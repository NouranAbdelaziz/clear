magic
tech sky130A
magscale 1 2
timestamp 1650625281
<< viali >>
rect 3985 20553 4019 20587
rect 7389 20553 7423 20587
rect 14289 20553 14323 20587
rect 15945 20553 15979 20587
rect 17969 20553 18003 20587
rect 19441 20553 19475 20587
rect 20545 20553 20579 20587
rect 2145 20485 2179 20519
rect 3249 20485 3283 20519
rect 4353 20485 4387 20519
rect 8493 20485 8527 20519
rect 9965 20485 9999 20519
rect 2605 20417 2639 20451
rect 3801 20417 3835 20451
rect 5273 20417 5307 20451
rect 5825 20417 5859 20451
rect 6653 20417 6687 20451
rect 6837 20417 6871 20451
rect 7205 20417 7239 20451
rect 7757 20417 7791 20451
rect 8309 20417 8343 20451
rect 9229 20417 9263 20451
rect 10517 20417 10551 20451
rect 11161 20417 11195 20451
rect 11529 20417 11563 20451
rect 12633 20417 12667 20451
rect 13553 20417 13587 20451
rect 14105 20417 14139 20451
rect 14657 20417 14691 20451
rect 15209 20417 15243 20451
rect 15761 20417 15795 20451
rect 16681 20417 16715 20451
rect 17233 20417 17267 20451
rect 17785 20417 17819 20451
rect 18337 20417 18371 20451
rect 19257 20417 19291 20451
rect 19809 20417 19843 20451
rect 20361 20417 20395 20451
rect 21097 20417 21131 20451
rect 1777 20349 1811 20383
rect 11805 20349 11839 20383
rect 2329 20281 2363 20315
rect 4537 20281 4571 20315
rect 4905 20281 4939 20315
rect 10977 20281 11011 20315
rect 14841 20281 14875 20315
rect 16865 20281 16899 20315
rect 18521 20281 18555 20315
rect 19993 20281 20027 20315
rect 2789 20213 2823 20247
rect 3341 20213 3375 20247
rect 5365 20213 5399 20247
rect 5917 20213 5951 20247
rect 7849 20213 7883 20247
rect 9321 20213 9355 20247
rect 10057 20213 10091 20247
rect 10609 20213 10643 20247
rect 13277 20213 13311 20247
rect 13737 20213 13771 20247
rect 15393 20213 15427 20247
rect 17417 20213 17451 20247
rect 21281 20213 21315 20247
rect 4353 20009 4387 20043
rect 4813 20009 4847 20043
rect 5273 20009 5307 20043
rect 6653 20009 6687 20043
rect 7573 20009 7607 20043
rect 14289 20009 14323 20043
rect 17233 20009 17267 20043
rect 17785 20009 17819 20043
rect 18337 20009 18371 20043
rect 18889 20009 18923 20043
rect 2421 19941 2455 19975
rect 5733 19941 5767 19975
rect 6193 19941 6227 19975
rect 7113 19941 7147 19975
rect 19441 19941 19475 19975
rect 10149 19873 10183 19907
rect 13001 19873 13035 19907
rect 14841 19873 14875 19907
rect 1685 19805 1719 19839
rect 2237 19805 2271 19839
rect 2697 19805 2731 19839
rect 3249 19805 3283 19839
rect 3893 19805 3927 19839
rect 4169 19805 4203 19839
rect 4629 19805 4663 19839
rect 5089 19805 5123 19839
rect 5549 19805 5583 19839
rect 6009 19805 6043 19839
rect 6469 19805 6503 19839
rect 6929 19805 6963 19839
rect 7389 19805 7423 19839
rect 7849 19805 7883 19839
rect 8309 19805 8343 19839
rect 9413 19805 9447 19839
rect 10977 19805 11011 19839
rect 11244 19805 11278 19839
rect 13185 19805 13219 19839
rect 14105 19805 14139 19839
rect 15025 19805 15059 19839
rect 16129 19805 16163 19839
rect 17049 19805 17083 19839
rect 17601 19805 17635 19839
rect 18153 19805 18187 19839
rect 18705 19805 18739 19839
rect 19257 19805 19291 19839
rect 20821 19805 20855 19839
rect 10333 19737 10367 19771
rect 15669 19737 15703 19771
rect 20177 19737 20211 19771
rect 21281 19737 21315 19771
rect 1777 19669 1811 19703
rect 2881 19669 2915 19703
rect 3341 19669 3375 19703
rect 8033 19669 8067 19703
rect 8493 19669 8527 19703
rect 9137 19669 9171 19703
rect 9597 19669 9631 19703
rect 10241 19669 10275 19703
rect 10701 19669 10735 19703
rect 12357 19669 12391 19703
rect 13093 19669 13127 19703
rect 13553 19669 13587 19703
rect 14933 19669 14967 19703
rect 15393 19669 15427 19703
rect 16773 19669 16807 19703
rect 3709 19465 3743 19499
rect 4169 19465 4203 19499
rect 6469 19465 6503 19499
rect 7113 19465 7147 19499
rect 7573 19465 7607 19499
rect 8493 19465 8527 19499
rect 8953 19465 8987 19499
rect 12725 19465 12759 19499
rect 16129 19465 16163 19499
rect 16865 19465 16899 19499
rect 17417 19465 17451 19499
rect 18521 19465 18555 19499
rect 19625 19465 19659 19499
rect 20177 19465 20211 19499
rect 21281 19465 21315 19499
rect 6009 19397 6043 19431
rect 3985 19329 4019 19363
rect 4445 19329 4479 19363
rect 4905 19329 4939 19363
rect 5549 19329 5583 19363
rect 6653 19329 6687 19363
rect 6929 19329 6963 19363
rect 7389 19329 7423 19363
rect 7849 19329 7883 19363
rect 8309 19329 8343 19363
rect 8769 19329 8803 19363
rect 9505 19329 9539 19363
rect 9781 19329 9815 19363
rect 10048 19329 10082 19363
rect 11897 19329 11931 19363
rect 11989 19329 12023 19363
rect 12541 19329 12575 19363
rect 13360 19329 13394 19363
rect 14749 19329 14783 19363
rect 15005 19329 15039 19363
rect 16681 19329 16715 19363
rect 17233 19329 17267 19363
rect 17785 19329 17819 19363
rect 18337 19329 18371 19363
rect 18889 19329 18923 19363
rect 19441 19329 19475 19363
rect 19993 19329 20027 19363
rect 20545 19329 20579 19363
rect 21097 19329 21131 19363
rect 2973 19261 3007 19295
rect 12081 19261 12115 19295
rect 13093 19261 13127 19295
rect 2237 19193 2271 19227
rect 3341 19193 3375 19227
rect 5089 19193 5123 19227
rect 8033 19193 8067 19227
rect 11161 19193 11195 19227
rect 17969 19193 18003 19227
rect 1501 19125 1535 19159
rect 1869 19125 1903 19159
rect 2605 19125 2639 19159
rect 4629 19125 4663 19159
rect 5365 19125 5399 19159
rect 9321 19125 9355 19159
rect 11529 19125 11563 19159
rect 14473 19125 14507 19159
rect 19073 19125 19107 19159
rect 20729 19125 20763 19159
rect 1593 18921 1627 18955
rect 2605 18921 2639 18955
rect 3065 18921 3099 18955
rect 4445 18921 4479 18955
rect 4905 18921 4939 18955
rect 5365 18921 5399 18955
rect 5825 18921 5859 18955
rect 6285 18921 6319 18955
rect 7205 18921 7239 18955
rect 8125 18921 8159 18955
rect 10609 18921 10643 18955
rect 13277 18921 13311 18955
rect 13737 18921 13771 18955
rect 18797 18921 18831 18955
rect 1961 18853 1995 18887
rect 4077 18785 4111 18819
rect 11529 18785 11563 18819
rect 14381 18785 14415 18819
rect 4721 18717 4755 18751
rect 5181 18717 5215 18751
rect 5641 18717 5675 18751
rect 6101 18717 6135 18751
rect 6561 18717 6595 18751
rect 7021 18717 7055 18751
rect 7481 18717 7515 18751
rect 7941 18717 7975 18751
rect 8585 18717 8619 18751
rect 9229 18717 9263 18751
rect 11897 18717 11931 18751
rect 13553 18717 13587 18751
rect 14473 18717 14507 18751
rect 15393 18717 15427 18751
rect 17233 18717 17267 18751
rect 18153 18717 18187 18751
rect 18613 18717 18647 18751
rect 19993 18717 20027 18751
rect 20453 18717 20487 18751
rect 21373 18717 21407 18751
rect 9496 18649 9530 18683
rect 11253 18649 11287 18683
rect 12164 18649 12198 18683
rect 15660 18649 15694 18683
rect 20729 18649 20763 18683
rect 2329 18581 2363 18615
rect 3433 18581 3467 18615
rect 6745 18581 6779 18615
rect 7665 18581 7699 18615
rect 8401 18581 8435 18615
rect 10885 18581 10919 18615
rect 11345 18581 11379 18615
rect 14565 18581 14599 18615
rect 14933 18581 14967 18615
rect 16773 18581 16807 18615
rect 17049 18581 17083 18615
rect 17509 18581 17543 18615
rect 19349 18581 19383 18615
rect 20269 18581 20303 18615
rect 2145 18377 2179 18411
rect 2881 18377 2915 18411
rect 6009 18377 6043 18411
rect 7297 18377 7331 18411
rect 8309 18377 8343 18411
rect 10517 18377 10551 18411
rect 11529 18377 11563 18411
rect 12909 18377 12943 18411
rect 13921 18377 13955 18411
rect 14749 18377 14783 18411
rect 15209 18377 15243 18411
rect 17141 18377 17175 18411
rect 19901 18377 19935 18411
rect 20729 18377 20763 18411
rect 1777 18309 1811 18343
rect 4353 18309 4387 18343
rect 5549 18309 5583 18343
rect 7941 18309 7975 18343
rect 9781 18309 9815 18343
rect 15117 18309 15151 18343
rect 19993 18309 20027 18343
rect 2513 18241 2547 18275
rect 5825 18241 5859 18275
rect 6653 18241 6687 18275
rect 7849 18241 7883 18275
rect 8953 18241 8987 18275
rect 11161 18241 11195 18275
rect 11897 18241 11931 18275
rect 12725 18241 12759 18275
rect 13277 18241 13311 18275
rect 14197 18241 14231 18275
rect 16037 18241 16071 18275
rect 18236 18241 18270 18275
rect 21373 18241 21407 18275
rect 3249 18173 3283 18207
rect 3985 18173 4019 18207
rect 7665 18173 7699 18207
rect 9597 18173 9631 18207
rect 9689 18173 9723 18207
rect 11989 18173 12023 18207
rect 12081 18173 12115 18207
rect 15301 18173 15335 18207
rect 16865 18173 16899 18207
rect 17049 18173 17083 18207
rect 17969 18173 18003 18207
rect 19717 18173 19751 18207
rect 3617 18105 3651 18139
rect 6837 18105 6871 18139
rect 16221 18105 16255 18139
rect 4721 18037 4755 18071
rect 5089 18037 5123 18071
rect 8677 18037 8711 18071
rect 9137 18037 9171 18071
rect 10149 18037 10183 18071
rect 14381 18037 14415 18071
rect 17509 18037 17543 18071
rect 19349 18037 19383 18071
rect 20361 18037 20395 18071
rect 5181 17833 5215 17867
rect 7113 17833 7147 17867
rect 10609 17833 10643 17867
rect 12265 17833 12299 17867
rect 12725 17833 12759 17867
rect 20269 17833 20303 17867
rect 4445 17765 4479 17799
rect 5549 17765 5583 17799
rect 17509 17765 17543 17799
rect 18521 17765 18555 17799
rect 19993 17765 20027 17799
rect 3065 17697 3099 17731
rect 11161 17697 11195 17731
rect 13185 17697 13219 17731
rect 13277 17697 13311 17731
rect 14289 17697 14323 17731
rect 17969 17697 18003 17731
rect 19349 17697 19383 17731
rect 20821 17697 20855 17731
rect 1685 17629 1719 17663
rect 3433 17629 3467 17663
rect 5825 17629 5859 17663
rect 6837 17629 6871 17663
rect 8493 17629 8527 17663
rect 8953 17629 8987 17663
rect 11621 17629 11655 17663
rect 12541 17629 12575 17663
rect 15761 17629 15795 17663
rect 16129 17629 16163 17663
rect 16396 17629 16430 17663
rect 18153 17629 18187 17663
rect 20637 17629 20671 17663
rect 8226 17561 8260 17595
rect 9220 17561 9254 17595
rect 11069 17561 11103 17595
rect 13369 17561 13403 17595
rect 15117 17561 15151 17595
rect 18797 17561 18831 17595
rect 19533 17561 19567 17595
rect 20729 17561 20763 17595
rect 1501 17493 1535 17527
rect 1961 17493 1995 17527
rect 2697 17493 2731 17527
rect 4077 17493 4111 17527
rect 4721 17493 4755 17527
rect 6193 17493 6227 17527
rect 10333 17493 10367 17527
rect 10977 17493 11011 17527
rect 13737 17493 13771 17527
rect 14381 17493 14415 17527
rect 14473 17493 14507 17527
rect 14841 17493 14875 17527
rect 18061 17493 18095 17527
rect 19625 17493 19659 17527
rect 21373 17493 21407 17527
rect 1409 17289 1443 17323
rect 1961 17289 1995 17323
rect 2237 17289 2271 17323
rect 3065 17289 3099 17323
rect 3433 17289 3467 17323
rect 3801 17289 3835 17323
rect 6009 17289 6043 17323
rect 9597 17289 9631 17323
rect 11161 17289 11195 17323
rect 14565 17289 14599 17323
rect 18429 17289 18463 17323
rect 2697 17221 2731 17255
rect 8116 17221 8150 17255
rect 9965 17221 9999 17255
rect 10057 17221 10091 17255
rect 16221 17221 16255 17255
rect 18972 17221 19006 17255
rect 4905 17153 4939 17187
rect 5273 17153 5307 17187
rect 6469 17153 6503 17187
rect 6929 17153 6963 17187
rect 7849 17153 7883 17187
rect 10977 17153 11011 17187
rect 11621 17153 11655 17187
rect 13176 17153 13210 17187
rect 15689 17153 15723 17187
rect 17316 17153 17350 17187
rect 18705 17153 18739 17187
rect 21005 17153 21039 17187
rect 4537 17085 4571 17119
rect 10241 17085 10275 17119
rect 12909 17085 12943 17119
rect 15945 17085 15979 17119
rect 17049 17085 17083 17119
rect 9229 17017 9263 17051
rect 14289 17017 14323 17051
rect 21281 17017 21315 17051
rect 4169 16949 4203 16983
rect 5641 16949 5675 16983
rect 6653 16949 6687 16983
rect 7573 16949 7607 16983
rect 10701 16949 10735 16983
rect 12265 16949 12299 16983
rect 12633 16949 12667 16983
rect 16681 16949 16715 16983
rect 20085 16949 20119 16983
rect 20361 16949 20395 16983
rect 1869 16745 1903 16779
rect 2513 16745 2547 16779
rect 4353 16745 4387 16779
rect 4997 16745 5031 16779
rect 5365 16745 5399 16779
rect 5641 16745 5675 16779
rect 6929 16745 6963 16779
rect 15945 16745 15979 16779
rect 19257 16745 19291 16779
rect 21281 16745 21315 16779
rect 13277 16677 13311 16711
rect 8309 16609 8343 16643
rect 9321 16609 9355 16643
rect 9505 16609 9539 16643
rect 10241 16609 10275 16643
rect 11897 16609 11931 16643
rect 14289 16609 14323 16643
rect 14381 16609 14415 16643
rect 15393 16609 15427 16643
rect 16773 16609 16807 16643
rect 17785 16609 17819 16643
rect 19809 16609 19843 16643
rect 20821 16609 20855 16643
rect 6193 16541 6227 16575
rect 12164 16541 12198 16575
rect 13553 16541 13587 16575
rect 15577 16541 15611 16575
rect 17693 16541 17727 16575
rect 18889 16541 18923 16575
rect 8064 16473 8098 16507
rect 10508 16473 10542 16507
rect 14473 16473 14507 16507
rect 16589 16473 16623 16507
rect 19717 16473 19751 16507
rect 20729 16473 20763 16507
rect 6009 16405 6043 16439
rect 6653 16405 6687 16439
rect 9597 16405 9631 16439
rect 9965 16405 9999 16439
rect 11621 16405 11655 16439
rect 13737 16405 13771 16439
rect 14841 16405 14875 16439
rect 15485 16405 15519 16439
rect 16221 16405 16255 16439
rect 16681 16405 16715 16439
rect 17233 16405 17267 16439
rect 17601 16405 17635 16439
rect 18245 16405 18279 16439
rect 19625 16405 19659 16439
rect 20269 16405 20303 16439
rect 20637 16405 20671 16439
rect 6745 16201 6779 16235
rect 9689 16201 9723 16235
rect 9781 16201 9815 16235
rect 10425 16201 10459 16235
rect 11713 16201 11747 16235
rect 12725 16201 12759 16235
rect 13369 16201 13403 16235
rect 19073 16201 19107 16235
rect 19625 16201 19659 16235
rect 20085 16201 20119 16235
rect 20361 16201 20395 16235
rect 12265 16133 12299 16167
rect 6837 16065 6871 16099
rect 7481 16065 7515 16099
rect 7737 16065 7771 16099
rect 10793 16065 10827 16099
rect 11529 16065 11563 16099
rect 12357 16065 12391 16099
rect 13461 16065 13495 16099
rect 14657 16065 14691 16099
rect 16057 16065 16091 16099
rect 17417 16065 17451 16099
rect 17960 16065 17994 16099
rect 19717 16065 19751 16099
rect 20729 16065 20763 16099
rect 5641 15997 5675 16031
rect 6653 15997 6687 16031
rect 9597 15997 9631 16031
rect 10885 15997 10919 16031
rect 10977 15997 11011 16031
rect 12081 15997 12115 16031
rect 13553 15997 13587 16031
rect 16313 15997 16347 16031
rect 17693 15997 17727 16031
rect 19441 15997 19475 16031
rect 20821 15997 20855 16031
rect 20913 15997 20947 16031
rect 5181 15929 5215 15963
rect 10149 15929 10183 15963
rect 4905 15861 4939 15895
rect 6009 15861 6043 15895
rect 7205 15861 7239 15895
rect 8861 15861 8895 15895
rect 13001 15861 13035 15895
rect 14013 15861 14047 15895
rect 14933 15861 14967 15895
rect 16773 15861 16807 15895
rect 6929 15657 6963 15691
rect 9965 15657 9999 15691
rect 10885 15657 10919 15691
rect 12449 15657 12483 15691
rect 14197 15657 14231 15691
rect 15393 15657 15427 15691
rect 17693 15657 17727 15691
rect 16957 15589 16991 15623
rect 18705 15589 18739 15623
rect 7941 15521 7975 15555
rect 8125 15521 8159 15555
rect 9137 15521 9171 15555
rect 13093 15521 13127 15555
rect 14749 15521 14783 15555
rect 18245 15521 18279 15555
rect 6469 15453 6503 15487
rect 7573 15453 7607 15487
rect 9321 15453 9355 15487
rect 10149 15453 10183 15487
rect 15209 15453 15243 15487
rect 18889 15453 18923 15487
rect 20370 15453 20404 15487
rect 20637 15453 20671 15487
rect 21097 15453 21131 15487
rect 6193 15385 6227 15419
rect 8217 15385 8251 15419
rect 12173 15385 12207 15419
rect 12817 15385 12851 15419
rect 13461 15385 13495 15419
rect 15669 15385 15703 15419
rect 5733 15317 5767 15351
rect 6653 15317 6687 15351
rect 8585 15317 8619 15351
rect 9229 15317 9263 15351
rect 9689 15317 9723 15351
rect 12909 15317 12943 15351
rect 14565 15317 14599 15351
rect 14657 15317 14691 15351
rect 18061 15317 18095 15351
rect 18153 15317 18187 15351
rect 19257 15317 19291 15351
rect 21281 15317 21315 15351
rect 9781 15113 9815 15147
rect 11529 15113 11563 15147
rect 13369 15113 13403 15147
rect 16313 15113 16347 15147
rect 18061 15113 18095 15147
rect 18797 15113 18831 15147
rect 20821 15113 20855 15147
rect 7481 15045 7515 15079
rect 8881 15045 8915 15079
rect 11897 15045 11931 15079
rect 14280 15045 14314 15079
rect 19708 15045 19742 15079
rect 6837 14977 6871 15011
rect 9137 14977 9171 15011
rect 10894 14977 10928 15011
rect 11161 14977 11195 15011
rect 12541 14977 12575 15011
rect 14013 14977 14047 15011
rect 15669 14977 15703 15011
rect 16681 14977 16715 15011
rect 17877 14977 17911 15011
rect 19441 14977 19475 15011
rect 21097 14977 21131 15011
rect 9505 14909 9539 14943
rect 11989 14909 12023 14943
rect 12081 14909 12115 14943
rect 13093 14909 13127 14943
rect 13277 14909 13311 14943
rect 18521 14909 18555 14943
rect 18705 14909 18739 14943
rect 6469 14773 6503 14807
rect 7021 14773 7055 14807
rect 7757 14773 7791 14807
rect 12725 14773 12759 14807
rect 13737 14773 13771 14807
rect 15393 14773 15427 14807
rect 17325 14773 17359 14807
rect 19165 14773 19199 14807
rect 21281 14773 21315 14807
rect 6745 14569 6779 14603
rect 16313 14569 16347 14603
rect 18797 14569 18831 14603
rect 19625 14569 19659 14603
rect 7481 14501 7515 14535
rect 11897 14501 11931 14535
rect 13737 14501 13771 14535
rect 7205 14433 7239 14467
rect 9689 14433 9723 14467
rect 9781 14433 9815 14467
rect 14197 14433 14231 14467
rect 14381 14433 14415 14467
rect 15577 14433 15611 14467
rect 15761 14433 15795 14467
rect 18153 14433 18187 14467
rect 20453 14433 20487 14467
rect 20637 14433 20671 14467
rect 7665 14365 7699 14399
rect 8574 14365 8608 14399
rect 9597 14365 9631 14399
rect 10241 14365 10275 14399
rect 12081 14365 12115 14399
rect 12357 14365 12391 14399
rect 16129 14365 16163 14399
rect 18613 14365 18647 14399
rect 19441 14365 19475 14399
rect 21005 14365 21039 14399
rect 10508 14297 10542 14331
rect 12624 14297 12658 14331
rect 17886 14297 17920 14331
rect 7941 14229 7975 14263
rect 9229 14229 9263 14263
rect 11621 14229 11655 14263
rect 14473 14229 14507 14263
rect 14841 14229 14875 14263
rect 15117 14229 15151 14263
rect 15485 14229 15519 14263
rect 16773 14229 16807 14263
rect 19993 14229 20027 14263
rect 20361 14229 20395 14263
rect 21189 14229 21223 14263
rect 8125 14025 8159 14059
rect 9505 14025 9539 14059
rect 11529 14025 11563 14059
rect 14381 14025 14415 14059
rect 14749 14025 14783 14059
rect 15393 14025 15427 14059
rect 18337 14025 18371 14059
rect 19349 14025 19383 14059
rect 20361 14025 20395 14059
rect 7849 13957 7883 13991
rect 10640 13957 10674 13991
rect 13737 13957 13771 13991
rect 19717 13957 19751 13991
rect 20729 13957 20763 13991
rect 8309 13889 8343 13923
rect 9229 13889 9263 13923
rect 10885 13889 10919 13923
rect 12642 13889 12676 13923
rect 12909 13889 12943 13923
rect 14289 13889 14323 13923
rect 16948 13889 16982 13923
rect 18705 13889 18739 13923
rect 19809 13889 19843 13923
rect 7389 13821 7423 13855
rect 8585 13821 8619 13855
rect 14105 13821 14139 13855
rect 15485 13821 15519 13855
rect 15577 13821 15611 13855
rect 16221 13821 16255 13855
rect 16681 13821 16715 13855
rect 18797 13821 18831 13855
rect 18889 13821 18923 13855
rect 19901 13821 19935 13855
rect 20821 13821 20855 13855
rect 21005 13821 21039 13855
rect 18061 13753 18095 13787
rect 13185 13685 13219 13719
rect 15025 13685 15059 13719
rect 7757 13481 7791 13515
rect 10885 13481 10919 13515
rect 12449 13481 12483 13515
rect 21281 13481 21315 13515
rect 9781 13413 9815 13447
rect 13461 13413 13495 13447
rect 15301 13413 15335 13447
rect 18797 13413 18831 13447
rect 8125 13345 8159 13379
rect 9229 13345 9263 13379
rect 12909 13345 12943 13379
rect 13001 13345 13035 13379
rect 14657 13345 14691 13379
rect 14841 13345 14875 13379
rect 19901 13345 19935 13379
rect 20453 13345 20487 13379
rect 8585 13277 8619 13311
rect 9413 13277 9447 13311
rect 12173 13277 12207 13311
rect 13645 13277 13679 13311
rect 14289 13277 14323 13311
rect 14933 13277 14967 13311
rect 17693 13277 17727 13311
rect 18613 13277 18647 13311
rect 19717 13277 19751 13311
rect 20545 13277 20579 13311
rect 9321 13209 9355 13243
rect 15669 13209 15703 13243
rect 17417 13209 17451 13243
rect 19625 13209 19659 13243
rect 7297 13141 7331 13175
rect 8401 13141 8435 13175
rect 10149 13141 10183 13175
rect 12817 13141 12851 13175
rect 14105 13141 14139 13175
rect 18337 13141 18371 13175
rect 19257 13141 19291 13175
rect 20637 13141 20671 13175
rect 21005 13141 21039 13175
rect 8033 12937 8067 12971
rect 8585 12937 8619 12971
rect 10333 12937 10367 12971
rect 10977 12937 11011 12971
rect 14565 12937 14599 12971
rect 15577 12937 15611 12971
rect 15945 12937 15979 12971
rect 18613 12937 18647 12971
rect 20269 12937 20303 12971
rect 20637 12937 20671 12971
rect 21373 12937 21407 12971
rect 14013 12869 14047 12903
rect 14933 12869 14967 12903
rect 16037 12869 16071 12903
rect 8953 12801 8987 12835
rect 9209 12801 9243 12835
rect 11805 12801 11839 12835
rect 12725 12801 12759 12835
rect 13369 12801 13403 12835
rect 17805 12801 17839 12835
rect 18061 12801 18095 12835
rect 19726 12801 19760 12835
rect 19993 12801 20027 12835
rect 12817 12733 12851 12767
rect 13001 12733 13035 12767
rect 15025 12733 15059 12767
rect 15117 12733 15151 12767
rect 16221 12733 16255 12767
rect 20729 12733 20763 12767
rect 20913 12733 20947 12767
rect 12357 12665 12391 12699
rect 11621 12597 11655 12631
rect 16681 12597 16715 12631
rect 8953 12393 8987 12427
rect 10609 12393 10643 12427
rect 12081 12393 12115 12427
rect 15761 12393 15795 12427
rect 17693 12393 17727 12427
rect 19257 12393 19291 12427
rect 21189 12393 21223 12427
rect 7665 12325 7699 12359
rect 13737 12325 13771 12359
rect 10333 12257 10367 12291
rect 11529 12257 11563 12291
rect 16313 12257 16347 12291
rect 17141 12257 17175 12291
rect 18613 12257 18647 12291
rect 19809 12257 19843 12291
rect 7481 12189 7515 12223
rect 8585 12189 8619 12223
rect 10793 12189 10827 12223
rect 12357 12189 12391 12223
rect 15218 12189 15252 12223
rect 15485 12189 15519 12223
rect 18337 12189 18371 12223
rect 19441 12189 19475 12223
rect 10066 12121 10100 12155
rect 11621 12121 11655 12155
rect 12602 12121 12636 12155
rect 16129 12121 16163 12155
rect 17233 12121 17267 12155
rect 20076 12121 20110 12155
rect 7941 12053 7975 12087
rect 11713 12053 11747 12087
rect 14105 12053 14139 12087
rect 16221 12053 16255 12087
rect 17325 12053 17359 12087
rect 17969 12053 18003 12087
rect 18429 12053 18463 12087
rect 6929 11849 6963 11883
rect 7849 11849 7883 11883
rect 10425 11849 10459 11883
rect 13829 11849 13863 11883
rect 18337 11849 18371 11883
rect 18797 11849 18831 11883
rect 19717 11849 19751 11883
rect 20361 11849 20395 11883
rect 8125 11781 8159 11815
rect 9290 11781 9324 11815
rect 15853 11781 15887 11815
rect 16948 11781 16982 11815
rect 18705 11781 18739 11815
rect 20821 11781 20855 11815
rect 7665 11713 7699 11747
rect 8769 11713 8803 11747
rect 9045 11713 9079 11747
rect 11713 11713 11747 11747
rect 11980 11713 12014 11747
rect 16129 11713 16163 11747
rect 20729 11713 20763 11747
rect 10977 11645 11011 11679
rect 16681 11645 16715 11679
rect 18889 11645 18923 11679
rect 19809 11645 19843 11679
rect 19993 11645 20027 11679
rect 20913 11645 20947 11679
rect 7297 11577 7331 11611
rect 13093 11509 13127 11543
rect 14565 11509 14599 11543
rect 16313 11509 16347 11543
rect 18061 11509 18095 11543
rect 19349 11509 19383 11543
rect 6837 11305 6871 11339
rect 7665 11305 7699 11339
rect 8585 11305 8619 11339
rect 11437 11305 11471 11339
rect 13185 11305 13219 11339
rect 14841 11305 14875 11339
rect 16497 11305 16531 11339
rect 21189 11305 21223 11339
rect 9321 11237 9355 11271
rect 14565 11237 14599 11271
rect 20729 11237 20763 11271
rect 7113 11169 7147 11203
rect 11989 11169 12023 11203
rect 12633 11169 12667 11203
rect 13461 11169 13495 11203
rect 17049 11169 17083 11203
rect 18061 11169 18095 11203
rect 18521 11169 18555 11203
rect 7481 11101 7515 11135
rect 7941 11101 7975 11135
rect 9505 11101 9539 11135
rect 11161 11101 11195 11135
rect 11897 11101 11931 11135
rect 14381 11101 14415 11135
rect 15954 11101 15988 11135
rect 16221 11101 16255 11135
rect 19349 11101 19383 11135
rect 9045 11033 9079 11067
rect 10894 11033 10928 11067
rect 16957 11033 16991 11067
rect 19594 11033 19628 11067
rect 21281 11033 21315 11067
rect 9781 10965 9815 10999
rect 11805 10965 11839 10999
rect 12725 10965 12759 10999
rect 12817 10965 12851 10999
rect 16865 10965 16899 10999
rect 17509 10965 17543 10999
rect 17877 10965 17911 10999
rect 17969 10965 18003 10999
rect 8217 10761 8251 10795
rect 9137 10761 9171 10795
rect 9781 10761 9815 10795
rect 10149 10761 10183 10795
rect 10793 10761 10827 10795
rect 11161 10761 11195 10795
rect 13093 10761 13127 10795
rect 14565 10761 14599 10795
rect 15209 10761 15243 10795
rect 15669 10761 15703 10795
rect 18337 10761 18371 10795
rect 6561 10693 6595 10727
rect 11980 10693 12014 10727
rect 14105 10693 14139 10727
rect 20260 10693 20294 10727
rect 7573 10625 7607 10659
rect 8493 10625 8527 10659
rect 14197 10625 14231 10659
rect 15301 10625 15335 10659
rect 15945 10625 15979 10659
rect 17805 10625 17839 10659
rect 19461 10625 19495 10659
rect 19717 10625 19751 10659
rect 19993 10625 20027 10659
rect 9597 10557 9631 10591
rect 9689 10557 9723 10591
rect 10609 10557 10643 10591
rect 10701 10557 10735 10591
rect 11713 10557 11747 10591
rect 13553 10557 13587 10591
rect 13921 10557 13955 10591
rect 15117 10557 15151 10591
rect 18061 10557 18095 10591
rect 7205 10489 7239 10523
rect 7757 10489 7791 10523
rect 6929 10421 6963 10455
rect 16129 10421 16163 10455
rect 16681 10421 16715 10455
rect 21373 10421 21407 10455
rect 7113 10217 7147 10251
rect 8953 10217 8987 10251
rect 12633 10217 12667 10251
rect 14105 10217 14139 10251
rect 16865 10217 16899 10251
rect 20637 10217 20671 10251
rect 10149 10149 10183 10183
rect 11989 10149 12023 10183
rect 6837 10081 6871 10115
rect 9505 10081 9539 10115
rect 13185 10081 13219 10115
rect 14657 10081 14691 10115
rect 15669 10081 15703 10115
rect 19257 10081 19291 10115
rect 7481 10013 7515 10047
rect 8585 10013 8619 10047
rect 9137 10013 9171 10047
rect 10609 10013 10643 10047
rect 15485 10013 15519 10047
rect 17978 10013 18012 10047
rect 18245 10013 18279 10047
rect 18613 10013 18647 10047
rect 19513 10013 19547 10047
rect 20913 10013 20947 10047
rect 7941 9945 7975 9979
rect 9689 9945 9723 9979
rect 10854 9945 10888 9979
rect 12357 9945 12391 9979
rect 13093 9945 13127 9979
rect 16589 9945 16623 9979
rect 6377 9877 6411 9911
rect 7665 9877 7699 9911
rect 9781 9877 9815 9911
rect 13001 9877 13035 9911
rect 13737 9877 13771 9911
rect 14473 9877 14507 9911
rect 14565 9877 14599 9911
rect 15117 9877 15151 9911
rect 15577 9877 15611 9911
rect 18797 9877 18831 9911
rect 21097 9877 21131 9911
rect 7481 9673 7515 9707
rect 13369 9673 13403 9707
rect 15945 9673 15979 9707
rect 7757 9605 7791 9639
rect 8677 9605 8711 9639
rect 10710 9605 10744 9639
rect 12173 9605 12207 9639
rect 12449 9605 12483 9639
rect 17233 9605 17267 9639
rect 18398 9605 18432 9639
rect 7113 9537 7147 9571
rect 8401 9537 8435 9571
rect 9321 9537 9355 9571
rect 11529 9537 11563 9571
rect 13093 9537 13127 9571
rect 13737 9537 13771 9571
rect 14749 9537 14783 9571
rect 16037 9537 16071 9571
rect 17141 9537 17175 9571
rect 17785 9537 17819 9571
rect 20177 9537 20211 9571
rect 21097 9537 21131 9571
rect 10977 9469 11011 9503
rect 13829 9469 13863 9503
rect 14013 9469 14047 9503
rect 14841 9469 14875 9503
rect 14933 9469 14967 9503
rect 16129 9469 16163 9503
rect 17325 9469 17359 9503
rect 18153 9469 18187 9503
rect 20269 9469 20303 9503
rect 20453 9469 20487 9503
rect 19533 9401 19567 9435
rect 19809 9401 19843 9435
rect 6653 9333 6687 9367
rect 9597 9333 9631 9367
rect 14381 9333 14415 9367
rect 15577 9333 15611 9367
rect 16773 9333 16807 9367
rect 21281 9333 21315 9367
rect 10425 9129 10459 9163
rect 11897 9129 11931 9163
rect 16037 9129 16071 9163
rect 20269 9129 20303 9163
rect 21281 9129 21315 9163
rect 7297 9061 7331 9095
rect 8125 9061 8159 9095
rect 6929 8993 6963 9027
rect 9505 8993 9539 9027
rect 10977 8993 11011 9027
rect 12173 8993 12207 9027
rect 16497 8993 16531 9027
rect 16589 8993 16623 9027
rect 17601 8993 17635 9027
rect 18245 8993 18279 9027
rect 19809 8993 19843 9027
rect 20821 8993 20855 9027
rect 7941 8925 7975 8959
rect 9689 8925 9723 8959
rect 11713 8925 11747 8959
rect 15772 8925 15806 8959
rect 17417 8925 17451 8959
rect 18429 8925 18463 8959
rect 20637 8925 20671 8959
rect 6561 8857 6595 8891
rect 9137 8857 9171 8891
rect 9781 8857 9815 8891
rect 10793 8857 10827 8891
rect 12440 8857 12474 8891
rect 15494 8857 15528 8891
rect 17509 8857 17543 8891
rect 18337 8857 18371 8891
rect 20729 8857 20763 8891
rect 7573 8789 7607 8823
rect 8585 8789 8619 8823
rect 10149 8789 10183 8823
rect 10885 8789 10919 8823
rect 13553 8789 13587 8823
rect 14381 8789 14415 8823
rect 16405 8789 16439 8823
rect 17049 8789 17083 8823
rect 18797 8789 18831 8823
rect 19257 8789 19291 8823
rect 19625 8789 19659 8823
rect 19717 8789 19751 8823
rect 7481 8585 7515 8619
rect 8309 8585 8343 8619
rect 9229 8585 9263 8619
rect 17049 8585 17083 8619
rect 18061 8585 18095 8619
rect 18429 8585 18463 8619
rect 21189 8585 21223 8619
rect 17417 8517 17451 8551
rect 20076 8517 20110 8551
rect 7113 8449 7147 8483
rect 8125 8449 8159 8483
rect 8769 8449 8803 8483
rect 10618 8449 10652 8483
rect 11897 8449 11931 8483
rect 12541 8449 12575 8483
rect 12797 8449 12831 8483
rect 14381 8449 14415 8483
rect 15189 8449 15223 8483
rect 16773 8449 16807 8483
rect 17509 8449 17543 8483
rect 18521 8449 18555 8483
rect 19073 8449 19107 8483
rect 19809 8449 19843 8483
rect 7757 8381 7791 8415
rect 10885 8381 10919 8415
rect 11621 8381 11655 8415
rect 11805 8381 11839 8415
rect 14933 8381 14967 8415
rect 17601 8381 17635 8415
rect 18613 8381 18647 8415
rect 8585 8313 8619 8347
rect 9505 8313 9539 8347
rect 12265 8313 12299 8347
rect 13921 8313 13955 8347
rect 16313 8313 16347 8347
rect 6745 8245 6779 8279
rect 14197 8245 14231 8279
rect 19257 8245 19291 8279
rect 9505 8041 9539 8075
rect 13645 8041 13679 8075
rect 14841 8041 14875 8075
rect 16957 8041 16991 8075
rect 18889 8041 18923 8075
rect 21281 8041 21315 8075
rect 19349 7973 19383 8007
rect 7297 7905 7331 7939
rect 8585 7905 8619 7939
rect 13001 7905 13035 7939
rect 14289 7905 14323 7939
rect 14381 7905 14415 7939
rect 18337 7905 18371 7939
rect 6561 7837 6595 7871
rect 7573 7837 7607 7871
rect 10149 7837 10183 7871
rect 13461 7837 13495 7871
rect 15117 7837 15151 7871
rect 18705 7837 18739 7871
rect 19625 7837 19659 7871
rect 19881 7837 19915 7871
rect 6193 7769 6227 7803
rect 10425 7769 10459 7803
rect 12173 7769 12207 7803
rect 12817 7769 12851 7803
rect 14473 7769 14507 7803
rect 15669 7769 15703 7803
rect 6929 7701 6963 7735
rect 8217 7701 8251 7735
rect 9229 7701 9263 7735
rect 12449 7701 12483 7735
rect 12909 7701 12943 7735
rect 15301 7701 15335 7735
rect 17693 7701 17727 7735
rect 18061 7701 18095 7735
rect 18153 7701 18187 7735
rect 21005 7701 21039 7735
rect 6561 7497 6595 7531
rect 10333 7497 10367 7531
rect 10701 7497 10735 7531
rect 11161 7497 11195 7531
rect 11529 7497 11563 7531
rect 13921 7497 13955 7531
rect 14013 7497 14047 7531
rect 14565 7497 14599 7531
rect 17141 7497 17175 7531
rect 18797 7497 18831 7531
rect 19257 7497 19291 7531
rect 20177 7497 20211 7531
rect 9198 7429 9232 7463
rect 20269 7429 20303 7463
rect 21189 7429 21223 7463
rect 8410 7361 8444 7395
rect 8677 7361 8711 7395
rect 8953 7361 8987 7395
rect 10977 7361 11011 7395
rect 12173 7361 12207 7395
rect 12817 7361 12851 7395
rect 16057 7361 16091 7395
rect 16313 7361 16347 7395
rect 16865 7361 16899 7395
rect 18265 7361 18299 7395
rect 18521 7361 18555 7395
rect 19165 7361 19199 7395
rect 12909 7293 12943 7327
rect 13001 7293 13035 7327
rect 14197 7293 14231 7327
rect 19349 7293 19383 7327
rect 20361 7293 20395 7327
rect 6929 7225 6963 7259
rect 14933 7225 14967 7259
rect 21373 7225 21407 7259
rect 5273 7157 5307 7191
rect 5549 7157 5583 7191
rect 5917 7157 5951 7191
rect 7297 7157 7331 7191
rect 12449 7157 12483 7191
rect 13553 7157 13587 7191
rect 16681 7157 16715 7191
rect 19809 7157 19843 7191
rect 5181 6953 5215 6987
rect 13001 6953 13035 6987
rect 15577 6953 15611 6987
rect 8585 6885 8619 6919
rect 9045 6885 9079 6919
rect 11345 6885 11379 6919
rect 17601 6885 17635 6919
rect 4813 6817 4847 6851
rect 5549 6817 5583 6851
rect 6929 6817 6963 6851
rect 8033 6817 8067 6851
rect 9413 6817 9447 6851
rect 10885 6817 10919 6851
rect 13645 6817 13679 6851
rect 14749 6817 14783 6851
rect 16129 6817 16163 6851
rect 17049 6817 17083 6851
rect 17141 6817 17175 6851
rect 18153 6817 18187 6851
rect 6193 6749 6227 6783
rect 7573 6749 7607 6783
rect 10701 6749 10735 6783
rect 12725 6749 12759 6783
rect 13369 6749 13403 6783
rect 13461 6749 13495 6783
rect 14289 6749 14323 6783
rect 15945 6749 15979 6783
rect 18613 6749 18647 6783
rect 19441 6749 19475 6783
rect 21097 6749 21131 6783
rect 5917 6681 5951 6715
rect 9597 6681 9631 6715
rect 10793 6681 10827 6715
rect 12480 6681 12514 6715
rect 14933 6681 14967 6715
rect 16037 6681 16071 6715
rect 17969 6681 18003 6715
rect 18061 6681 18095 6715
rect 19708 6681 19742 6715
rect 1409 6613 1443 6647
rect 4169 6613 4203 6647
rect 6653 6613 6687 6647
rect 8125 6613 8159 6647
rect 8217 6613 8251 6647
rect 9689 6613 9723 6647
rect 10057 6613 10091 6647
rect 10333 6613 10367 6647
rect 14841 6613 14875 6647
rect 15301 6613 15335 6647
rect 16589 6613 16623 6647
rect 16957 6613 16991 6647
rect 18797 6613 18831 6647
rect 20821 6613 20855 6647
rect 21281 6613 21315 6647
rect 3157 6409 3191 6443
rect 3893 6409 3927 6443
rect 4537 6409 4571 6443
rect 6009 6409 6043 6443
rect 7021 6409 7055 6443
rect 9137 6409 9171 6443
rect 10333 6409 10367 6443
rect 10701 6409 10735 6443
rect 11529 6409 11563 6443
rect 11897 6409 11931 6443
rect 11989 6409 12023 6443
rect 13093 6409 13127 6443
rect 20545 6409 20579 6443
rect 20913 6409 20947 6443
rect 8024 6341 8058 6375
rect 1409 6273 1443 6307
rect 1869 6273 1903 6307
rect 5641 6273 5675 6307
rect 7297 6273 7331 6307
rect 10057 6273 10091 6307
rect 12541 6273 12575 6307
rect 14217 6273 14251 6307
rect 14933 6273 14967 6307
rect 15200 6273 15234 6307
rect 16681 6273 16715 6307
rect 17141 6273 17175 6307
rect 17408 6273 17442 6307
rect 18797 6273 18831 6307
rect 19064 6273 19098 6307
rect 6561 6205 6595 6239
rect 7757 6205 7791 6239
rect 10793 6205 10827 6239
rect 10885 6205 10919 6239
rect 12081 6205 12115 6239
rect 14473 6205 14507 6239
rect 21005 6205 21039 6239
rect 21189 6205 21223 6239
rect 1593 6069 1627 6103
rect 2237 6069 2271 6103
rect 3433 6069 3467 6103
rect 4905 6069 4939 6103
rect 5273 6069 5307 6103
rect 7481 6069 7515 6103
rect 9413 6069 9447 6103
rect 12725 6069 12759 6103
rect 16313 6069 16347 6103
rect 16865 6069 16899 6103
rect 18521 6069 18555 6103
rect 20177 6069 20211 6103
rect 3433 5865 3467 5899
rect 6469 5865 6503 5899
rect 9045 5865 9079 5899
rect 10701 5865 10735 5899
rect 15301 5865 15335 5899
rect 17141 5865 17175 5899
rect 17877 5865 17911 5899
rect 20637 5865 20671 5899
rect 5917 5797 5951 5831
rect 6745 5729 6779 5763
rect 9689 5729 9723 5763
rect 12725 5729 12759 5763
rect 12817 5729 12851 5763
rect 14381 5729 14415 5763
rect 18337 5729 18371 5763
rect 18429 5729 18463 5763
rect 4445 5661 4479 5695
rect 5549 5661 5583 5695
rect 6285 5661 6319 5695
rect 7001 5661 7035 5695
rect 12173 5661 12207 5695
rect 13737 5661 13771 5695
rect 14565 5661 14599 5695
rect 19257 5661 19291 5695
rect 20913 5661 20947 5695
rect 21097 5661 21131 5695
rect 3065 5593 3099 5627
rect 4905 5593 4939 5627
rect 9413 5593 9447 5627
rect 9505 5593 9539 5627
rect 15669 5593 15703 5627
rect 19502 5593 19536 5627
rect 1501 5525 1535 5559
rect 1961 5525 1995 5559
rect 2329 5525 2363 5559
rect 2697 5525 2731 5559
rect 4169 5525 4203 5559
rect 5273 5525 5307 5559
rect 8125 5525 8159 5559
rect 8585 5525 8619 5559
rect 10149 5525 10183 5559
rect 12909 5525 12943 5559
rect 13277 5525 13311 5559
rect 13553 5525 13587 5559
rect 14657 5525 14691 5559
rect 15025 5525 15059 5559
rect 18245 5525 18279 5559
rect 1869 5321 1903 5355
rect 4077 5321 4111 5355
rect 7665 5321 7699 5355
rect 8401 5321 8435 5355
rect 14565 5321 14599 5355
rect 19441 5321 19475 5355
rect 19809 5321 19843 5355
rect 20637 5321 20671 5355
rect 4445 5253 4479 5287
rect 5549 5253 5583 5287
rect 9321 5253 9355 5287
rect 10701 5253 10735 5287
rect 15086 5253 15120 5287
rect 17202 5253 17236 5287
rect 2973 5185 3007 5219
rect 4813 5185 4847 5219
rect 6009 5185 6043 5219
rect 6561 5185 6595 5219
rect 7021 5185 7055 5219
rect 7481 5185 7515 5219
rect 7941 5185 7975 5219
rect 9045 5185 9079 5219
rect 9965 5185 9999 5219
rect 10609 5185 10643 5219
rect 11529 5185 11563 5219
rect 11785 5185 11819 5219
rect 13185 5185 13219 5219
rect 13441 5185 13475 5219
rect 16957 5185 16991 5219
rect 18613 5185 18647 5219
rect 21005 5185 21039 5219
rect 1501 5117 1535 5151
rect 10885 5117 10919 5151
rect 14841 5117 14875 5151
rect 19901 5117 19935 5151
rect 19993 5117 20027 5151
rect 21097 5117 21131 5151
rect 21281 5117 21315 5151
rect 2605 5049 2639 5083
rect 3709 5049 3743 5083
rect 6745 5049 6779 5083
rect 10241 5049 10275 5083
rect 18797 5049 18831 5083
rect 2237 4981 2271 5015
rect 3341 4981 3375 5015
rect 5089 4981 5123 5015
rect 5825 4981 5859 5015
rect 7205 4981 7239 5015
rect 8125 4981 8159 5015
rect 12909 4981 12943 5015
rect 16221 4981 16255 5015
rect 18337 4981 18371 5015
rect 4537 4777 4571 4811
rect 5365 4777 5399 4811
rect 5825 4777 5859 4811
rect 6745 4777 6779 4811
rect 7205 4777 7239 4811
rect 17877 4777 17911 4811
rect 3433 4709 3467 4743
rect 6285 4709 6319 4743
rect 13645 4709 13679 4743
rect 14289 4709 14323 4743
rect 16589 4709 16623 4743
rect 16865 4709 16899 4743
rect 4169 4641 4203 4675
rect 7665 4641 7699 4675
rect 9321 4641 9355 4675
rect 12357 4641 12391 4675
rect 13185 4641 13219 4675
rect 15025 4641 15059 4675
rect 15945 4641 15979 4675
rect 17417 4641 17451 4675
rect 18521 4641 18555 4675
rect 19257 4641 19291 4675
rect 2697 4573 2731 4607
rect 5181 4573 5215 4607
rect 5641 4573 5675 4607
rect 6101 4573 6135 4607
rect 6561 4573 6595 4607
rect 7021 4573 7055 4607
rect 8585 4573 8619 4607
rect 12090 4573 12124 4607
rect 13001 4573 13035 4607
rect 14105 4573 14139 4607
rect 15117 4573 15151 4607
rect 20913 4573 20947 4607
rect 7941 4505 7975 4539
rect 9588 4505 9622 4539
rect 16221 4505 16255 4539
rect 17325 4505 17359 4539
rect 19524 4505 19558 4539
rect 1593 4437 1627 4471
rect 1961 4437 1995 4471
rect 2329 4437 2363 4471
rect 2973 4437 3007 4471
rect 4905 4437 4939 4471
rect 9045 4437 9079 4471
rect 10701 4437 10735 4471
rect 10977 4437 11011 4471
rect 12633 4437 12667 4471
rect 13093 4437 13127 4471
rect 15209 4437 15243 4471
rect 15577 4437 15611 4471
rect 16129 4437 16163 4471
rect 17233 4437 17267 4471
rect 18245 4437 18279 4471
rect 18337 4437 18371 4471
rect 20637 4437 20671 4471
rect 21097 4437 21131 4471
rect 2605 4233 2639 4267
rect 11989 4233 12023 4267
rect 12633 4233 12667 4267
rect 14197 4233 14231 4267
rect 15209 4233 15243 4267
rect 15577 4233 15611 4267
rect 17509 4233 17543 4267
rect 17969 4233 18003 4267
rect 3709 4165 3743 4199
rect 6837 4165 6871 4199
rect 8953 4165 8987 4199
rect 9137 4165 9171 4199
rect 13001 4165 13035 4199
rect 16037 4165 16071 4199
rect 17601 4165 17635 4199
rect 20821 4165 20855 4199
rect 1501 4097 1535 4131
rect 2237 4097 2271 4131
rect 3985 4097 4019 4131
rect 4445 4097 4479 4131
rect 5081 4097 5115 4131
rect 5365 4097 5399 4131
rect 7297 4097 7331 4131
rect 7573 4097 7607 4131
rect 8217 4097 8251 4131
rect 8493 4097 8527 4131
rect 9505 4097 9539 4131
rect 10149 4097 10183 4131
rect 10793 4097 10827 4131
rect 10885 4097 10919 4131
rect 12081 4097 12115 4131
rect 16681 4097 16715 4131
rect 18245 4097 18279 4131
rect 18501 4097 18535 4131
rect 19901 4097 19935 4131
rect 3341 4029 3375 4063
rect 6009 4029 6043 4063
rect 10977 4029 11011 4063
rect 12173 4029 12207 4063
rect 13093 4029 13127 4063
rect 13185 4029 13219 4063
rect 14289 4029 14323 4063
rect 14473 4029 14507 4063
rect 15025 4029 15059 4063
rect 15117 4029 15151 4063
rect 15853 4029 15887 4063
rect 17325 4029 17359 4063
rect 20913 4029 20947 4063
rect 21097 4029 21131 4063
rect 4629 3961 4663 3995
rect 10425 3961 10459 3995
rect 20453 3961 20487 3995
rect 1869 3893 1903 3927
rect 2973 3893 3007 3927
rect 4169 3893 4203 3927
rect 4905 3893 4939 3927
rect 5549 3893 5583 3927
rect 7113 3893 7147 3927
rect 7757 3893 7791 3927
rect 8033 3893 8067 3927
rect 8677 3893 8711 3927
rect 11621 3893 11655 3927
rect 13829 3893 13863 3927
rect 16865 3893 16899 3927
rect 19625 3893 19659 3927
rect 20085 3893 20119 3927
rect 6469 3689 6503 3723
rect 7849 3689 7883 3723
rect 10793 3689 10827 3723
rect 15485 3689 15519 3723
rect 18797 3689 18831 3723
rect 21189 3689 21223 3723
rect 2605 3621 2639 3655
rect 3433 3621 3467 3655
rect 6009 3621 6043 3655
rect 6929 3621 6963 3655
rect 8493 3621 8527 3655
rect 10241 3553 10275 3587
rect 10333 3553 10367 3587
rect 13093 3553 13127 3587
rect 18153 3553 18187 3587
rect 19993 3553 20027 3587
rect 20637 3553 20671 3587
rect 1869 3485 1903 3519
rect 3249 3485 3283 3519
rect 3985 3485 4019 3519
rect 4629 3485 4663 3519
rect 4905 3485 4939 3519
rect 5365 3485 5399 3519
rect 5825 3485 5859 3519
rect 6285 3485 6319 3519
rect 6745 3485 6779 3519
rect 7205 3485 7239 3519
rect 8309 3485 8343 3519
rect 9781 3485 9815 3519
rect 10425 3485 10459 3519
rect 11069 3485 11103 3519
rect 11336 3485 11370 3519
rect 13369 3485 13403 3519
rect 14105 3485 14139 3519
rect 15945 3485 15979 3519
rect 17969 3485 18003 3519
rect 18613 3485 18647 3519
rect 19809 3485 19843 3519
rect 20821 3485 20855 3519
rect 2237 3417 2271 3451
rect 2973 3417 3007 3451
rect 7757 3417 7791 3451
rect 14350 3417 14384 3451
rect 16212 3417 16246 3451
rect 19901 3417 19935 3451
rect 20729 3417 20763 3451
rect 1501 3349 1535 3383
rect 4169 3349 4203 3383
rect 4445 3349 4479 3383
rect 5089 3349 5123 3383
rect 5549 3349 5583 3383
rect 7389 3349 7423 3383
rect 9137 3349 9171 3383
rect 12449 3349 12483 3383
rect 13277 3349 13311 3383
rect 13737 3349 13771 3383
rect 17325 3349 17359 3383
rect 17601 3349 17635 3383
rect 18061 3349 18095 3383
rect 19441 3349 19475 3383
rect 3433 3145 3467 3179
rect 5089 3145 5123 3179
rect 8309 3145 8343 3179
rect 11621 3145 11655 3179
rect 14289 3145 14323 3179
rect 20269 3145 20303 3179
rect 3801 3077 3835 3111
rect 10517 3077 10551 3111
rect 12909 3077 12943 3111
rect 14902 3077 14936 3111
rect 17294 3077 17328 3111
rect 1409 3009 1443 3043
rect 1869 3009 1903 3043
rect 2329 3009 2363 3043
rect 2789 3009 2823 3043
rect 3249 3009 3283 3043
rect 3985 3009 4019 3043
rect 4445 3009 4479 3043
rect 4905 3009 4939 3043
rect 5365 3009 5399 3043
rect 5825 3009 5859 3043
rect 6653 3009 6687 3043
rect 7297 3009 7331 3043
rect 7573 3009 7607 3043
rect 7757 3009 7791 3043
rect 8125 3009 8159 3043
rect 9321 3009 9355 3043
rect 9597 3009 9631 3043
rect 10241 3009 10275 3043
rect 11161 3009 11195 3043
rect 12265 3009 12299 3043
rect 12817 3009 12851 3043
rect 13921 3009 13955 3043
rect 14657 3009 14691 3043
rect 17049 3009 17083 3043
rect 18705 3009 18739 3043
rect 19901 3009 19935 3043
rect 20821 3009 20855 3043
rect 6837 2941 6871 2975
rect 12633 2941 12667 2975
rect 13645 2941 13679 2975
rect 13829 2941 13863 2975
rect 16773 2941 16807 2975
rect 19625 2941 19659 2975
rect 19809 2941 19843 2975
rect 20545 2941 20579 2975
rect 6009 2873 6043 2907
rect 16037 2873 16071 2907
rect 18889 2873 18923 2907
rect 1593 2805 1627 2839
rect 2053 2805 2087 2839
rect 2513 2805 2547 2839
rect 2973 2805 3007 2839
rect 4629 2805 4663 2839
rect 5549 2805 5583 2839
rect 7113 2805 7147 2839
rect 8677 2805 8711 2839
rect 13277 2805 13311 2839
rect 18429 2805 18463 2839
rect 3341 2601 3375 2635
rect 4813 2601 4847 2635
rect 5917 2601 5951 2635
rect 7297 2601 7331 2635
rect 9413 2601 9447 2635
rect 15577 2601 15611 2635
rect 17417 2601 17451 2635
rect 2789 2533 2823 2567
rect 4537 2533 4571 2567
rect 6653 2533 6687 2567
rect 8493 2533 8527 2567
rect 11713 2533 11747 2567
rect 19671 2533 19705 2567
rect 1409 2465 1443 2499
rect 1685 2465 1719 2499
rect 10149 2465 10183 2499
rect 13093 2465 13127 2499
rect 14749 2465 14783 2499
rect 16221 2465 16255 2499
rect 16773 2465 16807 2499
rect 16957 2465 16991 2499
rect 17877 2465 17911 2499
rect 18705 2465 18739 2499
rect 2605 2397 2639 2431
rect 3249 2397 3283 2431
rect 3801 2397 3835 2431
rect 7757 2397 7791 2431
rect 8309 2397 8343 2431
rect 9873 2397 9907 2431
rect 11161 2397 11195 2431
rect 11529 2397 11563 2431
rect 12725 2397 12759 2431
rect 14841 2397 14875 2431
rect 19441 2397 19475 2431
rect 21097 2397 21131 2431
rect 21373 2397 21407 2431
rect 4353 2329 4387 2363
rect 5365 2329 5399 2363
rect 5825 2329 5859 2363
rect 6837 2329 6871 2363
rect 7389 2329 7423 2363
rect 9505 2329 9539 2363
rect 14933 2329 14967 2363
rect 15945 2329 15979 2363
rect 16037 2329 16071 2363
rect 18613 2329 18647 2363
rect 3985 2261 4019 2295
rect 5273 2261 5307 2295
rect 7941 2261 7975 2295
rect 8953 2261 8987 2295
rect 10977 2261 11011 2295
rect 12081 2261 12115 2295
rect 13277 2261 13311 2295
rect 13369 2261 13403 2295
rect 13737 2261 13771 2295
rect 14289 2261 14323 2295
rect 15301 2261 15335 2295
rect 17049 2261 17083 2295
rect 18153 2261 18187 2295
rect 18521 2261 18555 2295
<< metal1 >>
rect 5994 21292 6000 21344
rect 6052 21332 6058 21344
rect 14642 21332 14648 21344
rect 6052 21304 14648 21332
rect 6052 21292 6058 21304
rect 14642 21292 14648 21304
rect 14700 21292 14706 21344
rect 8202 21224 8208 21276
rect 8260 21264 8266 21276
rect 12342 21264 12348 21276
rect 8260 21236 12348 21264
rect 8260 21224 8266 21236
rect 12342 21224 12348 21236
rect 12400 21224 12406 21276
rect 4890 21156 4896 21208
rect 4948 21196 4954 21208
rect 18414 21196 18420 21208
rect 4948 21168 18420 21196
rect 4948 21156 4954 21168
rect 18414 21156 18420 21168
rect 18472 21156 18478 21208
rect 4798 21088 4804 21140
rect 4856 21128 4862 21140
rect 20346 21128 20352 21140
rect 4856 21100 20352 21128
rect 4856 21088 4862 21100
rect 20346 21088 20352 21100
rect 20404 21088 20410 21140
rect 9306 21020 9312 21072
rect 9364 21060 9370 21072
rect 17586 21060 17592 21072
rect 9364 21032 17592 21060
rect 9364 21020 9370 21032
rect 17586 21020 17592 21032
rect 17644 21020 17650 21072
rect 7466 20952 7472 21004
rect 7524 20992 7530 21004
rect 17126 20992 17132 21004
rect 7524 20964 17132 20992
rect 7524 20952 7530 20964
rect 17126 20952 17132 20964
rect 17184 20952 17190 21004
rect 7098 20884 7104 20936
rect 7156 20924 7162 20936
rect 17218 20924 17224 20936
rect 7156 20896 17224 20924
rect 7156 20884 7162 20896
rect 17218 20884 17224 20896
rect 17276 20884 17282 20936
rect 7650 20816 7656 20868
rect 7708 20856 7714 20868
rect 11422 20856 11428 20868
rect 7708 20828 11428 20856
rect 7708 20816 7714 20828
rect 11422 20816 11428 20828
rect 11480 20816 11486 20868
rect 7374 20748 7380 20800
rect 7432 20788 7438 20800
rect 16206 20788 16212 20800
rect 7432 20760 16212 20788
rect 7432 20748 7438 20760
rect 16206 20748 16212 20760
rect 16264 20748 16270 20800
rect 1104 20698 21896 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21896 20698
rect 1104 20624 21896 20646
rect 3973 20587 4031 20593
rect 3973 20553 3985 20587
rect 4019 20584 4031 20587
rect 7190 20584 7196 20596
rect 4019 20556 7196 20584
rect 4019 20553 4031 20556
rect 3973 20547 4031 20553
rect 7190 20544 7196 20556
rect 7248 20544 7254 20596
rect 7377 20587 7435 20593
rect 7377 20553 7389 20587
rect 7423 20584 7435 20587
rect 7423 20556 12434 20584
rect 7423 20553 7435 20556
rect 7377 20547 7435 20553
rect 1946 20476 1952 20528
rect 2004 20516 2010 20528
rect 2133 20519 2191 20525
rect 2133 20516 2145 20519
rect 2004 20488 2145 20516
rect 2004 20476 2010 20488
rect 2133 20485 2145 20488
rect 2179 20485 2191 20519
rect 2133 20479 2191 20485
rect 3050 20476 3056 20528
rect 3108 20516 3114 20528
rect 3237 20519 3295 20525
rect 3237 20516 3249 20519
rect 3108 20488 3249 20516
rect 3108 20476 3114 20488
rect 3237 20485 3249 20488
rect 3283 20516 3295 20519
rect 3602 20516 3608 20528
rect 3283 20488 3608 20516
rect 3283 20485 3295 20488
rect 3237 20479 3295 20485
rect 3602 20476 3608 20488
rect 3660 20476 3666 20528
rect 4154 20476 4160 20528
rect 4212 20516 4218 20528
rect 4341 20519 4399 20525
rect 4341 20516 4353 20519
rect 4212 20488 4353 20516
rect 4212 20476 4218 20488
rect 4341 20485 4353 20488
rect 4387 20485 4399 20519
rect 7006 20516 7012 20528
rect 4341 20479 4399 20485
rect 4448 20488 7012 20516
rect 2498 20408 2504 20460
rect 2556 20448 2562 20460
rect 2593 20451 2651 20457
rect 2593 20448 2605 20451
rect 2556 20420 2605 20448
rect 2556 20408 2562 20420
rect 2593 20417 2605 20420
rect 2639 20417 2651 20451
rect 2593 20411 2651 20417
rect 3418 20408 3424 20460
rect 3476 20448 3482 20460
rect 3789 20451 3847 20457
rect 3789 20448 3801 20451
rect 3476 20420 3801 20448
rect 3476 20408 3482 20420
rect 3789 20417 3801 20420
rect 3835 20448 3847 20451
rect 4448 20448 4476 20488
rect 7006 20476 7012 20488
rect 7064 20476 7070 20528
rect 8481 20519 8539 20525
rect 8481 20485 8493 20519
rect 8527 20516 8539 20519
rect 9398 20516 9404 20528
rect 8527 20488 9404 20516
rect 8527 20485 8539 20488
rect 8481 20479 8539 20485
rect 9398 20476 9404 20488
rect 9456 20476 9462 20528
rect 9950 20516 9956 20528
rect 9911 20488 9956 20516
rect 9950 20476 9956 20488
rect 10008 20476 10014 20528
rect 11054 20476 11060 20528
rect 11112 20516 11118 20528
rect 12406 20516 12434 20556
rect 12618 20544 12624 20596
rect 12676 20584 12682 20596
rect 14277 20587 14335 20593
rect 14277 20584 14289 20587
rect 12676 20556 14289 20584
rect 12676 20544 12682 20556
rect 14277 20553 14289 20556
rect 14323 20553 14335 20587
rect 14277 20547 14335 20553
rect 14458 20544 14464 20596
rect 14516 20584 14522 20596
rect 14516 20556 15240 20584
rect 14516 20544 14522 20556
rect 11112 20488 11560 20516
rect 12406 20488 14136 20516
rect 11112 20476 11118 20488
rect 3835 20420 4476 20448
rect 5261 20451 5319 20457
rect 3835 20417 3847 20420
rect 3789 20411 3847 20417
rect 5261 20417 5273 20451
rect 5307 20417 5319 20451
rect 5261 20411 5319 20417
rect 1765 20383 1823 20389
rect 1765 20349 1777 20383
rect 1811 20380 1823 20383
rect 5166 20380 5172 20392
rect 1811 20352 5172 20380
rect 1811 20349 1823 20352
rect 1765 20343 1823 20349
rect 5166 20340 5172 20352
rect 5224 20340 5230 20392
rect 5278 20380 5306 20411
rect 5626 20408 5632 20460
rect 5684 20448 5690 20460
rect 5810 20448 5816 20460
rect 5684 20420 5816 20448
rect 5684 20408 5690 20420
rect 5810 20408 5816 20420
rect 5868 20408 5874 20460
rect 6638 20448 6644 20460
rect 6599 20420 6644 20448
rect 6638 20408 6644 20420
rect 6696 20408 6702 20460
rect 6822 20448 6828 20460
rect 6783 20420 6828 20448
rect 6822 20408 6828 20420
rect 6880 20408 6886 20460
rect 7193 20451 7251 20457
rect 7193 20417 7205 20451
rect 7239 20417 7251 20451
rect 7193 20411 7251 20417
rect 5350 20380 5356 20392
rect 5278 20352 5356 20380
rect 5350 20340 5356 20352
rect 5408 20340 5414 20392
rect 7208 20380 7236 20411
rect 7282 20408 7288 20460
rect 7340 20448 7346 20460
rect 7558 20448 7564 20460
rect 7340 20420 7564 20448
rect 7340 20408 7346 20420
rect 7558 20408 7564 20420
rect 7616 20448 7622 20460
rect 7745 20451 7803 20457
rect 7745 20448 7757 20451
rect 7616 20420 7757 20448
rect 7616 20408 7622 20420
rect 7745 20417 7757 20420
rect 7791 20417 7803 20451
rect 7745 20411 7803 20417
rect 7926 20408 7932 20460
rect 7984 20448 7990 20460
rect 8110 20448 8116 20460
rect 7984 20420 8116 20448
rect 7984 20408 7990 20420
rect 8110 20408 8116 20420
rect 8168 20448 8174 20460
rect 8297 20451 8355 20457
rect 8297 20448 8309 20451
rect 8168 20420 8309 20448
rect 8168 20408 8174 20420
rect 8297 20417 8309 20420
rect 8343 20417 8355 20451
rect 8297 20411 8355 20417
rect 8662 20408 8668 20460
rect 8720 20448 8726 20460
rect 9217 20451 9275 20457
rect 9217 20448 9229 20451
rect 8720 20420 9229 20448
rect 8720 20408 8726 20420
rect 9217 20417 9229 20420
rect 9263 20417 9275 20451
rect 9217 20411 9275 20417
rect 9674 20408 9680 20460
rect 9732 20448 9738 20460
rect 10318 20448 10324 20460
rect 9732 20420 10324 20448
rect 9732 20408 9738 20420
rect 10318 20408 10324 20420
rect 10376 20448 10382 20460
rect 10505 20451 10563 20457
rect 10505 20448 10517 20451
rect 10376 20420 10517 20448
rect 10376 20408 10382 20420
rect 10505 20417 10517 20420
rect 10551 20417 10563 20451
rect 11146 20448 11152 20460
rect 11107 20420 11152 20448
rect 10505 20411 10563 20417
rect 11146 20408 11152 20420
rect 11204 20408 11210 20460
rect 11532 20457 11560 20488
rect 11517 20451 11575 20457
rect 11517 20417 11529 20451
rect 11563 20417 11575 20451
rect 11517 20411 11575 20417
rect 12250 20408 12256 20460
rect 12308 20448 12314 20460
rect 12621 20451 12679 20457
rect 12621 20448 12633 20451
rect 12308 20420 12633 20448
rect 12308 20408 12314 20420
rect 12621 20417 12633 20420
rect 12667 20417 12679 20451
rect 12621 20411 12679 20417
rect 13354 20408 13360 20460
rect 13412 20448 13418 20460
rect 14108 20457 14136 20488
rect 14366 20476 14372 20528
rect 14424 20516 14430 20528
rect 14424 20488 15148 20516
rect 14424 20476 14430 20488
rect 13541 20451 13599 20457
rect 13541 20448 13553 20451
rect 13412 20420 13553 20448
rect 13412 20408 13418 20420
rect 13541 20417 13553 20420
rect 13587 20417 13599 20451
rect 13541 20411 13599 20417
rect 14093 20451 14151 20457
rect 14093 20417 14105 20451
rect 14139 20417 14151 20451
rect 14093 20411 14151 20417
rect 14645 20451 14703 20457
rect 14645 20417 14657 20451
rect 14691 20417 14703 20451
rect 14645 20411 14703 20417
rect 7834 20380 7840 20392
rect 7208 20352 7840 20380
rect 7834 20340 7840 20352
rect 7892 20340 7898 20392
rect 8018 20340 8024 20392
rect 8076 20380 8082 20392
rect 11793 20383 11851 20389
rect 8076 20352 11100 20380
rect 8076 20340 8082 20352
rect 2314 20312 2320 20324
rect 2275 20284 2320 20312
rect 2314 20272 2320 20284
rect 2372 20272 2378 20324
rect 4522 20312 4528 20324
rect 4483 20284 4528 20312
rect 4522 20272 4528 20284
rect 4580 20272 4586 20324
rect 4893 20315 4951 20321
rect 4893 20281 4905 20315
rect 4939 20312 4951 20315
rect 6822 20312 6828 20324
rect 4939 20284 6828 20312
rect 4939 20281 4951 20284
rect 4893 20275 4951 20281
rect 6822 20272 6828 20284
rect 6880 20272 6886 20324
rect 8294 20272 8300 20324
rect 8352 20312 8358 20324
rect 10965 20315 11023 20321
rect 10965 20312 10977 20315
rect 8352 20284 10977 20312
rect 8352 20272 8358 20284
rect 10965 20281 10977 20284
rect 11011 20281 11023 20315
rect 11072 20312 11100 20352
rect 11793 20349 11805 20383
rect 11839 20380 11851 20383
rect 11974 20380 11980 20392
rect 11839 20352 11980 20380
rect 11839 20349 11851 20352
rect 11793 20343 11851 20349
rect 11974 20340 11980 20352
rect 12032 20340 12038 20392
rect 14660 20380 14688 20411
rect 12406 20352 14688 20380
rect 12406 20312 12434 20352
rect 11072 20284 12434 20312
rect 10965 20275 11023 20281
rect 13170 20272 13176 20324
rect 13228 20312 13234 20324
rect 14829 20315 14887 20321
rect 14829 20312 14841 20315
rect 13228 20284 14841 20312
rect 13228 20272 13234 20284
rect 14829 20281 14841 20284
rect 14875 20281 14887 20315
rect 15120 20312 15148 20488
rect 15212 20457 15240 20556
rect 15378 20544 15384 20596
rect 15436 20584 15442 20596
rect 15933 20587 15991 20593
rect 15933 20584 15945 20587
rect 15436 20556 15945 20584
rect 15436 20544 15442 20556
rect 15933 20553 15945 20556
rect 15979 20553 15991 20587
rect 15933 20547 15991 20553
rect 16390 20544 16396 20596
rect 16448 20584 16454 20596
rect 17957 20587 18015 20593
rect 17957 20584 17969 20587
rect 16448 20556 17969 20584
rect 16448 20544 16454 20556
rect 17957 20553 17969 20556
rect 18003 20553 18015 20587
rect 17957 20547 18015 20553
rect 19429 20587 19487 20593
rect 19429 20553 19441 20587
rect 19475 20553 19487 20587
rect 19429 20547 19487 20553
rect 20533 20587 20591 20593
rect 20533 20553 20545 20587
rect 20579 20584 20591 20587
rect 21542 20584 21548 20596
rect 20579 20556 21548 20584
rect 20579 20553 20591 20556
rect 20533 20547 20591 20553
rect 15286 20476 15292 20528
rect 15344 20516 15350 20528
rect 15344 20488 17356 20516
rect 15344 20476 15350 20488
rect 15197 20451 15255 20457
rect 15197 20417 15209 20451
rect 15243 20417 15255 20451
rect 15746 20448 15752 20460
rect 15707 20420 15752 20448
rect 15197 20411 15255 20417
rect 15746 20408 15752 20420
rect 15804 20408 15810 20460
rect 16669 20451 16727 20457
rect 16669 20417 16681 20451
rect 16715 20448 16727 20451
rect 16942 20448 16948 20460
rect 16715 20420 16948 20448
rect 16715 20417 16727 20420
rect 16669 20411 16727 20417
rect 16942 20408 16948 20420
rect 17000 20408 17006 20460
rect 17218 20448 17224 20460
rect 17179 20420 17224 20448
rect 17218 20408 17224 20420
rect 17276 20408 17282 20460
rect 17328 20448 17356 20488
rect 17678 20476 17684 20528
rect 17736 20516 17742 20528
rect 19444 20516 19472 20547
rect 21542 20544 21548 20556
rect 21600 20544 21606 20596
rect 17736 20488 19472 20516
rect 17736 20476 17742 20488
rect 17773 20451 17831 20457
rect 17773 20448 17785 20451
rect 17328 20420 17785 20448
rect 17773 20417 17785 20420
rect 17819 20417 17831 20451
rect 17773 20411 17831 20417
rect 18046 20408 18052 20460
rect 18104 20448 18110 20460
rect 18325 20451 18383 20457
rect 18325 20448 18337 20451
rect 18104 20420 18337 20448
rect 18104 20408 18110 20420
rect 18325 20417 18337 20420
rect 18371 20417 18383 20451
rect 18325 20411 18383 20417
rect 18874 20408 18880 20460
rect 18932 20448 18938 20460
rect 19245 20451 19303 20457
rect 19245 20448 19257 20451
rect 18932 20420 19257 20448
rect 18932 20408 18938 20420
rect 19245 20417 19257 20420
rect 19291 20417 19303 20451
rect 19794 20448 19800 20460
rect 19755 20420 19800 20448
rect 19245 20411 19303 20417
rect 19794 20408 19800 20420
rect 19852 20408 19858 20460
rect 20346 20448 20352 20460
rect 20307 20420 20352 20448
rect 20346 20408 20352 20420
rect 20404 20408 20410 20460
rect 21082 20448 21088 20460
rect 21043 20420 21088 20448
rect 21082 20408 21088 20420
rect 21140 20408 21146 20460
rect 15286 20340 15292 20392
rect 15344 20380 15350 20392
rect 15344 20352 16988 20380
rect 15344 20340 15350 20352
rect 16853 20315 16911 20321
rect 16853 20312 16865 20315
rect 15120 20284 16865 20312
rect 14829 20275 14887 20281
rect 16853 20281 16865 20284
rect 16899 20281 16911 20315
rect 16853 20275 16911 20281
rect 2777 20247 2835 20253
rect 2777 20213 2789 20247
rect 2823 20244 2835 20247
rect 2958 20244 2964 20256
rect 2823 20216 2964 20244
rect 2823 20213 2835 20216
rect 2777 20207 2835 20213
rect 2958 20204 2964 20216
rect 3016 20204 3022 20256
rect 3326 20244 3332 20256
rect 3287 20216 3332 20244
rect 3326 20204 3332 20216
rect 3384 20204 3390 20256
rect 5353 20247 5411 20253
rect 5353 20213 5365 20247
rect 5399 20244 5411 20247
rect 5442 20244 5448 20256
rect 5399 20216 5448 20244
rect 5399 20213 5411 20216
rect 5353 20207 5411 20213
rect 5442 20204 5448 20216
rect 5500 20204 5506 20256
rect 5905 20247 5963 20253
rect 5905 20213 5917 20247
rect 5951 20244 5963 20247
rect 6270 20244 6276 20256
rect 5951 20216 6276 20244
rect 5951 20213 5963 20216
rect 5905 20207 5963 20213
rect 6270 20204 6276 20216
rect 6328 20204 6334 20256
rect 7742 20204 7748 20256
rect 7800 20244 7806 20256
rect 7837 20247 7895 20253
rect 7837 20244 7849 20247
rect 7800 20216 7849 20244
rect 7800 20204 7806 20216
rect 7837 20213 7849 20216
rect 7883 20213 7895 20247
rect 7837 20207 7895 20213
rect 9309 20247 9367 20253
rect 9309 20213 9321 20247
rect 9355 20244 9367 20247
rect 9490 20244 9496 20256
rect 9355 20216 9496 20244
rect 9355 20213 9367 20216
rect 9309 20207 9367 20213
rect 9490 20204 9496 20216
rect 9548 20204 9554 20256
rect 10042 20244 10048 20256
rect 10003 20216 10048 20244
rect 10042 20204 10048 20216
rect 10100 20204 10106 20256
rect 10597 20247 10655 20253
rect 10597 20213 10609 20247
rect 10643 20244 10655 20247
rect 10870 20244 10876 20256
rect 10643 20216 10876 20244
rect 10643 20213 10655 20216
rect 10597 20207 10655 20213
rect 10870 20204 10876 20216
rect 10928 20204 10934 20256
rect 13262 20244 13268 20256
rect 13223 20216 13268 20244
rect 13262 20204 13268 20216
rect 13320 20204 13326 20256
rect 13446 20204 13452 20256
rect 13504 20244 13510 20256
rect 13725 20247 13783 20253
rect 13725 20244 13737 20247
rect 13504 20216 13737 20244
rect 13504 20204 13510 20216
rect 13725 20213 13737 20216
rect 13771 20213 13783 20247
rect 13725 20207 13783 20213
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 15381 20247 15439 20253
rect 15381 20244 15393 20247
rect 13872 20216 15393 20244
rect 13872 20204 13878 20216
rect 15381 20213 15393 20216
rect 15427 20213 15439 20247
rect 16960 20244 16988 20352
rect 17034 20272 17040 20324
rect 17092 20312 17098 20324
rect 18509 20315 18567 20321
rect 18509 20312 18521 20315
rect 17092 20284 18521 20312
rect 17092 20272 17098 20284
rect 18509 20281 18521 20284
rect 18555 20281 18567 20315
rect 18509 20275 18567 20281
rect 19981 20315 20039 20321
rect 19981 20281 19993 20315
rect 20027 20312 20039 20315
rect 22094 20312 22100 20324
rect 20027 20284 22100 20312
rect 20027 20281 20039 20284
rect 19981 20275 20039 20281
rect 22094 20272 22100 20284
rect 22152 20272 22158 20324
rect 17405 20247 17463 20253
rect 17405 20244 17417 20247
rect 16960 20216 17417 20244
rect 15381 20207 15439 20213
rect 17405 20213 17417 20216
rect 17451 20213 17463 20247
rect 17405 20207 17463 20213
rect 18966 20204 18972 20256
rect 19024 20244 19030 20256
rect 21269 20247 21327 20253
rect 21269 20244 21281 20247
rect 19024 20216 21281 20244
rect 19024 20204 19030 20216
rect 21269 20213 21281 20216
rect 21315 20213 21327 20247
rect 21269 20207 21327 20213
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 4338 20040 4344 20052
rect 4299 20012 4344 20040
rect 4338 20000 4344 20012
rect 4396 20000 4402 20052
rect 4798 20040 4804 20052
rect 4759 20012 4804 20040
rect 4798 20000 4804 20012
rect 4856 20000 4862 20052
rect 5261 20043 5319 20049
rect 5261 20009 5273 20043
rect 5307 20040 5319 20043
rect 6641 20043 6699 20049
rect 5307 20012 5672 20040
rect 5307 20009 5319 20012
rect 5261 20003 5319 20009
rect 1394 19932 1400 19984
rect 1452 19932 1458 19984
rect 1670 19932 1676 19984
rect 1728 19972 1734 19984
rect 2409 19975 2467 19981
rect 2409 19972 2421 19975
rect 1728 19944 2421 19972
rect 1728 19932 1734 19944
rect 2409 19941 2421 19944
rect 2455 19941 2467 19975
rect 2409 19935 2467 19941
rect 3326 19932 3332 19984
rect 3384 19972 3390 19984
rect 5534 19972 5540 19984
rect 3384 19944 5540 19972
rect 3384 19932 3390 19944
rect 5534 19932 5540 19944
rect 5592 19932 5598 19984
rect 1412 19904 1440 19932
rect 2038 19904 2044 19916
rect 1412 19876 2044 19904
rect 2038 19864 2044 19876
rect 2096 19904 2102 19916
rect 5644 19904 5672 20012
rect 6641 20009 6653 20043
rect 6687 20040 6699 20043
rect 6914 20040 6920 20052
rect 6687 20012 6920 20040
rect 6687 20009 6699 20012
rect 6641 20003 6699 20009
rect 6914 20000 6920 20012
rect 6972 20000 6978 20052
rect 7561 20043 7619 20049
rect 7561 20009 7573 20043
rect 7607 20040 7619 20043
rect 7607 20012 12020 20040
rect 7607 20009 7619 20012
rect 7561 20003 7619 20009
rect 5718 19932 5724 19984
rect 5776 19972 5782 19984
rect 6181 19975 6239 19981
rect 5776 19944 5821 19972
rect 5776 19932 5782 19944
rect 6181 19941 6193 19975
rect 6227 19972 6239 19975
rect 6730 19972 6736 19984
rect 6227 19944 6736 19972
rect 6227 19941 6239 19944
rect 6181 19935 6239 19941
rect 6730 19932 6736 19944
rect 6788 19932 6794 19984
rect 7101 19975 7159 19981
rect 7101 19941 7113 19975
rect 7147 19972 7159 19975
rect 7147 19944 10640 19972
rect 7147 19941 7159 19944
rect 7101 19935 7159 19941
rect 2096 19876 2268 19904
rect 5644 19876 5856 19904
rect 2096 19864 2102 19876
rect 290 19796 296 19848
rect 348 19836 354 19848
rect 1394 19836 1400 19848
rect 348 19808 1400 19836
rect 348 19796 354 19808
rect 1394 19796 1400 19808
rect 1452 19836 1458 19848
rect 2240 19845 2268 19876
rect 1673 19839 1731 19845
rect 1673 19836 1685 19839
rect 1452 19808 1685 19836
rect 1452 19796 1458 19808
rect 1673 19805 1685 19808
rect 1719 19805 1731 19839
rect 1673 19799 1731 19805
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19805 2283 19839
rect 2225 19799 2283 19805
rect 2685 19839 2743 19845
rect 2685 19805 2697 19839
rect 2731 19805 2743 19839
rect 2685 19799 2743 19805
rect 842 19728 848 19780
rect 900 19768 906 19780
rect 2700 19768 2728 19799
rect 3142 19796 3148 19848
rect 3200 19836 3206 19848
rect 3237 19839 3295 19845
rect 3237 19836 3249 19839
rect 3200 19808 3249 19836
rect 3200 19796 3206 19808
rect 3237 19805 3249 19808
rect 3283 19805 3295 19839
rect 3237 19799 3295 19805
rect 3881 19839 3939 19845
rect 3881 19805 3893 19839
rect 3927 19836 3939 19839
rect 3970 19836 3976 19848
rect 3927 19808 3976 19836
rect 3927 19805 3939 19808
rect 3881 19799 3939 19805
rect 3970 19796 3976 19808
rect 4028 19796 4034 19848
rect 4157 19839 4215 19845
rect 4157 19805 4169 19839
rect 4203 19836 4215 19839
rect 4430 19836 4436 19848
rect 4203 19808 4436 19836
rect 4203 19805 4215 19808
rect 4157 19799 4215 19805
rect 4430 19796 4436 19808
rect 4488 19796 4494 19848
rect 4617 19839 4675 19845
rect 4617 19805 4629 19839
rect 4663 19836 4675 19839
rect 4798 19836 4804 19848
rect 4663 19808 4804 19836
rect 4663 19805 4675 19808
rect 4617 19799 4675 19805
rect 4798 19796 4804 19808
rect 4856 19796 4862 19848
rect 5077 19839 5135 19845
rect 5077 19805 5089 19839
rect 5123 19805 5135 19839
rect 5077 19799 5135 19805
rect 5537 19839 5595 19845
rect 5537 19805 5549 19839
rect 5583 19836 5595 19839
rect 5718 19836 5724 19848
rect 5583 19808 5724 19836
rect 5583 19805 5595 19808
rect 5537 19799 5595 19805
rect 900 19740 2728 19768
rect 900 19728 906 19740
rect 2240 19712 2268 19740
rect 2774 19728 2780 19780
rect 2832 19768 2838 19780
rect 2832 19740 3924 19768
rect 2832 19728 2838 19740
rect 1762 19700 1768 19712
rect 1723 19672 1768 19700
rect 1762 19660 1768 19672
rect 1820 19660 1826 19712
rect 2222 19660 2228 19712
rect 2280 19660 2286 19712
rect 2869 19703 2927 19709
rect 2869 19669 2881 19703
rect 2915 19700 2927 19703
rect 3234 19700 3240 19712
rect 2915 19672 3240 19700
rect 2915 19669 2927 19672
rect 2869 19663 2927 19669
rect 3234 19660 3240 19672
rect 3292 19660 3298 19712
rect 3329 19703 3387 19709
rect 3329 19669 3341 19703
rect 3375 19700 3387 19703
rect 3786 19700 3792 19712
rect 3375 19672 3792 19700
rect 3375 19669 3387 19672
rect 3329 19663 3387 19669
rect 3786 19660 3792 19672
rect 3844 19660 3850 19712
rect 3896 19700 3924 19740
rect 4246 19728 4252 19780
rect 4304 19768 4310 19780
rect 5092 19768 5120 19799
rect 5718 19796 5724 19808
rect 5776 19796 5782 19848
rect 4304 19740 5120 19768
rect 5828 19768 5856 19876
rect 6270 19864 6276 19916
rect 6328 19904 6334 19916
rect 7742 19904 7748 19916
rect 6328 19876 6776 19904
rect 6328 19864 6334 19876
rect 6748 19848 6776 19876
rect 6932 19876 7748 19904
rect 5994 19836 6000 19848
rect 5955 19808 6000 19836
rect 5994 19796 6000 19808
rect 6052 19796 6058 19848
rect 6086 19796 6092 19848
rect 6144 19836 6150 19848
rect 6457 19839 6515 19845
rect 6457 19836 6469 19839
rect 6144 19808 6469 19836
rect 6144 19796 6150 19808
rect 6457 19805 6469 19808
rect 6503 19805 6515 19839
rect 6457 19799 6515 19805
rect 6730 19796 6736 19848
rect 6788 19796 6794 19848
rect 6932 19845 6960 19876
rect 7742 19864 7748 19876
rect 7800 19864 7806 19916
rect 10134 19904 10140 19916
rect 10095 19876 10140 19904
rect 10134 19864 10140 19876
rect 10192 19864 10198 19916
rect 6917 19839 6975 19845
rect 6917 19805 6929 19839
rect 6963 19805 6975 19839
rect 6917 19799 6975 19805
rect 7377 19839 7435 19845
rect 7377 19805 7389 19839
rect 7423 19836 7435 19839
rect 7650 19836 7656 19848
rect 7423 19808 7656 19836
rect 7423 19805 7435 19808
rect 7377 19799 7435 19805
rect 7650 19796 7656 19808
rect 7708 19796 7714 19848
rect 7837 19839 7895 19845
rect 7837 19805 7849 19839
rect 7883 19836 7895 19839
rect 8202 19836 8208 19848
rect 7883 19808 8208 19836
rect 7883 19805 7895 19808
rect 7837 19799 7895 19805
rect 8202 19796 8208 19808
rect 8260 19796 8266 19848
rect 8297 19839 8355 19845
rect 8297 19805 8309 19839
rect 8343 19805 8355 19839
rect 8297 19799 8355 19805
rect 8312 19768 8340 19799
rect 8386 19796 8392 19848
rect 8444 19836 8450 19848
rect 9401 19839 9459 19845
rect 9401 19836 9413 19839
rect 8444 19808 9413 19836
rect 8444 19796 8450 19808
rect 9401 19805 9413 19808
rect 9447 19805 9459 19839
rect 9401 19799 9459 19805
rect 10321 19771 10379 19777
rect 10321 19768 10333 19771
rect 5828 19740 8340 19768
rect 8404 19740 10333 19768
rect 4304 19728 4310 19740
rect 7650 19700 7656 19712
rect 3896 19672 7656 19700
rect 7650 19660 7656 19672
rect 7708 19660 7714 19712
rect 8018 19700 8024 19712
rect 7979 19672 8024 19700
rect 8018 19660 8024 19672
rect 8076 19660 8082 19712
rect 8110 19660 8116 19712
rect 8168 19700 8174 19712
rect 8404 19700 8432 19740
rect 10321 19737 10333 19740
rect 10367 19737 10379 19771
rect 10612 19768 10640 19944
rect 10962 19836 10968 19848
rect 10923 19808 10968 19836
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 11238 19845 11244 19848
rect 11232 19836 11244 19845
rect 11199 19808 11244 19836
rect 11232 19799 11244 19808
rect 11238 19796 11244 19799
rect 11296 19796 11302 19848
rect 11992 19836 12020 20012
rect 12158 20000 12164 20052
rect 12216 20040 12222 20052
rect 14277 20043 14335 20049
rect 14277 20040 14289 20043
rect 12216 20012 14289 20040
rect 12216 20000 12222 20012
rect 14277 20009 14289 20012
rect 14323 20009 14335 20043
rect 14277 20003 14335 20009
rect 15930 20000 15936 20052
rect 15988 20040 15994 20052
rect 17221 20043 17279 20049
rect 17221 20040 17233 20043
rect 15988 20012 17233 20040
rect 15988 20000 15994 20012
rect 17221 20009 17233 20012
rect 17267 20009 17279 20043
rect 17221 20003 17279 20009
rect 17773 20043 17831 20049
rect 17773 20009 17785 20043
rect 17819 20040 17831 20043
rect 17862 20040 17868 20052
rect 17819 20012 17868 20040
rect 17819 20009 17831 20012
rect 17773 20003 17831 20009
rect 17862 20000 17868 20012
rect 17920 20000 17926 20052
rect 18322 20040 18328 20052
rect 18283 20012 18328 20040
rect 18322 20000 18328 20012
rect 18380 20000 18386 20052
rect 18874 20040 18880 20052
rect 18835 20012 18880 20040
rect 18874 20000 18880 20012
rect 18932 20000 18938 20052
rect 12066 19932 12072 19984
rect 12124 19972 12130 19984
rect 12124 19944 14136 19972
rect 12124 19932 12130 19944
rect 12986 19904 12992 19916
rect 12947 19876 12992 19904
rect 12986 19864 12992 19876
rect 13044 19864 13050 19916
rect 14108 19845 14136 19944
rect 18230 19932 18236 19984
rect 18288 19972 18294 19984
rect 19429 19975 19487 19981
rect 19429 19972 19441 19975
rect 18288 19944 19441 19972
rect 18288 19932 18294 19944
rect 19429 19941 19441 19944
rect 19475 19941 19487 19975
rect 19429 19935 19487 19941
rect 14826 19904 14832 19916
rect 14787 19876 14832 19904
rect 14826 19864 14832 19876
rect 14884 19864 14890 19916
rect 17494 19864 17500 19916
rect 17552 19904 17558 19916
rect 20530 19904 20536 19916
rect 17552 19876 20536 19904
rect 17552 19864 17558 19876
rect 20530 19864 20536 19876
rect 20588 19864 20594 19916
rect 13173 19839 13231 19845
rect 13173 19836 13185 19839
rect 11992 19808 13185 19836
rect 13173 19805 13185 19808
rect 13219 19805 13231 19839
rect 13173 19799 13231 19805
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19805 14151 19839
rect 15010 19836 15016 19848
rect 14971 19808 15016 19836
rect 14093 19799 14151 19805
rect 15010 19796 15016 19808
rect 15068 19796 15074 19848
rect 15102 19796 15108 19848
rect 15160 19836 15166 19848
rect 16114 19836 16120 19848
rect 15160 19808 16120 19836
rect 15160 19796 15166 19808
rect 16114 19796 16120 19808
rect 16172 19796 16178 19848
rect 16206 19796 16212 19848
rect 16264 19836 16270 19848
rect 17037 19839 17095 19845
rect 17037 19836 17049 19839
rect 16264 19808 17049 19836
rect 16264 19796 16270 19808
rect 17037 19805 17049 19808
rect 17083 19805 17095 19839
rect 17586 19836 17592 19848
rect 17547 19808 17592 19836
rect 17037 19799 17095 19805
rect 17586 19796 17592 19808
rect 17644 19796 17650 19848
rect 18138 19836 18144 19848
rect 18099 19808 18144 19836
rect 18138 19796 18144 19808
rect 18196 19796 18202 19848
rect 18598 19796 18604 19848
rect 18656 19836 18662 19848
rect 18693 19839 18751 19845
rect 18693 19836 18705 19839
rect 18656 19808 18705 19836
rect 18656 19796 18662 19808
rect 18693 19805 18705 19808
rect 18739 19805 18751 19839
rect 18693 19799 18751 19805
rect 19245 19839 19303 19845
rect 19245 19805 19257 19839
rect 19291 19805 19303 19839
rect 20806 19836 20812 19848
rect 20767 19808 20812 19836
rect 19245 19799 19303 19805
rect 10612 19740 11836 19768
rect 10321 19731 10379 19737
rect 8168 19672 8432 19700
rect 8168 19660 8174 19672
rect 8478 19660 8484 19712
rect 8536 19700 8542 19712
rect 9122 19700 9128 19712
rect 8536 19672 8581 19700
rect 9083 19672 9128 19700
rect 8536 19660 8542 19672
rect 9122 19660 9128 19672
rect 9180 19660 9186 19712
rect 9582 19700 9588 19712
rect 9543 19672 9588 19700
rect 9582 19660 9588 19672
rect 9640 19660 9646 19712
rect 10226 19700 10232 19712
rect 10187 19672 10232 19700
rect 10226 19660 10232 19672
rect 10284 19660 10290 19712
rect 10686 19700 10692 19712
rect 10647 19672 10692 19700
rect 10686 19660 10692 19672
rect 10744 19660 10750 19712
rect 11808 19700 11836 19740
rect 11882 19728 11888 19780
rect 11940 19768 11946 19780
rect 15657 19771 15715 19777
rect 15657 19768 15669 19771
rect 11940 19740 15669 19768
rect 11940 19728 11946 19740
rect 15657 19737 15669 19740
rect 15703 19737 15715 19771
rect 15657 19731 15715 19737
rect 16942 19728 16948 19780
rect 17000 19768 17006 19780
rect 19260 19768 19288 19799
rect 20806 19796 20812 19808
rect 20864 19796 20870 19848
rect 20162 19768 20168 19780
rect 17000 19740 19288 19768
rect 20123 19740 20168 19768
rect 17000 19728 17006 19740
rect 20162 19728 20168 19740
rect 20220 19728 20226 19780
rect 21266 19768 21272 19780
rect 21227 19740 21272 19768
rect 21266 19728 21272 19740
rect 21324 19728 21330 19780
rect 12066 19700 12072 19712
rect 11808 19672 12072 19700
rect 12066 19660 12072 19672
rect 12124 19660 12130 19712
rect 12250 19660 12256 19712
rect 12308 19700 12314 19712
rect 12345 19703 12403 19709
rect 12345 19700 12357 19703
rect 12308 19672 12357 19700
rect 12308 19660 12314 19672
rect 12345 19669 12357 19672
rect 12391 19669 12403 19703
rect 13078 19700 13084 19712
rect 13039 19672 13084 19700
rect 12345 19663 12403 19669
rect 13078 19660 13084 19672
rect 13136 19660 13142 19712
rect 13541 19703 13599 19709
rect 13541 19669 13553 19703
rect 13587 19700 13599 19703
rect 13722 19700 13728 19712
rect 13587 19672 13728 19700
rect 13587 19669 13599 19672
rect 13541 19663 13599 19669
rect 13722 19660 13728 19672
rect 13780 19660 13786 19712
rect 13814 19660 13820 19712
rect 13872 19700 13878 19712
rect 14921 19703 14979 19709
rect 14921 19700 14933 19703
rect 13872 19672 14933 19700
rect 13872 19660 13878 19672
rect 14921 19669 14933 19672
rect 14967 19669 14979 19703
rect 14921 19663 14979 19669
rect 15286 19660 15292 19712
rect 15344 19700 15350 19712
rect 15381 19703 15439 19709
rect 15381 19700 15393 19703
rect 15344 19672 15393 19700
rect 15344 19660 15350 19672
rect 15381 19669 15393 19672
rect 15427 19669 15439 19703
rect 15381 19663 15439 19669
rect 15746 19660 15752 19712
rect 15804 19700 15810 19712
rect 16761 19703 16819 19709
rect 16761 19700 16773 19703
rect 15804 19672 16773 19700
rect 15804 19660 15810 19672
rect 16761 19669 16773 19672
rect 16807 19669 16819 19703
rect 16761 19663 16819 19669
rect 18598 19660 18604 19712
rect 18656 19700 18662 19712
rect 18782 19700 18788 19712
rect 18656 19672 18788 19700
rect 18656 19660 18662 19672
rect 18782 19660 18788 19672
rect 18840 19660 18846 19712
rect 1104 19610 21896 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21896 19610
rect 1104 19536 21896 19558
rect 3697 19499 3755 19505
rect 3697 19465 3709 19499
rect 3743 19496 3755 19499
rect 3878 19496 3884 19508
rect 3743 19468 3884 19496
rect 3743 19465 3755 19468
rect 3697 19459 3755 19465
rect 3878 19456 3884 19468
rect 3936 19456 3942 19508
rect 4157 19499 4215 19505
rect 4157 19465 4169 19499
rect 4203 19496 4215 19499
rect 4522 19496 4528 19508
rect 4203 19468 4528 19496
rect 4203 19465 4215 19468
rect 4157 19459 4215 19465
rect 4522 19456 4528 19468
rect 4580 19456 4586 19508
rect 4706 19456 4712 19508
rect 4764 19496 4770 19508
rect 6457 19499 6515 19505
rect 6457 19496 6469 19499
rect 4764 19468 6469 19496
rect 4764 19456 4770 19468
rect 6457 19465 6469 19468
rect 6503 19465 6515 19499
rect 7098 19496 7104 19508
rect 7059 19468 7104 19496
rect 6457 19459 6515 19465
rect 7098 19456 7104 19468
rect 7156 19456 7162 19508
rect 7561 19499 7619 19505
rect 7561 19465 7573 19499
rect 7607 19496 7619 19499
rect 8386 19496 8392 19508
rect 7607 19468 8392 19496
rect 7607 19465 7619 19468
rect 7561 19459 7619 19465
rect 8386 19456 8392 19468
rect 8444 19456 8450 19508
rect 8481 19499 8539 19505
rect 8481 19465 8493 19499
rect 8527 19465 8539 19499
rect 8481 19459 8539 19465
rect 8941 19499 8999 19505
rect 8941 19465 8953 19499
rect 8987 19496 8999 19499
rect 12713 19499 12771 19505
rect 8987 19468 12664 19496
rect 8987 19465 8999 19468
rect 8941 19459 8999 19465
rect 4614 19428 4620 19440
rect 3988 19400 4620 19428
rect 3988 19369 4016 19400
rect 4614 19388 4620 19400
rect 4672 19388 4678 19440
rect 5997 19431 6055 19437
rect 5997 19397 6009 19431
rect 6043 19428 6055 19431
rect 7006 19428 7012 19440
rect 6043 19400 7012 19428
rect 6043 19397 6055 19400
rect 5997 19391 6055 19397
rect 7006 19388 7012 19400
rect 7064 19388 7070 19440
rect 8496 19428 8524 19459
rect 12636 19428 12664 19468
rect 12713 19465 12725 19499
rect 12759 19496 12771 19499
rect 16114 19496 16120 19508
rect 12759 19468 15976 19496
rect 16075 19468 16120 19496
rect 12759 19465 12771 19468
rect 12713 19459 12771 19465
rect 14458 19428 14464 19440
rect 7852 19400 8432 19428
rect 8496 19400 12434 19428
rect 12636 19400 14464 19428
rect 3973 19363 4031 19369
rect 3973 19329 3985 19363
rect 4019 19329 4031 19363
rect 3973 19323 4031 19329
rect 4338 19320 4344 19372
rect 4396 19360 4402 19372
rect 4433 19363 4491 19369
rect 4433 19360 4445 19363
rect 4396 19332 4445 19360
rect 4396 19320 4402 19332
rect 4433 19329 4445 19332
rect 4479 19329 4491 19363
rect 4433 19323 4491 19329
rect 4893 19363 4951 19369
rect 4893 19329 4905 19363
rect 4939 19360 4951 19363
rect 4982 19360 4988 19372
rect 4939 19332 4988 19360
rect 4939 19329 4951 19332
rect 4893 19323 4951 19329
rect 4982 19320 4988 19332
rect 5040 19320 5046 19372
rect 5166 19320 5172 19372
rect 5224 19360 5230 19372
rect 5350 19360 5356 19372
rect 5224 19332 5356 19360
rect 5224 19320 5230 19332
rect 5350 19320 5356 19332
rect 5408 19320 5414 19372
rect 5537 19363 5595 19369
rect 5537 19329 5549 19363
rect 5583 19360 5595 19363
rect 5810 19360 5816 19372
rect 5583 19332 5816 19360
rect 5583 19329 5595 19332
rect 5537 19323 5595 19329
rect 5810 19320 5816 19332
rect 5868 19320 5874 19372
rect 6086 19320 6092 19372
rect 6144 19360 6150 19372
rect 6641 19363 6699 19369
rect 6641 19360 6653 19363
rect 6144 19332 6653 19360
rect 6144 19320 6150 19332
rect 6641 19329 6653 19332
rect 6687 19329 6699 19363
rect 6914 19360 6920 19372
rect 6875 19332 6920 19360
rect 6641 19323 6699 19329
rect 6914 19320 6920 19332
rect 6972 19320 6978 19372
rect 7098 19320 7104 19372
rect 7156 19360 7162 19372
rect 7282 19360 7288 19372
rect 7156 19332 7288 19360
rect 7156 19320 7162 19332
rect 7282 19320 7288 19332
rect 7340 19320 7346 19372
rect 7377 19363 7435 19369
rect 7377 19329 7389 19363
rect 7423 19360 7435 19363
rect 7558 19360 7564 19372
rect 7423 19332 7564 19360
rect 7423 19329 7435 19332
rect 7377 19323 7435 19329
rect 7558 19320 7564 19332
rect 7616 19320 7622 19372
rect 7852 19369 7880 19400
rect 7837 19363 7895 19369
rect 7837 19329 7849 19363
rect 7883 19329 7895 19363
rect 8294 19360 8300 19372
rect 8255 19332 8300 19360
rect 7837 19323 7895 19329
rect 2961 19295 3019 19301
rect 2961 19261 2973 19295
rect 3007 19292 3019 19295
rect 7852 19292 7880 19323
rect 8294 19320 8300 19332
rect 8352 19320 8358 19372
rect 8404 19360 8432 19400
rect 8496 19360 8616 19364
rect 8754 19360 8760 19372
rect 8404 19336 8616 19360
rect 8404 19332 8524 19336
rect 3007 19264 7880 19292
rect 8588 19292 8616 19336
rect 8715 19332 8760 19360
rect 8754 19320 8760 19332
rect 8812 19320 8818 19372
rect 9214 19320 9220 19372
rect 9272 19360 9278 19372
rect 9493 19363 9551 19369
rect 9493 19360 9505 19363
rect 9272 19332 9505 19360
rect 9272 19320 9278 19332
rect 9493 19329 9505 19332
rect 9539 19329 9551 19363
rect 9766 19360 9772 19372
rect 9727 19332 9772 19360
rect 9493 19323 9551 19329
rect 9766 19320 9772 19332
rect 9824 19320 9830 19372
rect 10036 19363 10094 19369
rect 10036 19329 10048 19363
rect 10082 19360 10094 19363
rect 10502 19360 10508 19372
rect 10082 19332 10508 19360
rect 10082 19329 10094 19332
rect 10036 19323 10094 19329
rect 10502 19320 10508 19332
rect 10560 19320 10566 19372
rect 11882 19360 11888 19372
rect 11843 19332 11888 19360
rect 11882 19320 11888 19332
rect 11940 19320 11946 19372
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19360 12035 19363
rect 12158 19360 12164 19372
rect 12023 19332 12164 19360
rect 12023 19329 12035 19332
rect 11977 19323 12035 19329
rect 12158 19320 12164 19332
rect 12216 19320 12222 19372
rect 12406 19360 12434 19400
rect 14458 19388 14464 19400
rect 14516 19388 14522 19440
rect 15378 19428 15384 19440
rect 14752 19400 15384 19428
rect 12529 19363 12587 19369
rect 12529 19360 12541 19363
rect 12406 19332 12541 19360
rect 12529 19329 12541 19332
rect 12575 19329 12587 19363
rect 12529 19323 12587 19329
rect 13348 19363 13406 19369
rect 13348 19329 13360 19363
rect 13394 19360 13406 19363
rect 13630 19360 13636 19372
rect 13394 19332 13636 19360
rect 13394 19329 13406 19332
rect 13348 19323 13406 19329
rect 13630 19320 13636 19332
rect 13688 19320 13694 19372
rect 14752 19369 14780 19400
rect 15378 19388 15384 19400
rect 15436 19388 15442 19440
rect 15948 19428 15976 19468
rect 16114 19456 16120 19468
rect 16172 19456 16178 19508
rect 16853 19499 16911 19505
rect 16853 19465 16865 19499
rect 16899 19496 16911 19499
rect 17310 19496 17316 19508
rect 16899 19468 17316 19496
rect 16899 19465 16911 19468
rect 16853 19459 16911 19465
rect 17310 19456 17316 19468
rect 17368 19456 17374 19508
rect 17405 19499 17463 19505
rect 17405 19465 17417 19499
rect 17451 19496 17463 19499
rect 18046 19496 18052 19508
rect 17451 19468 18052 19496
rect 17451 19465 17463 19468
rect 17405 19459 17463 19465
rect 18046 19456 18052 19468
rect 18104 19456 18110 19508
rect 18506 19496 18512 19508
rect 18467 19468 18512 19496
rect 18506 19456 18512 19468
rect 18564 19456 18570 19508
rect 19242 19456 19248 19508
rect 19300 19496 19306 19508
rect 19613 19499 19671 19505
rect 19613 19496 19625 19499
rect 19300 19468 19625 19496
rect 19300 19456 19306 19468
rect 19613 19465 19625 19468
rect 19659 19465 19671 19499
rect 19613 19459 19671 19465
rect 20165 19499 20223 19505
rect 20165 19465 20177 19499
rect 20211 19465 20223 19499
rect 21266 19496 21272 19508
rect 21227 19468 21272 19496
rect 20165 19459 20223 19465
rect 17954 19428 17960 19440
rect 15948 19400 17960 19428
rect 17954 19388 17960 19400
rect 18012 19388 18018 19440
rect 18782 19388 18788 19440
rect 18840 19428 18846 19440
rect 20180 19428 20208 19459
rect 21266 19456 21272 19468
rect 21324 19456 21330 19508
rect 18840 19400 20208 19428
rect 18840 19388 18846 19400
rect 14737 19363 14795 19369
rect 14737 19329 14749 19363
rect 14783 19329 14795 19363
rect 14737 19323 14795 19329
rect 14826 19320 14832 19372
rect 14884 19360 14890 19372
rect 14993 19363 15051 19369
rect 14993 19360 15005 19363
rect 14884 19332 15005 19360
rect 14884 19320 14890 19332
rect 14993 19329 15005 19332
rect 15039 19329 15051 19363
rect 14993 19323 15051 19329
rect 16669 19363 16727 19369
rect 16669 19329 16681 19363
rect 16715 19360 16727 19363
rect 17034 19360 17040 19372
rect 16715 19332 17040 19360
rect 16715 19329 16727 19332
rect 16669 19323 16727 19329
rect 17034 19320 17040 19332
rect 17092 19320 17098 19372
rect 17126 19320 17132 19372
rect 17184 19360 17190 19372
rect 17221 19363 17279 19369
rect 17221 19360 17233 19363
rect 17184 19332 17233 19360
rect 17184 19320 17190 19332
rect 17221 19329 17233 19332
rect 17267 19329 17279 19363
rect 17770 19360 17776 19372
rect 17731 19332 17776 19360
rect 17221 19323 17279 19329
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 17862 19320 17868 19372
rect 17920 19360 17926 19372
rect 18325 19363 18383 19369
rect 18325 19360 18337 19363
rect 17920 19332 18337 19360
rect 17920 19320 17926 19332
rect 18325 19329 18337 19332
rect 18371 19329 18383 19363
rect 18874 19360 18880 19372
rect 18835 19332 18880 19360
rect 18325 19323 18383 19329
rect 18874 19320 18880 19332
rect 18932 19320 18938 19372
rect 19426 19360 19432 19372
rect 19387 19332 19432 19360
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 19610 19320 19616 19372
rect 19668 19360 19674 19372
rect 19981 19363 20039 19369
rect 19981 19360 19993 19363
rect 19668 19332 19993 19360
rect 19668 19320 19674 19332
rect 19981 19329 19993 19332
rect 20027 19329 20039 19363
rect 20530 19360 20536 19372
rect 20491 19332 20536 19360
rect 19981 19323 20039 19329
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 21085 19363 21143 19369
rect 21085 19329 21097 19363
rect 21131 19360 21143 19363
rect 21174 19360 21180 19372
rect 21131 19332 21180 19360
rect 21131 19329 21143 19332
rect 21085 19323 21143 19329
rect 21174 19320 21180 19332
rect 21232 19320 21238 19372
rect 9030 19292 9036 19304
rect 8588 19264 9036 19292
rect 3007 19261 3019 19264
rect 2961 19255 3019 19261
rect 9030 19252 9036 19264
rect 9088 19252 9094 19304
rect 9674 19292 9680 19304
rect 9140 19264 9680 19292
rect 2225 19227 2283 19233
rect 2225 19193 2237 19227
rect 2271 19224 2283 19227
rect 2682 19224 2688 19236
rect 2271 19196 2688 19224
rect 2271 19193 2283 19196
rect 2225 19187 2283 19193
rect 2682 19184 2688 19196
rect 2740 19184 2746 19236
rect 3329 19227 3387 19233
rect 3329 19193 3341 19227
rect 3375 19224 3387 19227
rect 5074 19224 5080 19236
rect 3375 19196 4936 19224
rect 5035 19196 5080 19224
rect 3375 19193 3387 19196
rect 3329 19187 3387 19193
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 1854 19156 1860 19168
rect 1815 19128 1860 19156
rect 1854 19116 1860 19128
rect 1912 19116 1918 19168
rect 2590 19156 2596 19168
rect 2551 19128 2596 19156
rect 2590 19116 2596 19128
rect 2648 19116 2654 19168
rect 4617 19159 4675 19165
rect 4617 19125 4629 19159
rect 4663 19156 4675 19159
rect 4798 19156 4804 19168
rect 4663 19128 4804 19156
rect 4663 19125 4675 19128
rect 4617 19119 4675 19125
rect 4798 19116 4804 19128
rect 4856 19116 4862 19168
rect 4908 19156 4936 19196
rect 5074 19184 5080 19196
rect 5132 19184 5138 19236
rect 8021 19227 8079 19233
rect 5184 19196 6500 19224
rect 5184 19156 5212 19196
rect 5350 19156 5356 19168
rect 4908 19128 5212 19156
rect 5311 19128 5356 19156
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 6472 19156 6500 19196
rect 8021 19193 8033 19227
rect 8067 19224 8079 19227
rect 8110 19224 8116 19236
rect 8067 19196 8116 19224
rect 8067 19193 8079 19196
rect 8021 19187 8079 19193
rect 8110 19184 8116 19196
rect 8168 19184 8174 19236
rect 9140 19224 9168 19264
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 11238 19252 11244 19304
rect 11296 19252 11302 19304
rect 12066 19252 12072 19304
rect 12124 19292 12130 19304
rect 13078 19292 13084 19304
rect 12124 19264 12169 19292
rect 13039 19264 13084 19292
rect 12124 19252 12130 19264
rect 13078 19252 13084 19264
rect 13136 19252 13142 19304
rect 14844 19292 14872 19320
rect 19334 19292 19340 19304
rect 14476 19264 14872 19292
rect 15764 19264 19340 19292
rect 8772 19196 9168 19224
rect 8772 19156 8800 19196
rect 9582 19184 9588 19236
rect 9640 19224 9646 19236
rect 11149 19227 11207 19233
rect 9640 19196 9812 19224
rect 9640 19184 9646 19196
rect 6472 19128 8800 19156
rect 9306 19116 9312 19168
rect 9364 19156 9370 19168
rect 9784 19156 9812 19196
rect 11149 19193 11161 19227
rect 11195 19224 11207 19227
rect 11256 19224 11284 19252
rect 12084 19224 12112 19252
rect 11195 19196 12112 19224
rect 11195 19193 11207 19196
rect 11149 19187 11207 19193
rect 11054 19156 11060 19168
rect 9364 19128 9409 19156
rect 9784 19128 11060 19156
rect 9364 19116 9370 19128
rect 11054 19116 11060 19128
rect 11112 19116 11118 19168
rect 11238 19116 11244 19168
rect 11296 19156 11302 19168
rect 11517 19159 11575 19165
rect 11517 19156 11529 19159
rect 11296 19128 11529 19156
rect 11296 19116 11302 19128
rect 11517 19125 11529 19128
rect 11563 19125 11575 19159
rect 11517 19119 11575 19125
rect 14366 19116 14372 19168
rect 14424 19156 14430 19168
rect 14476 19165 14504 19264
rect 14461 19159 14519 19165
rect 14461 19156 14473 19159
rect 14424 19128 14473 19156
rect 14424 19116 14430 19128
rect 14461 19125 14473 19128
rect 14507 19125 14519 19159
rect 14461 19119 14519 19125
rect 14550 19116 14556 19168
rect 14608 19156 14614 19168
rect 15764 19156 15792 19264
rect 19334 19252 19340 19264
rect 19392 19252 19398 19304
rect 19518 19252 19524 19304
rect 19576 19292 19582 19304
rect 22646 19292 22652 19304
rect 19576 19264 22652 19292
rect 19576 19252 19582 19264
rect 22646 19252 22652 19264
rect 22704 19252 22710 19304
rect 17957 19227 18015 19233
rect 17957 19193 17969 19227
rect 18003 19224 18015 19227
rect 20990 19224 20996 19236
rect 18003 19196 20996 19224
rect 18003 19193 18015 19196
rect 17957 19187 18015 19193
rect 20990 19184 20996 19196
rect 21048 19184 21054 19236
rect 14608 19128 15792 19156
rect 19061 19159 19119 19165
rect 14608 19116 14614 19128
rect 19061 19125 19073 19159
rect 19107 19156 19119 19159
rect 19518 19156 19524 19168
rect 19107 19128 19524 19156
rect 19107 19125 19119 19128
rect 19061 19119 19119 19125
rect 19518 19116 19524 19128
rect 19576 19116 19582 19168
rect 20714 19156 20720 19168
rect 20675 19128 20720 19156
rect 20714 19116 20720 19128
rect 20772 19116 20778 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1578 18952 1584 18964
rect 1539 18924 1584 18952
rect 1578 18912 1584 18924
rect 1636 18912 1642 18964
rect 2406 18912 2412 18964
rect 2464 18952 2470 18964
rect 2593 18955 2651 18961
rect 2593 18952 2605 18955
rect 2464 18924 2605 18952
rect 2464 18912 2470 18924
rect 2593 18921 2605 18924
rect 2639 18921 2651 18955
rect 2593 18915 2651 18921
rect 3053 18955 3111 18961
rect 3053 18921 3065 18955
rect 3099 18952 3111 18955
rect 4062 18952 4068 18964
rect 3099 18924 4068 18952
rect 3099 18921 3111 18924
rect 3053 18915 3111 18921
rect 4062 18912 4068 18924
rect 4120 18912 4126 18964
rect 4433 18955 4491 18961
rect 4433 18921 4445 18955
rect 4479 18952 4491 18955
rect 4798 18952 4804 18964
rect 4479 18924 4804 18952
rect 4479 18921 4491 18924
rect 4433 18915 4491 18921
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 4893 18955 4951 18961
rect 4893 18921 4905 18955
rect 4939 18952 4951 18955
rect 5074 18952 5080 18964
rect 4939 18924 5080 18952
rect 4939 18921 4951 18924
rect 4893 18915 4951 18921
rect 5074 18912 5080 18924
rect 5132 18912 5138 18964
rect 5350 18952 5356 18964
rect 5311 18924 5356 18952
rect 5350 18912 5356 18924
rect 5408 18912 5414 18964
rect 5810 18952 5816 18964
rect 5771 18924 5816 18952
rect 5810 18912 5816 18924
rect 5868 18912 5874 18964
rect 6273 18955 6331 18961
rect 6273 18921 6285 18955
rect 6319 18952 6331 18955
rect 6546 18952 6552 18964
rect 6319 18924 6552 18952
rect 6319 18921 6331 18924
rect 6273 18915 6331 18921
rect 6546 18912 6552 18924
rect 6604 18912 6610 18964
rect 7098 18952 7104 18964
rect 6748 18924 7104 18952
rect 1949 18887 2007 18893
rect 1949 18853 1961 18887
rect 1995 18884 2007 18887
rect 6638 18884 6644 18896
rect 1995 18856 6644 18884
rect 1995 18853 2007 18856
rect 1949 18847 2007 18853
rect 6638 18844 6644 18856
rect 6696 18844 6702 18896
rect 4062 18816 4068 18828
rect 4023 18788 4068 18816
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 4890 18776 4896 18828
rect 4948 18816 4954 18828
rect 6748 18816 6776 18924
rect 7098 18912 7104 18924
rect 7156 18912 7162 18964
rect 7193 18955 7251 18961
rect 7193 18921 7205 18955
rect 7239 18952 7251 18955
rect 7466 18952 7472 18964
rect 7239 18924 7472 18952
rect 7239 18921 7251 18924
rect 7193 18915 7251 18921
rect 7466 18912 7472 18924
rect 7524 18912 7530 18964
rect 8113 18955 8171 18961
rect 8113 18921 8125 18955
rect 8159 18952 8171 18955
rect 8202 18952 8208 18964
rect 8159 18924 8208 18952
rect 8159 18921 8171 18924
rect 8113 18915 8171 18921
rect 8202 18912 8208 18924
rect 8260 18912 8266 18964
rect 8570 18912 8576 18964
rect 8628 18952 8634 18964
rect 8628 18924 10180 18952
rect 8628 18912 8634 18924
rect 6822 18844 6828 18896
rect 6880 18884 6886 18896
rect 8478 18884 8484 18896
rect 6880 18856 8484 18884
rect 6880 18844 6886 18856
rect 8478 18844 8484 18856
rect 8536 18844 8542 18896
rect 10152 18884 10180 18924
rect 10226 18912 10232 18964
rect 10284 18952 10290 18964
rect 10594 18952 10600 18964
rect 10284 18924 10600 18952
rect 10284 18912 10290 18924
rect 10594 18912 10600 18924
rect 10652 18912 10658 18964
rect 12250 18952 12256 18964
rect 11532 18924 12256 18952
rect 10410 18884 10416 18896
rect 10152 18856 10416 18884
rect 10410 18844 10416 18856
rect 10468 18844 10474 18896
rect 11054 18816 11060 18828
rect 4948 18788 6776 18816
rect 7484 18788 9168 18816
rect 4948 18776 4954 18788
rect 4706 18748 4712 18760
rect 4667 18720 4712 18748
rect 4706 18708 4712 18720
rect 4764 18708 4770 18760
rect 5166 18748 5172 18760
rect 5127 18720 5172 18748
rect 5166 18708 5172 18720
rect 5224 18708 5230 18760
rect 5350 18708 5356 18760
rect 5408 18748 5414 18760
rect 5629 18751 5687 18757
rect 5629 18748 5641 18751
rect 5408 18720 5641 18748
rect 5408 18708 5414 18720
rect 5629 18717 5641 18720
rect 5675 18717 5687 18751
rect 6089 18751 6147 18757
rect 6089 18748 6101 18751
rect 5629 18711 5687 18717
rect 5736 18720 6101 18748
rect 1854 18640 1860 18692
rect 1912 18680 1918 18692
rect 4798 18680 4804 18692
rect 1912 18652 4804 18680
rect 1912 18640 1918 18652
rect 4798 18640 4804 18652
rect 4856 18640 4862 18692
rect 4890 18640 4896 18692
rect 4948 18680 4954 18692
rect 5736 18680 5764 18720
rect 6089 18717 6101 18720
rect 6135 18717 6147 18751
rect 6089 18711 6147 18717
rect 6454 18708 6460 18760
rect 6512 18748 6518 18760
rect 6549 18751 6607 18757
rect 6549 18748 6561 18751
rect 6512 18720 6561 18748
rect 6512 18708 6518 18720
rect 6549 18717 6561 18720
rect 6595 18748 6607 18751
rect 6638 18748 6644 18760
rect 6595 18720 6644 18748
rect 6595 18717 6607 18720
rect 6549 18711 6607 18717
rect 6638 18708 6644 18720
rect 6696 18708 6702 18760
rect 7484 18757 7512 18788
rect 7009 18751 7067 18757
rect 7009 18717 7021 18751
rect 7055 18717 7067 18751
rect 7009 18711 7067 18717
rect 7469 18751 7527 18757
rect 7469 18717 7481 18751
rect 7515 18717 7527 18751
rect 7469 18711 7527 18717
rect 7929 18751 7987 18757
rect 7929 18717 7941 18751
rect 7975 18748 7987 18751
rect 8570 18748 8576 18760
rect 7975 18720 8432 18748
rect 8531 18720 8576 18748
rect 7975 18717 7987 18720
rect 7929 18711 7987 18717
rect 4948 18652 5764 18680
rect 7024 18680 7052 18711
rect 8294 18680 8300 18692
rect 7024 18652 8300 18680
rect 4948 18640 4954 18652
rect 8294 18640 8300 18652
rect 8352 18640 8358 18692
rect 2317 18615 2375 18621
rect 2317 18581 2329 18615
rect 2363 18612 2375 18615
rect 2406 18612 2412 18624
rect 2363 18584 2412 18612
rect 2363 18581 2375 18584
rect 2317 18575 2375 18581
rect 2406 18572 2412 18584
rect 2464 18572 2470 18624
rect 3421 18615 3479 18621
rect 3421 18581 3433 18615
rect 3467 18612 3479 18615
rect 4706 18612 4712 18624
rect 3467 18584 4712 18612
rect 3467 18581 3479 18584
rect 3421 18575 3479 18581
rect 4706 18572 4712 18584
rect 4764 18572 4770 18624
rect 6733 18615 6791 18621
rect 6733 18581 6745 18615
rect 6779 18612 6791 18615
rect 7374 18612 7380 18624
rect 6779 18584 7380 18612
rect 6779 18581 6791 18584
rect 6733 18575 6791 18581
rect 7374 18572 7380 18584
rect 7432 18572 7438 18624
rect 7650 18612 7656 18624
rect 7611 18584 7656 18612
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 8404 18621 8432 18720
rect 8570 18708 8576 18720
rect 8628 18708 8634 18760
rect 8389 18615 8447 18621
rect 8389 18581 8401 18615
rect 8435 18581 8447 18615
rect 9140 18612 9168 18788
rect 10612 18788 11060 18816
rect 9217 18751 9275 18757
rect 9217 18717 9229 18751
rect 9263 18748 9275 18751
rect 9766 18748 9772 18760
rect 9263 18720 9772 18748
rect 9263 18717 9275 18720
rect 9217 18711 9275 18717
rect 9766 18708 9772 18720
rect 9824 18748 9830 18760
rect 9950 18748 9956 18760
rect 9824 18720 9956 18748
rect 9824 18708 9830 18720
rect 9950 18708 9956 18720
rect 10008 18708 10014 18760
rect 9484 18683 9542 18689
rect 9484 18649 9496 18683
rect 9530 18680 9542 18683
rect 10612 18680 10640 18788
rect 11054 18776 11060 18788
rect 11112 18776 11118 18828
rect 11532 18825 11560 18924
rect 12250 18912 12256 18924
rect 12308 18912 12314 18964
rect 12986 18912 12992 18964
rect 13044 18952 13050 18964
rect 13265 18955 13323 18961
rect 13265 18952 13277 18955
rect 13044 18924 13277 18952
rect 13044 18912 13050 18924
rect 13265 18921 13277 18924
rect 13311 18921 13323 18955
rect 13265 18915 13323 18921
rect 13725 18955 13783 18961
rect 13725 18921 13737 18955
rect 13771 18952 13783 18955
rect 16942 18952 16948 18964
rect 13771 18924 16948 18952
rect 13771 18921 13783 18924
rect 13725 18915 13783 18921
rect 16942 18912 16948 18924
rect 17000 18912 17006 18964
rect 18690 18912 18696 18964
rect 18748 18952 18754 18964
rect 18785 18955 18843 18961
rect 18785 18952 18797 18955
rect 18748 18924 18797 18952
rect 18748 18912 18754 18924
rect 18785 18921 18797 18924
rect 18831 18921 18843 18955
rect 18785 18915 18843 18921
rect 12894 18844 12900 18896
rect 12952 18884 12958 18896
rect 14550 18884 14556 18896
rect 12952 18856 14556 18884
rect 12952 18844 12958 18856
rect 14550 18844 14556 18856
rect 14608 18844 14614 18896
rect 11517 18819 11575 18825
rect 11517 18785 11529 18819
rect 11563 18785 11575 18819
rect 14366 18816 14372 18828
rect 14327 18788 14372 18816
rect 11517 18779 11575 18785
rect 14366 18776 14372 18788
rect 14424 18776 14430 18828
rect 16408 18788 20484 18816
rect 10962 18708 10968 18760
rect 11020 18748 11026 18760
rect 11882 18748 11888 18760
rect 11020 18720 11888 18748
rect 11020 18708 11026 18720
rect 11882 18708 11888 18720
rect 11940 18748 11946 18760
rect 13078 18748 13084 18760
rect 11940 18720 13084 18748
rect 11940 18708 11946 18720
rect 13078 18708 13084 18720
rect 13136 18708 13142 18760
rect 13538 18748 13544 18760
rect 13499 18720 13544 18748
rect 13538 18708 13544 18720
rect 13596 18708 13602 18760
rect 13722 18708 13728 18760
rect 13780 18748 13786 18760
rect 14461 18751 14519 18757
rect 14461 18748 14473 18751
rect 13780 18720 14473 18748
rect 13780 18708 13786 18720
rect 14461 18717 14473 18720
rect 14507 18717 14519 18751
rect 15378 18748 15384 18760
rect 15291 18720 15384 18748
rect 14461 18711 14519 18717
rect 15378 18708 15384 18720
rect 15436 18748 15442 18760
rect 16114 18748 16120 18760
rect 15436 18720 16120 18748
rect 15436 18708 15442 18720
rect 16114 18708 16120 18720
rect 16172 18708 16178 18760
rect 10778 18680 10784 18692
rect 9530 18652 10640 18680
rect 10704 18652 10784 18680
rect 9530 18649 9542 18652
rect 9484 18643 9542 18649
rect 10704 18612 10732 18652
rect 10778 18640 10784 18652
rect 10836 18640 10842 18692
rect 11238 18680 11244 18692
rect 11199 18652 11244 18680
rect 11238 18640 11244 18652
rect 11296 18640 11302 18692
rect 12152 18683 12210 18689
rect 12152 18649 12164 18683
rect 12198 18680 12210 18683
rect 13262 18680 13268 18692
rect 12198 18652 13268 18680
rect 12198 18649 12210 18652
rect 12152 18643 12210 18649
rect 13262 18640 13268 18652
rect 13320 18640 13326 18692
rect 15470 18680 15476 18692
rect 13648 18652 15476 18680
rect 10870 18612 10876 18624
rect 9140 18584 10732 18612
rect 10831 18584 10876 18612
rect 8389 18575 8447 18581
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 11333 18615 11391 18621
rect 11333 18581 11345 18615
rect 11379 18612 11391 18615
rect 11698 18612 11704 18624
rect 11379 18584 11704 18612
rect 11379 18581 11391 18584
rect 11333 18575 11391 18581
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 11790 18572 11796 18624
rect 11848 18612 11854 18624
rect 13648 18612 13676 18652
rect 15470 18640 15476 18652
rect 15528 18640 15534 18692
rect 15648 18683 15706 18689
rect 15648 18649 15660 18683
rect 15694 18680 15706 18683
rect 15746 18680 15752 18692
rect 15694 18652 15752 18680
rect 15694 18649 15706 18652
rect 15648 18643 15706 18649
rect 15746 18640 15752 18652
rect 15804 18640 15810 18692
rect 16408 18680 16436 18788
rect 17218 18748 17224 18760
rect 17179 18720 17224 18748
rect 17218 18708 17224 18720
rect 17276 18708 17282 18760
rect 18046 18708 18052 18760
rect 18104 18748 18110 18760
rect 18141 18751 18199 18757
rect 18141 18748 18153 18751
rect 18104 18720 18153 18748
rect 18104 18708 18110 18720
rect 18141 18717 18153 18720
rect 18187 18717 18199 18751
rect 18141 18711 18199 18717
rect 18414 18708 18420 18760
rect 18472 18748 18478 18760
rect 18601 18751 18659 18757
rect 18601 18748 18613 18751
rect 18472 18720 18613 18748
rect 18472 18708 18478 18720
rect 18601 18717 18613 18720
rect 18647 18717 18659 18751
rect 18601 18711 18659 18717
rect 19518 18708 19524 18760
rect 19576 18748 19582 18760
rect 20456 18757 20484 18788
rect 19981 18751 20039 18757
rect 19981 18748 19993 18751
rect 19576 18720 19993 18748
rect 19576 18708 19582 18720
rect 19981 18717 19993 18720
rect 20027 18717 20039 18751
rect 19981 18711 20039 18717
rect 20441 18751 20499 18757
rect 20441 18717 20453 18751
rect 20487 18717 20499 18751
rect 20441 18711 20499 18717
rect 20898 18708 20904 18760
rect 20956 18748 20962 18760
rect 21361 18751 21419 18757
rect 21361 18748 21373 18751
rect 20956 18720 21373 18748
rect 20956 18708 20962 18720
rect 21361 18717 21373 18720
rect 21407 18717 21419 18751
rect 21361 18711 21419 18717
rect 15856 18652 16436 18680
rect 11848 18584 13676 18612
rect 11848 18572 11854 18584
rect 14458 18572 14464 18624
rect 14516 18612 14522 18624
rect 14553 18615 14611 18621
rect 14553 18612 14565 18615
rect 14516 18584 14565 18612
rect 14516 18572 14522 18584
rect 14553 18581 14565 18584
rect 14599 18581 14611 18615
rect 14918 18612 14924 18624
rect 14879 18584 14924 18612
rect 14553 18575 14611 18581
rect 14918 18572 14924 18584
rect 14976 18572 14982 18624
rect 15010 18572 15016 18624
rect 15068 18612 15074 18624
rect 15856 18612 15884 18652
rect 16482 18640 16488 18692
rect 16540 18680 16546 18692
rect 18690 18680 18696 18692
rect 16540 18652 18696 18680
rect 16540 18640 16546 18652
rect 18690 18640 18696 18652
rect 18748 18640 18754 18692
rect 19702 18640 19708 18692
rect 19760 18680 19766 18692
rect 20717 18683 20775 18689
rect 20717 18680 20729 18683
rect 19760 18652 20729 18680
rect 19760 18640 19766 18652
rect 20717 18649 20729 18652
rect 20763 18649 20775 18683
rect 20717 18643 20775 18649
rect 15068 18584 15884 18612
rect 15068 18572 15074 18584
rect 16390 18572 16396 18624
rect 16448 18612 16454 18624
rect 16761 18615 16819 18621
rect 16761 18612 16773 18615
rect 16448 18584 16773 18612
rect 16448 18572 16454 18584
rect 16761 18581 16773 18584
rect 16807 18581 16819 18615
rect 16761 18575 16819 18581
rect 16942 18572 16948 18624
rect 17000 18612 17006 18624
rect 17037 18615 17095 18621
rect 17037 18612 17049 18615
rect 17000 18584 17049 18612
rect 17000 18572 17006 18584
rect 17037 18581 17049 18584
rect 17083 18581 17095 18615
rect 17037 18575 17095 18581
rect 17310 18572 17316 18624
rect 17368 18612 17374 18624
rect 17497 18615 17555 18621
rect 17497 18612 17509 18615
rect 17368 18584 17509 18612
rect 17368 18572 17374 18584
rect 17497 18581 17509 18584
rect 17543 18581 17555 18615
rect 17497 18575 17555 18581
rect 18966 18572 18972 18624
rect 19024 18612 19030 18624
rect 19337 18615 19395 18621
rect 19337 18612 19349 18615
rect 19024 18584 19349 18612
rect 19024 18572 19030 18584
rect 19337 18581 19349 18584
rect 19383 18581 19395 18615
rect 20254 18612 20260 18624
rect 20215 18584 20260 18612
rect 19337 18575 19395 18581
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 1104 18522 21896 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21896 18522
rect 1104 18448 21896 18470
rect 2130 18408 2136 18420
rect 2091 18380 2136 18408
rect 2130 18368 2136 18380
rect 2188 18368 2194 18420
rect 2866 18408 2872 18420
rect 2827 18380 2872 18408
rect 2866 18368 2872 18380
rect 2924 18408 2930 18420
rect 4062 18408 4068 18420
rect 2924 18380 4068 18408
rect 2924 18368 2930 18380
rect 4062 18368 4068 18380
rect 4120 18368 4126 18420
rect 5902 18408 5908 18420
rect 5552 18380 5908 18408
rect 1765 18343 1823 18349
rect 1765 18309 1777 18343
rect 1811 18340 1823 18343
rect 4154 18340 4160 18352
rect 1811 18312 4160 18340
rect 1811 18309 1823 18312
rect 1765 18303 1823 18309
rect 4154 18300 4160 18312
rect 4212 18300 4218 18352
rect 4341 18343 4399 18349
rect 4341 18309 4353 18343
rect 4387 18340 4399 18343
rect 5350 18340 5356 18352
rect 4387 18312 5356 18340
rect 4387 18309 4399 18312
rect 4341 18303 4399 18309
rect 5350 18300 5356 18312
rect 5408 18300 5414 18352
rect 5552 18349 5580 18380
rect 5902 18368 5908 18380
rect 5960 18368 5966 18420
rect 5997 18411 6055 18417
rect 5997 18377 6009 18411
rect 6043 18408 6055 18411
rect 6546 18408 6552 18420
rect 6043 18380 6552 18408
rect 6043 18377 6055 18380
rect 5997 18371 6055 18377
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 7282 18408 7288 18420
rect 7243 18380 7288 18408
rect 7282 18368 7288 18380
rect 7340 18368 7346 18420
rect 8297 18411 8355 18417
rect 8297 18377 8309 18411
rect 8343 18408 8355 18411
rect 9030 18408 9036 18420
rect 8343 18380 9036 18408
rect 8343 18377 8355 18380
rect 8297 18371 8355 18377
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 9306 18368 9312 18420
rect 9364 18408 9370 18420
rect 10226 18408 10232 18420
rect 9364 18380 10232 18408
rect 9364 18368 9370 18380
rect 10226 18368 10232 18380
rect 10284 18368 10290 18420
rect 10502 18408 10508 18420
rect 10463 18380 10508 18408
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 10778 18368 10784 18420
rect 10836 18408 10842 18420
rect 11517 18411 11575 18417
rect 10836 18380 11284 18408
rect 10836 18368 10842 18380
rect 5537 18343 5595 18349
rect 5537 18309 5549 18343
rect 5583 18309 5595 18343
rect 7006 18340 7012 18352
rect 5537 18303 5595 18309
rect 5736 18312 7012 18340
rect 2501 18275 2559 18281
rect 2501 18241 2513 18275
rect 2547 18272 2559 18275
rect 5626 18272 5632 18284
rect 2547 18244 5632 18272
rect 2547 18241 2559 18244
rect 2501 18235 2559 18241
rect 5626 18232 5632 18244
rect 5684 18232 5690 18284
rect 3234 18204 3240 18216
rect 3195 18176 3240 18204
rect 3234 18164 3240 18176
rect 3292 18164 3298 18216
rect 3973 18207 4031 18213
rect 3973 18173 3985 18207
rect 4019 18204 4031 18207
rect 5736 18204 5764 18312
rect 6656 18281 6684 18312
rect 7006 18300 7012 18312
rect 7064 18300 7070 18352
rect 7190 18300 7196 18352
rect 7248 18340 7254 18352
rect 7929 18343 7987 18349
rect 7929 18340 7941 18343
rect 7248 18312 7941 18340
rect 7248 18300 7254 18312
rect 7929 18309 7941 18312
rect 7975 18309 7987 18343
rect 7929 18303 7987 18309
rect 8202 18300 8208 18352
rect 8260 18340 8266 18352
rect 8662 18340 8668 18352
rect 8260 18312 8668 18340
rect 8260 18300 8266 18312
rect 8662 18300 8668 18312
rect 8720 18300 8726 18352
rect 8956 18312 9628 18340
rect 5813 18275 5871 18281
rect 5813 18241 5825 18275
rect 5859 18241 5871 18275
rect 5813 18235 5871 18241
rect 6641 18275 6699 18281
rect 6641 18241 6653 18275
rect 6687 18241 6699 18275
rect 6641 18235 6699 18241
rect 4019 18176 5764 18204
rect 5828 18204 5856 18235
rect 6730 18232 6736 18284
rect 6788 18272 6794 18284
rect 8956 18281 8984 18312
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 6788 18244 7849 18272
rect 6788 18232 6794 18244
rect 7837 18241 7849 18244
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 8941 18275 8999 18281
rect 8941 18241 8953 18275
rect 8987 18241 8999 18275
rect 8941 18235 8999 18241
rect 9030 18232 9036 18284
rect 9088 18272 9094 18284
rect 9490 18272 9496 18284
rect 9088 18244 9496 18272
rect 9088 18232 9094 18244
rect 9490 18232 9496 18244
rect 9548 18232 9554 18284
rect 9600 18272 9628 18312
rect 9674 18300 9680 18352
rect 9732 18340 9738 18352
rect 9769 18343 9827 18349
rect 9769 18340 9781 18343
rect 9732 18312 9781 18340
rect 9732 18300 9738 18312
rect 9769 18309 9781 18312
rect 9815 18309 9827 18343
rect 9769 18303 9827 18309
rect 10594 18300 10600 18352
rect 10652 18340 10658 18352
rect 11256 18340 11284 18380
rect 11517 18377 11529 18411
rect 11563 18408 11575 18411
rect 11698 18408 11704 18420
rect 11563 18380 11704 18408
rect 11563 18377 11575 18380
rect 11517 18371 11575 18377
rect 11698 18368 11704 18380
rect 11756 18368 11762 18420
rect 11882 18368 11888 18420
rect 11940 18408 11946 18420
rect 12250 18408 12256 18420
rect 11940 18380 12256 18408
rect 11940 18368 11946 18380
rect 12250 18368 12256 18380
rect 12308 18368 12314 18420
rect 12894 18408 12900 18420
rect 12855 18380 12900 18408
rect 12894 18368 12900 18380
rect 12952 18368 12958 18420
rect 13630 18368 13636 18420
rect 13688 18408 13694 18420
rect 13909 18411 13967 18417
rect 13909 18408 13921 18411
rect 13688 18380 13921 18408
rect 13688 18368 13694 18380
rect 13909 18377 13921 18380
rect 13955 18377 13967 18411
rect 13909 18371 13967 18377
rect 14737 18411 14795 18417
rect 14737 18377 14749 18411
rect 14783 18377 14795 18411
rect 14737 18371 14795 18377
rect 14752 18340 14780 18371
rect 14918 18368 14924 18420
rect 14976 18408 14982 18420
rect 15197 18411 15255 18417
rect 15197 18408 15209 18411
rect 14976 18380 15209 18408
rect 14976 18368 14982 18380
rect 15197 18377 15209 18380
rect 15243 18377 15255 18411
rect 15197 18371 15255 18377
rect 15470 18368 15476 18420
rect 15528 18408 15534 18420
rect 17129 18411 17187 18417
rect 17129 18408 17141 18411
rect 15528 18380 17141 18408
rect 15528 18368 15534 18380
rect 17129 18377 17141 18380
rect 17175 18377 17187 18411
rect 17129 18371 17187 18377
rect 17402 18368 17408 18420
rect 17460 18408 17466 18420
rect 18598 18408 18604 18420
rect 17460 18380 18604 18408
rect 17460 18368 17466 18380
rect 18598 18368 18604 18380
rect 18656 18368 18662 18420
rect 18690 18368 18696 18420
rect 18748 18408 18754 18420
rect 19889 18411 19947 18417
rect 19889 18408 19901 18411
rect 18748 18380 19901 18408
rect 18748 18368 18754 18380
rect 19889 18377 19901 18380
rect 19935 18377 19947 18411
rect 19889 18371 19947 18377
rect 20717 18411 20775 18417
rect 20717 18377 20729 18411
rect 20763 18408 20775 18411
rect 20806 18408 20812 18420
rect 20763 18380 20812 18408
rect 20763 18377 20775 18380
rect 20717 18371 20775 18377
rect 20806 18368 20812 18380
rect 20864 18368 20870 18420
rect 10652 18312 11192 18340
rect 11256 18312 14780 18340
rect 15105 18343 15163 18349
rect 10652 18300 10658 18312
rect 10870 18272 10876 18284
rect 9600 18244 10876 18272
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 11164 18281 11192 18312
rect 15105 18309 15117 18343
rect 15151 18340 15163 18343
rect 15286 18340 15292 18352
rect 15151 18312 15292 18340
rect 15151 18309 15163 18312
rect 15105 18303 15163 18309
rect 15286 18300 15292 18312
rect 15344 18300 15350 18352
rect 16298 18340 16304 18352
rect 15396 18312 16304 18340
rect 11149 18275 11207 18281
rect 11149 18241 11161 18275
rect 11195 18241 11207 18275
rect 11882 18272 11888 18284
rect 11843 18244 11888 18272
rect 11149 18235 11207 18241
rect 11882 18232 11888 18244
rect 11940 18232 11946 18284
rect 12710 18272 12716 18284
rect 12671 18244 12716 18272
rect 12710 18232 12716 18244
rect 12768 18232 12774 18284
rect 12986 18232 12992 18284
rect 13044 18272 13050 18284
rect 13265 18275 13323 18281
rect 13265 18272 13277 18275
rect 13044 18244 13277 18272
rect 13044 18232 13050 18244
rect 13265 18241 13277 18244
rect 13311 18241 13323 18275
rect 13265 18235 13323 18241
rect 14185 18275 14243 18281
rect 14185 18241 14197 18275
rect 14231 18272 14243 18275
rect 14274 18272 14280 18284
rect 14231 18244 14280 18272
rect 14231 18241 14243 18244
rect 14185 18235 14243 18241
rect 14274 18232 14280 18244
rect 14332 18232 14338 18284
rect 14918 18232 14924 18284
rect 14976 18272 14982 18284
rect 15396 18272 15424 18312
rect 16298 18300 16304 18312
rect 16356 18300 16362 18352
rect 16390 18300 16396 18352
rect 16448 18340 16454 18352
rect 19794 18340 19800 18352
rect 16448 18312 19800 18340
rect 16448 18300 16454 18312
rect 16022 18272 16028 18284
rect 14976 18244 15424 18272
rect 15983 18244 16028 18272
rect 14976 18232 14982 18244
rect 16022 18232 16028 18244
rect 16080 18232 16086 18284
rect 7098 18204 7104 18216
rect 5828 18176 7104 18204
rect 4019 18173 4031 18176
rect 3973 18167 4031 18173
rect 7098 18164 7104 18176
rect 7156 18164 7162 18216
rect 7282 18164 7288 18216
rect 7340 18204 7346 18216
rect 7653 18207 7711 18213
rect 7653 18204 7665 18207
rect 7340 18176 7665 18204
rect 7340 18164 7346 18176
rect 7653 18173 7665 18176
rect 7699 18173 7711 18207
rect 7653 18167 7711 18173
rect 8662 18164 8668 18216
rect 8720 18204 8726 18216
rect 9398 18204 9404 18216
rect 8720 18176 9404 18204
rect 8720 18164 8726 18176
rect 9398 18164 9404 18176
rect 9456 18164 9462 18216
rect 9585 18207 9643 18213
rect 9585 18173 9597 18207
rect 9631 18173 9643 18207
rect 9585 18167 9643 18173
rect 9677 18207 9735 18213
rect 9677 18173 9689 18207
rect 9723 18204 9735 18207
rect 10594 18204 10600 18216
rect 9723 18176 10600 18204
rect 9723 18173 9735 18176
rect 9677 18167 9735 18173
rect 2682 18096 2688 18148
rect 2740 18136 2746 18148
rect 2774 18136 2780 18148
rect 2740 18108 2780 18136
rect 2740 18096 2746 18108
rect 2774 18096 2780 18108
rect 2832 18096 2838 18148
rect 3605 18139 3663 18145
rect 3605 18105 3617 18139
rect 3651 18136 3663 18139
rect 6822 18136 6828 18148
rect 3651 18108 6684 18136
rect 6783 18108 6828 18136
rect 3651 18105 3663 18108
rect 3605 18099 3663 18105
rect 4709 18071 4767 18077
rect 4709 18037 4721 18071
rect 4755 18068 4767 18071
rect 4798 18068 4804 18080
rect 4755 18040 4804 18068
rect 4755 18037 4767 18040
rect 4709 18031 4767 18037
rect 4798 18028 4804 18040
rect 4856 18028 4862 18080
rect 5074 18068 5080 18080
rect 5035 18040 5080 18068
rect 5074 18028 5080 18040
rect 5132 18028 5138 18080
rect 6656 18068 6684 18108
rect 6822 18096 6828 18108
rect 6880 18096 6886 18148
rect 7006 18096 7012 18148
rect 7064 18136 7070 18148
rect 7190 18136 7196 18148
rect 7064 18108 7196 18136
rect 7064 18096 7070 18108
rect 7190 18096 7196 18108
rect 7248 18096 7254 18148
rect 9600 18136 9628 18167
rect 10594 18164 10600 18176
rect 10652 18164 10658 18216
rect 10686 18164 10692 18216
rect 10744 18204 10750 18216
rect 11977 18207 12035 18213
rect 11977 18204 11989 18207
rect 10744 18176 11989 18204
rect 10744 18164 10750 18176
rect 11977 18173 11989 18176
rect 12023 18173 12035 18207
rect 11977 18167 12035 18173
rect 12066 18164 12072 18216
rect 12124 18204 12130 18216
rect 14366 18204 14372 18216
rect 12124 18176 12169 18204
rect 12268 18176 14372 18204
rect 12124 18164 12130 18176
rect 9766 18136 9772 18148
rect 9600 18108 9772 18136
rect 9766 18096 9772 18108
rect 9824 18096 9830 18148
rect 10502 18096 10508 18148
rect 10560 18136 10566 18148
rect 12268 18136 12296 18176
rect 14366 18164 14372 18176
rect 14424 18164 14430 18216
rect 15102 18164 15108 18216
rect 15160 18204 15166 18216
rect 15289 18207 15347 18213
rect 15289 18204 15301 18207
rect 15160 18176 15301 18204
rect 15160 18164 15166 18176
rect 15289 18173 15301 18176
rect 15335 18173 15347 18207
rect 16758 18204 16764 18216
rect 15289 18167 15347 18173
rect 15396 18176 16764 18204
rect 10560 18108 12296 18136
rect 10560 18096 10566 18108
rect 12342 18096 12348 18148
rect 12400 18136 12406 18148
rect 15396 18136 15424 18176
rect 16758 18164 16764 18176
rect 16816 18164 16822 18216
rect 16868 18213 16896 18312
rect 19794 18300 19800 18312
rect 19852 18300 19858 18352
rect 19978 18340 19984 18352
rect 19939 18312 19984 18340
rect 19978 18300 19984 18312
rect 20036 18300 20042 18352
rect 18230 18281 18236 18284
rect 18224 18272 18236 18281
rect 18191 18244 18236 18272
rect 18224 18235 18236 18244
rect 18288 18272 18294 18284
rect 18288 18244 19748 18272
rect 18230 18232 18236 18235
rect 18288 18232 18294 18244
rect 16853 18207 16911 18213
rect 16853 18173 16865 18207
rect 16899 18173 16911 18207
rect 17034 18204 17040 18216
rect 16995 18176 17040 18204
rect 16853 18167 16911 18173
rect 17034 18164 17040 18176
rect 17092 18164 17098 18216
rect 17954 18204 17960 18216
rect 17915 18176 17960 18204
rect 17954 18164 17960 18176
rect 18012 18164 18018 18216
rect 19720 18213 19748 18244
rect 20806 18232 20812 18284
rect 20864 18272 20870 18284
rect 21361 18275 21419 18281
rect 21361 18272 21373 18275
rect 20864 18244 21373 18272
rect 20864 18232 20870 18244
rect 21361 18241 21373 18244
rect 21407 18241 21419 18275
rect 21361 18235 21419 18241
rect 19705 18207 19763 18213
rect 19705 18173 19717 18207
rect 19751 18173 19763 18207
rect 19705 18167 19763 18173
rect 12400 18108 15424 18136
rect 16209 18139 16267 18145
rect 12400 18096 12406 18108
rect 16209 18105 16221 18139
rect 16255 18136 16267 18139
rect 17862 18136 17868 18148
rect 16255 18108 17868 18136
rect 16255 18105 16267 18108
rect 16209 18099 16267 18105
rect 17862 18096 17868 18108
rect 17920 18096 17926 18148
rect 7926 18068 7932 18080
rect 6656 18040 7932 18068
rect 7926 18028 7932 18040
rect 7984 18028 7990 18080
rect 8386 18028 8392 18080
rect 8444 18068 8450 18080
rect 8662 18068 8668 18080
rect 8444 18040 8668 18068
rect 8444 18028 8450 18040
rect 8662 18028 8668 18040
rect 8720 18028 8726 18080
rect 9125 18071 9183 18077
rect 9125 18037 9137 18071
rect 9171 18068 9183 18071
rect 9582 18068 9588 18080
rect 9171 18040 9588 18068
rect 9171 18037 9183 18040
rect 9125 18031 9183 18037
rect 9582 18028 9588 18040
rect 9640 18028 9646 18080
rect 10134 18068 10140 18080
rect 10095 18040 10140 18068
rect 10134 18028 10140 18040
rect 10192 18028 10198 18080
rect 10226 18028 10232 18080
rect 10284 18068 10290 18080
rect 12066 18068 12072 18080
rect 10284 18040 12072 18068
rect 10284 18028 10290 18040
rect 12066 18028 12072 18040
rect 12124 18028 12130 18080
rect 14369 18071 14427 18077
rect 14369 18037 14381 18071
rect 14415 18068 14427 18071
rect 17402 18068 17408 18080
rect 14415 18040 17408 18068
rect 14415 18037 14427 18040
rect 14369 18031 14427 18037
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 17497 18071 17555 18077
rect 17497 18037 17509 18071
rect 17543 18068 17555 18071
rect 18138 18068 18144 18080
rect 17543 18040 18144 18068
rect 17543 18037 17555 18040
rect 17497 18031 17555 18037
rect 18138 18028 18144 18040
rect 18196 18028 18202 18080
rect 19337 18071 19395 18077
rect 19337 18037 19349 18071
rect 19383 18068 19395 18071
rect 19518 18068 19524 18080
rect 19383 18040 19524 18068
rect 19383 18037 19395 18040
rect 19337 18031 19395 18037
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 20346 18068 20352 18080
rect 20307 18040 20352 18068
rect 20346 18028 20352 18040
rect 20404 18028 20410 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 5166 17864 5172 17876
rect 5127 17836 5172 17864
rect 5166 17824 5172 17836
rect 5224 17824 5230 17876
rect 6914 17864 6920 17876
rect 5460 17836 6920 17864
rect 4433 17799 4491 17805
rect 4433 17765 4445 17799
rect 4479 17796 4491 17799
rect 5460 17796 5488 17836
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 7006 17824 7012 17876
rect 7064 17864 7070 17876
rect 7101 17867 7159 17873
rect 7101 17864 7113 17867
rect 7064 17836 7113 17864
rect 7064 17824 7070 17836
rect 7101 17833 7113 17836
rect 7147 17864 7159 17867
rect 7282 17864 7288 17876
rect 7147 17836 7288 17864
rect 7147 17833 7159 17836
rect 7101 17827 7159 17833
rect 7282 17824 7288 17836
rect 7340 17824 7346 17876
rect 10594 17864 10600 17876
rect 7576 17836 10180 17864
rect 10555 17836 10600 17864
rect 4479 17768 5488 17796
rect 5537 17799 5595 17805
rect 4479 17765 4491 17768
rect 4433 17759 4491 17765
rect 5537 17765 5549 17799
rect 5583 17796 5595 17799
rect 7576 17796 7604 17836
rect 5583 17768 7604 17796
rect 10152 17796 10180 17836
rect 10594 17824 10600 17836
rect 10652 17824 10658 17876
rect 11054 17824 11060 17876
rect 11112 17864 11118 17876
rect 12253 17867 12311 17873
rect 12253 17864 12265 17867
rect 11112 17836 12265 17864
rect 11112 17824 11118 17836
rect 12253 17833 12265 17836
rect 12299 17833 12311 17867
rect 12710 17864 12716 17876
rect 12671 17836 12716 17864
rect 12253 17827 12311 17833
rect 12710 17824 12716 17836
rect 12768 17824 12774 17876
rect 13354 17824 13360 17876
rect 13412 17864 13418 17876
rect 20257 17867 20315 17873
rect 20257 17864 20269 17867
rect 13412 17836 20269 17864
rect 13412 17824 13418 17836
rect 20257 17833 20269 17836
rect 20303 17833 20315 17867
rect 20257 17827 20315 17833
rect 10962 17796 10968 17808
rect 10152 17768 10968 17796
rect 5583 17765 5595 17768
rect 5537 17759 5595 17765
rect 10962 17756 10968 17768
rect 11020 17756 11026 17808
rect 11238 17756 11244 17808
rect 11296 17796 11302 17808
rect 11296 17768 13308 17796
rect 11296 17756 11302 17768
rect 3053 17731 3111 17737
rect 3053 17697 3065 17731
rect 3099 17728 3111 17731
rect 4338 17728 4344 17740
rect 3099 17700 4344 17728
rect 3099 17697 3111 17700
rect 3053 17691 3111 17697
rect 4338 17688 4344 17700
rect 4396 17728 4402 17740
rect 5166 17728 5172 17740
rect 4396 17700 5172 17728
rect 4396 17688 4402 17700
rect 5166 17688 5172 17700
rect 5224 17688 5230 17740
rect 5828 17700 7236 17728
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 3421 17663 3479 17669
rect 1719 17632 1992 17660
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 1964 17536 1992 17632
rect 3421 17629 3433 17663
rect 3467 17660 3479 17663
rect 3510 17660 3516 17672
rect 3467 17632 3516 17660
rect 3467 17629 3479 17632
rect 3421 17623 3479 17629
rect 3510 17620 3516 17632
rect 3568 17620 3574 17672
rect 3970 17620 3976 17672
rect 4028 17660 4034 17672
rect 5626 17660 5632 17672
rect 4028 17632 5632 17660
rect 4028 17620 4034 17632
rect 5626 17620 5632 17632
rect 5684 17660 5690 17672
rect 5828 17669 5856 17700
rect 5813 17663 5871 17669
rect 5813 17660 5825 17663
rect 5684 17632 5825 17660
rect 5684 17620 5690 17632
rect 5813 17629 5825 17632
rect 5859 17629 5871 17663
rect 5813 17623 5871 17629
rect 6825 17663 6883 17669
rect 6825 17629 6837 17663
rect 6871 17660 6883 17663
rect 6914 17660 6920 17672
rect 6871 17632 6920 17660
rect 6871 17629 6883 17632
rect 6825 17623 6883 17629
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 7208 17660 7236 17700
rect 10226 17688 10232 17740
rect 10284 17728 10290 17740
rect 11149 17731 11207 17737
rect 11149 17728 11161 17731
rect 10284 17700 11161 17728
rect 10284 17688 10290 17700
rect 11149 17697 11161 17700
rect 11195 17697 11207 17731
rect 13170 17728 13176 17740
rect 13131 17700 13176 17728
rect 11149 17691 11207 17697
rect 13170 17688 13176 17700
rect 13228 17688 13234 17740
rect 13280 17737 13308 17768
rect 13538 17756 13544 17808
rect 13596 17796 13602 17808
rect 15102 17796 15108 17808
rect 13596 17768 15108 17796
rect 13596 17756 13602 17768
rect 15102 17756 15108 17768
rect 15160 17756 15166 17808
rect 17497 17799 17555 17805
rect 17497 17765 17509 17799
rect 17543 17796 17555 17799
rect 18509 17799 18567 17805
rect 17543 17768 18000 17796
rect 17543 17765 17555 17768
rect 17497 17759 17555 17765
rect 13265 17731 13323 17737
rect 13265 17697 13277 17731
rect 13311 17697 13323 17731
rect 14274 17728 14280 17740
rect 14235 17700 14280 17728
rect 13265 17691 13323 17697
rect 14274 17688 14280 17700
rect 14332 17688 14338 17740
rect 17972 17737 18000 17768
rect 18509 17765 18521 17799
rect 18555 17796 18567 17799
rect 19886 17796 19892 17808
rect 18555 17768 19892 17796
rect 18555 17765 18567 17768
rect 18509 17759 18567 17765
rect 19886 17756 19892 17768
rect 19944 17756 19950 17808
rect 19978 17756 19984 17808
rect 20036 17796 20042 17808
rect 20036 17768 20081 17796
rect 20036 17756 20042 17768
rect 17957 17731 18015 17737
rect 17957 17697 17969 17731
rect 18003 17728 18015 17731
rect 18046 17728 18052 17740
rect 18003 17700 18052 17728
rect 18003 17697 18015 17700
rect 17957 17691 18015 17697
rect 18046 17688 18052 17700
rect 18104 17688 18110 17740
rect 18230 17688 18236 17740
rect 18288 17728 18294 17740
rect 19337 17731 19395 17737
rect 19337 17728 19349 17731
rect 18288 17700 19349 17728
rect 18288 17688 18294 17700
rect 19337 17697 19349 17700
rect 19383 17697 19395 17731
rect 19337 17691 19395 17697
rect 19518 17688 19524 17740
rect 19576 17728 19582 17740
rect 20809 17731 20867 17737
rect 20809 17728 20821 17731
rect 19576 17700 20821 17728
rect 19576 17688 19582 17700
rect 20809 17697 20821 17700
rect 20855 17697 20867 17731
rect 20809 17691 20867 17697
rect 8386 17660 8392 17672
rect 7208 17632 8392 17660
rect 8386 17620 8392 17632
rect 8444 17620 8450 17672
rect 8481 17663 8539 17669
rect 8481 17629 8493 17663
rect 8527 17660 8539 17663
rect 8941 17663 8999 17669
rect 8941 17660 8953 17663
rect 8527 17632 8953 17660
rect 8527 17629 8539 17632
rect 8481 17623 8539 17629
rect 8941 17629 8953 17632
rect 8987 17660 8999 17663
rect 9950 17660 9956 17672
rect 8987 17632 9956 17660
rect 8987 17629 8999 17632
rect 8941 17623 8999 17629
rect 9950 17620 9956 17632
rect 10008 17620 10014 17672
rect 10318 17620 10324 17672
rect 10376 17660 10382 17672
rect 11609 17663 11667 17669
rect 11609 17660 11621 17663
rect 10376 17632 11621 17660
rect 10376 17620 10382 17632
rect 11609 17629 11621 17632
rect 11655 17629 11667 17663
rect 11609 17623 11667 17629
rect 11698 17620 11704 17672
rect 11756 17660 11762 17672
rect 12529 17663 12587 17669
rect 12529 17660 12541 17663
rect 11756 17632 12541 17660
rect 11756 17620 11762 17632
rect 12529 17629 12541 17632
rect 12575 17660 12587 17663
rect 13814 17660 13820 17672
rect 12575 17632 13820 17660
rect 12575 17629 12587 17632
rect 12529 17623 12587 17629
rect 13814 17620 13820 17632
rect 13872 17620 13878 17672
rect 14550 17620 14556 17672
rect 14608 17660 14614 17672
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 14608 17632 15761 17660
rect 14608 17620 14614 17632
rect 15749 17629 15761 17632
rect 15795 17629 15807 17663
rect 16114 17660 16120 17672
rect 16075 17632 16120 17660
rect 15749 17623 15807 17629
rect 16114 17620 16120 17632
rect 16172 17620 16178 17672
rect 16390 17669 16396 17672
rect 16384 17660 16396 17669
rect 16351 17632 16396 17660
rect 16384 17623 16396 17632
rect 16390 17620 16396 17623
rect 16448 17620 16454 17672
rect 18138 17660 18144 17672
rect 18099 17632 18144 17660
rect 18138 17620 18144 17632
rect 18196 17620 18202 17672
rect 20346 17620 20352 17672
rect 20404 17660 20410 17672
rect 20625 17663 20683 17669
rect 20625 17660 20637 17663
rect 20404 17632 20637 17660
rect 20404 17620 20410 17632
rect 20625 17629 20637 17632
rect 20671 17629 20683 17663
rect 20625 17623 20683 17629
rect 6730 17592 6736 17604
rect 4724 17564 6736 17592
rect 4724 17536 4752 17564
rect 6730 17552 6736 17564
rect 6788 17552 6794 17604
rect 7006 17552 7012 17604
rect 7064 17592 7070 17604
rect 8214 17595 8272 17601
rect 8214 17592 8226 17595
rect 7064 17564 8226 17592
rect 7064 17552 7070 17564
rect 8214 17561 8226 17564
rect 8260 17561 8272 17595
rect 8214 17555 8272 17561
rect 9208 17595 9266 17601
rect 9208 17561 9220 17595
rect 9254 17592 9266 17595
rect 9254 17564 9444 17592
rect 9254 17561 9266 17564
rect 9208 17555 9266 17561
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 1946 17524 1952 17536
rect 1907 17496 1952 17524
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 2682 17524 2688 17536
rect 2643 17496 2688 17524
rect 2682 17484 2688 17496
rect 2740 17484 2746 17536
rect 4065 17527 4123 17533
rect 4065 17493 4077 17527
rect 4111 17524 4123 17527
rect 4246 17524 4252 17536
rect 4111 17496 4252 17524
rect 4111 17493 4123 17496
rect 4065 17487 4123 17493
rect 4246 17484 4252 17496
rect 4304 17484 4310 17536
rect 4706 17524 4712 17536
rect 4667 17496 4712 17524
rect 4706 17484 4712 17496
rect 4764 17484 4770 17536
rect 6181 17527 6239 17533
rect 6181 17493 6193 17527
rect 6227 17524 6239 17527
rect 8110 17524 8116 17536
rect 6227 17496 8116 17524
rect 6227 17493 6239 17496
rect 6181 17487 6239 17493
rect 8110 17484 8116 17496
rect 8168 17484 8174 17536
rect 9416 17524 9444 17564
rect 9490 17552 9496 17604
rect 9548 17592 9554 17604
rect 11057 17595 11115 17601
rect 11057 17592 11069 17595
rect 9548 17564 11069 17592
rect 9548 17552 9554 17564
rect 11057 17561 11069 17564
rect 11103 17561 11115 17595
rect 11057 17555 11115 17561
rect 11330 17552 11336 17604
rect 11388 17592 11394 17604
rect 13357 17595 13415 17601
rect 13357 17592 13369 17595
rect 11388 17564 13369 17592
rect 11388 17552 11394 17564
rect 13357 17561 13369 17564
rect 13403 17561 13415 17595
rect 13357 17555 13415 17561
rect 13630 17552 13636 17604
rect 13688 17592 13694 17604
rect 15105 17595 15163 17601
rect 15105 17592 15117 17595
rect 13688 17564 15117 17592
rect 13688 17552 13694 17564
rect 15105 17561 15117 17564
rect 15151 17561 15163 17595
rect 15105 17555 15163 17561
rect 16298 17552 16304 17604
rect 16356 17592 16362 17604
rect 18785 17595 18843 17601
rect 18785 17592 18797 17595
rect 16356 17564 18797 17592
rect 16356 17552 16362 17564
rect 18785 17561 18797 17564
rect 18831 17561 18843 17595
rect 19518 17592 19524 17604
rect 19479 17564 19524 17592
rect 18785 17555 18843 17561
rect 19518 17552 19524 17564
rect 19576 17552 19582 17604
rect 19978 17552 19984 17604
rect 20036 17592 20042 17604
rect 20717 17595 20775 17601
rect 20717 17592 20729 17595
rect 20036 17564 20729 17592
rect 20036 17552 20042 17564
rect 20717 17561 20729 17564
rect 20763 17561 20775 17595
rect 21542 17592 21548 17604
rect 20717 17555 20775 17561
rect 21192 17564 21548 17592
rect 10226 17524 10232 17536
rect 9416 17496 10232 17524
rect 10226 17484 10232 17496
rect 10284 17484 10290 17536
rect 10318 17484 10324 17536
rect 10376 17524 10382 17536
rect 10962 17524 10968 17536
rect 10376 17496 10421 17524
rect 10875 17496 10968 17524
rect 10376 17484 10382 17496
rect 10962 17484 10968 17496
rect 11020 17524 11026 17536
rect 13538 17524 13544 17536
rect 11020 17496 13544 17524
rect 11020 17484 11026 17496
rect 13538 17484 13544 17496
rect 13596 17484 13602 17536
rect 13725 17527 13783 17533
rect 13725 17493 13737 17527
rect 13771 17524 13783 17527
rect 14369 17527 14427 17533
rect 14369 17524 14381 17527
rect 13771 17496 14381 17524
rect 13771 17493 13783 17496
rect 13725 17487 13783 17493
rect 14369 17493 14381 17496
rect 14415 17493 14427 17527
rect 14369 17487 14427 17493
rect 14458 17484 14464 17536
rect 14516 17524 14522 17536
rect 14826 17524 14832 17536
rect 14516 17496 14561 17524
rect 14787 17496 14832 17524
rect 14516 17484 14522 17496
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 18046 17524 18052 17536
rect 18007 17496 18052 17524
rect 18046 17484 18052 17496
rect 18104 17484 18110 17536
rect 18138 17484 18144 17536
rect 18196 17524 18202 17536
rect 19613 17527 19671 17533
rect 19613 17524 19625 17527
rect 18196 17496 19625 17524
rect 18196 17484 18202 17496
rect 19613 17493 19625 17496
rect 19659 17524 19671 17527
rect 21192 17524 21220 17564
rect 21542 17552 21548 17564
rect 21600 17552 21606 17604
rect 19659 17496 21220 17524
rect 21361 17527 21419 17533
rect 19659 17493 19671 17496
rect 19613 17487 19671 17493
rect 21361 17493 21373 17527
rect 21407 17524 21419 17527
rect 21450 17524 21456 17536
rect 21407 17496 21456 17524
rect 21407 17493 21419 17496
rect 21361 17487 21419 17493
rect 21450 17484 21456 17496
rect 21508 17484 21514 17536
rect 1104 17434 21896 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21896 17434
rect 1104 17360 21896 17382
rect 1394 17320 1400 17332
rect 1355 17292 1400 17320
rect 1394 17280 1400 17292
rect 1452 17280 1458 17332
rect 1949 17323 2007 17329
rect 1949 17289 1961 17323
rect 1995 17320 2007 17323
rect 2038 17320 2044 17332
rect 1995 17292 2044 17320
rect 1995 17289 2007 17292
rect 1949 17283 2007 17289
rect 2038 17280 2044 17292
rect 2096 17280 2102 17332
rect 2222 17320 2228 17332
rect 2183 17292 2228 17320
rect 2222 17280 2228 17292
rect 2280 17280 2286 17332
rect 3050 17320 3056 17332
rect 3011 17292 3056 17320
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 3418 17320 3424 17332
rect 3379 17292 3424 17320
rect 3418 17280 3424 17292
rect 3476 17280 3482 17332
rect 3789 17323 3847 17329
rect 3789 17289 3801 17323
rect 3835 17320 3847 17323
rect 5258 17320 5264 17332
rect 3835 17292 5264 17320
rect 3835 17289 3847 17292
rect 3789 17283 3847 17289
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 5997 17323 6055 17329
rect 5997 17289 6009 17323
rect 6043 17320 6055 17323
rect 6546 17320 6552 17332
rect 6043 17292 6552 17320
rect 6043 17289 6055 17292
rect 5997 17283 6055 17289
rect 2685 17255 2743 17261
rect 2685 17221 2697 17255
rect 2731 17252 2743 17255
rect 3142 17252 3148 17264
rect 2731 17224 3148 17252
rect 2731 17221 2743 17224
rect 2685 17215 2743 17221
rect 3142 17212 3148 17224
rect 3200 17212 3206 17264
rect 5902 17252 5908 17264
rect 3896 17224 5908 17252
rect 1578 17076 1584 17128
rect 1636 17116 1642 17128
rect 3896 17116 3924 17224
rect 5902 17212 5908 17224
rect 5960 17252 5966 17264
rect 6012 17252 6040 17283
rect 6546 17280 6552 17292
rect 6604 17280 6610 17332
rect 7650 17280 7656 17332
rect 7708 17320 7714 17332
rect 9585 17323 9643 17329
rect 7708 17292 9076 17320
rect 7708 17280 7714 17292
rect 5960 17224 6040 17252
rect 5960 17212 5966 17224
rect 6086 17212 6092 17264
rect 6144 17252 6150 17264
rect 8110 17261 8116 17264
rect 6144 17224 8064 17252
rect 6144 17212 6150 17224
rect 4890 17184 4896 17196
rect 4851 17156 4896 17184
rect 4890 17144 4896 17156
rect 4948 17144 4954 17196
rect 5261 17187 5319 17193
rect 5261 17153 5273 17187
rect 5307 17184 5319 17187
rect 6457 17187 6515 17193
rect 5307 17156 6408 17184
rect 5307 17153 5319 17156
rect 5261 17147 5319 17153
rect 1636 17088 3924 17116
rect 4525 17119 4583 17125
rect 1636 17076 1642 17088
rect 4525 17085 4537 17119
rect 4571 17116 4583 17119
rect 5350 17116 5356 17128
rect 4571 17088 5356 17116
rect 4571 17085 4583 17088
rect 4525 17079 4583 17085
rect 5350 17076 5356 17088
rect 5408 17076 5414 17128
rect 6380 17116 6408 17156
rect 6457 17153 6469 17187
rect 6503 17184 6515 17187
rect 6730 17184 6736 17196
rect 6503 17156 6736 17184
rect 6503 17153 6515 17156
rect 6457 17147 6515 17153
rect 6730 17144 6736 17156
rect 6788 17144 6794 17196
rect 6914 17184 6920 17196
rect 6875 17156 6920 17184
rect 6914 17144 6920 17156
rect 6972 17144 6978 17196
rect 7837 17187 7895 17193
rect 7837 17153 7849 17187
rect 7883 17184 7895 17187
rect 7926 17184 7932 17196
rect 7883 17156 7932 17184
rect 7883 17153 7895 17156
rect 7837 17147 7895 17153
rect 7926 17144 7932 17156
rect 7984 17144 7990 17196
rect 8036 17184 8064 17224
rect 8104 17215 8116 17261
rect 8168 17252 8174 17264
rect 8168 17224 8204 17252
rect 8110 17212 8116 17215
rect 8168 17212 8174 17224
rect 9048 17184 9076 17292
rect 9585 17289 9597 17323
rect 9631 17320 9643 17323
rect 9674 17320 9680 17332
rect 9631 17292 9680 17320
rect 9631 17289 9643 17292
rect 9585 17283 9643 17289
rect 9674 17280 9680 17292
rect 9732 17280 9738 17332
rect 9766 17280 9772 17332
rect 9824 17320 9830 17332
rect 9824 17292 10088 17320
rect 9824 17280 9830 17292
rect 9122 17212 9128 17264
rect 9180 17252 9186 17264
rect 10060 17261 10088 17292
rect 10962 17280 10968 17332
rect 11020 17280 11026 17332
rect 11149 17323 11207 17329
rect 11149 17289 11161 17323
rect 11195 17320 11207 17323
rect 14550 17320 14556 17332
rect 11195 17292 12756 17320
rect 14511 17292 14556 17320
rect 11195 17289 11207 17292
rect 11149 17283 11207 17289
rect 9953 17255 10011 17261
rect 9953 17252 9965 17255
rect 9180 17224 9965 17252
rect 9180 17212 9186 17224
rect 9953 17221 9965 17224
rect 9999 17221 10011 17255
rect 9953 17215 10011 17221
rect 10045 17255 10103 17261
rect 10045 17221 10057 17255
rect 10091 17252 10103 17255
rect 10870 17252 10876 17264
rect 10091 17224 10876 17252
rect 10091 17221 10103 17224
rect 10045 17215 10103 17221
rect 10870 17212 10876 17224
rect 10928 17212 10934 17264
rect 10980 17252 11008 17280
rect 12434 17252 12440 17264
rect 10980 17224 12440 17252
rect 12434 17212 12440 17224
rect 12492 17212 12498 17264
rect 10965 17187 11023 17193
rect 10965 17184 10977 17187
rect 8036 17156 8892 17184
rect 9048 17156 10977 17184
rect 7098 17116 7104 17128
rect 6380 17088 7104 17116
rect 7098 17076 7104 17088
rect 7156 17076 7162 17128
rect 8864 17116 8892 17156
rect 10965 17153 10977 17156
rect 11011 17153 11023 17187
rect 10965 17147 11023 17153
rect 11514 17144 11520 17196
rect 11572 17184 11578 17196
rect 11609 17187 11667 17193
rect 11609 17184 11621 17187
rect 11572 17156 11621 17184
rect 11572 17144 11578 17156
rect 11609 17153 11621 17156
rect 11655 17153 11667 17187
rect 12728 17184 12756 17292
rect 14550 17280 14556 17292
rect 14608 17280 14614 17332
rect 17494 17320 17500 17332
rect 14660 17292 17500 17320
rect 14660 17252 14688 17292
rect 17494 17280 17500 17292
rect 17552 17280 17558 17332
rect 17678 17280 17684 17332
rect 17736 17320 17742 17332
rect 18138 17320 18144 17332
rect 17736 17292 18144 17320
rect 17736 17280 17742 17292
rect 18138 17280 18144 17292
rect 18196 17280 18202 17332
rect 18230 17280 18236 17332
rect 18288 17320 18294 17332
rect 18417 17323 18475 17329
rect 18417 17320 18429 17323
rect 18288 17292 18429 17320
rect 18288 17280 18294 17292
rect 18417 17289 18429 17292
rect 18463 17289 18475 17323
rect 18417 17283 18475 17289
rect 13004 17224 14688 17252
rect 13004 17184 13032 17224
rect 15102 17212 15108 17264
rect 15160 17252 15166 17264
rect 16209 17255 16267 17261
rect 16209 17252 16221 17255
rect 15160 17224 16221 17252
rect 15160 17212 15166 17224
rect 16209 17221 16221 17224
rect 16255 17252 16267 17255
rect 16298 17252 16304 17264
rect 16255 17224 16304 17252
rect 16255 17221 16267 17224
rect 16209 17215 16267 17221
rect 16298 17212 16304 17224
rect 16356 17212 16362 17264
rect 17954 17252 17960 17264
rect 17052 17224 17960 17252
rect 13170 17193 13176 17196
rect 13164 17184 13176 17193
rect 12728 17156 13032 17184
rect 13131 17156 13176 17184
rect 11609 17147 11667 17153
rect 13164 17147 13176 17156
rect 13170 17144 13176 17147
rect 13228 17144 13234 17196
rect 14274 17184 14280 17196
rect 14187 17156 14280 17184
rect 14274 17144 14280 17156
rect 14332 17184 14338 17196
rect 15677 17187 15735 17193
rect 15677 17184 15689 17187
rect 14332 17156 15689 17184
rect 14332 17144 14338 17156
rect 15677 17153 15689 17156
rect 15723 17184 15735 17187
rect 16758 17184 16764 17196
rect 15723 17156 16764 17184
rect 15723 17153 15735 17156
rect 15677 17147 15735 17153
rect 16758 17144 16764 17156
rect 16816 17144 16822 17196
rect 9306 17116 9312 17128
rect 8864 17088 9312 17116
rect 9306 17076 9312 17088
rect 9364 17076 9370 17128
rect 10226 17116 10232 17128
rect 10187 17088 10232 17116
rect 10226 17076 10232 17088
rect 10284 17076 10290 17128
rect 11698 17116 11704 17128
rect 10612 17088 11704 17116
rect 1670 17008 1676 17060
rect 1728 17048 1734 17060
rect 9217 17051 9275 17057
rect 1728 17020 7880 17048
rect 1728 17008 1734 17020
rect 4157 16983 4215 16989
rect 4157 16949 4169 16983
rect 4203 16980 4215 16983
rect 4246 16980 4252 16992
rect 4203 16952 4252 16980
rect 4203 16949 4215 16952
rect 4157 16943 4215 16949
rect 4246 16940 4252 16952
rect 4304 16940 4310 16992
rect 5629 16983 5687 16989
rect 5629 16949 5641 16983
rect 5675 16980 5687 16983
rect 6086 16980 6092 16992
rect 5675 16952 6092 16980
rect 5675 16949 5687 16952
rect 5629 16943 5687 16949
rect 6086 16940 6092 16952
rect 6144 16940 6150 16992
rect 6641 16983 6699 16989
rect 6641 16949 6653 16983
rect 6687 16980 6699 16983
rect 6822 16980 6828 16992
rect 6687 16952 6828 16980
rect 6687 16949 6699 16952
rect 6641 16943 6699 16949
rect 6822 16940 6828 16952
rect 6880 16940 6886 16992
rect 7558 16980 7564 16992
rect 7519 16952 7564 16980
rect 7558 16940 7564 16952
rect 7616 16940 7622 16992
rect 7852 16980 7880 17020
rect 9217 17017 9229 17051
rect 9263 17048 9275 17051
rect 10244 17048 10272 17076
rect 9263 17020 10272 17048
rect 9263 17017 9275 17020
rect 9217 17011 9275 17017
rect 9490 16980 9496 16992
rect 7852 16952 9496 16980
rect 9490 16940 9496 16952
rect 9548 16940 9554 16992
rect 9674 16940 9680 16992
rect 9732 16980 9738 16992
rect 10612 16980 10640 17088
rect 11698 17076 11704 17088
rect 11756 17076 11762 17128
rect 12250 17076 12256 17128
rect 12308 17116 12314 17128
rect 12897 17119 12955 17125
rect 12897 17116 12909 17119
rect 12308 17088 12909 17116
rect 12308 17076 12314 17088
rect 12897 17085 12909 17088
rect 12943 17085 12955 17119
rect 12897 17079 12955 17085
rect 10870 17008 10876 17060
rect 10928 17048 10934 17060
rect 12802 17048 12808 17060
rect 10928 17020 12808 17048
rect 10928 17008 10934 17020
rect 12802 17008 12808 17020
rect 12860 17008 12866 17060
rect 14292 17057 14320 17144
rect 15933 17119 15991 17125
rect 15933 17085 15945 17119
rect 15979 17116 15991 17119
rect 16114 17116 16120 17128
rect 15979 17088 16120 17116
rect 15979 17085 15991 17088
rect 15933 17079 15991 17085
rect 16114 17076 16120 17088
rect 16172 17116 16178 17128
rect 16298 17116 16304 17128
rect 16172 17088 16304 17116
rect 16172 17076 16178 17088
rect 16298 17076 16304 17088
rect 16356 17116 16362 17128
rect 17052 17125 17080 17224
rect 17954 17212 17960 17224
rect 18012 17252 18018 17264
rect 18966 17261 18972 17264
rect 18960 17252 18972 17261
rect 18012 17224 18736 17252
rect 18927 17224 18972 17252
rect 18012 17212 18018 17224
rect 17310 17193 17316 17196
rect 17304 17184 17316 17193
rect 17271 17156 17316 17184
rect 17304 17147 17316 17156
rect 17310 17144 17316 17147
rect 17368 17144 17374 17196
rect 18708 17193 18736 17224
rect 18960 17215 18972 17224
rect 18966 17212 18972 17215
rect 19024 17212 19030 17264
rect 18693 17187 18751 17193
rect 18693 17153 18705 17187
rect 18739 17153 18751 17187
rect 20622 17184 20628 17196
rect 18693 17147 18751 17153
rect 18800 17156 20628 17184
rect 17037 17119 17095 17125
rect 17037 17116 17049 17119
rect 16356 17088 17049 17116
rect 16356 17076 16362 17088
rect 17037 17085 17049 17088
rect 17083 17085 17095 17119
rect 17037 17079 17095 17085
rect 18138 17076 18144 17128
rect 18196 17116 18202 17128
rect 18800 17116 18828 17156
rect 20622 17144 20628 17156
rect 20680 17144 20686 17196
rect 20990 17184 20996 17196
rect 20951 17156 20996 17184
rect 20990 17144 20996 17156
rect 21048 17144 21054 17196
rect 18196 17088 18828 17116
rect 18196 17076 18202 17088
rect 14277 17051 14335 17057
rect 14277 17017 14289 17051
rect 14323 17017 14335 17051
rect 21269 17051 21327 17057
rect 21269 17048 21281 17051
rect 14277 17011 14335 17017
rect 15948 17020 16804 17048
rect 9732 16952 10640 16980
rect 10689 16983 10747 16989
rect 9732 16940 9738 16952
rect 10689 16949 10701 16983
rect 10735 16980 10747 16983
rect 10778 16980 10784 16992
rect 10735 16952 10784 16980
rect 10735 16949 10747 16952
rect 10689 16943 10747 16949
rect 10778 16940 10784 16952
rect 10836 16980 10842 16992
rect 11882 16980 11888 16992
rect 10836 16952 11888 16980
rect 10836 16940 10842 16952
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 12158 16940 12164 16992
rect 12216 16980 12222 16992
rect 12253 16983 12311 16989
rect 12253 16980 12265 16983
rect 12216 16952 12265 16980
rect 12216 16940 12222 16952
rect 12253 16949 12265 16952
rect 12299 16949 12311 16983
rect 12253 16943 12311 16949
rect 12621 16983 12679 16989
rect 12621 16949 12633 16983
rect 12667 16980 12679 16983
rect 13814 16980 13820 16992
rect 12667 16952 13820 16980
rect 12667 16949 12679 16952
rect 12621 16943 12679 16949
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 15654 16940 15660 16992
rect 15712 16980 15718 16992
rect 15948 16980 15976 17020
rect 16666 16980 16672 16992
rect 15712 16952 15976 16980
rect 16627 16952 16672 16980
rect 15712 16940 15718 16952
rect 16666 16940 16672 16952
rect 16724 16940 16730 16992
rect 16776 16980 16804 17020
rect 19628 17020 21281 17048
rect 19628 16980 19656 17020
rect 21269 17017 21281 17020
rect 21315 17017 21327 17051
rect 21269 17011 21327 17017
rect 16776 16952 19656 16980
rect 19978 16940 19984 16992
rect 20036 16980 20042 16992
rect 20073 16983 20131 16989
rect 20073 16980 20085 16983
rect 20036 16952 20085 16980
rect 20036 16940 20042 16952
rect 20073 16949 20085 16952
rect 20119 16949 20131 16983
rect 20073 16943 20131 16949
rect 20349 16983 20407 16989
rect 20349 16949 20361 16983
rect 20395 16980 20407 16983
rect 20438 16980 20444 16992
rect 20395 16952 20444 16980
rect 20395 16949 20407 16952
rect 20349 16943 20407 16949
rect 20438 16940 20444 16952
rect 20496 16940 20502 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 1854 16776 1860 16788
rect 1815 16748 1860 16776
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 2498 16776 2504 16788
rect 2459 16748 2504 16776
rect 2498 16736 2504 16748
rect 2556 16736 2562 16788
rect 4341 16779 4399 16785
rect 4341 16745 4353 16779
rect 4387 16776 4399 16779
rect 4614 16776 4620 16788
rect 4387 16748 4620 16776
rect 4387 16745 4399 16748
rect 4341 16739 4399 16745
rect 4614 16736 4620 16748
rect 4672 16736 4678 16788
rect 4982 16776 4988 16788
rect 4943 16748 4988 16776
rect 4982 16736 4988 16748
rect 5040 16736 5046 16788
rect 5350 16776 5356 16788
rect 5311 16748 5356 16776
rect 5350 16736 5356 16748
rect 5408 16736 5414 16788
rect 5534 16736 5540 16788
rect 5592 16776 5598 16788
rect 5629 16779 5687 16785
rect 5629 16776 5641 16779
rect 5592 16748 5641 16776
rect 5592 16736 5598 16748
rect 5629 16745 5641 16748
rect 5675 16745 5687 16779
rect 6914 16776 6920 16788
rect 6875 16748 6920 16776
rect 5629 16739 5687 16745
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 7926 16736 7932 16788
rect 7984 16776 7990 16788
rect 7984 16748 8340 16776
rect 7984 16736 7990 16748
rect 5000 16708 5028 16736
rect 5994 16708 6000 16720
rect 5000 16680 6000 16708
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 8312 16708 8340 16748
rect 8386 16736 8392 16788
rect 8444 16776 8450 16788
rect 9674 16776 9680 16788
rect 8444 16748 9680 16776
rect 8444 16736 8450 16748
rect 9674 16736 9680 16748
rect 9732 16736 9738 16788
rect 9950 16736 9956 16788
rect 10008 16776 10014 16788
rect 11146 16776 11152 16788
rect 10008 16748 11152 16776
rect 10008 16736 10014 16748
rect 9968 16708 9996 16736
rect 8312 16680 9996 16708
rect 5350 16600 5356 16652
rect 5408 16640 5414 16652
rect 5626 16640 5632 16652
rect 5408 16612 5632 16640
rect 5408 16600 5414 16612
rect 5626 16600 5632 16612
rect 5684 16600 5690 16652
rect 8312 16649 8340 16680
rect 8297 16643 8355 16649
rect 8297 16609 8309 16643
rect 8343 16609 8355 16643
rect 9306 16640 9312 16652
rect 9267 16612 9312 16640
rect 8297 16603 8355 16609
rect 9306 16600 9312 16612
rect 9364 16600 9370 16652
rect 9490 16640 9496 16652
rect 9451 16612 9496 16640
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 9582 16600 9588 16652
rect 9640 16640 9646 16652
rect 10244 16649 10272 16748
rect 11146 16736 11152 16748
rect 11204 16776 11210 16788
rect 12250 16776 12256 16788
rect 11204 16748 12256 16776
rect 11204 16736 11210 16748
rect 11900 16649 11928 16748
rect 12250 16736 12256 16748
rect 12308 16736 12314 16788
rect 12802 16736 12808 16788
rect 12860 16776 12866 16788
rect 15194 16776 15200 16788
rect 12860 16748 15200 16776
rect 12860 16736 12866 16748
rect 15194 16736 15200 16748
rect 15252 16736 15258 16788
rect 15930 16776 15936 16788
rect 15891 16748 15936 16776
rect 15930 16736 15936 16748
rect 15988 16736 15994 16788
rect 18046 16736 18052 16788
rect 18104 16776 18110 16788
rect 19245 16779 19303 16785
rect 19245 16776 19257 16779
rect 18104 16748 19257 16776
rect 18104 16736 18110 16748
rect 19245 16745 19257 16748
rect 19291 16745 19303 16779
rect 19245 16739 19303 16745
rect 20622 16736 20628 16788
rect 20680 16776 20686 16788
rect 21269 16779 21327 16785
rect 21269 16776 21281 16779
rect 20680 16748 21281 16776
rect 20680 16736 20686 16748
rect 21269 16745 21281 16748
rect 21315 16745 21327 16779
rect 21269 16739 21327 16745
rect 13170 16668 13176 16720
rect 13228 16708 13234 16720
rect 13265 16711 13323 16717
rect 13265 16708 13277 16711
rect 13228 16680 13277 16708
rect 13228 16668 13234 16680
rect 13265 16677 13277 16680
rect 13311 16708 13323 16711
rect 14550 16708 14556 16720
rect 13311 16680 14228 16708
rect 13311 16677 13323 16680
rect 13265 16671 13323 16677
rect 10229 16643 10287 16649
rect 9640 16612 10088 16640
rect 9640 16600 9646 16612
rect 6181 16575 6239 16581
rect 6181 16541 6193 16575
rect 6227 16572 6239 16575
rect 9950 16572 9956 16584
rect 6227 16544 9956 16572
rect 6227 16541 6239 16544
rect 6181 16535 6239 16541
rect 9950 16532 9956 16544
rect 10008 16532 10014 16584
rect 10060 16572 10088 16612
rect 10229 16609 10241 16643
rect 10275 16609 10287 16643
rect 10229 16603 10287 16609
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16609 11943 16643
rect 11885 16603 11943 16609
rect 12158 16581 12164 16584
rect 12152 16572 12164 16581
rect 10060 16544 12020 16572
rect 12119 16544 12164 16572
rect 8052 16507 8110 16513
rect 8052 16473 8064 16507
rect 8098 16504 8110 16507
rect 10226 16504 10232 16516
rect 8098 16476 10232 16504
rect 8098 16473 8110 16476
rect 8052 16467 8110 16473
rect 10226 16464 10232 16476
rect 10284 16464 10290 16516
rect 10496 16507 10554 16513
rect 10496 16473 10508 16507
rect 10542 16504 10554 16507
rect 10686 16504 10692 16516
rect 10542 16476 10692 16504
rect 10542 16473 10554 16476
rect 10496 16467 10554 16473
rect 10686 16464 10692 16476
rect 10744 16464 10750 16516
rect 11514 16464 11520 16516
rect 11572 16464 11578 16516
rect 11992 16504 12020 16544
rect 12152 16535 12164 16544
rect 12158 16532 12164 16535
rect 12216 16532 12222 16584
rect 13541 16575 13599 16581
rect 13541 16572 13553 16575
rect 12406 16544 13553 16572
rect 12406 16504 12434 16544
rect 13541 16541 13553 16544
rect 13587 16541 13599 16575
rect 14200 16572 14228 16680
rect 14292 16680 14556 16708
rect 14292 16649 14320 16680
rect 14550 16668 14556 16680
rect 14608 16668 14614 16720
rect 15838 16668 15844 16720
rect 15896 16708 15902 16720
rect 20162 16708 20168 16720
rect 15896 16680 20168 16708
rect 15896 16668 15902 16680
rect 20162 16668 20168 16680
rect 20220 16668 20226 16720
rect 14277 16643 14335 16649
rect 14277 16609 14289 16643
rect 14323 16609 14335 16643
rect 14277 16603 14335 16609
rect 14369 16643 14427 16649
rect 14369 16609 14381 16643
rect 14415 16640 14427 16643
rect 14826 16640 14832 16652
rect 14415 16612 14832 16640
rect 14415 16609 14427 16612
rect 14369 16603 14427 16609
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 15381 16643 15439 16649
rect 15381 16640 15393 16643
rect 14936 16612 15393 16640
rect 14734 16572 14740 16584
rect 14200 16544 14740 16572
rect 13541 16535 13599 16541
rect 14734 16532 14740 16544
rect 14792 16572 14798 16584
rect 14936 16572 14964 16612
rect 15381 16609 15393 16612
rect 15427 16640 15439 16643
rect 16758 16640 16764 16652
rect 15427 16612 16620 16640
rect 16719 16612 16764 16640
rect 15427 16609 15439 16612
rect 15381 16603 15439 16609
rect 15562 16572 15568 16584
rect 14792 16544 14964 16572
rect 15523 16544 15568 16572
rect 14792 16532 14798 16544
rect 15562 16532 15568 16544
rect 15620 16532 15626 16584
rect 16592 16572 16620 16612
rect 16758 16600 16764 16612
rect 16816 16600 16822 16652
rect 17773 16643 17831 16649
rect 17773 16640 17785 16643
rect 16868 16612 17785 16640
rect 16868 16572 16896 16612
rect 17773 16609 17785 16612
rect 17819 16609 17831 16643
rect 17773 16603 17831 16609
rect 19242 16600 19248 16652
rect 19300 16640 19306 16652
rect 19300 16612 19748 16640
rect 19300 16600 19306 16612
rect 16592 16544 16896 16572
rect 17678 16532 17684 16584
rect 17736 16572 17742 16584
rect 18874 16572 18880 16584
rect 17736 16544 17781 16572
rect 18835 16544 18880 16572
rect 17736 16532 17742 16544
rect 18874 16532 18880 16544
rect 18932 16532 18938 16584
rect 19610 16572 19616 16584
rect 18984 16544 19616 16572
rect 11992 16476 12434 16504
rect 14461 16507 14519 16513
rect 14461 16473 14473 16507
rect 14507 16504 14519 16507
rect 14507 16476 15700 16504
rect 14507 16473 14519 16476
rect 14461 16467 14519 16473
rect 2682 16396 2688 16448
rect 2740 16436 2746 16448
rect 5997 16439 6055 16445
rect 5997 16436 6009 16439
rect 2740 16408 6009 16436
rect 2740 16396 2746 16408
rect 5997 16405 6009 16408
rect 6043 16436 6055 16439
rect 6546 16436 6552 16448
rect 6043 16408 6552 16436
rect 6043 16405 6055 16408
rect 5997 16399 6055 16405
rect 6546 16396 6552 16408
rect 6604 16396 6610 16448
rect 6641 16439 6699 16445
rect 6641 16405 6653 16439
rect 6687 16436 6699 16439
rect 9306 16436 9312 16448
rect 6687 16408 9312 16436
rect 6687 16405 6699 16408
rect 6641 16399 6699 16405
rect 9306 16396 9312 16408
rect 9364 16396 9370 16448
rect 9582 16436 9588 16448
rect 9543 16408 9588 16436
rect 9582 16396 9588 16408
rect 9640 16396 9646 16448
rect 9674 16396 9680 16448
rect 9732 16436 9738 16448
rect 9953 16439 10011 16445
rect 9953 16436 9965 16439
rect 9732 16408 9965 16436
rect 9732 16396 9738 16408
rect 9953 16405 9965 16408
rect 9999 16405 10011 16439
rect 11532 16436 11560 16464
rect 11609 16439 11667 16445
rect 11609 16436 11621 16439
rect 11532 16408 11621 16436
rect 9953 16399 10011 16405
rect 11609 16405 11621 16408
rect 11655 16436 11667 16439
rect 13538 16436 13544 16448
rect 11655 16408 13544 16436
rect 11655 16405 11667 16408
rect 11609 16399 11667 16405
rect 13538 16396 13544 16408
rect 13596 16396 13602 16448
rect 13725 16439 13783 16445
rect 13725 16405 13737 16439
rect 13771 16436 13783 16439
rect 13906 16436 13912 16448
rect 13771 16408 13912 16436
rect 13771 16405 13783 16408
rect 13725 16399 13783 16405
rect 13906 16396 13912 16408
rect 13964 16396 13970 16448
rect 14366 16396 14372 16448
rect 14424 16436 14430 16448
rect 14550 16436 14556 16448
rect 14424 16408 14556 16436
rect 14424 16396 14430 16408
rect 14550 16396 14556 16408
rect 14608 16396 14614 16448
rect 14829 16439 14887 16445
rect 14829 16405 14841 16439
rect 14875 16436 14887 16439
rect 15010 16436 15016 16448
rect 14875 16408 15016 16436
rect 14875 16405 14887 16408
rect 14829 16399 14887 16405
rect 15010 16396 15016 16408
rect 15068 16396 15074 16448
rect 15473 16439 15531 16445
rect 15473 16405 15485 16439
rect 15519 16436 15531 16439
rect 15562 16436 15568 16448
rect 15519 16408 15568 16436
rect 15519 16405 15531 16408
rect 15473 16399 15531 16405
rect 15562 16396 15568 16408
rect 15620 16396 15626 16448
rect 15672 16436 15700 16476
rect 15930 16464 15936 16516
rect 15988 16504 15994 16516
rect 16577 16507 16635 16513
rect 16577 16504 16589 16507
rect 15988 16476 16589 16504
rect 15988 16464 15994 16476
rect 16577 16473 16589 16476
rect 16623 16473 16635 16507
rect 16577 16467 16635 16473
rect 16942 16464 16948 16516
rect 17000 16504 17006 16516
rect 18984 16504 19012 16544
rect 19610 16532 19616 16544
rect 19668 16532 19674 16584
rect 19720 16572 19748 16612
rect 19794 16600 19800 16652
rect 19852 16640 19858 16652
rect 20809 16643 20867 16649
rect 20809 16640 20821 16643
rect 19852 16612 19897 16640
rect 19996 16612 20821 16640
rect 19852 16600 19858 16612
rect 19996 16572 20024 16612
rect 20809 16609 20821 16612
rect 20855 16640 20867 16643
rect 20990 16640 20996 16652
rect 20855 16612 20996 16640
rect 20855 16609 20867 16612
rect 20809 16603 20867 16609
rect 20990 16600 20996 16612
rect 21048 16600 21054 16652
rect 19720 16544 20024 16572
rect 17000 16476 19012 16504
rect 17000 16464 17006 16476
rect 19518 16464 19524 16516
rect 19576 16504 19582 16516
rect 19705 16507 19763 16513
rect 19705 16504 19717 16507
rect 19576 16476 19717 16504
rect 19576 16464 19582 16476
rect 19705 16473 19717 16476
rect 19751 16473 19763 16507
rect 19705 16467 19763 16473
rect 20070 16464 20076 16516
rect 20128 16504 20134 16516
rect 20717 16507 20775 16513
rect 20717 16504 20729 16507
rect 20128 16476 20729 16504
rect 20128 16464 20134 16476
rect 20717 16473 20729 16476
rect 20763 16473 20775 16507
rect 20717 16467 20775 16473
rect 16209 16439 16267 16445
rect 16209 16436 16221 16439
rect 15672 16408 16221 16436
rect 16209 16405 16221 16408
rect 16255 16405 16267 16439
rect 16209 16399 16267 16405
rect 16669 16439 16727 16445
rect 16669 16405 16681 16439
rect 16715 16436 16727 16439
rect 17221 16439 17279 16445
rect 17221 16436 17233 16439
rect 16715 16408 17233 16436
rect 16715 16405 16727 16408
rect 16669 16399 16727 16405
rect 17221 16405 17233 16408
rect 17267 16405 17279 16439
rect 17586 16436 17592 16448
rect 17547 16408 17592 16436
rect 17221 16399 17279 16405
rect 17586 16396 17592 16408
rect 17644 16396 17650 16448
rect 17770 16396 17776 16448
rect 17828 16436 17834 16448
rect 18233 16439 18291 16445
rect 18233 16436 18245 16439
rect 17828 16408 18245 16436
rect 17828 16396 17834 16408
rect 18233 16405 18245 16408
rect 18279 16405 18291 16439
rect 18233 16399 18291 16405
rect 19613 16439 19671 16445
rect 19613 16405 19625 16439
rect 19659 16436 19671 16439
rect 19794 16436 19800 16448
rect 19659 16408 19800 16436
rect 19659 16405 19671 16408
rect 19613 16399 19671 16405
rect 19794 16396 19800 16408
rect 19852 16396 19858 16448
rect 20254 16436 20260 16448
rect 20215 16408 20260 16436
rect 20254 16396 20260 16408
rect 20312 16396 20318 16448
rect 20346 16396 20352 16448
rect 20404 16436 20410 16448
rect 20625 16439 20683 16445
rect 20625 16436 20637 16439
rect 20404 16408 20637 16436
rect 20404 16396 20410 16408
rect 20625 16405 20637 16408
rect 20671 16405 20683 16439
rect 20625 16399 20683 16405
rect 1104 16346 21896 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21896 16346
rect 1104 16272 21896 16294
rect 4522 16192 4528 16244
rect 4580 16232 4586 16244
rect 6733 16235 6791 16241
rect 6733 16232 6745 16235
rect 4580 16204 6745 16232
rect 4580 16192 4586 16204
rect 6733 16201 6745 16204
rect 6779 16201 6791 16235
rect 9674 16232 9680 16244
rect 6733 16195 6791 16201
rect 7392 16204 9536 16232
rect 9635 16204 9680 16232
rect 5810 16124 5816 16176
rect 5868 16164 5874 16176
rect 7392 16164 7420 16204
rect 7926 16164 7932 16176
rect 5868 16136 7420 16164
rect 7484 16136 7932 16164
rect 5868 16124 5874 16136
rect 5442 16096 5448 16108
rect 5184 16068 5448 16096
rect 4614 15920 4620 15972
rect 4672 15960 4678 15972
rect 5184 15969 5212 16068
rect 5442 16056 5448 16068
rect 5500 16096 5506 16108
rect 7484 16105 7512 16136
rect 7926 16124 7932 16136
rect 7984 16124 7990 16176
rect 9508 16164 9536 16204
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 9769 16235 9827 16241
rect 9769 16201 9781 16235
rect 9815 16232 9827 16235
rect 10413 16235 10471 16241
rect 10413 16232 10425 16235
rect 9815 16204 10425 16232
rect 9815 16201 9827 16204
rect 9769 16195 9827 16201
rect 10413 16201 10425 16204
rect 10459 16201 10471 16235
rect 11698 16232 11704 16244
rect 10413 16195 10471 16201
rect 10520 16204 11560 16232
rect 11659 16204 11704 16232
rect 10520 16164 10548 16204
rect 10686 16164 10692 16176
rect 9508 16136 10548 16164
rect 10612 16136 10692 16164
rect 6825 16099 6883 16105
rect 6825 16096 6837 16099
rect 5500 16068 6837 16096
rect 5500 16056 5506 16068
rect 6825 16065 6837 16068
rect 6871 16065 6883 16099
rect 6825 16059 6883 16065
rect 7469 16099 7527 16105
rect 7469 16065 7481 16099
rect 7515 16065 7527 16099
rect 7469 16059 7527 16065
rect 7558 16056 7564 16108
rect 7616 16096 7622 16108
rect 7725 16099 7783 16105
rect 7725 16096 7737 16099
rect 7616 16068 7737 16096
rect 7616 16056 7622 16068
rect 7725 16065 7737 16068
rect 7771 16065 7783 16099
rect 7725 16059 7783 16065
rect 5258 15988 5264 16040
rect 5316 16028 5322 16040
rect 5626 16028 5632 16040
rect 5316 16000 5632 16028
rect 5316 15988 5322 16000
rect 5626 15988 5632 16000
rect 5684 15988 5690 16040
rect 6641 16031 6699 16037
rect 6641 15997 6653 16031
rect 6687 15997 6699 16031
rect 6641 15991 6699 15997
rect 9585 16031 9643 16037
rect 9585 15997 9597 16031
rect 9631 16028 9643 16031
rect 9766 16028 9772 16040
rect 9631 16000 9772 16028
rect 9631 15997 9643 16000
rect 9585 15991 9643 15997
rect 5169 15963 5227 15969
rect 5169 15960 5181 15963
rect 4672 15932 5181 15960
rect 4672 15920 4678 15932
rect 5169 15929 5181 15932
rect 5215 15929 5227 15963
rect 6656 15960 6684 15991
rect 9766 15988 9772 16000
rect 9824 16028 9830 16040
rect 10612 16028 10640 16136
rect 10686 16124 10692 16136
rect 10744 16164 10750 16176
rect 10744 16136 11192 16164
rect 10744 16124 10750 16136
rect 10778 16096 10784 16108
rect 10739 16068 10784 16096
rect 10778 16056 10784 16068
rect 10836 16056 10842 16108
rect 10870 16028 10876 16040
rect 9824 16000 10640 16028
rect 10831 16000 10876 16028
rect 9824 15988 9830 16000
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 10962 15988 10968 16040
rect 11020 16028 11026 16040
rect 11164 16028 11192 16136
rect 11532 16105 11560 16204
rect 11698 16192 11704 16204
rect 11756 16192 11762 16244
rect 12713 16235 12771 16241
rect 12713 16201 12725 16235
rect 12759 16232 12771 16235
rect 13357 16235 13415 16241
rect 13357 16232 13369 16235
rect 12759 16204 13369 16232
rect 12759 16201 12771 16204
rect 12713 16195 12771 16201
rect 13357 16201 13369 16204
rect 13403 16201 13415 16235
rect 13357 16195 13415 16201
rect 13722 16192 13728 16244
rect 13780 16232 13786 16244
rect 19061 16235 19119 16241
rect 13780 16204 17816 16232
rect 13780 16192 13786 16204
rect 12253 16167 12311 16173
rect 12253 16133 12265 16167
rect 12299 16164 12311 16167
rect 17678 16164 17684 16176
rect 12299 16136 17684 16164
rect 12299 16133 12311 16136
rect 12253 16127 12311 16133
rect 17678 16124 17684 16136
rect 17736 16124 17742 16176
rect 17788 16164 17816 16204
rect 19061 16201 19073 16235
rect 19107 16232 19119 16235
rect 19242 16232 19248 16244
rect 19107 16204 19248 16232
rect 19107 16201 19119 16204
rect 19061 16195 19119 16201
rect 19242 16192 19248 16204
rect 19300 16192 19306 16244
rect 19613 16235 19671 16241
rect 19613 16232 19625 16235
rect 19352 16204 19625 16232
rect 19352 16164 19380 16204
rect 19613 16201 19625 16204
rect 19659 16201 19671 16235
rect 20070 16232 20076 16244
rect 20031 16204 20076 16232
rect 19613 16195 19671 16201
rect 20070 16192 20076 16204
rect 20128 16192 20134 16244
rect 20346 16232 20352 16244
rect 20307 16204 20352 16232
rect 20346 16192 20352 16204
rect 20404 16192 20410 16244
rect 19978 16164 19984 16176
rect 17788 16136 19380 16164
rect 19444 16136 19984 16164
rect 11517 16099 11575 16105
rect 11517 16065 11529 16099
rect 11563 16065 11575 16099
rect 11517 16059 11575 16065
rect 12345 16099 12403 16105
rect 12345 16065 12357 16099
rect 12391 16096 12403 16099
rect 12434 16096 12440 16108
rect 12391 16068 12440 16096
rect 12391 16065 12403 16068
rect 12345 16059 12403 16065
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 13449 16099 13507 16105
rect 13449 16065 13461 16099
rect 13495 16096 13507 16099
rect 13495 16068 13676 16096
rect 13495 16065 13507 16068
rect 13449 16059 13507 16065
rect 12069 16031 12127 16037
rect 12069 16028 12081 16031
rect 11020 16000 11065 16028
rect 11164 16000 12081 16028
rect 11020 15988 11026 16000
rect 12069 15997 12081 16000
rect 12115 15997 12127 16031
rect 13538 16028 13544 16040
rect 13499 16000 13544 16028
rect 12069 15991 12127 15997
rect 13538 15988 13544 16000
rect 13596 15988 13602 16040
rect 6914 15960 6920 15972
rect 6656 15932 6920 15960
rect 5169 15923 5227 15929
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 7282 15960 7288 15972
rect 7116 15932 7288 15960
rect 4893 15895 4951 15901
rect 4893 15861 4905 15895
rect 4939 15892 4951 15895
rect 4982 15892 4988 15904
rect 4939 15864 4988 15892
rect 4939 15861 4951 15864
rect 4893 15855 4951 15861
rect 4982 15852 4988 15864
rect 5040 15852 5046 15904
rect 5997 15895 6055 15901
rect 5997 15861 6009 15895
rect 6043 15892 6055 15895
rect 7116 15892 7144 15932
rect 7282 15920 7288 15932
rect 7340 15920 7346 15972
rect 10137 15963 10195 15969
rect 10137 15929 10149 15963
rect 10183 15960 10195 15963
rect 13648 15960 13676 16068
rect 14366 16056 14372 16108
rect 14424 16096 14430 16108
rect 14645 16099 14703 16105
rect 14645 16096 14657 16099
rect 14424 16068 14657 16096
rect 14424 16056 14430 16068
rect 14645 16065 14657 16068
rect 14691 16065 14703 16099
rect 14645 16059 14703 16065
rect 16045 16099 16103 16105
rect 16045 16065 16057 16099
rect 16091 16096 16103 16099
rect 16206 16096 16212 16108
rect 16091 16068 16212 16096
rect 16091 16065 16103 16068
rect 16045 16059 16103 16065
rect 16206 16056 16212 16068
rect 16264 16056 16270 16108
rect 17402 16096 17408 16108
rect 17363 16068 17408 16096
rect 17402 16056 17408 16068
rect 17460 16056 17466 16108
rect 17948 16099 18006 16105
rect 17948 16065 17960 16099
rect 17994 16096 18006 16099
rect 19444 16096 19472 16136
rect 19978 16124 19984 16136
rect 20036 16164 20042 16176
rect 20036 16136 20944 16164
rect 20036 16124 20042 16136
rect 19705 16099 19763 16105
rect 19705 16096 19717 16099
rect 17994 16068 19472 16096
rect 17994 16065 18006 16068
rect 17948 16059 18006 16065
rect 16298 16028 16304 16040
rect 16259 16000 16304 16028
rect 16298 15988 16304 16000
rect 16356 16028 16362 16040
rect 19444 16037 19472 16068
rect 19536 16068 19717 16096
rect 17681 16031 17739 16037
rect 17681 16028 17693 16031
rect 16356 16000 17693 16028
rect 16356 15988 16362 16000
rect 17681 15997 17693 16000
rect 17727 15997 17739 16031
rect 17681 15991 17739 15997
rect 19429 16031 19487 16037
rect 19429 15997 19441 16031
rect 19475 15997 19487 16031
rect 19429 15991 19487 15997
rect 10183 15932 13676 15960
rect 10183 15929 10195 15932
rect 10137 15923 10195 15929
rect 13906 15920 13912 15972
rect 13964 15960 13970 15972
rect 16942 15960 16948 15972
rect 13964 15932 15056 15960
rect 13964 15920 13970 15932
rect 6043 15864 7144 15892
rect 7193 15895 7251 15901
rect 6043 15861 6055 15864
rect 5997 15855 6055 15861
rect 7193 15861 7205 15895
rect 7239 15892 7251 15895
rect 8110 15892 8116 15904
rect 7239 15864 8116 15892
rect 7239 15861 7251 15864
rect 7193 15855 7251 15861
rect 8110 15852 8116 15864
rect 8168 15852 8174 15904
rect 8849 15895 8907 15901
rect 8849 15861 8861 15895
rect 8895 15892 8907 15895
rect 9122 15892 9128 15904
rect 8895 15864 9128 15892
rect 8895 15861 8907 15864
rect 8849 15855 8907 15861
rect 9122 15852 9128 15864
rect 9180 15852 9186 15904
rect 9398 15852 9404 15904
rect 9456 15892 9462 15904
rect 10962 15892 10968 15904
rect 9456 15864 10968 15892
rect 9456 15852 9462 15864
rect 10962 15852 10968 15864
rect 11020 15852 11026 15904
rect 12526 15852 12532 15904
rect 12584 15892 12590 15904
rect 12989 15895 13047 15901
rect 12989 15892 13001 15895
rect 12584 15864 13001 15892
rect 12584 15852 12590 15864
rect 12989 15861 13001 15864
rect 13035 15861 13047 15895
rect 12989 15855 13047 15861
rect 14001 15895 14059 15901
rect 14001 15861 14013 15895
rect 14047 15892 14059 15895
rect 14274 15892 14280 15904
rect 14047 15864 14280 15892
rect 14047 15861 14059 15864
rect 14001 15855 14059 15861
rect 14274 15852 14280 15864
rect 14332 15852 14338 15904
rect 14918 15892 14924 15904
rect 14879 15864 14924 15892
rect 14918 15852 14924 15864
rect 14976 15852 14982 15904
rect 15028 15892 15056 15932
rect 16316 15932 16948 15960
rect 16316 15892 16344 15932
rect 16942 15920 16948 15932
rect 17000 15920 17006 15972
rect 18966 15920 18972 15972
rect 19024 15960 19030 15972
rect 19536 15960 19564 16068
rect 19705 16065 19717 16068
rect 19751 16065 19763 16099
rect 20714 16096 20720 16108
rect 20675 16068 20720 16096
rect 19705 16059 19763 16065
rect 20714 16056 20720 16068
rect 20772 16056 20778 16108
rect 20916 16037 20944 16136
rect 20809 16031 20867 16037
rect 20809 15997 20821 16031
rect 20855 15997 20867 16031
rect 20809 15991 20867 15997
rect 20901 16031 20959 16037
rect 20901 15997 20913 16031
rect 20947 15997 20959 16031
rect 20901 15991 20959 15997
rect 19024 15932 19564 15960
rect 19024 15920 19030 15932
rect 15028 15864 16344 15892
rect 16761 15895 16819 15901
rect 16761 15861 16773 15895
rect 16807 15892 16819 15895
rect 18414 15892 18420 15904
rect 16807 15864 18420 15892
rect 16807 15861 16819 15864
rect 16761 15855 16819 15861
rect 18414 15852 18420 15864
rect 18472 15852 18478 15904
rect 18598 15852 18604 15904
rect 18656 15892 18662 15904
rect 20824 15892 20852 15991
rect 18656 15864 20852 15892
rect 18656 15852 18662 15864
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 6917 15691 6975 15697
rect 6917 15657 6929 15691
rect 6963 15688 6975 15691
rect 7006 15688 7012 15700
rect 6963 15660 7012 15688
rect 6963 15657 6975 15660
rect 6917 15651 6975 15657
rect 7006 15648 7012 15660
rect 7064 15648 7070 15700
rect 9582 15688 9588 15700
rect 7852 15660 9588 15688
rect 5534 15580 5540 15632
rect 5592 15620 5598 15632
rect 6730 15620 6736 15632
rect 5592 15592 6736 15620
rect 5592 15580 5598 15592
rect 6730 15580 6736 15592
rect 6788 15620 6794 15632
rect 7852 15620 7880 15660
rect 9582 15648 9588 15660
rect 9640 15648 9646 15700
rect 9950 15688 9956 15700
rect 9911 15660 9956 15688
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 10873 15691 10931 15697
rect 10873 15657 10885 15691
rect 10919 15688 10931 15691
rect 11146 15688 11152 15700
rect 10919 15660 11152 15688
rect 10919 15657 10931 15660
rect 10873 15651 10931 15657
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 12434 15648 12440 15700
rect 12492 15688 12498 15700
rect 14185 15691 14243 15697
rect 12492 15660 12537 15688
rect 12492 15648 12498 15660
rect 14185 15657 14197 15691
rect 14231 15688 14243 15691
rect 14458 15688 14464 15700
rect 14231 15660 14464 15688
rect 14231 15657 14243 15660
rect 14185 15651 14243 15657
rect 14458 15648 14464 15660
rect 14516 15648 14522 15700
rect 15381 15691 15439 15697
rect 15381 15657 15393 15691
rect 15427 15688 15439 15691
rect 16022 15688 16028 15700
rect 15427 15660 16028 15688
rect 15427 15657 15439 15660
rect 15381 15651 15439 15657
rect 16022 15648 16028 15660
rect 16080 15648 16086 15700
rect 17678 15688 17684 15700
rect 17639 15660 17684 15688
rect 17678 15648 17684 15660
rect 17736 15648 17742 15700
rect 20254 15688 20260 15700
rect 18524 15660 20260 15688
rect 6788 15592 7880 15620
rect 7944 15592 9168 15620
rect 6788 15580 6794 15592
rect 7944 15561 7972 15592
rect 9140 15564 9168 15592
rect 10226 15580 10232 15632
rect 10284 15620 10290 15632
rect 13630 15620 13636 15632
rect 10284 15592 13636 15620
rect 10284 15580 10290 15592
rect 13630 15580 13636 15592
rect 13688 15580 13694 15632
rect 13998 15580 14004 15632
rect 14056 15620 14062 15632
rect 16298 15620 16304 15632
rect 14056 15592 16304 15620
rect 14056 15580 14062 15592
rect 16298 15580 16304 15592
rect 16356 15620 16362 15632
rect 16945 15623 17003 15629
rect 16945 15620 16957 15623
rect 16356 15592 16957 15620
rect 16356 15580 16362 15592
rect 16945 15589 16957 15592
rect 16991 15589 17003 15623
rect 16945 15583 17003 15589
rect 17402 15580 17408 15632
rect 17460 15620 17466 15632
rect 18524 15620 18552 15660
rect 20254 15648 20260 15660
rect 20312 15648 20318 15700
rect 18690 15620 18696 15632
rect 17460 15592 18552 15620
rect 18651 15592 18696 15620
rect 17460 15580 17466 15592
rect 18690 15580 18696 15592
rect 18748 15580 18754 15632
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15521 7987 15555
rect 8110 15552 8116 15564
rect 8071 15524 8116 15552
rect 7929 15515 7987 15521
rect 8110 15512 8116 15524
rect 8168 15512 8174 15564
rect 9122 15552 9128 15564
rect 9083 15524 9128 15552
rect 9122 15512 9128 15524
rect 9180 15512 9186 15564
rect 10962 15512 10968 15564
rect 11020 15552 11026 15564
rect 13081 15555 13139 15561
rect 13081 15552 13093 15555
rect 11020 15524 13093 15552
rect 11020 15512 11026 15524
rect 13081 15521 13093 15524
rect 13127 15521 13139 15555
rect 13081 15515 13139 15521
rect 6454 15484 6460 15496
rect 6415 15456 6460 15484
rect 6454 15444 6460 15456
rect 6512 15444 6518 15496
rect 7561 15487 7619 15493
rect 7561 15453 7573 15487
rect 7607 15484 7619 15487
rect 7742 15484 7748 15496
rect 7607 15456 7748 15484
rect 7607 15453 7619 15456
rect 7561 15447 7619 15453
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 9306 15484 9312 15496
rect 9267 15456 9312 15484
rect 9306 15444 9312 15456
rect 9364 15444 9370 15496
rect 10134 15484 10140 15496
rect 10095 15456 10140 15484
rect 10134 15444 10140 15456
rect 10192 15444 10198 15496
rect 13096 15484 13124 15515
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 14458 15552 14464 15564
rect 13872 15524 14464 15552
rect 13872 15512 13878 15524
rect 14458 15512 14464 15524
rect 14516 15512 14522 15564
rect 14734 15552 14740 15564
rect 14695 15524 14740 15552
rect 14734 15512 14740 15524
rect 14792 15512 14798 15564
rect 14918 15512 14924 15564
rect 14976 15552 14982 15564
rect 18233 15555 18291 15561
rect 18233 15552 18245 15555
rect 14976 15524 18245 15552
rect 14976 15512 14982 15524
rect 18233 15521 18245 15524
rect 18279 15521 18291 15555
rect 18233 15515 18291 15521
rect 14936 15484 14964 15512
rect 13096 15456 14964 15484
rect 15197 15487 15255 15493
rect 15197 15453 15209 15487
rect 15243 15453 15255 15487
rect 15197 15447 15255 15453
rect 6178 15416 6184 15428
rect 6139 15388 6184 15416
rect 6178 15376 6184 15388
rect 6236 15376 6242 15428
rect 6914 15416 6920 15428
rect 6472 15388 6920 15416
rect 5721 15351 5779 15357
rect 5721 15317 5733 15351
rect 5767 15348 5779 15351
rect 5810 15348 5816 15360
rect 5767 15320 5816 15348
rect 5767 15317 5779 15320
rect 5721 15311 5779 15317
rect 5810 15308 5816 15320
rect 5868 15348 5874 15360
rect 6472 15348 6500 15388
rect 6914 15376 6920 15388
rect 6972 15376 6978 15428
rect 7282 15376 7288 15428
rect 7340 15416 7346 15428
rect 8202 15416 8208 15428
rect 7340 15388 8208 15416
rect 7340 15376 7346 15388
rect 8202 15376 8208 15388
rect 8260 15416 8266 15428
rect 10870 15416 10876 15428
rect 8260 15388 10876 15416
rect 8260 15376 8266 15388
rect 10870 15376 10876 15388
rect 10928 15376 10934 15428
rect 12158 15416 12164 15428
rect 12119 15388 12164 15416
rect 12158 15376 12164 15388
rect 12216 15376 12222 15428
rect 12805 15419 12863 15425
rect 12805 15385 12817 15419
rect 12851 15416 12863 15419
rect 13449 15419 13507 15425
rect 13449 15416 13461 15419
rect 12851 15388 13461 15416
rect 12851 15385 12863 15388
rect 12805 15379 12863 15385
rect 13449 15385 13461 15388
rect 13495 15385 13507 15419
rect 13449 15379 13507 15385
rect 13538 15376 13544 15428
rect 13596 15416 13602 15428
rect 15212 15416 15240 15447
rect 18046 15444 18052 15496
rect 18104 15484 18110 15496
rect 18877 15487 18935 15493
rect 18877 15484 18889 15487
rect 18104 15456 18889 15484
rect 18104 15444 18110 15456
rect 18877 15453 18889 15456
rect 18923 15453 18935 15487
rect 18877 15447 18935 15453
rect 20358 15487 20416 15493
rect 20358 15453 20370 15487
rect 20404 15453 20416 15487
rect 20622 15484 20628 15496
rect 20583 15456 20628 15484
rect 20358 15447 20416 15453
rect 15654 15416 15660 15428
rect 13596 15388 15240 15416
rect 15615 15388 15660 15416
rect 13596 15376 13602 15388
rect 15654 15376 15660 15388
rect 15712 15376 15718 15428
rect 18230 15416 18236 15428
rect 18064 15388 18236 15416
rect 6638 15348 6644 15360
rect 5868 15320 6500 15348
rect 6599 15320 6644 15348
rect 5868 15308 5874 15320
rect 6638 15308 6644 15320
rect 6696 15308 6702 15360
rect 8573 15351 8631 15357
rect 8573 15317 8585 15351
rect 8619 15348 8631 15351
rect 8662 15348 8668 15360
rect 8619 15320 8668 15348
rect 8619 15317 8631 15320
rect 8573 15311 8631 15317
rect 8662 15308 8668 15320
rect 8720 15308 8726 15360
rect 8754 15308 8760 15360
rect 8812 15348 8818 15360
rect 9217 15351 9275 15357
rect 9217 15348 9229 15351
rect 8812 15320 9229 15348
rect 8812 15308 8818 15320
rect 9217 15317 9229 15320
rect 9263 15317 9275 15351
rect 9217 15311 9275 15317
rect 9582 15308 9588 15360
rect 9640 15348 9646 15360
rect 9677 15351 9735 15357
rect 9677 15348 9689 15351
rect 9640 15320 9689 15348
rect 9640 15308 9646 15320
rect 9677 15317 9689 15320
rect 9723 15317 9735 15351
rect 9677 15311 9735 15317
rect 9858 15308 9864 15360
rect 9916 15348 9922 15360
rect 12250 15348 12256 15360
rect 9916 15320 12256 15348
rect 9916 15308 9922 15320
rect 12250 15308 12256 15320
rect 12308 15308 12314 15360
rect 12897 15351 12955 15357
rect 12897 15317 12909 15351
rect 12943 15348 12955 15351
rect 13814 15348 13820 15360
rect 12943 15320 13820 15348
rect 12943 15317 12955 15320
rect 12897 15311 12955 15317
rect 13814 15308 13820 15320
rect 13872 15308 13878 15360
rect 14550 15348 14556 15360
rect 14511 15320 14556 15348
rect 14550 15308 14556 15320
rect 14608 15308 14614 15360
rect 14645 15351 14703 15357
rect 14645 15317 14657 15351
rect 14691 15348 14703 15351
rect 15102 15348 15108 15360
rect 14691 15320 15108 15348
rect 14691 15317 14703 15320
rect 14645 15311 14703 15317
rect 15102 15308 15108 15320
rect 15160 15308 15166 15360
rect 18064 15357 18092 15388
rect 18230 15376 18236 15388
rect 18288 15416 18294 15428
rect 18966 15416 18972 15428
rect 18288 15388 18972 15416
rect 18288 15376 18294 15388
rect 18966 15376 18972 15388
rect 19024 15376 19030 15428
rect 19794 15416 19800 15428
rect 19076 15388 19800 15416
rect 18049 15351 18107 15357
rect 18049 15317 18061 15351
rect 18095 15317 18107 15351
rect 18049 15311 18107 15317
rect 18141 15351 18199 15357
rect 18141 15317 18153 15351
rect 18187 15348 18199 15351
rect 19076 15348 19104 15388
rect 19794 15376 19800 15388
rect 19852 15376 19858 15428
rect 20364 15416 20392 15447
rect 20622 15444 20628 15456
rect 20680 15444 20686 15496
rect 21085 15487 21143 15493
rect 21085 15453 21097 15487
rect 21131 15453 21143 15487
rect 21085 15447 21143 15453
rect 20438 15416 20444 15428
rect 20364 15388 20444 15416
rect 20438 15376 20444 15388
rect 20496 15376 20502 15428
rect 19242 15348 19248 15360
rect 18187 15320 19104 15348
rect 19203 15320 19248 15348
rect 18187 15317 18199 15320
rect 18141 15311 18199 15317
rect 19242 15308 19248 15320
rect 19300 15308 19306 15360
rect 20070 15308 20076 15360
rect 20128 15348 20134 15360
rect 21100 15348 21128 15447
rect 20128 15320 21128 15348
rect 21269 15351 21327 15357
rect 20128 15308 20134 15320
rect 21269 15317 21281 15351
rect 21315 15348 21327 15351
rect 21358 15348 21364 15360
rect 21315 15320 21364 15348
rect 21315 15317 21327 15320
rect 21269 15311 21327 15317
rect 21358 15308 21364 15320
rect 21416 15308 21422 15360
rect 1104 15258 21896 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21896 15258
rect 1104 15184 21896 15206
rect 7190 15104 7196 15156
rect 7248 15144 7254 15156
rect 8754 15144 8760 15156
rect 7248 15116 8760 15144
rect 7248 15104 7254 15116
rect 8754 15104 8760 15116
rect 8812 15104 8818 15156
rect 9122 15144 9128 15156
rect 8956 15116 9128 15144
rect 7469 15079 7527 15085
rect 7469 15045 7481 15079
rect 7515 15076 7527 15079
rect 8869 15079 8927 15085
rect 7515 15048 8800 15076
rect 7515 15045 7527 15048
rect 7469 15039 7527 15045
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 15008 6883 15011
rect 8110 15008 8116 15020
rect 6871 14980 8116 15008
rect 6871 14977 6883 14980
rect 6825 14971 6883 14977
rect 8110 14968 8116 14980
rect 8168 14968 8174 15020
rect 8772 15008 8800 15048
rect 8869 15045 8881 15079
rect 8915 15076 8927 15079
rect 8956 15076 8984 15116
rect 9122 15104 9128 15116
rect 9180 15104 9186 15156
rect 9766 15144 9772 15156
rect 9727 15116 9772 15144
rect 9766 15104 9772 15116
rect 9824 15104 9830 15156
rect 9968 15116 11192 15144
rect 9968 15076 9996 15116
rect 11164 15076 11192 15116
rect 11238 15104 11244 15156
rect 11296 15144 11302 15156
rect 11517 15147 11575 15153
rect 11517 15144 11529 15147
rect 11296 15116 11529 15144
rect 11296 15104 11302 15116
rect 11517 15113 11529 15116
rect 11563 15113 11575 15147
rect 11517 15107 11575 15113
rect 11698 15104 11704 15156
rect 11756 15144 11762 15156
rect 12066 15144 12072 15156
rect 11756 15116 12072 15144
rect 11756 15104 11762 15116
rect 12066 15104 12072 15116
rect 12124 15104 12130 15156
rect 12250 15104 12256 15156
rect 12308 15144 12314 15156
rect 13357 15147 13415 15153
rect 13357 15144 13369 15147
rect 12308 15116 13369 15144
rect 12308 15104 12314 15116
rect 13357 15113 13369 15116
rect 13403 15144 13415 15147
rect 13403 15116 14412 15144
rect 13403 15113 13415 15116
rect 13357 15107 13415 15113
rect 11790 15076 11796 15088
rect 8915 15048 8984 15076
rect 9048 15048 9996 15076
rect 10060 15048 11100 15076
rect 11164 15048 11796 15076
rect 8915 15045 8927 15048
rect 8869 15039 8927 15045
rect 9048 15008 9076 15048
rect 8772 14980 9076 15008
rect 9125 15011 9183 15017
rect 9125 14977 9137 15011
rect 9171 15008 9183 15011
rect 10060 15008 10088 15048
rect 9171 14980 10088 15008
rect 9171 14977 9183 14980
rect 9125 14971 9183 14977
rect 10870 14968 10876 15020
rect 10928 15017 10934 15020
rect 10928 15008 10940 15017
rect 11072 15008 11100 15048
rect 11790 15036 11796 15048
rect 11848 15036 11854 15088
rect 11885 15079 11943 15085
rect 11885 15045 11897 15079
rect 11931 15076 11943 15079
rect 12434 15076 12440 15088
rect 11931 15048 12440 15076
rect 11931 15045 11943 15048
rect 11885 15039 11943 15045
rect 12434 15036 12440 15048
rect 12492 15036 12498 15088
rect 14274 15085 14280 15088
rect 14268 15076 14280 15085
rect 14235 15048 14280 15076
rect 14268 15039 14280 15048
rect 14274 15036 14280 15039
rect 14332 15036 14338 15088
rect 14384 15076 14412 15116
rect 16206 15104 16212 15156
rect 16264 15144 16270 15156
rect 16301 15147 16359 15153
rect 16301 15144 16313 15147
rect 16264 15116 16313 15144
rect 16264 15104 16270 15116
rect 16301 15113 16313 15116
rect 16347 15113 16359 15147
rect 16301 15107 16359 15113
rect 18049 15147 18107 15153
rect 18049 15113 18061 15147
rect 18095 15144 18107 15147
rect 18322 15144 18328 15156
rect 18095 15116 18328 15144
rect 18095 15113 18107 15116
rect 18049 15107 18107 15113
rect 18322 15104 18328 15116
rect 18380 15104 18386 15156
rect 18506 15144 18512 15156
rect 18432 15116 18512 15144
rect 17034 15076 17040 15088
rect 14384 15048 17040 15076
rect 17034 15036 17040 15048
rect 17092 15036 17098 15088
rect 17586 15036 17592 15088
rect 17644 15076 17650 15088
rect 18432 15076 18460 15116
rect 18506 15104 18512 15116
rect 18564 15144 18570 15156
rect 18785 15147 18843 15153
rect 18785 15144 18797 15147
rect 18564 15116 18797 15144
rect 18564 15104 18570 15116
rect 18785 15113 18797 15116
rect 18831 15113 18843 15147
rect 18785 15107 18843 15113
rect 19426 15104 19432 15156
rect 19484 15144 19490 15156
rect 20622 15144 20628 15156
rect 19484 15116 20628 15144
rect 19484 15104 19490 15116
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 20806 15144 20812 15156
rect 20767 15116 20812 15144
rect 20806 15104 20812 15116
rect 20864 15104 20870 15156
rect 19242 15076 19248 15088
rect 17644 15048 18460 15076
rect 18524 15048 19248 15076
rect 17644 15036 17650 15048
rect 11146 15008 11152 15020
rect 10928 14980 10973 15008
rect 11072 14980 11152 15008
rect 10928 14971 10940 14980
rect 10928 14968 10934 14971
rect 11146 14968 11152 14980
rect 11204 14968 11210 15020
rect 12526 15008 12532 15020
rect 12487 14980 12532 15008
rect 12526 14968 12532 14980
rect 12584 14968 12590 15020
rect 13998 15008 14004 15020
rect 13959 14980 14004 15008
rect 13998 14968 14004 14980
rect 14056 14968 14062 15020
rect 14550 14968 14556 15020
rect 14608 15008 14614 15020
rect 14734 15008 14740 15020
rect 14608 14980 14740 15008
rect 14608 14968 14614 14980
rect 14734 14968 14740 14980
rect 14792 14968 14798 15020
rect 15657 15011 15715 15017
rect 15657 15008 15669 15011
rect 15396 14980 15669 15008
rect 9493 14943 9551 14949
rect 9493 14909 9505 14943
rect 9539 14940 9551 14943
rect 9858 14940 9864 14952
rect 9539 14912 9864 14940
rect 9539 14909 9551 14912
rect 9493 14903 9551 14909
rect 9858 14900 9864 14912
rect 9916 14900 9922 14952
rect 11974 14940 11980 14952
rect 11935 14912 11980 14940
rect 11974 14900 11980 14912
rect 12032 14900 12038 14952
rect 12069 14943 12127 14949
rect 12069 14909 12081 14943
rect 12115 14909 12127 14943
rect 12069 14903 12127 14909
rect 13081 14943 13139 14949
rect 13081 14909 13093 14943
rect 13127 14909 13139 14943
rect 13262 14940 13268 14952
rect 13223 14912 13268 14940
rect 13081 14903 13139 14909
rect 6822 14832 6828 14884
rect 6880 14872 6886 14884
rect 6880 14844 8248 14872
rect 6880 14832 6886 14844
rect 6454 14804 6460 14816
rect 6415 14776 6460 14804
rect 6454 14764 6460 14776
rect 6512 14764 6518 14816
rect 7006 14804 7012 14816
rect 6967 14776 7012 14804
rect 7006 14764 7012 14776
rect 7064 14764 7070 14816
rect 7742 14804 7748 14816
rect 7703 14776 7748 14804
rect 7742 14764 7748 14776
rect 7800 14764 7806 14816
rect 8220 14804 8248 14844
rect 9324 14844 9674 14872
rect 9324 14804 9352 14844
rect 8220 14776 9352 14804
rect 9646 14804 9674 14844
rect 11146 14832 11152 14884
rect 11204 14872 11210 14884
rect 12084 14872 12112 14903
rect 11204 14844 12112 14872
rect 13096 14872 13124 14903
rect 13262 14900 13268 14912
rect 13320 14900 13326 14952
rect 13814 14872 13820 14884
rect 13096 14844 13820 14872
rect 11204 14832 11210 14844
rect 13814 14832 13820 14844
rect 13872 14832 13878 14884
rect 11238 14804 11244 14816
rect 9646 14776 11244 14804
rect 11238 14764 11244 14776
rect 11296 14764 11302 14816
rect 12713 14807 12771 14813
rect 12713 14773 12725 14807
rect 12759 14804 12771 14807
rect 13630 14804 13636 14816
rect 12759 14776 13636 14804
rect 12759 14773 12771 14776
rect 12713 14767 12771 14773
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 13725 14807 13783 14813
rect 13725 14773 13737 14807
rect 13771 14804 13783 14807
rect 14366 14804 14372 14816
rect 13771 14776 14372 14804
rect 13771 14773 13783 14776
rect 13725 14767 13783 14773
rect 14366 14764 14372 14776
rect 14424 14764 14430 14816
rect 14642 14764 14648 14816
rect 14700 14804 14706 14816
rect 15396 14813 15424 14980
rect 15657 14977 15669 14980
rect 15703 14977 15715 15011
rect 15657 14971 15715 14977
rect 16669 15011 16727 15017
rect 16669 14977 16681 15011
rect 16715 15008 16727 15011
rect 16942 15008 16948 15020
rect 16715 14980 16948 15008
rect 16715 14977 16727 14980
rect 16669 14971 16727 14977
rect 16942 14968 16948 14980
rect 17000 14968 17006 15020
rect 17862 15008 17868 15020
rect 17823 14980 17868 15008
rect 17862 14968 17868 14980
rect 17920 14968 17926 15020
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 17586 14940 17592 14952
rect 15528 14912 17592 14940
rect 15528 14900 15534 14912
rect 17586 14900 17592 14912
rect 17644 14900 17650 14952
rect 18524 14949 18552 15048
rect 19242 15036 19248 15048
rect 19300 15076 19306 15088
rect 19696 15079 19754 15085
rect 19696 15076 19708 15079
rect 19300 15048 19708 15076
rect 19300 15036 19306 15048
rect 19696 15045 19708 15048
rect 19742 15076 19754 15079
rect 20990 15076 20996 15088
rect 19742 15048 20996 15076
rect 19742 15045 19754 15048
rect 19696 15039 19754 15045
rect 20990 15036 20996 15048
rect 21048 15036 21054 15088
rect 19426 15008 19432 15020
rect 19387 14980 19432 15008
rect 19426 14968 19432 14980
rect 19484 14968 19490 15020
rect 20714 15008 20720 15020
rect 19536 14980 20720 15008
rect 18509 14943 18567 14949
rect 18509 14909 18521 14943
rect 18555 14909 18567 14943
rect 18690 14940 18696 14952
rect 18651 14912 18696 14940
rect 18509 14903 18567 14909
rect 18690 14900 18696 14912
rect 18748 14900 18754 14952
rect 19536 14940 19564 14980
rect 20714 14968 20720 14980
rect 20772 14968 20778 15020
rect 21082 15008 21088 15020
rect 21043 14980 21088 15008
rect 21082 14968 21088 14980
rect 21140 14968 21146 15020
rect 18800 14912 19564 14940
rect 15562 14832 15568 14884
rect 15620 14872 15626 14884
rect 18800 14872 18828 14912
rect 15620 14844 18828 14872
rect 15620 14832 15626 14844
rect 15381 14807 15439 14813
rect 15381 14804 15393 14807
rect 14700 14776 15393 14804
rect 14700 14764 14706 14776
rect 15381 14773 15393 14776
rect 15427 14773 15439 14807
rect 17310 14804 17316 14816
rect 17271 14776 17316 14804
rect 15381 14767 15439 14773
rect 17310 14764 17316 14776
rect 17368 14764 17374 14816
rect 19153 14807 19211 14813
rect 19153 14773 19165 14807
rect 19199 14804 19211 14807
rect 20438 14804 20444 14816
rect 19199 14776 20444 14804
rect 19199 14773 19211 14776
rect 19153 14767 19211 14773
rect 20438 14764 20444 14776
rect 20496 14764 20502 14816
rect 21266 14804 21272 14816
rect 21227 14776 21272 14804
rect 21266 14764 21272 14776
rect 21324 14764 21330 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 6546 14560 6552 14612
rect 6604 14600 6610 14612
rect 6733 14603 6791 14609
rect 6733 14600 6745 14603
rect 6604 14572 6745 14600
rect 6604 14560 6610 14572
rect 6733 14569 6745 14572
rect 6779 14569 6791 14603
rect 6733 14563 6791 14569
rect 7006 14560 7012 14612
rect 7064 14600 7070 14612
rect 16301 14603 16359 14609
rect 7064 14572 16252 14600
rect 7064 14560 7070 14572
rect 4430 14492 4436 14544
rect 4488 14532 4494 14544
rect 7469 14535 7527 14541
rect 7469 14532 7481 14535
rect 4488 14504 7481 14532
rect 4488 14492 4494 14504
rect 7469 14501 7481 14504
rect 7515 14501 7527 14535
rect 7469 14495 7527 14501
rect 7742 14492 7748 14544
rect 7800 14532 7806 14544
rect 11882 14532 11888 14544
rect 7800 14504 9812 14532
rect 11843 14504 11888 14532
rect 7800 14492 7806 14504
rect 7006 14424 7012 14476
rect 7064 14464 7070 14476
rect 7190 14464 7196 14476
rect 7064 14436 7196 14464
rect 7064 14424 7070 14436
rect 7190 14424 7196 14436
rect 7248 14424 7254 14476
rect 7668 14436 9076 14464
rect 5534 14356 5540 14408
rect 5592 14396 5598 14408
rect 5994 14396 6000 14408
rect 5592 14368 6000 14396
rect 5592 14356 5598 14368
rect 5994 14356 6000 14368
rect 6052 14356 6058 14408
rect 7668 14405 7696 14436
rect 7653 14399 7711 14405
rect 7653 14365 7665 14399
rect 7699 14365 7711 14399
rect 7653 14359 7711 14365
rect 8562 14399 8620 14405
rect 8562 14365 8574 14399
rect 8608 14365 8620 14399
rect 9048 14396 9076 14436
rect 9122 14424 9128 14476
rect 9180 14464 9186 14476
rect 9784 14473 9812 14504
rect 11882 14492 11888 14504
rect 11940 14492 11946 14544
rect 13725 14535 13783 14541
rect 13725 14501 13737 14535
rect 13771 14501 13783 14535
rect 13725 14495 13783 14501
rect 9677 14467 9735 14473
rect 9677 14464 9689 14467
rect 9180 14436 9689 14464
rect 9180 14424 9186 14436
rect 9677 14433 9689 14436
rect 9723 14433 9735 14467
rect 9677 14427 9735 14433
rect 9769 14467 9827 14473
rect 9769 14433 9781 14467
rect 9815 14433 9827 14467
rect 9769 14427 9827 14433
rect 11238 14424 11244 14476
rect 11296 14464 11302 14476
rect 13740 14464 13768 14495
rect 13998 14492 14004 14544
rect 14056 14532 14062 14544
rect 14056 14504 15608 14532
rect 14056 14492 14062 14504
rect 15580 14476 15608 14504
rect 15663 14504 16160 14532
rect 14182 14464 14188 14476
rect 11296 14436 12480 14464
rect 13740 14436 14188 14464
rect 11296 14424 11302 14436
rect 9582 14396 9588 14408
rect 9048 14368 9444 14396
rect 9543 14368 9588 14396
rect 8562 14359 8620 14365
rect 8588 14328 8616 14359
rect 9306 14328 9312 14340
rect 8588 14300 9312 14328
rect 9306 14288 9312 14300
rect 9364 14288 9370 14340
rect 9416 14328 9444 14368
rect 9582 14356 9588 14368
rect 9640 14356 9646 14408
rect 10229 14399 10287 14405
rect 10229 14365 10241 14399
rect 10275 14396 10287 14399
rect 10870 14396 10876 14408
rect 10275 14368 10876 14396
rect 10275 14365 10287 14368
rect 10229 14359 10287 14365
rect 10870 14356 10876 14368
rect 10928 14356 10934 14408
rect 12069 14399 12127 14405
rect 12069 14365 12081 14399
rect 12115 14365 12127 14399
rect 12342 14396 12348 14408
rect 12303 14368 12348 14396
rect 12069 14359 12127 14365
rect 10042 14328 10048 14340
rect 9416 14300 10048 14328
rect 10042 14288 10048 14300
rect 10100 14288 10106 14340
rect 10496 14331 10554 14337
rect 10496 14297 10508 14331
rect 10542 14328 10554 14331
rect 10962 14328 10968 14340
rect 10542 14300 10968 14328
rect 10542 14297 10554 14300
rect 10496 14291 10554 14297
rect 10962 14288 10968 14300
rect 11020 14288 11026 14340
rect 12084 14328 12112 14359
rect 12342 14356 12348 14368
rect 12400 14356 12406 14408
rect 12452 14392 12480 14436
rect 14182 14424 14188 14436
rect 14240 14424 14246 14476
rect 14366 14464 14372 14476
rect 14327 14436 14372 14464
rect 14366 14424 14372 14436
rect 14424 14424 14430 14476
rect 15562 14464 15568 14476
rect 15523 14436 15568 14464
rect 15562 14424 15568 14436
rect 15620 14424 15626 14476
rect 15663 14396 15691 14504
rect 15749 14467 15807 14473
rect 15749 14433 15761 14467
rect 15795 14433 15807 14467
rect 15749 14427 15807 14433
rect 12544 14392 15691 14396
rect 12452 14368 15691 14392
rect 12452 14364 12572 14368
rect 12250 14328 12256 14340
rect 12084 14300 12256 14328
rect 12250 14288 12256 14300
rect 12308 14288 12314 14340
rect 12612 14331 12670 14337
rect 12612 14297 12624 14331
rect 12658 14328 12670 14331
rect 13814 14328 13820 14340
rect 12658 14300 13820 14328
rect 12658 14297 12670 14300
rect 12612 14291 12670 14297
rect 13814 14288 13820 14300
rect 13872 14328 13878 14340
rect 14090 14328 14096 14340
rect 13872 14300 14096 14328
rect 13872 14288 13878 14300
rect 14090 14288 14096 14300
rect 14148 14328 14154 14340
rect 15764 14328 15792 14427
rect 16132 14405 16160 14504
rect 16117 14399 16175 14405
rect 16117 14365 16129 14399
rect 16163 14365 16175 14399
rect 16224 14396 16252 14572
rect 16301 14569 16313 14603
rect 16347 14600 16359 14603
rect 17862 14600 17868 14612
rect 16347 14572 17868 14600
rect 16347 14569 16359 14572
rect 16301 14563 16359 14569
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 18782 14600 18788 14612
rect 18743 14572 18788 14600
rect 18782 14560 18788 14572
rect 18840 14560 18846 14612
rect 19610 14600 19616 14612
rect 19571 14572 19616 14600
rect 19610 14560 19616 14572
rect 19668 14560 19674 14612
rect 18141 14467 18199 14473
rect 18141 14433 18153 14467
rect 18187 14464 18199 14467
rect 19518 14464 19524 14476
rect 18187 14436 19524 14464
rect 18187 14433 18199 14436
rect 18141 14427 18199 14433
rect 19518 14424 19524 14436
rect 19576 14424 19582 14476
rect 20438 14464 20444 14476
rect 20399 14436 20444 14464
rect 20438 14424 20444 14436
rect 20496 14424 20502 14476
rect 20625 14467 20683 14473
rect 20625 14433 20637 14467
rect 20671 14464 20683 14467
rect 20806 14464 20812 14476
rect 20671 14436 20812 14464
rect 20671 14433 20683 14436
rect 20625 14427 20683 14433
rect 20806 14424 20812 14436
rect 20864 14424 20870 14476
rect 18601 14399 18659 14405
rect 18601 14396 18613 14399
rect 16224 14368 18613 14396
rect 16117 14359 16175 14365
rect 18601 14365 18613 14368
rect 18647 14365 18659 14399
rect 19426 14396 19432 14408
rect 19387 14368 19432 14396
rect 18601 14359 18659 14365
rect 19426 14356 19432 14368
rect 19484 14356 19490 14408
rect 20993 14399 21051 14405
rect 20993 14365 21005 14399
rect 21039 14365 21051 14399
rect 20993 14359 21051 14365
rect 14148 14300 16252 14328
rect 14148 14288 14154 14300
rect 16224 14272 16252 14300
rect 17770 14288 17776 14340
rect 17828 14328 17834 14340
rect 17874 14331 17932 14337
rect 17874 14328 17886 14331
rect 17828 14300 17886 14328
rect 17828 14288 17834 14300
rect 17874 14297 17886 14300
rect 17920 14297 17932 14331
rect 17874 14291 17932 14297
rect 18230 14288 18236 14340
rect 18288 14328 18294 14340
rect 21008 14328 21036 14359
rect 18288 14300 21036 14328
rect 18288 14288 18294 14300
rect 7742 14220 7748 14272
rect 7800 14260 7806 14272
rect 7929 14263 7987 14269
rect 7929 14260 7941 14263
rect 7800 14232 7941 14260
rect 7800 14220 7806 14232
rect 7929 14229 7941 14232
rect 7975 14229 7987 14263
rect 7929 14223 7987 14229
rect 8294 14220 8300 14272
rect 8352 14260 8358 14272
rect 9217 14263 9275 14269
rect 9217 14260 9229 14263
rect 8352 14232 9229 14260
rect 8352 14220 8358 14232
rect 9217 14229 9229 14232
rect 9263 14229 9275 14263
rect 9217 14223 9275 14229
rect 11609 14263 11667 14269
rect 11609 14229 11621 14263
rect 11655 14260 11667 14263
rect 11698 14260 11704 14272
rect 11655 14232 11704 14260
rect 11655 14229 11667 14232
rect 11609 14223 11667 14229
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 13998 14260 14004 14272
rect 11940 14232 14004 14260
rect 11940 14220 11946 14232
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 14458 14220 14464 14272
rect 14516 14260 14522 14272
rect 14826 14260 14832 14272
rect 14516 14232 14561 14260
rect 14787 14232 14832 14260
rect 14516 14220 14522 14232
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 14918 14220 14924 14272
rect 14976 14260 14982 14272
rect 15105 14263 15163 14269
rect 15105 14260 15117 14263
rect 14976 14232 15117 14260
rect 14976 14220 14982 14232
rect 15105 14229 15117 14232
rect 15151 14229 15163 14263
rect 15470 14260 15476 14272
rect 15431 14232 15476 14260
rect 15105 14223 15163 14229
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 16206 14220 16212 14272
rect 16264 14260 16270 14272
rect 16761 14263 16819 14269
rect 16761 14260 16773 14263
rect 16264 14232 16773 14260
rect 16264 14220 16270 14232
rect 16761 14229 16773 14232
rect 16807 14229 16819 14263
rect 16761 14223 16819 14229
rect 17218 14220 17224 14272
rect 17276 14260 17282 14272
rect 19981 14263 20039 14269
rect 19981 14260 19993 14263
rect 17276 14232 19993 14260
rect 17276 14220 17282 14232
rect 19981 14229 19993 14232
rect 20027 14229 20039 14263
rect 20346 14260 20352 14272
rect 20307 14232 20352 14260
rect 19981 14223 20039 14229
rect 20346 14220 20352 14232
rect 20404 14220 20410 14272
rect 21174 14260 21180 14272
rect 21135 14232 21180 14260
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 1104 14170 21896 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21896 14170
rect 1104 14096 21896 14118
rect 8110 14056 8116 14068
rect 8071 14028 8116 14056
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 9306 14016 9312 14068
rect 9364 14056 9370 14068
rect 9493 14059 9551 14065
rect 9493 14056 9505 14059
rect 9364 14028 9505 14056
rect 9364 14016 9370 14028
rect 9493 14025 9505 14028
rect 9539 14056 9551 14059
rect 11146 14056 11152 14068
rect 9539 14028 11152 14056
rect 9539 14025 9551 14028
rect 9493 14019 9551 14025
rect 11146 14016 11152 14028
rect 11204 14016 11210 14068
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14056 11575 14059
rect 12986 14056 12992 14068
rect 11563 14028 12992 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 7837 13991 7895 13997
rect 7837 13957 7849 13991
rect 7883 13988 7895 13991
rect 8202 13988 8208 14000
rect 7883 13960 8208 13988
rect 7883 13957 7895 13960
rect 7837 13951 7895 13957
rect 8202 13948 8208 13960
rect 8260 13948 8266 14000
rect 9858 13988 9864 14000
rect 8496 13960 9864 13988
rect 3878 13880 3884 13932
rect 3936 13920 3942 13932
rect 8294 13920 8300 13932
rect 3936 13892 8156 13920
rect 8255 13892 8300 13920
rect 3936 13880 3942 13892
rect 7098 13812 7104 13864
rect 7156 13852 7162 13864
rect 7377 13855 7435 13861
rect 7377 13852 7389 13855
rect 7156 13824 7389 13852
rect 7156 13812 7162 13824
rect 7377 13821 7389 13824
rect 7423 13821 7435 13855
rect 8128 13852 8156 13892
rect 8294 13880 8300 13892
rect 8352 13880 8358 13932
rect 8496 13852 8524 13960
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 10628 13991 10686 13997
rect 10628 13957 10640 13991
rect 10674 13988 10686 13991
rect 11532 13988 11560 14019
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 14274 14016 14280 14068
rect 14332 14056 14338 14068
rect 14369 14059 14427 14065
rect 14369 14056 14381 14059
rect 14332 14028 14381 14056
rect 14332 14016 14338 14028
rect 14369 14025 14381 14028
rect 14415 14025 14427 14059
rect 14369 14019 14427 14025
rect 14458 14016 14464 14068
rect 14516 14056 14522 14068
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 14516 14028 14749 14056
rect 14516 14016 14522 14028
rect 14737 14025 14749 14028
rect 14783 14025 14795 14059
rect 14737 14019 14795 14025
rect 14918 14016 14924 14068
rect 14976 14056 14982 14068
rect 15381 14059 15439 14065
rect 15381 14056 15393 14059
rect 14976 14028 15393 14056
rect 14976 14016 14982 14028
rect 15381 14025 15393 14028
rect 15427 14025 15439 14059
rect 15381 14019 15439 14025
rect 15562 14016 15568 14068
rect 15620 14056 15626 14068
rect 18325 14059 18383 14065
rect 18325 14056 18337 14059
rect 15620 14028 18337 14056
rect 15620 14016 15626 14028
rect 18325 14025 18337 14028
rect 18371 14025 18383 14059
rect 18325 14019 18383 14025
rect 19337 14059 19395 14065
rect 19337 14025 19349 14059
rect 19383 14056 19395 14059
rect 19610 14056 19616 14068
rect 19383 14028 19616 14056
rect 19383 14025 19395 14028
rect 19337 14019 19395 14025
rect 19610 14016 19616 14028
rect 19668 14016 19674 14068
rect 19794 14016 19800 14068
rect 19852 14016 19858 14068
rect 20346 14056 20352 14068
rect 20307 14028 20352 14056
rect 20346 14016 20352 14028
rect 20404 14016 20410 14068
rect 10674 13960 11560 13988
rect 10674 13957 10686 13960
rect 10628 13951 10686 13957
rect 12342 13948 12348 14000
rect 12400 13988 12406 14000
rect 13725 13991 13783 13997
rect 12400 13960 12940 13988
rect 12400 13948 12406 13960
rect 9217 13923 9275 13929
rect 9217 13889 9229 13923
rect 9263 13920 9275 13923
rect 10318 13920 10324 13932
rect 9263 13892 10324 13920
rect 9263 13889 9275 13892
rect 9217 13883 9275 13889
rect 10318 13880 10324 13892
rect 10376 13880 10382 13932
rect 10870 13920 10876 13932
rect 10783 13892 10876 13920
rect 10870 13880 10876 13892
rect 10928 13920 10934 13932
rect 12360 13920 12388 13948
rect 12618 13920 12624 13932
rect 12676 13929 12682 13932
rect 12912 13929 12940 13960
rect 13725 13957 13737 13991
rect 13771 13988 13783 13991
rect 15470 13988 15476 14000
rect 13771 13960 15476 13988
rect 13771 13957 13783 13960
rect 13725 13951 13783 13957
rect 15470 13948 15476 13960
rect 15528 13948 15534 14000
rect 19705 13991 19763 13997
rect 15580 13960 17724 13988
rect 10928 13892 12388 13920
rect 12588 13892 12624 13920
rect 10928 13880 10934 13892
rect 12618 13880 12624 13892
rect 12676 13883 12688 13929
rect 12897 13923 12955 13929
rect 12897 13889 12909 13923
rect 12943 13889 12955 13923
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 12897 13883 12955 13889
rect 13740 13892 14289 13920
rect 12676 13880 12682 13883
rect 13740 13864 13768 13892
rect 14277 13889 14289 13892
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 8128 13824 8524 13852
rect 8573 13855 8631 13861
rect 7377 13815 7435 13821
rect 8573 13821 8585 13855
rect 8619 13852 8631 13855
rect 9858 13852 9864 13864
rect 8619 13824 9864 13852
rect 8619 13821 8631 13824
rect 8573 13815 8631 13821
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 13722 13812 13728 13864
rect 13780 13812 13786 13864
rect 14090 13852 14096 13864
rect 14051 13824 14096 13852
rect 14090 13812 14096 13824
rect 14148 13812 14154 13864
rect 14292 13852 14320 13883
rect 14734 13880 14740 13932
rect 14792 13920 14798 13932
rect 15580 13920 15608 13960
rect 14792 13892 15608 13920
rect 16936 13923 16994 13929
rect 14792 13880 14798 13892
rect 16936 13889 16948 13923
rect 16982 13920 16994 13923
rect 17218 13920 17224 13932
rect 16982 13892 17224 13920
rect 16982 13889 16994 13892
rect 16936 13883 16994 13889
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 15102 13852 15108 13864
rect 14292 13824 15108 13852
rect 15102 13812 15108 13824
rect 15160 13812 15166 13864
rect 15470 13852 15476 13864
rect 15431 13824 15476 13852
rect 15470 13812 15476 13824
rect 15528 13812 15534 13864
rect 15565 13855 15623 13861
rect 15565 13821 15577 13855
rect 15611 13821 15623 13855
rect 15565 13815 15623 13821
rect 8202 13744 8208 13796
rect 8260 13784 8266 13796
rect 9490 13784 9496 13796
rect 8260 13756 9496 13784
rect 8260 13744 8266 13756
rect 9490 13744 9496 13756
rect 9548 13744 9554 13796
rect 14182 13744 14188 13796
rect 14240 13784 14246 13796
rect 15580 13784 15608 13815
rect 16114 13812 16120 13864
rect 16172 13852 16178 13864
rect 16209 13855 16267 13861
rect 16209 13852 16221 13855
rect 16172 13824 16221 13852
rect 16172 13812 16178 13824
rect 16209 13821 16221 13824
rect 16255 13821 16267 13855
rect 16209 13815 16267 13821
rect 16669 13855 16727 13861
rect 16669 13821 16681 13855
rect 16715 13821 16727 13855
rect 17696 13852 17724 13960
rect 19705 13957 19717 13991
rect 19751 13988 19763 13991
rect 19812 13988 19840 14016
rect 19978 13988 19984 14000
rect 19751 13960 19984 13988
rect 19751 13957 19763 13960
rect 19705 13951 19763 13957
rect 19978 13948 19984 13960
rect 20036 13948 20042 14000
rect 20162 13948 20168 14000
rect 20220 13988 20226 14000
rect 20717 13991 20775 13997
rect 20717 13988 20729 13991
rect 20220 13960 20729 13988
rect 20220 13948 20226 13960
rect 20717 13957 20729 13960
rect 20763 13957 20775 13991
rect 20717 13951 20775 13957
rect 17862 13880 17868 13932
rect 17920 13920 17926 13932
rect 18693 13923 18751 13929
rect 18693 13920 18705 13923
rect 17920 13892 18705 13920
rect 17920 13880 17926 13892
rect 18693 13889 18705 13892
rect 18739 13889 18751 13923
rect 18693 13883 18751 13889
rect 19797 13923 19855 13929
rect 19797 13889 19809 13923
rect 19843 13920 19855 13923
rect 20346 13920 20352 13932
rect 19843 13892 20352 13920
rect 19843 13889 19855 13892
rect 19797 13883 19855 13889
rect 20346 13880 20352 13892
rect 20404 13880 20410 13932
rect 18230 13852 18236 13864
rect 17696 13824 18236 13852
rect 16669 13815 16727 13821
rect 14240 13756 15608 13784
rect 14240 13744 14246 13756
rect 9306 13676 9312 13728
rect 9364 13716 9370 13728
rect 12710 13716 12716 13728
rect 9364 13688 12716 13716
rect 9364 13676 9370 13688
rect 12710 13676 12716 13688
rect 12768 13676 12774 13728
rect 12894 13676 12900 13728
rect 12952 13716 12958 13728
rect 13173 13719 13231 13725
rect 13173 13716 13185 13719
rect 12952 13688 13185 13716
rect 12952 13676 12958 13688
rect 13173 13685 13185 13688
rect 13219 13685 13231 13719
rect 15010 13716 15016 13728
rect 14971 13688 15016 13716
rect 13173 13679 13231 13685
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 16684 13716 16712 13815
rect 18230 13812 18236 13824
rect 18288 13812 18294 13864
rect 18322 13812 18328 13864
rect 18380 13852 18386 13864
rect 18785 13855 18843 13861
rect 18785 13852 18797 13855
rect 18380 13824 18797 13852
rect 18380 13812 18386 13824
rect 18785 13821 18797 13824
rect 18831 13821 18843 13855
rect 18785 13815 18843 13821
rect 18874 13812 18880 13864
rect 18932 13852 18938 13864
rect 19886 13852 19892 13864
rect 18932 13824 18977 13852
rect 19306 13824 19748 13852
rect 19847 13824 19892 13852
rect 18932 13812 18938 13824
rect 18049 13787 18107 13793
rect 18049 13753 18061 13787
rect 18095 13784 18107 13787
rect 18892 13784 18920 13812
rect 18095 13756 18920 13784
rect 18095 13753 18107 13756
rect 18049 13747 18107 13753
rect 17402 13716 17408 13728
rect 16684 13688 17408 13716
rect 17402 13676 17408 13688
rect 17460 13676 17466 13728
rect 17770 13676 17776 13728
rect 17828 13716 17834 13728
rect 19306 13716 19334 13824
rect 19720 13784 19748 13824
rect 19886 13812 19892 13824
rect 19944 13812 19950 13864
rect 20809 13855 20867 13861
rect 20809 13852 20821 13855
rect 19996 13824 20821 13852
rect 19996 13784 20024 13824
rect 20809 13821 20821 13824
rect 20855 13821 20867 13855
rect 20990 13852 20996 13864
rect 20951 13824 20996 13852
rect 20809 13815 20867 13821
rect 20990 13812 20996 13824
rect 21048 13812 21054 13864
rect 19720 13756 20024 13784
rect 17828 13688 19334 13716
rect 17828 13676 17834 13688
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 5442 13472 5448 13524
rect 5500 13512 5506 13524
rect 7745 13515 7803 13521
rect 7745 13512 7757 13515
rect 5500 13484 7757 13512
rect 5500 13472 5506 13484
rect 7745 13481 7757 13484
rect 7791 13512 7803 13515
rect 9674 13512 9680 13524
rect 7791 13484 9680 13512
rect 7791 13481 7803 13484
rect 7745 13475 7803 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 10870 13512 10876 13524
rect 10831 13484 10876 13512
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12492 13484 12537 13512
rect 12492 13472 12498 13484
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 17954 13512 17960 13524
rect 12768 13484 17960 13512
rect 12768 13472 12774 13484
rect 17954 13472 17960 13484
rect 18012 13472 18018 13524
rect 20714 13472 20720 13524
rect 20772 13512 20778 13524
rect 21269 13515 21327 13521
rect 21269 13512 21281 13515
rect 20772 13484 21281 13512
rect 20772 13472 20778 13484
rect 21269 13481 21281 13484
rect 21315 13481 21327 13515
rect 21269 13475 21327 13481
rect 5166 13404 5172 13456
rect 5224 13444 5230 13456
rect 9769 13447 9827 13453
rect 5224 13416 9536 13444
rect 5224 13404 5230 13416
rect 8113 13379 8171 13385
rect 8113 13345 8125 13379
rect 8159 13376 8171 13379
rect 8202 13376 8208 13388
rect 8159 13348 8208 13376
rect 8159 13345 8171 13348
rect 8113 13339 8171 13345
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 9214 13376 9220 13388
rect 9175 13348 9220 13376
rect 9214 13336 9220 13348
rect 9272 13336 9278 13388
rect 9508 13376 9536 13416
rect 9769 13413 9781 13447
rect 9815 13444 9827 13447
rect 10778 13444 10784 13456
rect 9815 13416 10784 13444
rect 9815 13413 9827 13416
rect 9769 13407 9827 13413
rect 10778 13404 10784 13416
rect 10836 13404 10842 13456
rect 11790 13404 11796 13456
rect 11848 13444 11854 13456
rect 13449 13447 13507 13453
rect 13449 13444 13461 13447
rect 11848 13416 13461 13444
rect 11848 13404 11854 13416
rect 13449 13413 13461 13416
rect 13495 13413 13507 13447
rect 13449 13407 13507 13413
rect 14274 13404 14280 13456
rect 14332 13444 14338 13456
rect 15289 13447 15347 13453
rect 14332 13416 14964 13444
rect 14332 13404 14338 13416
rect 12894 13376 12900 13388
rect 9508 13348 12900 13376
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 12986 13336 12992 13388
rect 13044 13376 13050 13388
rect 14642 13376 14648 13388
rect 13044 13348 13089 13376
rect 14603 13348 14648 13376
rect 13044 13336 13050 13348
rect 14642 13336 14648 13348
rect 14700 13336 14706 13388
rect 14826 13376 14832 13388
rect 14787 13348 14832 13376
rect 14826 13336 14832 13348
rect 14884 13336 14890 13388
rect 14936 13376 14964 13416
rect 15289 13413 15301 13447
rect 15335 13444 15347 13447
rect 18046 13444 18052 13456
rect 15335 13416 18052 13444
rect 15335 13413 15347 13416
rect 15289 13407 15347 13413
rect 18046 13404 18052 13416
rect 18104 13404 18110 13456
rect 18785 13447 18843 13453
rect 18785 13413 18797 13447
rect 18831 13444 18843 13447
rect 21082 13444 21088 13456
rect 18831 13416 21088 13444
rect 18831 13413 18843 13416
rect 18785 13407 18843 13413
rect 21082 13404 21088 13416
rect 21140 13404 21146 13456
rect 14936 13348 17816 13376
rect 2314 13268 2320 13320
rect 2372 13308 2378 13320
rect 5442 13308 5448 13320
rect 2372 13280 5448 13308
rect 2372 13268 2378 13280
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 8570 13308 8576 13320
rect 8531 13280 8576 13308
rect 8570 13268 8576 13280
rect 8628 13268 8634 13320
rect 9398 13308 9404 13320
rect 9359 13280 9404 13308
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 12158 13308 12164 13320
rect 12071 13280 12164 13308
rect 12158 13268 12164 13280
rect 12216 13308 12222 13320
rect 13630 13308 13636 13320
rect 12216 13280 13492 13308
rect 13591 13280 13636 13308
rect 12216 13268 12222 13280
rect 6914 13200 6920 13252
rect 6972 13240 6978 13252
rect 9309 13243 9367 13249
rect 6972 13212 8524 13240
rect 6972 13200 6978 13212
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 7285 13175 7343 13181
rect 7285 13172 7297 13175
rect 7248 13144 7297 13172
rect 7248 13132 7254 13144
rect 7285 13141 7297 13144
rect 7331 13141 7343 13175
rect 7285 13135 7343 13141
rect 8202 13132 8208 13184
rect 8260 13172 8266 13184
rect 8389 13175 8447 13181
rect 8389 13172 8401 13175
rect 8260 13144 8401 13172
rect 8260 13132 8266 13144
rect 8389 13141 8401 13144
rect 8435 13141 8447 13175
rect 8496 13172 8524 13212
rect 9309 13209 9321 13243
rect 9355 13240 9367 13243
rect 11238 13240 11244 13252
rect 9355 13212 11244 13240
rect 9355 13209 9367 13212
rect 9309 13203 9367 13209
rect 11238 13200 11244 13212
rect 11296 13200 11302 13252
rect 13464 13240 13492 13280
rect 13630 13268 13636 13280
rect 13688 13268 13694 13320
rect 14277 13311 14335 13317
rect 14277 13277 14289 13311
rect 14323 13308 14335 13311
rect 14550 13308 14556 13320
rect 14323 13280 14556 13308
rect 14323 13277 14335 13280
rect 14277 13271 14335 13277
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 14921 13311 14979 13317
rect 14921 13277 14933 13311
rect 14967 13308 14979 13311
rect 15010 13308 15016 13320
rect 14967 13280 15016 13308
rect 14967 13277 14979 13280
rect 14921 13271 14979 13277
rect 15010 13268 15016 13280
rect 15068 13268 15074 13320
rect 16298 13268 16304 13320
rect 16356 13308 16362 13320
rect 17681 13311 17739 13317
rect 17681 13308 17693 13311
rect 16356 13280 17693 13308
rect 16356 13268 16362 13280
rect 17681 13277 17693 13280
rect 17727 13277 17739 13311
rect 17681 13271 17739 13277
rect 15654 13240 15660 13252
rect 13464 13212 15660 13240
rect 15654 13200 15660 13212
rect 15712 13200 15718 13252
rect 17402 13240 17408 13252
rect 17363 13212 17408 13240
rect 17402 13200 17408 13212
rect 17460 13200 17466 13252
rect 17788 13240 17816 13348
rect 18690 13336 18696 13388
rect 18748 13376 18754 13388
rect 19886 13376 19892 13388
rect 18748 13348 19892 13376
rect 18748 13336 18754 13348
rect 19886 13336 19892 13348
rect 19944 13336 19950 13388
rect 20441 13379 20499 13385
rect 20441 13345 20453 13379
rect 20487 13376 20499 13379
rect 20714 13376 20720 13388
rect 20487 13348 20720 13376
rect 20487 13345 20499 13348
rect 20441 13339 20499 13345
rect 20714 13336 20720 13348
rect 20772 13336 20778 13388
rect 18598 13308 18604 13320
rect 18559 13280 18604 13308
rect 18598 13268 18604 13280
rect 18656 13268 18662 13320
rect 19058 13268 19064 13320
rect 19116 13308 19122 13320
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19116 13280 19717 13308
rect 19116 13268 19122 13280
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 20530 13308 20536 13320
rect 20491 13280 20536 13308
rect 19705 13271 19763 13277
rect 20530 13268 20536 13280
rect 20588 13308 20594 13320
rect 21450 13308 21456 13320
rect 20588 13280 21456 13308
rect 20588 13268 20594 13280
rect 21450 13268 21456 13280
rect 21508 13268 21514 13320
rect 19613 13243 19671 13249
rect 19613 13240 19625 13243
rect 17788 13212 19625 13240
rect 19613 13209 19625 13212
rect 19659 13209 19671 13243
rect 19613 13203 19671 13209
rect 10137 13175 10195 13181
rect 10137 13172 10149 13175
rect 8496 13144 10149 13172
rect 8389 13135 8447 13141
rect 10137 13141 10149 13144
rect 10183 13172 10195 13175
rect 12342 13172 12348 13184
rect 10183 13144 12348 13172
rect 10183 13141 10195 13144
rect 10137 13135 10195 13141
rect 12342 13132 12348 13144
rect 12400 13132 12406 13184
rect 12802 13172 12808 13184
rect 12763 13144 12808 13172
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 14093 13175 14151 13181
rect 14093 13141 14105 13175
rect 14139 13172 14151 13175
rect 14458 13172 14464 13184
rect 14139 13144 14464 13172
rect 14139 13141 14151 13144
rect 14093 13135 14151 13141
rect 14458 13132 14464 13144
rect 14516 13132 14522 13184
rect 14642 13132 14648 13184
rect 14700 13172 14706 13184
rect 14918 13172 14924 13184
rect 14700 13144 14924 13172
rect 14700 13132 14706 13144
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 15930 13132 15936 13184
rect 15988 13172 15994 13184
rect 18325 13175 18383 13181
rect 18325 13172 18337 13175
rect 15988 13144 18337 13172
rect 15988 13132 15994 13144
rect 18325 13141 18337 13144
rect 18371 13141 18383 13175
rect 18325 13135 18383 13141
rect 18874 13132 18880 13184
rect 18932 13172 18938 13184
rect 19245 13175 19303 13181
rect 19245 13172 19257 13175
rect 18932 13144 19257 13172
rect 18932 13132 18938 13144
rect 19245 13141 19257 13144
rect 19291 13141 19303 13175
rect 19245 13135 19303 13141
rect 19978 13132 19984 13184
rect 20036 13172 20042 13184
rect 20254 13172 20260 13184
rect 20036 13144 20260 13172
rect 20036 13132 20042 13144
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 20622 13132 20628 13184
rect 20680 13172 20686 13184
rect 20990 13172 20996 13184
rect 20680 13144 20725 13172
rect 20951 13144 20996 13172
rect 20680 13132 20686 13144
rect 20990 13132 20996 13144
rect 21048 13132 21054 13184
rect 1104 13082 21896 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21896 13082
rect 1104 13008 21896 13030
rect 7466 12928 7472 12980
rect 7524 12968 7530 12980
rect 8021 12971 8079 12977
rect 8021 12968 8033 12971
rect 7524 12940 8033 12968
rect 7524 12928 7530 12940
rect 8021 12937 8033 12940
rect 8067 12968 8079 12971
rect 8110 12968 8116 12980
rect 8067 12940 8116 12968
rect 8067 12937 8079 12940
rect 8021 12931 8079 12937
rect 8110 12928 8116 12940
rect 8168 12928 8174 12980
rect 8573 12971 8631 12977
rect 8573 12937 8585 12971
rect 8619 12968 8631 12971
rect 9398 12968 9404 12980
rect 8619 12940 9404 12968
rect 8619 12937 8631 12940
rect 8573 12931 8631 12937
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 10318 12968 10324 12980
rect 10279 12940 10324 12968
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 10965 12971 11023 12977
rect 10965 12937 10977 12971
rect 11011 12968 11023 12971
rect 12802 12968 12808 12980
rect 11011 12940 12808 12968
rect 11011 12937 11023 12940
rect 10965 12931 11023 12937
rect 12802 12928 12808 12940
rect 12860 12928 12866 12980
rect 14550 12968 14556 12980
rect 14511 12940 14556 12968
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 15194 12928 15200 12980
rect 15252 12928 15258 12980
rect 15470 12928 15476 12980
rect 15528 12968 15534 12980
rect 15565 12971 15623 12977
rect 15565 12968 15577 12971
rect 15528 12940 15577 12968
rect 15528 12928 15534 12940
rect 15565 12937 15577 12940
rect 15611 12937 15623 12971
rect 15565 12931 15623 12937
rect 15746 12928 15752 12980
rect 15804 12968 15810 12980
rect 15933 12971 15991 12977
rect 15933 12968 15945 12971
rect 15804 12940 15945 12968
rect 15804 12928 15810 12940
rect 15933 12937 15945 12940
rect 15979 12937 15991 12971
rect 15933 12931 15991 12937
rect 18601 12971 18659 12977
rect 18601 12937 18613 12971
rect 18647 12968 18659 12971
rect 18690 12968 18696 12980
rect 18647 12940 18696 12968
rect 18647 12937 18659 12940
rect 18601 12931 18659 12937
rect 18690 12928 18696 12940
rect 18748 12928 18754 12980
rect 20254 12968 20260 12980
rect 20215 12940 20260 12968
rect 20254 12928 20260 12940
rect 20312 12928 20318 12980
rect 20625 12971 20683 12977
rect 20625 12937 20637 12971
rect 20671 12968 20683 12971
rect 20990 12968 20996 12980
rect 20671 12940 20996 12968
rect 20671 12937 20683 12940
rect 20625 12931 20683 12937
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 21361 12971 21419 12977
rect 21361 12937 21373 12971
rect 21407 12968 21419 12971
rect 21542 12968 21548 12980
rect 21407 12940 21548 12968
rect 21407 12937 21419 12940
rect 21361 12931 21419 12937
rect 21542 12928 21548 12940
rect 21600 12928 21606 12980
rect 4982 12860 4988 12912
rect 5040 12900 5046 12912
rect 10410 12900 10416 12912
rect 5040 12872 10416 12900
rect 5040 12860 5046 12872
rect 10410 12860 10416 12872
rect 10468 12900 10474 12912
rect 12526 12900 12532 12912
rect 10468 12872 12532 12900
rect 10468 12860 10474 12872
rect 12526 12860 12532 12872
rect 12584 12860 12590 12912
rect 12618 12860 12624 12912
rect 12676 12900 12682 12912
rect 14001 12903 14059 12909
rect 14001 12900 14013 12903
rect 12676 12872 14013 12900
rect 12676 12860 12682 12872
rect 14001 12869 14013 12872
rect 14047 12869 14059 12903
rect 14001 12863 14059 12869
rect 14921 12903 14979 12909
rect 14921 12869 14933 12903
rect 14967 12900 14979 12903
rect 15102 12900 15108 12912
rect 14967 12872 15108 12900
rect 14967 12869 14979 12872
rect 14921 12863 14979 12869
rect 15102 12860 15108 12872
rect 15160 12860 15166 12912
rect 15212 12900 15240 12928
rect 16025 12903 16083 12909
rect 16025 12900 16037 12903
rect 15212 12872 16037 12900
rect 16025 12869 16037 12872
rect 16071 12869 16083 12903
rect 16025 12863 16083 12869
rect 17402 12860 17408 12912
rect 17460 12900 17466 12912
rect 19518 12900 19524 12912
rect 17460 12872 19524 12900
rect 17460 12860 17466 12872
rect 7742 12792 7748 12844
rect 7800 12792 7806 12844
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 8904 12804 8953 12832
rect 8904 12792 8910 12804
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 9197 12835 9255 12841
rect 9197 12832 9209 12835
rect 8941 12795 8999 12801
rect 9048 12804 9209 12832
rect 7760 12764 7788 12792
rect 9048 12764 9076 12804
rect 9197 12801 9209 12804
rect 9243 12801 9255 12835
rect 9197 12795 9255 12801
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 11793 12835 11851 12841
rect 11793 12832 11805 12835
rect 10284 12804 11805 12832
rect 10284 12792 10290 12804
rect 11793 12801 11805 12804
rect 11839 12801 11851 12835
rect 11793 12795 11851 12801
rect 12342 12792 12348 12844
rect 12400 12832 12406 12844
rect 12713 12835 12771 12841
rect 12713 12832 12725 12835
rect 12400 12804 12725 12832
rect 12400 12792 12406 12804
rect 12713 12801 12725 12804
rect 12759 12832 12771 12835
rect 12759 12804 13308 12832
rect 12759 12801 12771 12804
rect 12713 12795 12771 12801
rect 7760 12736 9076 12764
rect 12066 12724 12072 12776
rect 12124 12764 12130 12776
rect 12805 12767 12863 12773
rect 12805 12764 12817 12767
rect 12124 12736 12817 12764
rect 12124 12724 12130 12736
rect 12805 12733 12817 12736
rect 12851 12733 12863 12767
rect 12986 12764 12992 12776
rect 12947 12736 12992 12764
rect 12805 12727 12863 12733
rect 12986 12724 12992 12736
rect 13044 12724 13050 12776
rect 11974 12656 11980 12708
rect 12032 12696 12038 12708
rect 12345 12699 12403 12705
rect 12345 12696 12357 12699
rect 12032 12668 12357 12696
rect 12032 12656 12038 12668
rect 12345 12665 12357 12668
rect 12391 12665 12403 12699
rect 13280 12696 13308 12804
rect 13354 12792 13360 12844
rect 13412 12832 13418 12844
rect 16942 12832 16948 12844
rect 13412 12804 13457 12832
rect 15580 12804 16948 12832
rect 13412 12792 13418 12804
rect 13538 12724 13544 12776
rect 13596 12764 13602 12776
rect 14734 12764 14740 12776
rect 13596 12736 14740 12764
rect 13596 12724 13602 12736
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 15010 12764 15016 12776
rect 14971 12736 15016 12764
rect 15010 12724 15016 12736
rect 15068 12724 15074 12776
rect 15105 12767 15163 12773
rect 15105 12733 15117 12767
rect 15151 12764 15163 12767
rect 15580 12764 15608 12804
rect 16942 12792 16948 12804
rect 17000 12792 17006 12844
rect 18064 12841 18092 12872
rect 19518 12860 19524 12872
rect 19576 12900 19582 12912
rect 19576 12872 20024 12900
rect 19576 12860 19582 12872
rect 17793 12835 17851 12841
rect 17793 12801 17805 12835
rect 17839 12832 17851 12835
rect 18049 12835 18107 12841
rect 17839 12804 18000 12832
rect 17839 12801 17851 12804
rect 17793 12795 17851 12801
rect 16206 12764 16212 12776
rect 15151 12736 15608 12764
rect 16167 12736 16212 12764
rect 15151 12733 15163 12736
rect 15105 12727 15163 12733
rect 14550 12696 14556 12708
rect 13280 12668 14556 12696
rect 12345 12659 12403 12665
rect 14550 12656 14556 12668
rect 14608 12656 14614 12708
rect 14826 12656 14832 12708
rect 14884 12696 14890 12708
rect 15120 12696 15148 12727
rect 16206 12724 16212 12736
rect 16264 12724 16270 12776
rect 17972 12764 18000 12804
rect 18049 12801 18061 12835
rect 18095 12801 18107 12835
rect 18049 12795 18107 12801
rect 19702 12792 19708 12844
rect 19760 12841 19766 12844
rect 19996 12841 20024 12872
rect 19760 12832 19772 12841
rect 19981 12835 20039 12841
rect 19760 12804 19805 12832
rect 19760 12795 19772 12804
rect 19981 12801 19993 12835
rect 20027 12801 20039 12835
rect 19981 12795 20039 12801
rect 19760 12792 19766 12795
rect 18782 12764 18788 12776
rect 16316 12736 17080 12764
rect 17972 12736 18788 12764
rect 14884 12668 15148 12696
rect 14884 12656 14890 12668
rect 8110 12588 8116 12640
rect 8168 12628 8174 12640
rect 11609 12631 11667 12637
rect 11609 12628 11621 12631
rect 8168 12600 11621 12628
rect 8168 12588 8174 12600
rect 11609 12597 11621 12600
rect 11655 12597 11667 12631
rect 11609 12591 11667 12597
rect 11698 12588 11704 12640
rect 11756 12628 11762 12640
rect 13354 12628 13360 12640
rect 11756 12600 13360 12628
rect 11756 12588 11762 12600
rect 13354 12588 13360 12600
rect 13412 12588 13418 12640
rect 13814 12588 13820 12640
rect 13872 12628 13878 12640
rect 16316 12628 16344 12736
rect 16666 12628 16672 12640
rect 13872 12600 16344 12628
rect 16627 12600 16672 12628
rect 13872 12588 13878 12600
rect 16666 12588 16672 12600
rect 16724 12588 16730 12640
rect 17052 12628 17080 12736
rect 18782 12724 18788 12736
rect 18840 12724 18846 12776
rect 20530 12724 20536 12776
rect 20588 12764 20594 12776
rect 20717 12767 20775 12773
rect 20717 12764 20729 12767
rect 20588 12736 20729 12764
rect 20588 12724 20594 12736
rect 20717 12733 20729 12736
rect 20763 12733 20775 12767
rect 20898 12764 20904 12776
rect 20859 12736 20904 12764
rect 20717 12727 20775 12733
rect 20898 12724 20904 12736
rect 20956 12724 20962 12776
rect 18506 12656 18512 12708
rect 18564 12696 18570 12708
rect 18690 12696 18696 12708
rect 18564 12668 18696 12696
rect 18564 12656 18570 12668
rect 18690 12656 18696 12668
rect 18748 12656 18754 12708
rect 20622 12628 20628 12640
rect 17052 12600 20628 12628
rect 20622 12588 20628 12600
rect 20680 12588 20686 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 8941 12427 8999 12433
rect 8941 12393 8953 12427
rect 8987 12424 8999 12427
rect 9214 12424 9220 12436
rect 8987 12396 9220 12424
rect 8987 12393 8999 12396
rect 8941 12387 8999 12393
rect 7650 12356 7656 12368
rect 7611 12328 7656 12356
rect 7650 12316 7656 12328
rect 7708 12316 7714 12368
rect 8754 12316 8760 12368
rect 8812 12356 8818 12368
rect 8956 12356 8984 12387
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 10597 12427 10655 12433
rect 10597 12424 10609 12427
rect 9324 12396 10609 12424
rect 8812 12328 8984 12356
rect 8812 12316 8818 12328
rect 8386 12248 8392 12300
rect 8444 12288 8450 12300
rect 9324 12288 9352 12396
rect 10597 12393 10609 12396
rect 10643 12393 10655 12427
rect 12066 12424 12072 12436
rect 12027 12396 12072 12424
rect 10597 12387 10655 12393
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 15102 12384 15108 12436
rect 15160 12424 15166 12436
rect 15749 12427 15807 12433
rect 15749 12424 15761 12427
rect 15160 12396 15761 12424
rect 15160 12384 15166 12396
rect 15749 12393 15761 12396
rect 15795 12393 15807 12427
rect 17678 12424 17684 12436
rect 17639 12396 17684 12424
rect 15749 12387 15807 12393
rect 17678 12384 17684 12396
rect 17736 12384 17742 12436
rect 18598 12384 18604 12436
rect 18656 12424 18662 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 18656 12396 19257 12424
rect 18656 12384 18662 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 19245 12387 19303 12393
rect 20898 12384 20904 12436
rect 20956 12424 20962 12436
rect 21177 12427 21235 12433
rect 21177 12424 21189 12427
rect 20956 12396 21189 12424
rect 20956 12384 20962 12396
rect 21177 12393 21189 12396
rect 21223 12393 21235 12427
rect 21177 12387 21235 12393
rect 13725 12359 13783 12365
rect 13725 12325 13737 12359
rect 13771 12325 13783 12359
rect 13725 12319 13783 12325
rect 8444 12260 9352 12288
rect 10321 12291 10379 12297
rect 8444 12248 8450 12260
rect 10321 12257 10333 12291
rect 10367 12288 10379 12291
rect 10870 12288 10876 12300
rect 10367 12260 10876 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 7469 12223 7527 12229
rect 7469 12189 7481 12223
rect 7515 12220 7527 12223
rect 8110 12220 8116 12232
rect 7515 12192 8116 12220
rect 7515 12189 7527 12192
rect 7469 12183 7527 12189
rect 8110 12180 8116 12192
rect 8168 12180 8174 12232
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12220 8631 12223
rect 8938 12220 8944 12232
rect 8619 12192 8944 12220
rect 8619 12189 8631 12192
rect 8573 12183 8631 12189
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 9030 12180 9036 12232
rect 9088 12220 9094 12232
rect 10336 12220 10364 12251
rect 10870 12248 10876 12260
rect 10928 12248 10934 12300
rect 11517 12291 11575 12297
rect 11517 12257 11529 12291
rect 11563 12288 11575 12291
rect 11698 12288 11704 12300
rect 11563 12260 11704 12288
rect 11563 12257 11575 12260
rect 11517 12251 11575 12257
rect 11698 12248 11704 12260
rect 11756 12248 11762 12300
rect 10778 12220 10784 12232
rect 9088 12192 10364 12220
rect 10739 12192 10784 12220
rect 9088 12180 9094 12192
rect 10778 12180 10784 12192
rect 10836 12180 10842 12232
rect 10888 12220 10916 12248
rect 11790 12220 11796 12232
rect 10888 12192 11796 12220
rect 11790 12180 11796 12192
rect 11848 12220 11854 12232
rect 12345 12223 12403 12229
rect 12345 12220 12357 12223
rect 11848 12192 12357 12220
rect 11848 12180 11854 12192
rect 12345 12189 12357 12192
rect 12391 12189 12403 12223
rect 13740 12220 13768 12319
rect 15470 12316 15476 12368
rect 15528 12356 15534 12368
rect 17770 12356 17776 12368
rect 15528 12328 17776 12356
rect 15528 12316 15534 12328
rect 17770 12316 17776 12328
rect 17828 12316 17834 12368
rect 16298 12288 16304 12300
rect 15396 12260 16304 12288
rect 15194 12220 15200 12232
rect 15252 12229 15258 12232
rect 13740 12192 15200 12220
rect 12345 12183 12403 12189
rect 15194 12180 15200 12192
rect 15252 12183 15264 12229
rect 15252 12180 15258 12183
rect 9858 12112 9864 12164
rect 9916 12152 9922 12164
rect 10054 12155 10112 12161
rect 10054 12152 10066 12155
rect 9916 12124 10066 12152
rect 9916 12112 9922 12124
rect 10054 12121 10066 12124
rect 10100 12121 10112 12155
rect 11606 12152 11612 12164
rect 11519 12124 11612 12152
rect 10054 12115 10112 12121
rect 11606 12112 11612 12124
rect 11664 12152 11670 12164
rect 12158 12152 12164 12164
rect 11664 12124 12164 12152
rect 11664 12112 11670 12124
rect 12158 12112 12164 12124
rect 12216 12112 12222 12164
rect 12434 12112 12440 12164
rect 12492 12152 12498 12164
rect 12590 12155 12648 12161
rect 12590 12152 12602 12155
rect 12492 12124 12602 12152
rect 12492 12112 12498 12124
rect 12590 12121 12602 12124
rect 12636 12121 12648 12155
rect 14274 12152 14280 12164
rect 12590 12115 12648 12121
rect 13372 12124 14280 12152
rect 7929 12087 7987 12093
rect 7929 12053 7941 12087
rect 7975 12084 7987 12087
rect 10502 12084 10508 12096
rect 7975 12056 10508 12084
rect 7975 12053 7987 12056
rect 7929 12047 7987 12053
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 11146 12044 11152 12096
rect 11204 12084 11210 12096
rect 11701 12087 11759 12093
rect 11701 12084 11713 12087
rect 11204 12056 11713 12084
rect 11204 12044 11210 12056
rect 11701 12053 11713 12056
rect 11747 12084 11759 12087
rect 13372 12084 13400 12124
rect 14274 12112 14280 12124
rect 14332 12112 14338 12164
rect 11747 12056 13400 12084
rect 11747 12053 11759 12056
rect 11701 12047 11759 12053
rect 13906 12044 13912 12096
rect 13964 12084 13970 12096
rect 14093 12087 14151 12093
rect 14093 12084 14105 12087
rect 13964 12056 14105 12084
rect 13964 12044 13970 12056
rect 14093 12053 14105 12056
rect 14139 12084 14151 12087
rect 15396 12084 15424 12260
rect 16298 12248 16304 12260
rect 16356 12248 16362 12300
rect 16666 12248 16672 12300
rect 16724 12288 16730 12300
rect 17129 12291 17187 12297
rect 17129 12288 17141 12291
rect 16724 12260 17141 12288
rect 16724 12248 16730 12260
rect 17129 12257 17141 12260
rect 17175 12288 17187 12291
rect 17218 12288 17224 12300
rect 17175 12260 17224 12288
rect 17175 12257 17187 12260
rect 17129 12251 17187 12257
rect 17218 12248 17224 12260
rect 17276 12288 17282 12300
rect 17678 12288 17684 12300
rect 17276 12260 17684 12288
rect 17276 12248 17282 12260
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 18601 12291 18659 12297
rect 18601 12257 18613 12291
rect 18647 12288 18659 12291
rect 18782 12288 18788 12300
rect 18647 12260 18788 12288
rect 18647 12257 18659 12260
rect 18601 12251 18659 12257
rect 18782 12248 18788 12260
rect 18840 12248 18846 12300
rect 19518 12248 19524 12300
rect 19576 12288 19582 12300
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 19576 12260 19809 12288
rect 19576 12248 19582 12260
rect 19797 12257 19809 12260
rect 19843 12257 19855 12291
rect 19797 12251 19855 12257
rect 15473 12223 15531 12229
rect 15473 12189 15485 12223
rect 15519 12220 15531 12223
rect 17402 12220 17408 12232
rect 15519 12192 17408 12220
rect 15519 12189 15531 12192
rect 15473 12183 15531 12189
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 18230 12180 18236 12232
rect 18288 12220 18294 12232
rect 18325 12223 18383 12229
rect 18325 12220 18337 12223
rect 18288 12192 18337 12220
rect 18288 12180 18294 12192
rect 18325 12189 18337 12192
rect 18371 12189 18383 12223
rect 18325 12183 18383 12189
rect 19429 12223 19487 12229
rect 19429 12189 19441 12223
rect 19475 12220 19487 12223
rect 19702 12220 19708 12232
rect 19475 12192 19708 12220
rect 19475 12189 19487 12192
rect 19429 12183 19487 12189
rect 19702 12180 19708 12192
rect 19760 12180 19766 12232
rect 16114 12152 16120 12164
rect 16075 12124 16120 12152
rect 16114 12112 16120 12124
rect 16172 12112 16178 12164
rect 17221 12155 17279 12161
rect 17221 12121 17233 12155
rect 17267 12152 17279 12155
rect 20064 12155 20122 12161
rect 17267 12124 18000 12152
rect 17267 12121 17279 12124
rect 17221 12115 17279 12121
rect 16206 12084 16212 12096
rect 14139 12056 15424 12084
rect 16167 12056 16212 12084
rect 14139 12053 14151 12056
rect 14093 12047 14151 12053
rect 16206 12044 16212 12056
rect 16264 12044 16270 12096
rect 17313 12087 17371 12093
rect 17313 12053 17325 12087
rect 17359 12084 17371 12087
rect 17862 12084 17868 12096
rect 17359 12056 17868 12084
rect 17359 12053 17371 12056
rect 17313 12047 17371 12053
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 17972 12093 18000 12124
rect 20064 12121 20076 12155
rect 20110 12152 20122 12155
rect 20714 12152 20720 12164
rect 20110 12124 20720 12152
rect 20110 12121 20122 12124
rect 20064 12115 20122 12121
rect 20714 12112 20720 12124
rect 20772 12112 20778 12164
rect 17957 12087 18015 12093
rect 17957 12053 17969 12087
rect 18003 12053 18015 12087
rect 17957 12047 18015 12053
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 18417 12087 18475 12093
rect 18417 12084 18429 12087
rect 18196 12056 18429 12084
rect 18196 12044 18202 12056
rect 18417 12053 18429 12056
rect 18463 12084 18475 12087
rect 18506 12084 18512 12096
rect 18463 12056 18512 12084
rect 18463 12053 18475 12056
rect 18417 12047 18475 12053
rect 18506 12044 18512 12056
rect 18564 12044 18570 12096
rect 19886 12044 19892 12096
rect 19944 12084 19950 12096
rect 20438 12084 20444 12096
rect 19944 12056 20444 12084
rect 19944 12044 19950 12056
rect 20438 12044 20444 12056
rect 20496 12044 20502 12096
rect 1104 11994 21896 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21896 11994
rect 1104 11920 21896 11942
rect 4890 11840 4896 11892
rect 4948 11880 4954 11892
rect 6914 11880 6920 11892
rect 4948 11852 6920 11880
rect 4948 11840 4954 11852
rect 6914 11840 6920 11852
rect 6972 11880 6978 11892
rect 7190 11880 7196 11892
rect 6972 11852 7196 11880
rect 6972 11840 6978 11852
rect 7190 11840 7196 11852
rect 7248 11840 7254 11892
rect 7837 11883 7895 11889
rect 7837 11849 7849 11883
rect 7883 11880 7895 11883
rect 8478 11880 8484 11892
rect 7883 11852 8484 11880
rect 7883 11849 7895 11852
rect 7837 11843 7895 11849
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 8938 11840 8944 11892
rect 8996 11880 9002 11892
rect 9674 11880 9680 11892
rect 8996 11852 9680 11880
rect 8996 11840 9002 11852
rect 9674 11840 9680 11852
rect 9732 11880 9738 11892
rect 10413 11883 10471 11889
rect 10413 11880 10425 11883
rect 9732 11852 10425 11880
rect 9732 11840 9738 11852
rect 10413 11849 10425 11852
rect 10459 11849 10471 11883
rect 11790 11880 11796 11892
rect 10413 11843 10471 11849
rect 11716 11852 11796 11880
rect 8113 11815 8171 11821
rect 8113 11781 8125 11815
rect 8159 11812 8171 11815
rect 9278 11815 9336 11821
rect 9278 11812 9290 11815
rect 8159 11784 9290 11812
rect 8159 11781 8171 11784
rect 8113 11775 8171 11781
rect 9278 11781 9290 11784
rect 9324 11781 9336 11815
rect 9278 11775 9336 11781
rect 9490 11772 9496 11824
rect 9548 11812 9554 11824
rect 11146 11812 11152 11824
rect 9548 11784 11152 11812
rect 9548 11772 9554 11784
rect 11146 11772 11152 11784
rect 11204 11772 11210 11824
rect 7653 11747 7711 11753
rect 7653 11713 7665 11747
rect 7699 11744 7711 11747
rect 8018 11744 8024 11756
rect 7699 11716 8024 11744
rect 7699 11713 7711 11716
rect 7653 11707 7711 11713
rect 8018 11704 8024 11716
rect 8076 11704 8082 11756
rect 8754 11744 8760 11756
rect 8715 11716 8760 11744
rect 8754 11704 8760 11716
rect 8812 11704 8818 11756
rect 9030 11744 9036 11756
rect 8991 11716 9036 11744
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 11716 11753 11744 11852
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 13814 11880 13820 11892
rect 13775 11852 13820 11880
rect 13814 11840 13820 11852
rect 13872 11840 13878 11892
rect 18046 11880 18052 11892
rect 16224 11852 18052 11880
rect 14734 11812 14740 11824
rect 11808 11784 14740 11812
rect 11701 11747 11759 11753
rect 9140 11716 11100 11744
rect 6546 11636 6552 11688
rect 6604 11676 6610 11688
rect 9140 11676 9168 11716
rect 6604 11648 9168 11676
rect 6604 11636 6610 11648
rect 10042 11636 10048 11688
rect 10100 11676 10106 11688
rect 10965 11679 11023 11685
rect 10965 11676 10977 11679
rect 10100 11648 10977 11676
rect 10100 11636 10106 11648
rect 10965 11645 10977 11648
rect 11011 11645 11023 11679
rect 11072 11676 11100 11716
rect 11701 11713 11713 11747
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 11808 11676 11836 11784
rect 14734 11772 14740 11784
rect 14792 11772 14798 11824
rect 15838 11812 15844 11824
rect 15799 11784 15844 11812
rect 15838 11772 15844 11784
rect 15896 11772 15902 11824
rect 16224 11812 16252 11852
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 18322 11880 18328 11892
rect 18283 11852 18328 11880
rect 18322 11840 18328 11852
rect 18380 11840 18386 11892
rect 18785 11883 18843 11889
rect 18785 11849 18797 11883
rect 18831 11880 18843 11883
rect 18874 11880 18880 11892
rect 18831 11852 18880 11880
rect 18831 11849 18843 11852
rect 18785 11843 18843 11849
rect 18874 11840 18880 11852
rect 18932 11840 18938 11892
rect 19705 11883 19763 11889
rect 19705 11849 19717 11883
rect 19751 11880 19763 11883
rect 20349 11883 20407 11889
rect 20349 11880 20361 11883
rect 19751 11852 20361 11880
rect 19751 11849 19763 11852
rect 19705 11843 19763 11849
rect 20349 11849 20361 11852
rect 20395 11849 20407 11883
rect 20349 11843 20407 11849
rect 16132 11784 16252 11812
rect 16936 11815 16994 11821
rect 11974 11753 11980 11756
rect 11968 11707 11980 11753
rect 12032 11744 12038 11756
rect 16132 11753 16160 11784
rect 16936 11781 16948 11815
rect 16982 11812 16994 11815
rect 17310 11812 17316 11824
rect 16982 11784 17316 11812
rect 16982 11781 16994 11784
rect 16936 11775 16994 11781
rect 17310 11772 17316 11784
rect 17368 11772 17374 11824
rect 18693 11815 18751 11821
rect 18693 11781 18705 11815
rect 18739 11812 18751 11815
rect 19610 11812 19616 11824
rect 18739 11784 19616 11812
rect 18739 11781 18751 11784
rect 18693 11775 18751 11781
rect 19610 11772 19616 11784
rect 19668 11772 19674 11824
rect 20809 11815 20867 11821
rect 20809 11812 20821 11815
rect 20088 11784 20821 11812
rect 16117 11747 16175 11753
rect 12032 11716 12068 11744
rect 11974 11704 11980 11707
rect 12032 11704 12038 11716
rect 16117 11713 16129 11747
rect 16163 11713 16175 11747
rect 18598 11744 18604 11756
rect 16117 11707 16175 11713
rect 16224 11716 18604 11744
rect 11072 11648 11836 11676
rect 10965 11639 11023 11645
rect 15102 11636 15108 11688
rect 15160 11676 15166 11688
rect 16224 11676 16252 11716
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 18966 11704 18972 11756
rect 19024 11744 19030 11756
rect 20088 11744 20116 11784
rect 20809 11781 20821 11784
rect 20855 11781 20867 11815
rect 20809 11775 20867 11781
rect 20714 11744 20720 11756
rect 19024 11716 20116 11744
rect 20675 11716 20720 11744
rect 19024 11704 19030 11716
rect 20714 11704 20720 11716
rect 20772 11704 20778 11756
rect 16666 11676 16672 11688
rect 15160 11648 16252 11676
rect 16627 11648 16672 11676
rect 15160 11636 15166 11648
rect 16666 11636 16672 11648
rect 16724 11636 16730 11688
rect 17678 11636 17684 11688
rect 17736 11676 17742 11688
rect 18877 11679 18935 11685
rect 18877 11676 18889 11679
rect 17736 11648 18889 11676
rect 17736 11636 17742 11648
rect 18877 11645 18889 11648
rect 18923 11645 18935 11679
rect 19794 11676 19800 11688
rect 19755 11648 19800 11676
rect 18877 11639 18935 11645
rect 19794 11636 19800 11648
rect 19852 11636 19858 11688
rect 19978 11676 19984 11688
rect 19939 11648 19984 11676
rect 19978 11636 19984 11648
rect 20036 11636 20042 11688
rect 20901 11679 20959 11685
rect 20901 11645 20913 11679
rect 20947 11645 20959 11679
rect 20901 11639 20959 11645
rect 5074 11568 5080 11620
rect 5132 11608 5138 11620
rect 7285 11611 7343 11617
rect 7285 11608 7297 11611
rect 5132 11580 7297 11608
rect 5132 11568 5138 11580
rect 7285 11577 7297 11580
rect 7331 11608 7343 11611
rect 7650 11608 7656 11620
rect 7331 11580 7656 11608
rect 7331 11577 7343 11580
rect 7285 11571 7343 11577
rect 7650 11568 7656 11580
rect 7708 11568 7714 11620
rect 10318 11568 10324 11620
rect 10376 11608 10382 11620
rect 11330 11608 11336 11620
rect 10376 11580 11336 11608
rect 10376 11568 10382 11580
rect 11330 11568 11336 11580
rect 11388 11568 11394 11620
rect 12912 11580 16427 11608
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 12912 11540 12940 11580
rect 13078 11540 13084 11552
rect 7524 11512 12940 11540
rect 13039 11512 13084 11540
rect 7524 11500 7530 11512
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 14553 11543 14611 11549
rect 14553 11509 14565 11543
rect 14599 11540 14611 11543
rect 15654 11540 15660 11552
rect 14599 11512 15660 11540
rect 14599 11509 14611 11512
rect 14553 11503 14611 11509
rect 15654 11500 15660 11512
rect 15712 11500 15718 11552
rect 16298 11540 16304 11552
rect 16259 11512 16304 11540
rect 16298 11500 16304 11512
rect 16356 11500 16362 11552
rect 16399 11540 16427 11580
rect 20622 11568 20628 11620
rect 20680 11608 20686 11620
rect 20916 11608 20944 11639
rect 20680 11580 20944 11608
rect 20680 11568 20686 11580
rect 16850 11540 16856 11552
rect 16399 11512 16856 11540
rect 16850 11500 16856 11512
rect 16908 11500 16914 11552
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 18104 11512 18149 11540
rect 18104 11500 18110 11512
rect 18230 11500 18236 11552
rect 18288 11540 18294 11552
rect 19337 11543 19395 11549
rect 19337 11540 19349 11543
rect 18288 11512 19349 11540
rect 18288 11500 18294 11512
rect 19337 11509 19349 11512
rect 19383 11509 19395 11543
rect 19337 11503 19395 11509
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 6822 11336 6828 11348
rect 6783 11308 6828 11336
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7653 11339 7711 11345
rect 7653 11305 7665 11339
rect 7699 11336 7711 11339
rect 7742 11336 7748 11348
rect 7699 11308 7748 11336
rect 7699 11305 7711 11308
rect 7653 11299 7711 11305
rect 7742 11296 7748 11308
rect 7800 11296 7806 11348
rect 8570 11336 8576 11348
rect 8531 11308 8576 11336
rect 8570 11296 8576 11308
rect 8628 11296 8634 11348
rect 9214 11296 9220 11348
rect 9272 11336 9278 11348
rect 9490 11336 9496 11348
rect 9272 11308 9496 11336
rect 9272 11296 9278 11308
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 10778 11296 10784 11348
rect 10836 11336 10842 11348
rect 10836 11308 11192 11336
rect 10836 11296 10842 11308
rect 1762 11228 1768 11280
rect 1820 11268 1826 11280
rect 1820 11240 2774 11268
rect 1820 11228 1826 11240
rect 2746 11200 2774 11240
rect 5718 11228 5724 11280
rect 5776 11268 5782 11280
rect 9309 11271 9367 11277
rect 9309 11268 9321 11271
rect 5776 11240 9321 11268
rect 5776 11228 5782 11240
rect 9309 11237 9321 11240
rect 9355 11237 9367 11271
rect 11164 11268 11192 11308
rect 11238 11296 11244 11348
rect 11296 11336 11302 11348
rect 11425 11339 11483 11345
rect 11425 11336 11437 11339
rect 11296 11308 11437 11336
rect 11296 11296 11302 11308
rect 11425 11305 11437 11308
rect 11471 11305 11483 11339
rect 11425 11299 11483 11305
rect 13173 11339 13231 11345
rect 13173 11305 13185 11339
rect 13219 11336 13231 11339
rect 13630 11336 13636 11348
rect 13219 11308 13636 11336
rect 13219 11305 13231 11308
rect 13173 11299 13231 11305
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 14826 11336 14832 11348
rect 14787 11308 14832 11336
rect 14826 11296 14832 11308
rect 14884 11296 14890 11348
rect 14918 11296 14924 11348
rect 14976 11336 14982 11348
rect 16485 11339 16543 11345
rect 16485 11336 16497 11339
rect 14976 11308 16497 11336
rect 14976 11296 14982 11308
rect 16485 11305 16497 11308
rect 16531 11305 16543 11339
rect 16485 11299 16543 11305
rect 16574 11296 16580 11348
rect 16632 11336 16638 11348
rect 17126 11336 17132 11348
rect 16632 11308 17132 11336
rect 16632 11296 16638 11308
rect 17126 11296 17132 11308
rect 17184 11296 17190 11348
rect 18690 11296 18696 11348
rect 18748 11336 18754 11348
rect 21177 11339 21235 11345
rect 21177 11336 21189 11339
rect 18748 11308 21189 11336
rect 18748 11296 18754 11308
rect 21177 11305 21189 11308
rect 21223 11305 21235 11339
rect 21177 11299 21235 11305
rect 14553 11271 14611 11277
rect 11164 11240 13492 11268
rect 9309 11231 9367 11237
rect 5534 11200 5540 11212
rect 2746 11172 5540 11200
rect 5534 11160 5540 11172
rect 5592 11200 5598 11212
rect 7101 11203 7159 11209
rect 7101 11200 7113 11203
rect 5592 11172 7113 11200
rect 5592 11160 5598 11172
rect 7101 11169 7113 11172
rect 7147 11169 7159 11203
rect 8202 11200 8208 11212
rect 7101 11163 7159 11169
rect 7484 11172 8208 11200
rect 7484 11141 7512 11172
rect 8202 11160 8208 11172
rect 8260 11160 8266 11212
rect 11330 11160 11336 11212
rect 11388 11200 11394 11212
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 11388 11172 11989 11200
rect 11388 11160 11394 11172
rect 11977 11169 11989 11172
rect 12023 11169 12035 11203
rect 11977 11163 12035 11169
rect 12621 11203 12679 11209
rect 12621 11169 12633 11203
rect 12667 11200 12679 11203
rect 13078 11200 13084 11212
rect 12667 11172 13084 11200
rect 12667 11169 12679 11172
rect 12621 11163 12679 11169
rect 13078 11160 13084 11172
rect 13136 11160 13142 11212
rect 13464 11209 13492 11240
rect 14553 11237 14565 11271
rect 14599 11237 14611 11271
rect 14553 11231 14611 11237
rect 13449 11203 13507 11209
rect 13449 11169 13461 11203
rect 13495 11169 13507 11203
rect 14568 11200 14596 11231
rect 16298 11228 16304 11280
rect 16356 11268 16362 11280
rect 17678 11268 17684 11280
rect 16356 11240 17684 11268
rect 16356 11228 16362 11240
rect 17678 11228 17684 11240
rect 17736 11228 17742 11280
rect 17862 11228 17868 11280
rect 17920 11268 17926 11280
rect 20717 11271 20775 11277
rect 17920 11240 18552 11268
rect 17920 11228 17926 11240
rect 17034 11200 17040 11212
rect 14568 11172 15240 11200
rect 16995 11172 17040 11200
rect 13449 11163 13507 11169
rect 7469 11135 7527 11141
rect 7469 11101 7481 11135
rect 7515 11101 7527 11135
rect 7469 11095 7527 11101
rect 7650 11092 7656 11144
rect 7708 11132 7714 11144
rect 7929 11135 7987 11141
rect 7929 11132 7941 11135
rect 7708 11104 7941 11132
rect 7708 11092 7714 11104
rect 7929 11101 7941 11104
rect 7975 11101 7987 11135
rect 7929 11095 7987 11101
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 11149 11135 11207 11141
rect 9539 11104 11100 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 3142 11024 3148 11076
rect 3200 11064 3206 11076
rect 5810 11064 5816 11076
rect 3200 11036 5816 11064
rect 3200 11024 3206 11036
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 9033 11067 9091 11073
rect 9033 11033 9045 11067
rect 9079 11064 9091 11067
rect 9214 11064 9220 11076
rect 9079 11036 9220 11064
rect 9079 11033 9091 11036
rect 9033 11027 9091 11033
rect 9214 11024 9220 11036
rect 9272 11024 9278 11076
rect 9398 11024 9404 11076
rect 9456 11064 9462 11076
rect 9456 11036 9904 11064
rect 9456 11024 9462 11036
rect 9766 10996 9772 11008
rect 9727 10968 9772 10996
rect 9766 10956 9772 10968
rect 9824 10956 9830 11008
rect 9876 10996 9904 11036
rect 10502 11024 10508 11076
rect 10560 11064 10566 11076
rect 10882 11067 10940 11073
rect 10882 11064 10894 11067
rect 10560 11036 10894 11064
rect 10560 11024 10566 11036
rect 10882 11033 10894 11036
rect 10928 11033 10940 11067
rect 11072 11064 11100 11104
rect 11149 11101 11161 11135
rect 11195 11132 11207 11135
rect 11790 11132 11796 11144
rect 11195 11104 11796 11132
rect 11195 11101 11207 11104
rect 11149 11095 11207 11101
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 11885 11135 11943 11141
rect 11885 11101 11897 11135
rect 11931 11132 11943 11135
rect 13722 11132 13728 11144
rect 11931 11104 13728 11132
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 13722 11092 13728 11104
rect 13780 11132 13786 11144
rect 14274 11132 14280 11144
rect 13780 11104 14280 11132
rect 13780 11092 13786 11104
rect 14274 11092 14280 11104
rect 14332 11092 14338 11144
rect 14369 11135 14427 11141
rect 14369 11101 14381 11135
rect 14415 11132 14427 11135
rect 15102 11132 15108 11144
rect 14415 11104 15108 11132
rect 14415 11101 14427 11104
rect 14369 11095 14427 11101
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 15212 11132 15240 11172
rect 17034 11160 17040 11172
rect 17092 11200 17098 11212
rect 18524 11209 18552 11240
rect 20717 11237 20729 11271
rect 20763 11268 20775 11271
rect 20990 11268 20996 11280
rect 20763 11240 20996 11268
rect 20763 11237 20775 11240
rect 20717 11231 20775 11237
rect 20990 11228 20996 11240
rect 21048 11268 21054 11280
rect 21450 11268 21456 11280
rect 21048 11240 21456 11268
rect 21048 11228 21054 11240
rect 21450 11228 21456 11240
rect 21508 11228 21514 11280
rect 18049 11203 18107 11209
rect 18049 11200 18061 11203
rect 17092 11172 18061 11200
rect 17092 11160 17098 11172
rect 18049 11169 18061 11172
rect 18095 11169 18107 11203
rect 18049 11163 18107 11169
rect 18509 11203 18567 11209
rect 18509 11169 18521 11203
rect 18555 11169 18567 11203
rect 18509 11163 18567 11169
rect 15470 11132 15476 11144
rect 15212 11104 15476 11132
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 15930 11132 15936 11144
rect 15988 11141 15994 11144
rect 15900 11104 15936 11132
rect 15930 11092 15936 11104
rect 15988 11095 16000 11141
rect 16209 11135 16267 11141
rect 16209 11101 16221 11135
rect 16255 11132 16267 11135
rect 16666 11132 16672 11144
rect 16255 11104 16672 11132
rect 16255 11101 16267 11104
rect 16209 11095 16267 11101
rect 15988 11092 15994 11095
rect 16666 11092 16672 11104
rect 16724 11132 16730 11144
rect 18138 11132 18144 11144
rect 16724 11104 18144 11132
rect 16724 11092 16730 11104
rect 18138 11092 18144 11104
rect 18196 11132 18202 11144
rect 19242 11132 19248 11144
rect 18196 11104 19248 11132
rect 18196 11092 18202 11104
rect 19242 11092 19248 11104
rect 19300 11132 19306 11144
rect 19337 11135 19395 11141
rect 19337 11132 19349 11135
rect 19300 11104 19349 11132
rect 19300 11092 19306 11104
rect 19337 11101 19349 11104
rect 19383 11101 19395 11135
rect 19337 11095 19395 11101
rect 16574 11064 16580 11076
rect 11072 11036 16580 11064
rect 10882 11027 10940 11033
rect 16574 11024 16580 11036
rect 16632 11024 16638 11076
rect 16945 11067 17003 11073
rect 16945 11033 16957 11067
rect 16991 11064 17003 11067
rect 16991 11036 17080 11064
rect 16991 11033 17003 11036
rect 16945 11027 17003 11033
rect 11793 10999 11851 11005
rect 11793 10996 11805 10999
rect 9876 10968 11805 10996
rect 11793 10965 11805 10968
rect 11839 10965 11851 10999
rect 12710 10996 12716 11008
rect 12671 10968 12716 10996
rect 11793 10959 11851 10965
rect 12710 10956 12716 10968
rect 12768 10956 12774 11008
rect 12802 10956 12808 11008
rect 12860 10996 12866 11008
rect 12860 10968 12905 10996
rect 12860 10956 12866 10968
rect 16390 10956 16396 11008
rect 16448 10996 16454 11008
rect 16853 10999 16911 11005
rect 16853 10996 16865 10999
rect 16448 10968 16865 10996
rect 16448 10956 16454 10968
rect 16853 10965 16865 10968
rect 16899 10965 16911 10999
rect 17052 10996 17080 11036
rect 17126 11024 17132 11076
rect 17184 11064 17190 11076
rect 18230 11064 18236 11076
rect 17184 11036 18236 11064
rect 17184 11024 17190 11036
rect 18230 11024 18236 11036
rect 18288 11024 18294 11076
rect 18414 11024 18420 11076
rect 18472 11064 18478 11076
rect 19582 11067 19640 11073
rect 19582 11064 19594 11067
rect 18472 11036 19594 11064
rect 18472 11024 18478 11036
rect 19582 11033 19594 11036
rect 19628 11033 19640 11067
rect 19582 11027 19640 11033
rect 21269 11067 21327 11073
rect 21269 11033 21281 11067
rect 21315 11064 21327 11067
rect 21634 11064 21640 11076
rect 21315 11036 21640 11064
rect 21315 11033 21327 11036
rect 21269 11027 21327 11033
rect 21634 11024 21640 11036
rect 21692 11024 21698 11076
rect 17218 10996 17224 11008
rect 17052 10968 17224 10996
rect 16853 10959 16911 10965
rect 17218 10956 17224 10968
rect 17276 10956 17282 11008
rect 17494 10996 17500 11008
rect 17455 10968 17500 10996
rect 17494 10956 17500 10968
rect 17552 10956 17558 11008
rect 17678 10956 17684 11008
rect 17736 10996 17742 11008
rect 17865 10999 17923 11005
rect 17865 10996 17877 10999
rect 17736 10968 17877 10996
rect 17736 10956 17742 10968
rect 17865 10965 17877 10968
rect 17911 10965 17923 10999
rect 17865 10959 17923 10965
rect 17954 10956 17960 11008
rect 18012 10996 18018 11008
rect 18012 10968 18057 10996
rect 18012 10956 18018 10968
rect 1104 10906 21896 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21896 10906
rect 1104 10832 21896 10854
rect 8110 10752 8116 10804
rect 8168 10792 8174 10804
rect 8205 10795 8263 10801
rect 8205 10792 8217 10795
rect 8168 10764 8217 10792
rect 8168 10752 8174 10764
rect 8205 10761 8217 10764
rect 8251 10761 8263 10795
rect 8205 10755 8263 10761
rect 9125 10795 9183 10801
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 9769 10795 9827 10801
rect 9171 10764 9720 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 6549 10727 6607 10733
rect 6549 10693 6561 10727
rect 6595 10724 6607 10727
rect 9306 10724 9312 10736
rect 6595 10696 9312 10724
rect 6595 10693 6607 10696
rect 6549 10687 6607 10693
rect 7576 10665 7604 10696
rect 9306 10684 9312 10696
rect 9364 10684 9370 10736
rect 9692 10724 9720 10764
rect 9769 10761 9781 10795
rect 9815 10792 9827 10795
rect 10042 10792 10048 10804
rect 9815 10764 10048 10792
rect 9815 10761 9827 10764
rect 9769 10755 9827 10761
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 10137 10795 10195 10801
rect 10137 10761 10149 10795
rect 10183 10792 10195 10795
rect 10226 10792 10232 10804
rect 10183 10764 10232 10792
rect 10183 10761 10195 10764
rect 10137 10755 10195 10761
rect 10226 10752 10232 10764
rect 10284 10752 10290 10804
rect 10778 10792 10784 10804
rect 10739 10764 10784 10792
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 11149 10795 11207 10801
rect 11149 10761 11161 10795
rect 11195 10792 11207 10795
rect 12802 10792 12808 10804
rect 11195 10764 12808 10792
rect 11195 10761 11207 10764
rect 11149 10755 11207 10761
rect 12802 10752 12808 10764
rect 12860 10752 12866 10804
rect 13081 10795 13139 10801
rect 13081 10761 13093 10795
rect 13127 10761 13139 10795
rect 13081 10755 13139 10761
rect 14553 10795 14611 10801
rect 14553 10761 14565 10795
rect 14599 10792 14611 10795
rect 15010 10792 15016 10804
rect 14599 10764 15016 10792
rect 14599 10761 14611 10764
rect 14553 10755 14611 10761
rect 11790 10724 11796 10736
rect 9692 10696 11796 10724
rect 11790 10684 11796 10696
rect 11848 10684 11854 10736
rect 11968 10727 12026 10733
rect 11968 10693 11980 10727
rect 12014 10724 12026 10727
rect 12066 10724 12072 10736
rect 12014 10696 12072 10724
rect 12014 10693 12026 10696
rect 11968 10687 12026 10693
rect 12066 10684 12072 10696
rect 12124 10684 12130 10736
rect 12250 10684 12256 10736
rect 12308 10724 12314 10736
rect 13096 10724 13124 10755
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 15197 10795 15255 10801
rect 15197 10761 15209 10795
rect 15243 10792 15255 10795
rect 15286 10792 15292 10804
rect 15243 10764 15292 10792
rect 15243 10761 15255 10764
rect 15197 10755 15255 10761
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 15657 10795 15715 10801
rect 15657 10761 15669 10795
rect 15703 10792 15715 10795
rect 16206 10792 16212 10804
rect 15703 10764 16212 10792
rect 15703 10761 15715 10764
rect 15657 10755 15715 10761
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 18325 10795 18383 10801
rect 18325 10761 18337 10795
rect 18371 10792 18383 10795
rect 19978 10792 19984 10804
rect 18371 10764 19984 10792
rect 18371 10761 18383 10764
rect 18325 10755 18383 10761
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 12308 10696 13124 10724
rect 14093 10727 14151 10733
rect 12308 10684 12314 10696
rect 14093 10693 14105 10727
rect 14139 10724 14151 10727
rect 14918 10724 14924 10736
rect 14139 10696 14924 10724
rect 14139 10693 14151 10696
rect 14093 10687 14151 10693
rect 14918 10684 14924 10696
rect 14976 10684 14982 10736
rect 17494 10724 17500 10736
rect 15212 10696 17500 10724
rect 7561 10659 7619 10665
rect 7561 10625 7573 10659
rect 7607 10625 7619 10659
rect 7561 10619 7619 10625
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10656 8539 10659
rect 9766 10656 9772 10668
rect 8527 10628 9772 10656
rect 8527 10625 8539 10628
rect 8481 10619 8539 10625
rect 9306 10548 9312 10600
rect 9364 10588 9370 10600
rect 9490 10588 9496 10600
rect 9364 10560 9496 10588
rect 9364 10548 9370 10560
rect 9490 10548 9496 10560
rect 9548 10548 9554 10600
rect 9600 10597 9628 10628
rect 9766 10616 9772 10628
rect 9824 10616 9830 10668
rect 11146 10616 11152 10668
rect 11204 10656 11210 10668
rect 12342 10656 12348 10668
rect 11204 10628 12348 10656
rect 11204 10616 11210 10628
rect 12342 10616 12348 10628
rect 12400 10616 12406 10668
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10656 14243 10659
rect 15212 10656 15240 10696
rect 17494 10684 17500 10696
rect 17552 10684 17558 10736
rect 17954 10724 17960 10736
rect 17604 10696 17960 10724
rect 14231 10628 15240 10656
rect 14231 10625 14243 10628
rect 14185 10619 14243 10625
rect 15286 10616 15292 10668
rect 15344 10656 15350 10668
rect 15930 10656 15936 10668
rect 15344 10628 15389 10656
rect 15843 10628 15936 10656
rect 15344 10616 15350 10628
rect 15930 10616 15936 10628
rect 15988 10656 15994 10668
rect 17604 10656 17632 10696
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 18046 10684 18052 10736
rect 18104 10684 18110 10736
rect 19242 10684 19248 10736
rect 19300 10724 19306 10736
rect 20254 10733 20260 10736
rect 19300 10696 19748 10724
rect 19300 10684 19306 10696
rect 15988 10628 17632 10656
rect 17793 10659 17851 10665
rect 15988 10616 15994 10628
rect 17793 10625 17805 10659
rect 17839 10656 17851 10659
rect 18064 10656 18092 10684
rect 18230 10656 18236 10668
rect 17839 10628 18236 10656
rect 17839 10625 17851 10628
rect 17793 10619 17851 10625
rect 18230 10616 18236 10628
rect 18288 10616 18294 10668
rect 19720 10665 19748 10696
rect 20248 10687 20260 10733
rect 20312 10724 20318 10736
rect 20312 10696 20348 10724
rect 20254 10684 20260 10687
rect 20312 10684 20318 10696
rect 19449 10659 19507 10665
rect 19449 10625 19461 10659
rect 19495 10656 19507 10659
rect 19705 10659 19763 10665
rect 19495 10628 19656 10656
rect 19495 10625 19507 10628
rect 19449 10619 19507 10625
rect 9585 10591 9643 10597
rect 9585 10557 9597 10591
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10588 9735 10591
rect 10134 10588 10140 10600
rect 9723 10560 10140 10588
rect 9723 10557 9735 10560
rect 9677 10551 9735 10557
rect 10134 10548 10140 10560
rect 10192 10548 10198 10600
rect 10597 10591 10655 10597
rect 10597 10557 10609 10591
rect 10643 10557 10655 10591
rect 10597 10551 10655 10557
rect 10689 10591 10747 10597
rect 10689 10557 10701 10591
rect 10735 10557 10747 10591
rect 10689 10551 10747 10557
rect 5626 10480 5632 10532
rect 5684 10520 5690 10532
rect 7193 10523 7251 10529
rect 7193 10520 7205 10523
rect 5684 10492 7205 10520
rect 5684 10480 5690 10492
rect 7193 10489 7205 10492
rect 7239 10489 7251 10523
rect 7742 10520 7748 10532
rect 7703 10492 7748 10520
rect 7193 10483 7251 10489
rect 7742 10480 7748 10492
rect 7800 10480 7806 10532
rect 8386 10480 8392 10532
rect 8444 10520 8450 10532
rect 9122 10520 9128 10532
rect 8444 10492 9128 10520
rect 8444 10480 8450 10492
rect 9122 10480 9128 10492
rect 9180 10480 9186 10532
rect 6638 10412 6644 10464
rect 6696 10452 6702 10464
rect 6822 10452 6828 10464
rect 6696 10424 6828 10452
rect 6696 10412 6702 10424
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 6917 10455 6975 10461
rect 6917 10421 6929 10455
rect 6963 10452 6975 10455
rect 10226 10452 10232 10464
rect 6963 10424 10232 10452
rect 6963 10421 6975 10424
rect 6917 10415 6975 10421
rect 10226 10412 10232 10424
rect 10284 10412 10290 10464
rect 10612 10452 10640 10551
rect 10704 10520 10732 10551
rect 11054 10548 11060 10600
rect 11112 10588 11118 10600
rect 11701 10591 11759 10597
rect 11701 10588 11713 10591
rect 11112 10560 11713 10588
rect 11112 10548 11118 10560
rect 11701 10557 11713 10560
rect 11747 10557 11759 10591
rect 11701 10551 11759 10557
rect 13262 10548 13268 10600
rect 13320 10588 13326 10600
rect 13541 10591 13599 10597
rect 13541 10588 13553 10591
rect 13320 10560 13553 10588
rect 13320 10548 13326 10560
rect 13541 10557 13553 10560
rect 13587 10557 13599 10591
rect 13541 10551 13599 10557
rect 13814 10548 13820 10600
rect 13872 10588 13878 10600
rect 13909 10591 13967 10597
rect 13909 10588 13921 10591
rect 13872 10560 13921 10588
rect 13872 10548 13878 10560
rect 13909 10557 13921 10560
rect 13955 10557 13967 10591
rect 13909 10551 13967 10557
rect 15105 10591 15163 10597
rect 15105 10557 15117 10591
rect 15151 10588 15163 10591
rect 15194 10588 15200 10600
rect 15151 10560 15200 10588
rect 15151 10557 15163 10560
rect 15105 10551 15163 10557
rect 15194 10548 15200 10560
rect 15252 10588 15258 10600
rect 17034 10588 17040 10600
rect 15252 10560 17040 10588
rect 15252 10548 15258 10560
rect 17034 10548 17040 10560
rect 17092 10548 17098 10600
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 18138 10588 18144 10600
rect 18095 10560 18144 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 18138 10548 18144 10560
rect 18196 10548 18202 10600
rect 19628 10588 19656 10628
rect 19705 10625 19717 10659
rect 19751 10656 19763 10659
rect 19981 10659 20039 10665
rect 19981 10656 19993 10659
rect 19751 10628 19993 10656
rect 19751 10625 19763 10628
rect 19705 10619 19763 10625
rect 19981 10625 19993 10628
rect 20027 10625 20039 10659
rect 19981 10619 20039 10625
rect 19628 10560 19748 10588
rect 10704 10492 11560 10520
rect 11238 10452 11244 10464
rect 10612 10424 11244 10452
rect 11238 10412 11244 10424
rect 11296 10412 11302 10464
rect 11532 10452 11560 10492
rect 12802 10480 12808 10532
rect 12860 10520 12866 10532
rect 15562 10520 15568 10532
rect 12860 10492 15568 10520
rect 12860 10480 12866 10492
rect 15562 10480 15568 10492
rect 15620 10480 15626 10532
rect 15663 10492 16804 10520
rect 13814 10452 13820 10464
rect 11532 10424 13820 10452
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 14274 10412 14280 10464
rect 14332 10452 14338 10464
rect 15663 10452 15691 10492
rect 14332 10424 15691 10452
rect 16117 10455 16175 10461
rect 14332 10412 14338 10424
rect 16117 10421 16129 10455
rect 16163 10452 16175 10455
rect 16206 10452 16212 10464
rect 16163 10424 16212 10452
rect 16163 10421 16175 10424
rect 16117 10415 16175 10421
rect 16206 10412 16212 10424
rect 16264 10412 16270 10464
rect 16666 10452 16672 10464
rect 16627 10424 16672 10452
rect 16666 10412 16672 10424
rect 16724 10412 16730 10464
rect 16776 10452 16804 10492
rect 18046 10452 18052 10464
rect 16776 10424 18052 10452
rect 18046 10412 18052 10424
rect 18104 10412 18110 10464
rect 19720 10452 19748 10560
rect 20622 10452 20628 10464
rect 19720 10424 20628 10452
rect 20622 10412 20628 10424
rect 20680 10412 20686 10464
rect 20898 10412 20904 10464
rect 20956 10452 20962 10464
rect 21174 10452 21180 10464
rect 20956 10424 21180 10452
rect 20956 10412 20962 10424
rect 21174 10412 21180 10424
rect 21232 10452 21238 10464
rect 21361 10455 21419 10461
rect 21361 10452 21373 10455
rect 21232 10424 21373 10452
rect 21232 10412 21238 10424
rect 21361 10421 21373 10424
rect 21407 10421 21419 10455
rect 21361 10415 21419 10421
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 4246 10208 4252 10260
rect 4304 10248 4310 10260
rect 7101 10251 7159 10257
rect 7101 10248 7113 10251
rect 4304 10220 7113 10248
rect 4304 10208 4310 10220
rect 7101 10217 7113 10220
rect 7147 10248 7159 10251
rect 7650 10248 7656 10260
rect 7147 10220 7656 10248
rect 7147 10217 7159 10220
rect 7101 10211 7159 10217
rect 7650 10208 7656 10220
rect 7708 10208 7714 10260
rect 7926 10208 7932 10260
rect 7984 10248 7990 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 7984 10220 8953 10248
rect 7984 10208 7990 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 8941 10211 8999 10217
rect 9140 10220 10097 10248
rect 8386 10180 8392 10192
rect 7300 10152 8392 10180
rect 7300 10124 7328 10152
rect 8386 10140 8392 10152
rect 8444 10140 8450 10192
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 7282 10112 7288 10124
rect 6871 10084 7288 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 7282 10072 7288 10084
rect 7340 10072 7346 10124
rect 5810 10004 5816 10056
rect 5868 10044 5874 10056
rect 6730 10044 6736 10056
rect 5868 10016 6736 10044
rect 5868 10004 5874 10016
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 7466 10044 7472 10056
rect 7427 10016 7472 10044
rect 7466 10004 7472 10016
rect 7524 10004 7530 10056
rect 8570 10044 8576 10056
rect 8531 10016 8576 10044
rect 8570 10004 8576 10016
rect 8628 10004 8634 10056
rect 9140 10053 9168 10220
rect 9490 10072 9496 10124
rect 9548 10112 9554 10124
rect 10069 10112 10097 10220
rect 10226 10208 10232 10260
rect 10284 10248 10290 10260
rect 12621 10251 12679 10257
rect 10284 10220 12434 10248
rect 10284 10208 10290 10220
rect 10134 10140 10140 10192
rect 10192 10180 10198 10192
rect 11977 10183 12035 10189
rect 10192 10152 10237 10180
rect 10192 10140 10198 10152
rect 11977 10149 11989 10183
rect 12023 10180 12035 10183
rect 12066 10180 12072 10192
rect 12023 10152 12072 10180
rect 12023 10149 12035 10152
rect 11977 10143 12035 10149
rect 12066 10140 12072 10152
rect 12124 10140 12130 10192
rect 12406 10180 12434 10220
rect 12621 10217 12633 10251
rect 12667 10248 12679 10251
rect 12710 10248 12716 10260
rect 12667 10220 12716 10248
rect 12667 10217 12679 10220
rect 12621 10211 12679 10217
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 13872 10220 14105 10248
rect 13872 10208 13878 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 15562 10208 15568 10260
rect 15620 10248 15626 10260
rect 15620 10220 16068 10248
rect 15620 10208 15626 10220
rect 15930 10180 15936 10192
rect 12406 10152 15936 10180
rect 15930 10140 15936 10152
rect 15988 10140 15994 10192
rect 16040 10180 16068 10220
rect 16114 10208 16120 10260
rect 16172 10248 16178 10260
rect 16853 10251 16911 10257
rect 16853 10248 16865 10251
rect 16172 10220 16865 10248
rect 16172 10208 16178 10220
rect 16853 10217 16865 10220
rect 16899 10217 16911 10251
rect 20346 10248 20352 10260
rect 16853 10211 16911 10217
rect 16951 10220 20352 10248
rect 16951 10180 16979 10220
rect 20346 10208 20352 10220
rect 20404 10208 20410 10260
rect 20622 10248 20628 10260
rect 20583 10220 20628 10248
rect 20622 10208 20628 10220
rect 20680 10208 20686 10260
rect 16040 10152 16979 10180
rect 9548 10084 9593 10112
rect 10069 10084 10456 10112
rect 9548 10072 9554 10084
rect 10428 10056 10456 10084
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 10410 10004 10416 10056
rect 10468 10004 10474 10056
rect 10597 10047 10655 10053
rect 10597 10013 10609 10047
rect 10643 10044 10655 10047
rect 12084 10044 12112 10140
rect 12250 10072 12256 10124
rect 12308 10112 12314 10124
rect 13173 10115 13231 10121
rect 13173 10112 13185 10115
rect 12308 10084 13185 10112
rect 12308 10072 12314 10084
rect 13173 10081 13185 10084
rect 13219 10081 13231 10115
rect 13173 10075 13231 10081
rect 13538 10072 13544 10124
rect 13596 10112 13602 10124
rect 14550 10112 14556 10124
rect 13596 10084 14556 10112
rect 13596 10072 13602 10084
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 14645 10115 14703 10121
rect 14645 10081 14657 10115
rect 14691 10112 14703 10115
rect 15657 10115 15715 10121
rect 15657 10112 15669 10115
rect 14691 10084 15669 10112
rect 14691 10081 14703 10084
rect 14645 10075 14703 10081
rect 15657 10081 15669 10084
rect 15703 10081 15715 10115
rect 17218 10112 17224 10124
rect 15657 10075 15715 10081
rect 16592 10084 17224 10112
rect 13998 10044 14004 10056
rect 10643 10016 11100 10044
rect 12084 10016 14004 10044
rect 10643 10013 10655 10016
rect 10597 10007 10655 10013
rect 11072 9988 11100 10016
rect 13998 10004 14004 10016
rect 14056 10044 14062 10056
rect 14660 10044 14688 10075
rect 14056 10016 14688 10044
rect 14056 10004 14062 10016
rect 14734 10004 14740 10056
rect 14792 10044 14798 10056
rect 15473 10047 15531 10053
rect 15473 10044 15485 10047
rect 14792 10016 15485 10044
rect 14792 10004 14798 10016
rect 15473 10013 15485 10016
rect 15519 10013 15531 10047
rect 16592 10044 16620 10084
rect 17218 10072 17224 10084
rect 17276 10072 17282 10124
rect 19245 10115 19303 10121
rect 19245 10112 19257 10115
rect 18248 10084 19257 10112
rect 15473 10007 15531 10013
rect 15580 10016 16620 10044
rect 6638 9936 6644 9988
rect 6696 9976 6702 9988
rect 7926 9976 7932 9988
rect 6696 9948 7788 9976
rect 7887 9948 7932 9976
rect 6696 9936 6702 9948
rect 5902 9868 5908 9920
rect 5960 9908 5966 9920
rect 6365 9911 6423 9917
rect 6365 9908 6377 9911
rect 5960 9880 6377 9908
rect 5960 9868 5966 9880
rect 6365 9877 6377 9880
rect 6411 9908 6423 9911
rect 6546 9908 6552 9920
rect 6411 9880 6552 9908
rect 6411 9877 6423 9880
rect 6365 9871 6423 9877
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 7650 9908 7656 9920
rect 7611 9880 7656 9908
rect 7650 9868 7656 9880
rect 7708 9868 7714 9920
rect 7760 9908 7788 9948
rect 7926 9936 7932 9948
rect 7984 9936 7990 9988
rect 8386 9936 8392 9988
rect 8444 9976 8450 9988
rect 9677 9979 9735 9985
rect 9677 9976 9689 9979
rect 8444 9948 9689 9976
rect 8444 9936 8450 9948
rect 9677 9945 9689 9948
rect 9723 9945 9735 9979
rect 9677 9939 9735 9945
rect 10318 9936 10324 9988
rect 10376 9976 10382 9988
rect 10842 9979 10900 9985
rect 10842 9976 10854 9979
rect 10376 9948 10854 9976
rect 10376 9936 10382 9948
rect 10842 9945 10854 9948
rect 10888 9945 10900 9979
rect 10842 9939 10900 9945
rect 11054 9936 11060 9988
rect 11112 9936 11118 9988
rect 11698 9936 11704 9988
rect 11756 9976 11762 9988
rect 12158 9976 12164 9988
rect 11756 9948 12164 9976
rect 11756 9936 11762 9948
rect 12158 9936 12164 9948
rect 12216 9976 12222 9988
rect 12345 9979 12403 9985
rect 12345 9976 12357 9979
rect 12216 9948 12357 9976
rect 12216 9936 12222 9948
rect 12345 9945 12357 9948
rect 12391 9945 12403 9979
rect 12345 9939 12403 9945
rect 13081 9979 13139 9985
rect 13081 9945 13093 9979
rect 13127 9976 13139 9979
rect 13127 9948 15148 9976
rect 13127 9945 13139 9948
rect 13081 9939 13139 9945
rect 9769 9911 9827 9917
rect 9769 9908 9781 9911
rect 7760 9880 9781 9908
rect 9769 9877 9781 9880
rect 9815 9877 9827 9911
rect 12986 9908 12992 9920
rect 12947 9880 12992 9908
rect 9769 9871 9827 9877
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 13725 9911 13783 9917
rect 13725 9877 13737 9911
rect 13771 9908 13783 9911
rect 14274 9908 14280 9920
rect 13771 9880 14280 9908
rect 13771 9877 13783 9880
rect 13725 9871 13783 9877
rect 14274 9868 14280 9880
rect 14332 9868 14338 9920
rect 14458 9908 14464 9920
rect 14419 9880 14464 9908
rect 14458 9868 14464 9880
rect 14516 9868 14522 9920
rect 14550 9868 14556 9920
rect 14608 9908 14614 9920
rect 15120 9917 15148 9948
rect 15105 9911 15163 9917
rect 14608 9880 14653 9908
rect 14608 9868 14614 9880
rect 15105 9877 15117 9911
rect 15151 9877 15163 9911
rect 15105 9871 15163 9877
rect 15194 9868 15200 9920
rect 15252 9908 15258 9920
rect 15580 9917 15608 10016
rect 16666 10004 16672 10056
rect 16724 10044 16730 10056
rect 17678 10044 17684 10056
rect 16724 10016 17684 10044
rect 16724 10004 16730 10016
rect 17678 10004 17684 10016
rect 17736 10044 17742 10056
rect 17966 10047 18024 10053
rect 17966 10044 17978 10047
rect 17736 10016 17978 10044
rect 17736 10004 17742 10016
rect 17966 10013 17978 10016
rect 18012 10013 18024 10047
rect 17966 10007 18024 10013
rect 18138 10004 18144 10056
rect 18196 10044 18202 10056
rect 18248 10053 18276 10084
rect 19245 10081 19257 10084
rect 19291 10081 19303 10115
rect 19245 10075 19303 10081
rect 18233 10047 18291 10053
rect 18233 10044 18245 10047
rect 18196 10016 18245 10044
rect 18196 10004 18202 10016
rect 18233 10013 18245 10016
rect 18279 10013 18291 10047
rect 18598 10044 18604 10056
rect 18559 10016 18604 10044
rect 18233 10007 18291 10013
rect 18598 10004 18604 10016
rect 18656 10004 18662 10056
rect 19334 10004 19340 10056
rect 19392 10044 19398 10056
rect 19501 10047 19559 10053
rect 19501 10044 19513 10047
rect 19392 10016 19513 10044
rect 19392 10004 19398 10016
rect 19501 10013 19513 10016
rect 19547 10013 19559 10047
rect 19501 10007 19559 10013
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 20901 10047 20959 10053
rect 20901 10044 20913 10047
rect 20772 10016 20913 10044
rect 20772 10004 20778 10016
rect 20901 10013 20913 10016
rect 20947 10013 20959 10047
rect 20901 10007 20959 10013
rect 16577 9979 16635 9985
rect 16577 9945 16589 9979
rect 16623 9976 16635 9979
rect 20162 9976 20168 9988
rect 16623 9948 20168 9976
rect 16623 9945 16635 9948
rect 16577 9939 16635 9945
rect 20162 9936 20168 9948
rect 20220 9936 20226 9988
rect 15565 9911 15623 9917
rect 15565 9908 15577 9911
rect 15252 9880 15577 9908
rect 15252 9868 15258 9880
rect 15565 9877 15577 9880
rect 15611 9877 15623 9911
rect 15565 9871 15623 9877
rect 15838 9868 15844 9920
rect 15896 9908 15902 9920
rect 17862 9908 17868 9920
rect 15896 9880 17868 9908
rect 15896 9868 15902 9880
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 18785 9911 18843 9917
rect 18785 9877 18797 9911
rect 18831 9908 18843 9911
rect 19886 9908 19892 9920
rect 18831 9880 19892 9908
rect 18831 9877 18843 9880
rect 18785 9871 18843 9877
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 20806 9868 20812 9920
rect 20864 9908 20870 9920
rect 21085 9911 21143 9917
rect 21085 9908 21097 9911
rect 20864 9880 21097 9908
rect 20864 9868 20870 9880
rect 21085 9877 21097 9880
rect 21131 9877 21143 9911
rect 21085 9871 21143 9877
rect 1104 9818 21896 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21896 9818
rect 1104 9744 21896 9766
rect 7466 9704 7472 9716
rect 7427 9676 7472 9704
rect 7466 9664 7472 9676
rect 7524 9664 7530 9716
rect 7650 9664 7656 9716
rect 7708 9704 7714 9716
rect 12066 9704 12072 9716
rect 7708 9676 12072 9704
rect 7708 9664 7714 9676
rect 12066 9664 12072 9676
rect 12124 9664 12130 9716
rect 12986 9664 12992 9716
rect 13044 9704 13050 9716
rect 13357 9707 13415 9713
rect 13357 9704 13369 9707
rect 13044 9676 13369 9704
rect 13044 9664 13050 9676
rect 13357 9673 13369 9676
rect 13403 9673 13415 9707
rect 13357 9667 13415 9673
rect 14550 9664 14556 9716
rect 14608 9704 14614 9716
rect 15102 9704 15108 9716
rect 14608 9676 15108 9704
rect 14608 9664 14614 9676
rect 15102 9664 15108 9676
rect 15160 9664 15166 9716
rect 15838 9704 15844 9716
rect 15221 9676 15844 9704
rect 1854 9596 1860 9648
rect 1912 9636 1918 9648
rect 6822 9636 6828 9648
rect 1912 9608 6828 9636
rect 1912 9596 1918 9608
rect 6822 9596 6828 9608
rect 6880 9636 6886 9648
rect 7282 9636 7288 9648
rect 6880 9608 7288 9636
rect 6880 9596 6886 9608
rect 7282 9596 7288 9608
rect 7340 9596 7346 9648
rect 7745 9639 7803 9645
rect 7745 9605 7757 9639
rect 7791 9636 7803 9639
rect 8294 9636 8300 9648
rect 7791 9608 8300 9636
rect 7791 9605 7803 9608
rect 7745 9599 7803 9605
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 8662 9636 8668 9648
rect 8623 9608 8668 9636
rect 8662 9596 8668 9608
rect 8720 9596 8726 9648
rect 9122 9596 9128 9648
rect 9180 9636 9186 9648
rect 9180 9608 9444 9636
rect 9180 9596 9186 9608
rect 7098 9568 7104 9580
rect 7059 9540 7104 9568
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 8386 9568 8392 9580
rect 8347 9540 8392 9568
rect 8386 9528 8392 9540
rect 8444 9528 8450 9580
rect 9309 9571 9367 9577
rect 9309 9537 9321 9571
rect 9355 9537 9367 9571
rect 9416 9568 9444 9608
rect 9490 9596 9496 9648
rect 9548 9636 9554 9648
rect 10698 9639 10756 9645
rect 10698 9636 10710 9639
rect 9548 9608 10710 9636
rect 9548 9596 9554 9608
rect 10698 9605 10710 9608
rect 10744 9636 10756 9639
rect 11698 9636 11704 9648
rect 10744 9608 11704 9636
rect 10744 9605 10756 9608
rect 10698 9599 10756 9605
rect 11698 9596 11704 9608
rect 11756 9596 11762 9648
rect 11974 9596 11980 9648
rect 12032 9636 12038 9648
rect 12161 9639 12219 9645
rect 12161 9636 12173 9639
rect 12032 9608 12173 9636
rect 12032 9596 12038 9608
rect 12161 9605 12173 9608
rect 12207 9605 12219 9639
rect 12161 9599 12219 9605
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 12492 9608 12537 9636
rect 12492 9596 12498 9608
rect 14366 9596 14372 9648
rect 14424 9636 14430 9648
rect 15221 9636 15249 9676
rect 15838 9664 15844 9676
rect 15896 9704 15902 9716
rect 15933 9707 15991 9713
rect 15933 9704 15945 9707
rect 15896 9676 15945 9704
rect 15896 9664 15902 9676
rect 15933 9673 15945 9676
rect 15979 9673 15991 9707
rect 15933 9667 15991 9673
rect 16206 9664 16212 9716
rect 16264 9704 16270 9716
rect 20898 9704 20904 9716
rect 16264 9676 20904 9704
rect 16264 9664 16270 9676
rect 20898 9664 20904 9676
rect 20956 9664 20962 9716
rect 14424 9608 15249 9636
rect 14424 9596 14430 9608
rect 16114 9596 16120 9648
rect 16172 9636 16178 9648
rect 16172 9608 16804 9636
rect 16172 9596 16178 9608
rect 9858 9568 9864 9580
rect 9416 9540 9864 9568
rect 9309 9531 9367 9537
rect 5718 9324 5724 9376
rect 5776 9364 5782 9376
rect 6641 9367 6699 9373
rect 6641 9364 6653 9367
rect 5776 9336 6653 9364
rect 5776 9324 5782 9336
rect 6641 9333 6653 9336
rect 6687 9364 6699 9367
rect 6822 9364 6828 9376
rect 6687 9336 6828 9364
rect 6687 9333 6699 9336
rect 6641 9327 6699 9333
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 9324 9364 9352 9531
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 11238 9528 11244 9580
rect 11296 9568 11302 9580
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 11296 9540 11529 9568
rect 11296 9528 11302 9540
rect 11517 9537 11529 9540
rect 11563 9568 11575 9571
rect 12250 9568 12256 9580
rect 11563 9540 12256 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 13078 9568 13084 9580
rect 13039 9540 13084 9568
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 13725 9571 13783 9577
rect 13725 9568 13737 9571
rect 13188 9540 13737 9568
rect 10965 9503 11023 9509
rect 10965 9469 10977 9503
rect 11011 9500 11023 9503
rect 11054 9500 11060 9512
rect 11011 9472 11060 9500
rect 11011 9469 11023 9472
rect 10965 9463 11023 9469
rect 11054 9460 11060 9472
rect 11112 9460 11118 9512
rect 11606 9460 11612 9512
rect 11664 9500 11670 9512
rect 13188 9500 13216 9540
rect 13725 9537 13737 9540
rect 13771 9568 13783 9571
rect 14274 9568 14280 9580
rect 13771 9540 14280 9568
rect 13771 9537 13783 9540
rect 13725 9531 13783 9537
rect 14274 9528 14280 9540
rect 14332 9528 14338 9580
rect 14737 9571 14795 9577
rect 14737 9537 14749 9571
rect 14783 9568 14795 9571
rect 15930 9568 15936 9580
rect 14783 9540 15936 9568
rect 14783 9537 14795 9540
rect 14737 9531 14795 9537
rect 15930 9528 15936 9540
rect 15988 9528 15994 9580
rect 16025 9571 16083 9577
rect 16025 9537 16037 9571
rect 16071 9568 16083 9571
rect 16390 9568 16396 9580
rect 16071 9540 16396 9568
rect 16071 9537 16083 9540
rect 16025 9531 16083 9537
rect 11664 9472 13216 9500
rect 11664 9460 11670 9472
rect 13630 9460 13636 9512
rect 13688 9500 13694 9512
rect 13817 9503 13875 9509
rect 13817 9500 13829 9503
rect 13688 9472 13829 9500
rect 13688 9460 13694 9472
rect 13817 9469 13829 9472
rect 13863 9469 13875 9503
rect 13998 9500 14004 9512
rect 13959 9472 14004 9500
rect 13817 9463 13875 9469
rect 13998 9460 14004 9472
rect 14056 9460 14062 9512
rect 14826 9500 14832 9512
rect 14787 9472 14832 9500
rect 14826 9460 14832 9472
rect 14884 9460 14890 9512
rect 14921 9503 14979 9509
rect 14921 9469 14933 9503
rect 14967 9469 14979 9503
rect 14921 9463 14979 9469
rect 13538 9432 13544 9444
rect 12268 9404 13544 9432
rect 9582 9364 9588 9376
rect 9324 9336 9588 9364
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 10226 9324 10232 9376
rect 10284 9364 10290 9376
rect 12268 9364 12296 9404
rect 13538 9392 13544 9404
rect 13596 9392 13602 9444
rect 14936 9432 14964 9463
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 15746 9500 15752 9512
rect 15344 9472 15752 9500
rect 15344 9460 15350 9472
rect 15746 9460 15752 9472
rect 15804 9460 15810 9512
rect 16114 9500 16120 9512
rect 16075 9472 16120 9500
rect 16114 9460 16120 9472
rect 16172 9460 16178 9512
rect 16224 9432 16252 9540
rect 16390 9528 16396 9540
rect 16448 9528 16454 9580
rect 16776 9568 16804 9608
rect 16850 9596 16856 9648
rect 16908 9636 16914 9648
rect 17221 9639 17279 9645
rect 17221 9636 17233 9639
rect 16908 9608 17233 9636
rect 16908 9596 16914 9608
rect 17221 9605 17233 9608
rect 17267 9605 17279 9639
rect 17221 9599 17279 9605
rect 17954 9596 17960 9648
rect 18012 9636 18018 9648
rect 18386 9639 18444 9645
rect 18386 9636 18398 9639
rect 18012 9608 18398 9636
rect 18012 9596 18018 9608
rect 18386 9605 18398 9608
rect 18432 9605 18444 9639
rect 18386 9599 18444 9605
rect 16942 9568 16948 9580
rect 16776 9540 16948 9568
rect 16942 9528 16948 9540
rect 17000 9528 17006 9580
rect 17034 9528 17040 9580
rect 17092 9568 17098 9580
rect 17129 9571 17187 9577
rect 17129 9568 17141 9571
rect 17092 9540 17141 9568
rect 17092 9528 17098 9540
rect 17129 9537 17141 9540
rect 17175 9537 17187 9571
rect 17129 9531 17187 9537
rect 17773 9571 17831 9577
rect 17773 9537 17785 9571
rect 17819 9568 17831 9571
rect 18690 9568 18696 9580
rect 17819 9540 18696 9568
rect 17819 9537 17831 9540
rect 17773 9531 17831 9537
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 20162 9568 20168 9580
rect 20123 9540 20168 9568
rect 20162 9528 20168 9540
rect 20220 9528 20226 9580
rect 21082 9568 21088 9580
rect 21043 9540 21088 9568
rect 21082 9528 21088 9540
rect 21140 9528 21146 9580
rect 17313 9503 17371 9509
rect 17313 9469 17325 9503
rect 17359 9469 17371 9503
rect 18138 9500 18144 9512
rect 18099 9472 18144 9500
rect 17313 9463 17371 9469
rect 13740 9404 14964 9432
rect 15221 9404 16252 9432
rect 10284 9336 12296 9364
rect 10284 9324 10290 9336
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 13740 9364 13768 9404
rect 13504 9336 13768 9364
rect 13504 9324 13510 9336
rect 13814 9324 13820 9376
rect 13872 9364 13878 9376
rect 14369 9367 14427 9373
rect 14369 9364 14381 9367
rect 13872 9336 14381 9364
rect 13872 9324 13878 9336
rect 14369 9333 14381 9336
rect 14415 9333 14427 9367
rect 14369 9327 14427 9333
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 15221 9364 15249 9404
rect 14792 9336 15249 9364
rect 14792 9324 14798 9336
rect 15286 9324 15292 9376
rect 15344 9364 15350 9376
rect 15565 9367 15623 9373
rect 15565 9364 15577 9367
rect 15344 9336 15577 9364
rect 15344 9324 15350 9336
rect 15565 9333 15577 9336
rect 15611 9333 15623 9367
rect 15565 9327 15623 9333
rect 15838 9324 15844 9376
rect 15896 9364 15902 9376
rect 16574 9364 16580 9376
rect 15896 9336 16580 9364
rect 15896 9324 15902 9336
rect 16574 9324 16580 9336
rect 16632 9324 16638 9376
rect 16666 9324 16672 9376
rect 16724 9364 16730 9376
rect 16761 9367 16819 9373
rect 16761 9364 16773 9367
rect 16724 9336 16773 9364
rect 16724 9324 16730 9336
rect 16761 9333 16773 9336
rect 16807 9333 16819 9367
rect 16761 9327 16819 9333
rect 16942 9324 16948 9376
rect 17000 9364 17006 9376
rect 17328 9364 17356 9463
rect 18138 9460 18144 9472
rect 18196 9460 18202 9512
rect 20254 9500 20260 9512
rect 20215 9472 20260 9500
rect 20254 9460 20260 9472
rect 20312 9460 20318 9512
rect 20346 9460 20352 9512
rect 20404 9460 20410 9512
rect 20441 9503 20499 9509
rect 20441 9469 20453 9503
rect 20487 9500 20499 9503
rect 20622 9500 20628 9512
rect 20487 9472 20628 9500
rect 20487 9469 20499 9472
rect 20441 9463 20499 9469
rect 20622 9460 20628 9472
rect 20680 9460 20686 9512
rect 19518 9432 19524 9444
rect 19479 9404 19524 9432
rect 19518 9392 19524 9404
rect 19576 9392 19582 9444
rect 19794 9432 19800 9444
rect 19755 9404 19800 9432
rect 19794 9392 19800 9404
rect 19852 9392 19858 9444
rect 20364 9432 20392 9460
rect 20364 9404 20668 9432
rect 20640 9376 20668 9404
rect 17000 9336 17356 9364
rect 17000 9324 17006 9336
rect 17402 9324 17408 9376
rect 17460 9364 17466 9376
rect 20346 9364 20352 9376
rect 17460 9336 20352 9364
rect 17460 9324 17466 9336
rect 20346 9324 20352 9336
rect 20404 9324 20410 9376
rect 20622 9324 20628 9376
rect 20680 9324 20686 9376
rect 21266 9364 21272 9376
rect 21227 9336 21272 9364
rect 21266 9324 21272 9336
rect 21324 9324 21330 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 10226 9160 10232 9172
rect 7116 9132 10232 9160
rect 7116 9036 7144 9132
rect 10226 9120 10232 9132
rect 10284 9120 10290 9172
rect 10410 9160 10416 9172
rect 10371 9132 10416 9160
rect 10410 9120 10416 9132
rect 10468 9120 10474 9172
rect 11885 9163 11943 9169
rect 11885 9129 11897 9163
rect 11931 9160 11943 9163
rect 14366 9160 14372 9172
rect 11931 9132 14372 9160
rect 11931 9129 11943 9132
rect 11885 9123 11943 9129
rect 14366 9120 14372 9132
rect 14424 9120 14430 9172
rect 15378 9160 15384 9172
rect 14752 9132 15384 9160
rect 7282 9092 7288 9104
rect 7243 9064 7288 9092
rect 7282 9052 7288 9064
rect 7340 9052 7346 9104
rect 8113 9095 8171 9101
rect 8113 9061 8125 9095
rect 8159 9092 8171 9095
rect 11606 9092 11612 9104
rect 8159 9064 11612 9092
rect 8159 9061 8171 9064
rect 8113 9055 8171 9061
rect 11606 9052 11612 9064
rect 11664 9052 11670 9104
rect 13538 9052 13544 9104
rect 13596 9092 13602 9104
rect 14458 9092 14464 9104
rect 13596 9064 14464 9092
rect 13596 9052 13602 9064
rect 14458 9052 14464 9064
rect 14516 9052 14522 9104
rect 6914 9024 6920 9036
rect 6827 8996 6920 9024
rect 6914 8984 6920 8996
rect 6972 9024 6978 9036
rect 7098 9024 7104 9036
rect 6972 8996 7104 9024
rect 6972 8984 6978 8996
rect 7098 8984 7104 8996
rect 7156 8984 7162 9036
rect 8478 9024 8484 9036
rect 7208 8996 8484 9024
rect 6822 8916 6828 8968
rect 6880 8956 6886 8968
rect 7208 8956 7236 8996
rect 8478 8984 8484 8996
rect 8536 8984 8542 9036
rect 9490 9024 9496 9036
rect 9451 8996 9496 9024
rect 9490 8984 9496 8996
rect 9548 8984 9554 9036
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 10965 9027 11023 9033
rect 10965 9024 10977 9027
rect 9640 8996 10977 9024
rect 9640 8984 9646 8996
rect 10965 8993 10977 8996
rect 11011 8993 11023 9027
rect 10965 8987 11023 8993
rect 11054 8984 11060 9036
rect 11112 9024 11118 9036
rect 12158 9024 12164 9036
rect 11112 8996 12164 9024
rect 11112 8984 11118 8996
rect 12158 8984 12164 8996
rect 12216 8984 12222 9036
rect 13722 8984 13728 9036
rect 13780 9024 13786 9036
rect 14752 9024 14780 9132
rect 15378 9120 15384 9132
rect 15436 9160 15442 9172
rect 15436 9132 15884 9160
rect 15436 9120 15442 9132
rect 13780 8996 14780 9024
rect 15856 9024 15884 9132
rect 15930 9120 15936 9172
rect 15988 9160 15994 9172
rect 16025 9163 16083 9169
rect 16025 9160 16037 9163
rect 15988 9132 16037 9160
rect 15988 9120 15994 9132
rect 16025 9129 16037 9132
rect 16071 9129 16083 9163
rect 16025 9123 16083 9129
rect 16574 9120 16580 9172
rect 16632 9160 16638 9172
rect 16632 9132 16804 9160
rect 16632 9120 16638 9132
rect 16776 9092 16804 9132
rect 17218 9120 17224 9172
rect 17276 9160 17282 9172
rect 17402 9160 17408 9172
rect 17276 9132 17408 9160
rect 17276 9120 17282 9132
rect 17402 9120 17408 9132
rect 17460 9160 17466 9172
rect 17460 9132 17724 9160
rect 17460 9120 17466 9132
rect 17126 9092 17132 9104
rect 16776 9064 17132 9092
rect 17126 9052 17132 9064
rect 17184 9052 17190 9104
rect 15856 8996 16160 9024
rect 13780 8984 13786 8996
rect 16132 8968 16160 8996
rect 16298 8984 16304 9036
rect 16356 9024 16362 9036
rect 16485 9027 16543 9033
rect 16485 9024 16497 9027
rect 16356 8996 16497 9024
rect 16356 8984 16362 8996
rect 16485 8993 16497 8996
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 16632 8996 16677 9024
rect 16632 8984 16638 8996
rect 17494 8984 17500 9036
rect 17552 9024 17558 9036
rect 17589 9027 17647 9033
rect 17589 9024 17601 9027
rect 17552 8996 17601 9024
rect 17552 8984 17558 8996
rect 17589 8993 17601 8996
rect 17635 8993 17647 9027
rect 17589 8987 17647 8993
rect 6880 8928 7236 8956
rect 7929 8959 7987 8965
rect 6880 8916 6886 8928
rect 7929 8925 7941 8959
rect 7975 8956 7987 8959
rect 8018 8956 8024 8968
rect 7975 8928 8024 8956
rect 7975 8925 7987 8928
rect 7929 8919 7987 8925
rect 8018 8916 8024 8928
rect 8076 8916 8082 8968
rect 9677 8959 9735 8965
rect 9677 8956 9689 8959
rect 8128 8928 9689 8956
rect 6546 8888 6552 8900
rect 6507 8860 6552 8888
rect 6546 8848 6552 8860
rect 6604 8848 6610 8900
rect 8128 8888 8156 8928
rect 9677 8925 9689 8928
rect 9723 8925 9735 8959
rect 9677 8919 9735 8925
rect 10686 8916 10692 8968
rect 10744 8956 10750 8968
rect 11701 8959 11759 8965
rect 11701 8956 11713 8959
rect 10744 8928 11713 8956
rect 10744 8916 10750 8928
rect 11701 8925 11713 8928
rect 11747 8956 11759 8959
rect 14274 8956 14280 8968
rect 11747 8928 14280 8956
rect 11747 8925 11759 8928
rect 11701 8919 11759 8925
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 15760 8959 15818 8965
rect 15028 8928 15608 8956
rect 7576 8860 8156 8888
rect 9125 8891 9183 8897
rect 7576 8832 7604 8860
rect 9125 8857 9137 8891
rect 9171 8888 9183 8891
rect 9769 8891 9827 8897
rect 9769 8888 9781 8891
rect 9171 8860 9781 8888
rect 9171 8857 9183 8860
rect 9125 8851 9183 8857
rect 9769 8857 9781 8860
rect 9815 8857 9827 8891
rect 10781 8891 10839 8897
rect 10781 8888 10793 8891
rect 9769 8851 9827 8857
rect 10152 8860 10793 8888
rect 7558 8820 7564 8832
rect 7519 8792 7564 8820
rect 7558 8780 7564 8792
rect 7616 8780 7622 8832
rect 8570 8820 8576 8832
rect 8531 8792 8576 8820
rect 8570 8780 8576 8792
rect 8628 8780 8634 8832
rect 10152 8829 10180 8860
rect 10781 8857 10793 8860
rect 10827 8857 10839 8891
rect 10781 8851 10839 8857
rect 12428 8891 12486 8897
rect 12428 8857 12440 8891
rect 12474 8888 12486 8891
rect 13078 8888 13084 8900
rect 12474 8860 13084 8888
rect 12474 8857 12486 8860
rect 12428 8851 12486 8857
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 10137 8823 10195 8829
rect 10137 8789 10149 8823
rect 10183 8789 10195 8823
rect 10137 8783 10195 8789
rect 10873 8823 10931 8829
rect 10873 8789 10885 8823
rect 10919 8820 10931 8823
rect 11146 8820 11152 8832
rect 10919 8792 11152 8820
rect 10919 8789 10931 8792
rect 10873 8783 10931 8789
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 12342 8780 12348 8832
rect 12400 8820 12406 8832
rect 13446 8820 13452 8832
rect 12400 8792 13452 8820
rect 12400 8780 12406 8792
rect 13446 8780 13452 8792
rect 13504 8820 13510 8832
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 13504 8792 13553 8820
rect 13504 8780 13510 8792
rect 13541 8789 13553 8792
rect 13587 8789 13599 8823
rect 14366 8820 14372 8832
rect 14327 8792 14372 8820
rect 13541 8783 13599 8789
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 14458 8780 14464 8832
rect 14516 8820 14522 8832
rect 15028 8820 15056 8928
rect 15482 8891 15540 8897
rect 15482 8857 15494 8891
rect 15528 8857 15540 8891
rect 15580 8888 15608 8928
rect 15760 8925 15772 8959
rect 15806 8956 15818 8959
rect 15930 8956 15936 8968
rect 15806 8928 15936 8956
rect 15806 8925 15818 8928
rect 15760 8919 15818 8925
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 16114 8916 16120 8968
rect 16172 8916 16178 8968
rect 16666 8916 16672 8968
rect 16724 8956 16730 8968
rect 16942 8956 16948 8968
rect 16724 8928 16948 8956
rect 16724 8916 16730 8928
rect 16942 8916 16948 8928
rect 17000 8916 17006 8968
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 17405 8959 17463 8965
rect 17405 8956 17417 8959
rect 17368 8928 17417 8956
rect 17368 8916 17374 8928
rect 17405 8925 17417 8928
rect 17451 8925 17463 8959
rect 17405 8919 17463 8925
rect 15580 8860 16528 8888
rect 15482 8851 15540 8857
rect 14516 8792 15056 8820
rect 15497 8820 15525 8851
rect 15838 8820 15844 8832
rect 15497 8792 15844 8820
rect 14516 8780 14522 8792
rect 15838 8780 15844 8792
rect 15896 8780 15902 8832
rect 16022 8780 16028 8832
rect 16080 8820 16086 8832
rect 16393 8823 16451 8829
rect 16393 8820 16405 8823
rect 16080 8792 16405 8820
rect 16080 8780 16086 8792
rect 16393 8789 16405 8792
rect 16439 8789 16451 8823
rect 16500 8820 16528 8860
rect 16850 8848 16856 8900
rect 16908 8888 16914 8900
rect 17218 8888 17224 8900
rect 16908 8860 17224 8888
rect 16908 8848 16914 8860
rect 17218 8848 17224 8860
rect 17276 8848 17282 8900
rect 17497 8891 17555 8897
rect 17497 8857 17509 8891
rect 17543 8888 17555 8891
rect 17696 8888 17724 9132
rect 18046 9120 18052 9172
rect 18104 9160 18110 9172
rect 18506 9160 18512 9172
rect 18104 9132 18512 9160
rect 18104 9120 18110 9132
rect 18506 9120 18512 9132
rect 18564 9120 18570 9172
rect 20254 9160 20260 9172
rect 20215 9132 20260 9160
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 20346 9120 20352 9172
rect 20404 9160 20410 9172
rect 21269 9163 21327 9169
rect 21269 9160 21281 9163
rect 20404 9132 21281 9160
rect 20404 9120 20410 9132
rect 21269 9129 21281 9132
rect 21315 9129 21327 9163
rect 21269 9123 21327 9129
rect 19150 9052 19156 9104
rect 19208 9092 19214 9104
rect 19426 9092 19432 9104
rect 19208 9064 19432 9092
rect 19208 9052 19214 9064
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 19518 9052 19524 9104
rect 19576 9092 19582 9104
rect 19576 9064 19932 9092
rect 19576 9052 19582 9064
rect 18230 9024 18236 9036
rect 18143 8996 18236 9024
rect 18230 8984 18236 8996
rect 18288 9024 18294 9036
rect 19797 9027 19855 9033
rect 19797 9024 19809 9027
rect 18288 8996 19809 9024
rect 18288 8984 18294 8996
rect 19797 8993 19809 8996
rect 19843 8993 19855 9027
rect 19904 9024 19932 9064
rect 20809 9027 20867 9033
rect 20809 9024 20821 9027
rect 19904 8996 20821 9024
rect 19797 8987 19855 8993
rect 20809 8993 20821 8996
rect 20855 8993 20867 9027
rect 20809 8987 20867 8993
rect 17862 8916 17868 8968
rect 17920 8956 17926 8968
rect 18417 8959 18475 8965
rect 18417 8956 18429 8959
rect 17920 8928 18429 8956
rect 17920 8916 17926 8928
rect 18417 8925 18429 8928
rect 18463 8925 18475 8959
rect 18417 8919 18475 8925
rect 19426 8916 19432 8968
rect 19484 8956 19490 8968
rect 20162 8956 20168 8968
rect 19484 8928 20168 8956
rect 19484 8916 19490 8928
rect 20162 8916 20168 8928
rect 20220 8956 20226 8968
rect 20625 8959 20683 8965
rect 20625 8956 20637 8959
rect 20220 8928 20637 8956
rect 20220 8916 20226 8928
rect 20625 8925 20637 8928
rect 20671 8925 20683 8959
rect 20625 8919 20683 8925
rect 18322 8888 18328 8900
rect 17543 8860 17724 8888
rect 18283 8860 18328 8888
rect 17543 8857 17555 8860
rect 17497 8851 17555 8857
rect 18322 8848 18328 8860
rect 18380 8888 18386 8900
rect 18690 8888 18696 8900
rect 18380 8860 18696 8888
rect 18380 8848 18386 8860
rect 18690 8848 18696 8860
rect 18748 8848 18754 8900
rect 18966 8848 18972 8900
rect 19024 8888 19030 8900
rect 20717 8891 20775 8897
rect 20717 8888 20729 8891
rect 19024 8860 20729 8888
rect 19024 8848 19030 8860
rect 20717 8857 20729 8860
rect 20763 8888 20775 8891
rect 21358 8888 21364 8900
rect 20763 8860 21364 8888
rect 20763 8857 20775 8860
rect 20717 8851 20775 8857
rect 21358 8848 21364 8860
rect 21416 8848 21422 8900
rect 17037 8823 17095 8829
rect 17037 8820 17049 8823
rect 16500 8792 17049 8820
rect 16393 8783 16451 8789
rect 17037 8789 17049 8792
rect 17083 8789 17095 8823
rect 18782 8820 18788 8832
rect 18743 8792 18788 8820
rect 17037 8783 17095 8789
rect 18782 8780 18788 8792
rect 18840 8780 18846 8832
rect 18874 8780 18880 8832
rect 18932 8820 18938 8832
rect 19245 8823 19303 8829
rect 19245 8820 19257 8823
rect 18932 8792 19257 8820
rect 18932 8780 18938 8792
rect 19245 8789 19257 8792
rect 19291 8789 19303 8823
rect 19610 8820 19616 8832
rect 19571 8792 19616 8820
rect 19245 8783 19303 8789
rect 19610 8780 19616 8792
rect 19668 8780 19674 8832
rect 19705 8823 19763 8829
rect 19705 8789 19717 8823
rect 19751 8820 19763 8823
rect 19794 8820 19800 8832
rect 19751 8792 19800 8820
rect 19751 8789 19763 8792
rect 19705 8783 19763 8789
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 1104 8730 21896 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21896 8730
rect 1104 8656 21896 8678
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 8018 8616 8024 8628
rect 7515 8588 8024 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 8018 8576 8024 8588
rect 8076 8576 8082 8628
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8585 8355 8619
rect 8297 8579 8355 8585
rect 9217 8619 9275 8625
rect 9217 8585 9229 8619
rect 9263 8616 9275 8619
rect 16022 8616 16028 8628
rect 9263 8588 16028 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 7101 8483 7159 8489
rect 7101 8449 7113 8483
rect 7147 8480 7159 8483
rect 8110 8480 8116 8492
rect 7147 8452 8116 8480
rect 7147 8449 7159 8452
rect 7101 8443 7159 8449
rect 8110 8440 8116 8452
rect 8168 8440 8174 8492
rect 3326 8372 3332 8424
rect 3384 8412 3390 8424
rect 7742 8412 7748 8424
rect 3384 8384 7748 8412
rect 3384 8372 3390 8384
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 8312 8412 8340 8579
rect 16022 8576 16028 8588
rect 16080 8576 16086 8628
rect 17034 8616 17040 8628
rect 16995 8588 17040 8616
rect 17034 8576 17040 8588
rect 17092 8576 17098 8628
rect 17218 8576 17224 8628
rect 17276 8616 17282 8628
rect 18049 8619 18107 8625
rect 18049 8616 18061 8619
rect 17276 8588 18061 8616
rect 17276 8576 17282 8588
rect 18049 8585 18061 8588
rect 18095 8585 18107 8619
rect 18049 8579 18107 8585
rect 18417 8619 18475 8625
rect 18417 8585 18429 8619
rect 18463 8616 18475 8619
rect 18782 8616 18788 8628
rect 18463 8588 18788 8616
rect 18463 8585 18475 8588
rect 18417 8579 18475 8585
rect 18782 8576 18788 8588
rect 18840 8576 18846 8628
rect 21082 8576 21088 8628
rect 21140 8616 21146 8628
rect 21177 8619 21235 8625
rect 21177 8616 21189 8619
rect 21140 8588 21189 8616
rect 21140 8576 21146 8588
rect 21177 8585 21189 8588
rect 21223 8585 21235 8619
rect 21177 8579 21235 8585
rect 8570 8508 8576 8560
rect 8628 8548 8634 8560
rect 17405 8551 17463 8557
rect 17405 8548 17417 8551
rect 8628 8520 17417 8548
rect 8628 8508 8634 8520
rect 17405 8517 17417 8520
rect 17451 8517 17463 8551
rect 17405 8511 17463 8517
rect 18138 8508 18144 8560
rect 18196 8548 18202 8560
rect 20064 8551 20122 8557
rect 18196 8520 19840 8548
rect 18196 8508 18202 8520
rect 8757 8483 8815 8489
rect 8757 8449 8769 8483
rect 8803 8480 8815 8483
rect 10318 8480 10324 8492
rect 8803 8452 10324 8480
rect 8803 8449 8815 8452
rect 8757 8443 8815 8449
rect 10318 8440 10324 8452
rect 10376 8440 10382 8492
rect 10594 8440 10600 8492
rect 10652 8489 10658 8492
rect 10652 8480 10664 8489
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 10652 8452 11652 8480
rect 10652 8443 10664 8452
rect 10652 8440 10658 8443
rect 9858 8412 9864 8424
rect 8312 8384 9864 8412
rect 9858 8372 9864 8384
rect 9916 8372 9922 8424
rect 10873 8415 10931 8421
rect 10873 8381 10885 8415
rect 10919 8412 10931 8415
rect 11054 8412 11060 8424
rect 10919 8384 11060 8412
rect 10919 8381 10931 8384
rect 10873 8375 10931 8381
rect 11054 8372 11060 8384
rect 11112 8372 11118 8424
rect 11624 8421 11652 8452
rect 11716 8452 11897 8480
rect 11609 8415 11667 8421
rect 11609 8381 11621 8415
rect 11655 8381 11667 8415
rect 11609 8375 11667 8381
rect 7834 8304 7840 8356
rect 7892 8344 7898 8356
rect 8573 8347 8631 8353
rect 8573 8344 8585 8347
rect 7892 8316 8585 8344
rect 7892 8304 7898 8316
rect 8573 8313 8585 8316
rect 8619 8313 8631 8347
rect 9490 8344 9496 8356
rect 9451 8316 9496 8344
rect 8573 8307 8631 8313
rect 9490 8304 9496 8316
rect 9548 8304 9554 8356
rect 10962 8304 10968 8356
rect 11020 8344 11026 8356
rect 11716 8344 11744 8452
rect 11885 8449 11897 8452
rect 11931 8480 11943 8483
rect 11974 8480 11980 8492
rect 11931 8452 11980 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 11974 8440 11980 8452
rect 12032 8440 12038 8492
rect 12158 8440 12164 8492
rect 12216 8480 12222 8492
rect 12529 8483 12587 8489
rect 12529 8480 12541 8483
rect 12216 8452 12541 8480
rect 12216 8440 12222 8452
rect 12529 8449 12541 8452
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 12618 8440 12624 8492
rect 12676 8480 12682 8492
rect 12785 8483 12843 8489
rect 12785 8480 12797 8483
rect 12676 8452 12797 8480
rect 12676 8440 12682 8452
rect 12785 8449 12797 8452
rect 12831 8449 12843 8483
rect 12785 8443 12843 8449
rect 13538 8440 13544 8492
rect 13596 8480 13602 8492
rect 14366 8484 14372 8492
rect 14292 8480 14372 8484
rect 13596 8456 14372 8480
rect 13596 8452 14320 8456
rect 13596 8440 13602 8452
rect 14366 8440 14372 8456
rect 14424 8480 14430 8492
rect 15177 8483 15235 8489
rect 15177 8480 15189 8483
rect 14424 8452 14469 8480
rect 14568 8452 15189 8480
rect 14424 8440 14430 8452
rect 11793 8415 11851 8421
rect 11793 8381 11805 8415
rect 11839 8412 11851 8415
rect 12066 8412 12072 8424
rect 11839 8384 12072 8412
rect 11839 8381 11851 8384
rect 11793 8375 11851 8381
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 14568 8412 14596 8452
rect 15177 8449 15189 8452
rect 15223 8449 15235 8483
rect 15177 8443 15235 8449
rect 15930 8440 15936 8492
rect 15988 8480 15994 8492
rect 16666 8480 16672 8492
rect 15988 8452 16672 8480
rect 15988 8440 15994 8452
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 16761 8483 16819 8489
rect 16761 8449 16773 8483
rect 16807 8480 16819 8483
rect 17126 8480 17132 8492
rect 16807 8452 17132 8480
rect 16807 8449 16819 8452
rect 16761 8443 16819 8449
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 17497 8483 17555 8489
rect 17497 8449 17509 8483
rect 17543 8449 17555 8483
rect 17497 8443 17555 8449
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8480 18567 8483
rect 18874 8480 18880 8492
rect 18555 8452 18880 8480
rect 18555 8449 18567 8452
rect 18509 8443 18567 8449
rect 14918 8412 14924 8424
rect 13556 8384 14596 8412
rect 14879 8384 14924 8412
rect 11020 8316 11744 8344
rect 11020 8304 11026 8316
rect 11882 8304 11888 8356
rect 11940 8344 11946 8356
rect 12253 8347 12311 8353
rect 12253 8344 12265 8347
rect 11940 8316 12265 8344
rect 11940 8304 11946 8316
rect 12253 8313 12265 8316
rect 12299 8313 12311 8347
rect 13556 8344 13584 8384
rect 14918 8372 14924 8384
rect 14976 8372 14982 8424
rect 16114 8372 16120 8424
rect 16172 8412 16178 8424
rect 17512 8412 17540 8443
rect 18874 8440 18880 8452
rect 18932 8440 18938 8492
rect 18966 8440 18972 8492
rect 19024 8480 19030 8492
rect 19812 8489 19840 8520
rect 20064 8517 20076 8551
rect 20110 8548 20122 8551
rect 20714 8548 20720 8560
rect 20110 8520 20720 8548
rect 20110 8517 20122 8520
rect 20064 8511 20122 8517
rect 20714 8508 20720 8520
rect 20772 8508 20778 8560
rect 19061 8483 19119 8489
rect 19061 8480 19073 8483
rect 19024 8452 19073 8480
rect 19024 8440 19030 8452
rect 19061 8449 19073 8452
rect 19107 8449 19119 8483
rect 19061 8443 19119 8449
rect 19797 8483 19855 8489
rect 19797 8449 19809 8483
rect 19843 8449 19855 8483
rect 19797 8443 19855 8449
rect 16172 8384 17540 8412
rect 17589 8415 17647 8421
rect 16172 8372 16178 8384
rect 17589 8381 17601 8415
rect 17635 8412 17647 8415
rect 18601 8415 18659 8421
rect 18601 8412 18613 8415
rect 17635 8384 18613 8412
rect 17635 8381 17647 8384
rect 17589 8375 17647 8381
rect 18601 8381 18613 8384
rect 18647 8381 18659 8415
rect 18601 8375 18659 8381
rect 12253 8307 12311 8313
rect 13464 8316 13584 8344
rect 6733 8279 6791 8285
rect 6733 8245 6745 8279
rect 6779 8276 6791 8279
rect 7282 8276 7288 8288
rect 6779 8248 7288 8276
rect 6779 8245 6791 8248
rect 6733 8239 6791 8245
rect 7282 8236 7288 8248
rect 7340 8236 7346 8288
rect 9582 8236 9588 8288
rect 9640 8276 9646 8288
rect 13464 8276 13492 8316
rect 13722 8304 13728 8356
rect 13780 8344 13786 8356
rect 13909 8347 13967 8353
rect 13909 8344 13921 8347
rect 13780 8316 13921 8344
rect 13780 8304 13786 8316
rect 13909 8313 13921 8316
rect 13955 8313 13967 8347
rect 13909 8307 13967 8313
rect 13998 8304 14004 8356
rect 14056 8344 14062 8356
rect 14056 8316 14228 8344
rect 14056 8304 14062 8316
rect 14200 8285 14228 8316
rect 15930 8304 15936 8356
rect 15988 8344 15994 8356
rect 16301 8347 16359 8353
rect 16301 8344 16313 8347
rect 15988 8316 16313 8344
rect 15988 8304 15994 8316
rect 16301 8313 16313 8316
rect 16347 8344 16359 8347
rect 17494 8344 17500 8356
rect 16347 8316 17500 8344
rect 16347 8313 16359 8316
rect 16301 8307 16359 8313
rect 17494 8304 17500 8316
rect 17552 8304 17558 8356
rect 17604 8344 17632 8375
rect 17678 8344 17684 8356
rect 17604 8316 17684 8344
rect 17678 8304 17684 8316
rect 17736 8304 17742 8356
rect 19150 8344 19156 8356
rect 17788 8316 19156 8344
rect 9640 8248 13492 8276
rect 14185 8279 14243 8285
rect 9640 8236 9646 8248
rect 14185 8245 14197 8279
rect 14231 8245 14243 8279
rect 14185 8239 14243 8245
rect 16114 8236 16120 8288
rect 16172 8276 16178 8288
rect 17788 8276 17816 8316
rect 19150 8304 19156 8316
rect 19208 8304 19214 8356
rect 16172 8248 17816 8276
rect 16172 8236 16178 8248
rect 18414 8236 18420 8288
rect 18472 8276 18478 8288
rect 18874 8276 18880 8288
rect 18472 8248 18880 8276
rect 18472 8236 18478 8248
rect 18874 8236 18880 8248
rect 18932 8236 18938 8288
rect 18966 8236 18972 8288
rect 19024 8276 19030 8288
rect 19245 8279 19303 8285
rect 19245 8276 19257 8279
rect 19024 8248 19257 8276
rect 19024 8236 19030 8248
rect 19245 8245 19257 8248
rect 19291 8245 19303 8279
rect 19245 8239 19303 8245
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 7006 8032 7012 8084
rect 7064 8072 7070 8084
rect 9493 8075 9551 8081
rect 7064 8044 7328 8072
rect 7064 8032 7070 8044
rect 7300 7945 7328 8044
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9582 8072 9588 8084
rect 9539 8044 9588 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 9766 8032 9772 8084
rect 9824 8072 9830 8084
rect 13630 8072 13636 8084
rect 9824 8044 13492 8072
rect 13591 8044 13636 8072
rect 9824 8032 9830 8044
rect 9950 7964 9956 8016
rect 10008 8004 10014 8016
rect 10502 8004 10508 8016
rect 10008 7976 10508 8004
rect 10008 7964 10014 7976
rect 10502 7964 10508 7976
rect 10560 7964 10566 8016
rect 10594 7964 10600 8016
rect 10652 8004 10658 8016
rect 13464 8004 13492 8044
rect 13630 8032 13636 8044
rect 13688 8032 13694 8084
rect 14826 8072 14832 8084
rect 14787 8044 14832 8072
rect 14826 8032 14832 8044
rect 14884 8032 14890 8084
rect 15378 8032 15384 8084
rect 15436 8072 15442 8084
rect 16114 8072 16120 8084
rect 15436 8044 16120 8072
rect 15436 8032 15442 8044
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 16666 8032 16672 8084
rect 16724 8072 16730 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16724 8044 16957 8072
rect 16724 8032 16730 8044
rect 16945 8041 16957 8044
rect 16991 8072 17003 8075
rect 18138 8072 18144 8084
rect 16991 8044 18144 8072
rect 16991 8041 17003 8044
rect 16945 8035 17003 8041
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 18877 8075 18935 8081
rect 18877 8041 18889 8075
rect 18923 8072 18935 8075
rect 19978 8072 19984 8084
rect 18923 8044 19984 8072
rect 18923 8041 18935 8044
rect 18877 8035 18935 8041
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 20622 8032 20628 8084
rect 20680 8072 20686 8084
rect 21269 8075 21327 8081
rect 21269 8072 21281 8075
rect 20680 8044 21281 8072
rect 20680 8032 20686 8044
rect 21269 8041 21281 8044
rect 21315 8041 21327 8075
rect 21269 8035 21327 8041
rect 14734 8004 14740 8016
rect 10652 7976 13032 8004
rect 13464 7976 14740 8004
rect 10652 7964 10658 7976
rect 7285 7939 7343 7945
rect 7285 7905 7297 7939
rect 7331 7936 7343 7939
rect 8478 7936 8484 7948
rect 7331 7908 8484 7936
rect 7331 7905 7343 7908
rect 7285 7899 7343 7905
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 13004 7945 13032 7976
rect 14734 7964 14740 7976
rect 14792 7964 14798 8016
rect 18506 7964 18512 8016
rect 18564 8004 18570 8016
rect 18966 8004 18972 8016
rect 18564 7976 18972 8004
rect 18564 7964 18570 7976
rect 18966 7964 18972 7976
rect 19024 7964 19030 8016
rect 19337 8007 19395 8013
rect 19337 7973 19349 8007
rect 19383 8004 19395 8007
rect 19518 8004 19524 8016
rect 19383 7976 19524 8004
rect 19383 7973 19395 7976
rect 19337 7967 19395 7973
rect 19518 7964 19524 7976
rect 19576 7964 19582 8016
rect 8573 7939 8631 7945
rect 8573 7905 8585 7939
rect 8619 7936 8631 7939
rect 12989 7939 13047 7945
rect 8619 7908 12940 7936
rect 8619 7905 8631 7908
rect 8573 7899 8631 7905
rect 6546 7868 6552 7880
rect 6507 7840 6552 7868
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 7558 7868 7564 7880
rect 7519 7840 7564 7868
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 10137 7871 10195 7877
rect 10137 7837 10149 7871
rect 10183 7868 10195 7871
rect 12710 7868 12716 7880
rect 10183 7840 12716 7868
rect 10183 7837 10195 7840
rect 10137 7831 10195 7837
rect 12710 7828 12716 7840
rect 12768 7828 12774 7880
rect 12912 7868 12940 7908
rect 12989 7905 13001 7939
rect 13035 7905 13047 7939
rect 12989 7899 13047 7905
rect 13078 7896 13084 7948
rect 13136 7936 13142 7948
rect 14277 7939 14335 7945
rect 14277 7936 14289 7939
rect 13136 7908 14289 7936
rect 13136 7896 13142 7908
rect 14277 7905 14289 7908
rect 14323 7905 14335 7939
rect 14277 7899 14335 7905
rect 14369 7939 14427 7945
rect 14369 7905 14381 7939
rect 14415 7936 14427 7939
rect 14458 7936 14464 7948
rect 14415 7908 14464 7936
rect 14415 7905 14427 7908
rect 14369 7899 14427 7905
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 17954 7936 17960 7948
rect 14936 7908 17960 7936
rect 13449 7871 13507 7877
rect 13449 7868 13461 7871
rect 12912 7840 13461 7868
rect 13449 7837 13461 7840
rect 13495 7868 13507 7871
rect 14936 7868 14964 7908
rect 17954 7896 17960 7908
rect 18012 7896 18018 7948
rect 18325 7939 18383 7945
rect 18325 7905 18337 7939
rect 18371 7936 18383 7939
rect 18414 7936 18420 7948
rect 18371 7908 18420 7936
rect 18371 7905 18383 7908
rect 18325 7899 18383 7905
rect 18414 7896 18420 7908
rect 18472 7896 18478 7948
rect 15102 7868 15108 7880
rect 13495 7840 14964 7868
rect 15063 7840 15108 7868
rect 13495 7837 13507 7840
rect 13449 7831 13507 7837
rect 15102 7828 15108 7840
rect 15160 7828 15166 7880
rect 15286 7828 15292 7880
rect 15344 7868 15350 7880
rect 15344 7840 15792 7868
rect 15344 7828 15350 7840
rect 6181 7803 6239 7809
rect 6181 7769 6193 7803
rect 6227 7800 6239 7803
rect 7834 7800 7840 7812
rect 6227 7772 7840 7800
rect 6227 7769 6239 7772
rect 6181 7763 6239 7769
rect 7834 7760 7840 7772
rect 7892 7760 7898 7812
rect 8938 7760 8944 7812
rect 8996 7800 9002 7812
rect 10413 7803 10471 7809
rect 10413 7800 10425 7803
rect 8996 7772 10425 7800
rect 8996 7760 9002 7772
rect 10413 7769 10425 7772
rect 10459 7800 10471 7803
rect 11054 7800 11060 7812
rect 10459 7772 11060 7800
rect 10459 7769 10471 7772
rect 10413 7763 10471 7769
rect 11054 7760 11060 7772
rect 11112 7760 11118 7812
rect 12158 7800 12164 7812
rect 12119 7772 12164 7800
rect 12158 7760 12164 7772
rect 12216 7760 12222 7812
rect 12802 7800 12808 7812
rect 12763 7772 12808 7800
rect 12802 7760 12808 7772
rect 12860 7760 12866 7812
rect 13722 7760 13728 7812
rect 13780 7800 13786 7812
rect 14182 7800 14188 7812
rect 13780 7772 14188 7800
rect 13780 7760 13786 7772
rect 14182 7760 14188 7772
rect 14240 7760 14246 7812
rect 14461 7803 14519 7809
rect 14461 7769 14473 7803
rect 14507 7800 14519 7803
rect 15194 7800 15200 7812
rect 14507 7772 15200 7800
rect 14507 7769 14519 7772
rect 14461 7763 14519 7769
rect 15194 7760 15200 7772
rect 15252 7760 15258 7812
rect 15654 7800 15660 7812
rect 15615 7772 15660 7800
rect 15654 7760 15660 7772
rect 15712 7760 15718 7812
rect 15764 7800 15792 7840
rect 17770 7828 17776 7880
rect 17828 7868 17834 7880
rect 18693 7871 18751 7877
rect 18693 7868 18705 7871
rect 17828 7840 18705 7868
rect 17828 7828 17834 7840
rect 18693 7837 18705 7840
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 19518 7828 19524 7880
rect 19576 7868 19582 7880
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 19576 7840 19625 7868
rect 19576 7828 19582 7840
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 19702 7828 19708 7880
rect 19760 7868 19766 7880
rect 19869 7871 19927 7877
rect 19869 7868 19881 7871
rect 19760 7840 19881 7868
rect 19760 7828 19766 7840
rect 19869 7837 19881 7840
rect 19915 7837 19927 7871
rect 19869 7831 19927 7837
rect 20162 7800 20168 7812
rect 15764 7772 20168 7800
rect 20162 7760 20168 7772
rect 20220 7760 20226 7812
rect 6917 7735 6975 7741
rect 6917 7701 6929 7735
rect 6963 7732 6975 7735
rect 7098 7732 7104 7744
rect 6963 7704 7104 7732
rect 6963 7701 6975 7704
rect 6917 7695 6975 7701
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 8202 7732 8208 7744
rect 8163 7704 8208 7732
rect 8202 7692 8208 7704
rect 8260 7692 8266 7744
rect 9217 7735 9275 7741
rect 9217 7701 9229 7735
rect 9263 7732 9275 7735
rect 10134 7732 10140 7744
rect 9263 7704 10140 7732
rect 9263 7701 9275 7704
rect 9217 7695 9275 7701
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 12437 7735 12495 7741
rect 12437 7701 12449 7735
rect 12483 7732 12495 7735
rect 12526 7732 12532 7744
rect 12483 7704 12532 7732
rect 12483 7701 12495 7704
rect 12437 7695 12495 7701
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 12897 7735 12955 7741
rect 12897 7701 12909 7735
rect 12943 7732 12955 7735
rect 12986 7732 12992 7744
rect 12943 7704 12992 7732
rect 12943 7701 12955 7704
rect 12897 7695 12955 7701
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 15289 7735 15347 7741
rect 15289 7701 15301 7735
rect 15335 7732 15347 7735
rect 16390 7732 16396 7744
rect 15335 7704 16396 7732
rect 15335 7701 15347 7704
rect 15289 7695 15347 7701
rect 16390 7692 16396 7704
rect 16448 7692 16454 7744
rect 17034 7692 17040 7744
rect 17092 7732 17098 7744
rect 17681 7735 17739 7741
rect 17681 7732 17693 7735
rect 17092 7704 17693 7732
rect 17092 7692 17098 7704
rect 17681 7701 17693 7704
rect 17727 7701 17739 7735
rect 18046 7732 18052 7744
rect 18007 7704 18052 7732
rect 17681 7695 17739 7701
rect 18046 7692 18052 7704
rect 18104 7692 18110 7744
rect 18141 7735 18199 7741
rect 18141 7701 18153 7735
rect 18187 7732 18199 7735
rect 18782 7732 18788 7744
rect 18187 7704 18788 7732
rect 18187 7701 18199 7704
rect 18141 7695 18199 7701
rect 18782 7692 18788 7704
rect 18840 7692 18846 7744
rect 20714 7692 20720 7744
rect 20772 7732 20778 7744
rect 20993 7735 21051 7741
rect 20993 7732 21005 7735
rect 20772 7704 21005 7732
rect 20772 7692 20778 7704
rect 20993 7701 21005 7704
rect 21039 7701 21051 7735
rect 20993 7695 21051 7701
rect 1104 7642 21896 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21896 7642
rect 1104 7568 21896 7590
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 5500 7500 6561 7528
rect 5500 7488 5506 7500
rect 6549 7497 6561 7500
rect 6595 7497 6607 7531
rect 6549 7491 6607 7497
rect 7742 7488 7748 7540
rect 7800 7528 7806 7540
rect 10321 7531 10379 7537
rect 7800 7500 9674 7528
rect 7800 7488 7806 7500
rect 8202 7420 8208 7472
rect 8260 7460 8266 7472
rect 9186 7463 9244 7469
rect 9186 7460 9198 7463
rect 8260 7432 9198 7460
rect 8260 7420 8266 7432
rect 9186 7429 9198 7432
rect 9232 7429 9244 7463
rect 9646 7460 9674 7500
rect 10321 7497 10333 7531
rect 10367 7528 10379 7531
rect 10594 7528 10600 7540
rect 10367 7500 10600 7528
rect 10367 7497 10379 7500
rect 10321 7491 10379 7497
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 10686 7488 10692 7540
rect 10744 7528 10750 7540
rect 11149 7531 11207 7537
rect 10744 7500 10789 7528
rect 10744 7488 10750 7500
rect 11149 7497 11161 7531
rect 11195 7528 11207 7531
rect 11238 7528 11244 7540
rect 11195 7500 11244 7528
rect 11195 7497 11207 7500
rect 11149 7491 11207 7497
rect 11238 7488 11244 7500
rect 11296 7488 11302 7540
rect 11517 7531 11575 7537
rect 11517 7497 11529 7531
rect 11563 7528 11575 7531
rect 12618 7528 12624 7540
rect 11563 7500 12624 7528
rect 11563 7497 11575 7500
rect 11517 7491 11575 7497
rect 12618 7488 12624 7500
rect 12676 7488 12682 7540
rect 13630 7488 13636 7540
rect 13688 7528 13694 7540
rect 13909 7531 13967 7537
rect 13909 7528 13921 7531
rect 13688 7500 13921 7528
rect 13688 7488 13694 7500
rect 13909 7497 13921 7500
rect 13955 7497 13967 7531
rect 13909 7491 13967 7497
rect 14001 7531 14059 7537
rect 14001 7497 14013 7531
rect 14047 7497 14059 7531
rect 14001 7491 14059 7497
rect 14553 7531 14611 7537
rect 14553 7497 14565 7531
rect 14599 7528 14611 7531
rect 15010 7528 15016 7540
rect 14599 7500 15016 7528
rect 14599 7497 14611 7500
rect 14553 7491 14611 7497
rect 14016 7460 14044 7491
rect 15010 7488 15016 7500
rect 15068 7488 15074 7540
rect 16206 7488 16212 7540
rect 16264 7528 16270 7540
rect 17129 7531 17187 7537
rect 17129 7528 17141 7531
rect 16264 7500 17141 7528
rect 16264 7488 16270 7500
rect 17129 7497 17141 7500
rect 17175 7528 17187 7531
rect 18414 7528 18420 7540
rect 17175 7500 18420 7528
rect 17175 7497 17187 7500
rect 17129 7491 17187 7497
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 18782 7528 18788 7540
rect 18743 7500 18788 7528
rect 18782 7488 18788 7500
rect 18840 7488 18846 7540
rect 19058 7488 19064 7540
rect 19116 7528 19122 7540
rect 19245 7531 19303 7537
rect 19245 7528 19257 7531
rect 19116 7500 19257 7528
rect 19116 7488 19122 7500
rect 19245 7497 19257 7500
rect 19291 7497 19303 7531
rect 20162 7528 20168 7540
rect 20123 7500 20168 7528
rect 19245 7491 19303 7497
rect 20162 7488 20168 7500
rect 20220 7488 20226 7540
rect 14642 7460 14648 7472
rect 9646 7432 14648 7460
rect 9186 7423 9244 7429
rect 14642 7420 14648 7432
rect 14700 7420 14706 7472
rect 14918 7420 14924 7472
rect 14976 7460 14982 7472
rect 14976 7432 18552 7460
rect 14976 7420 14982 7432
rect 8386 7352 8392 7404
rect 8444 7401 8450 7404
rect 8444 7392 8456 7401
rect 8665 7395 8723 7401
rect 8444 7364 8489 7392
rect 8444 7355 8456 7364
rect 8665 7361 8677 7395
rect 8711 7392 8723 7395
rect 8938 7392 8944 7404
rect 8711 7364 8944 7392
rect 8711 7361 8723 7364
rect 8665 7355 8723 7361
rect 8444 7352 8450 7355
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 10962 7392 10968 7404
rect 10923 7364 10968 7392
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 12161 7395 12219 7401
rect 12161 7361 12173 7395
rect 12207 7392 12219 7395
rect 12342 7392 12348 7404
rect 12207 7364 12348 7392
rect 12207 7361 12219 7364
rect 12161 7355 12219 7361
rect 12342 7352 12348 7364
rect 12400 7352 12406 7404
rect 12805 7395 12863 7401
rect 12805 7361 12817 7395
rect 12851 7392 12863 7395
rect 15102 7392 15108 7404
rect 12851 7364 15108 7392
rect 12851 7361 12863 7364
rect 12805 7355 12863 7361
rect 15102 7352 15108 7364
rect 15160 7352 15166 7404
rect 16045 7395 16103 7401
rect 16045 7361 16057 7395
rect 16091 7392 16103 7395
rect 16206 7392 16212 7404
rect 16091 7364 16212 7392
rect 16091 7361 16103 7364
rect 16045 7355 16103 7361
rect 16206 7352 16212 7364
rect 16264 7352 16270 7404
rect 16316 7401 16344 7432
rect 16301 7395 16359 7401
rect 16301 7361 16313 7395
rect 16347 7361 16359 7395
rect 16301 7355 16359 7361
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7392 16911 7395
rect 16942 7392 16948 7404
rect 16899 7364 16948 7392
rect 16899 7361 16911 7364
rect 16853 7355 16911 7361
rect 16942 7352 16948 7364
rect 17000 7352 17006 7404
rect 18524 7401 18552 7432
rect 18690 7420 18696 7472
rect 18748 7460 18754 7472
rect 20257 7463 20315 7469
rect 20257 7460 20269 7463
rect 18748 7432 20269 7460
rect 18748 7420 18754 7432
rect 20257 7429 20269 7432
rect 20303 7429 20315 7463
rect 20257 7423 20315 7429
rect 20990 7420 20996 7472
rect 21048 7460 21054 7472
rect 21177 7463 21235 7469
rect 21177 7460 21189 7463
rect 21048 7432 21189 7460
rect 21048 7420 21054 7432
rect 21177 7429 21189 7432
rect 21223 7460 21235 7463
rect 22002 7460 22008 7472
rect 21223 7432 22008 7460
rect 21223 7429 21235 7432
rect 21177 7423 21235 7429
rect 22002 7420 22008 7432
rect 22060 7420 22066 7472
rect 18253 7395 18311 7401
rect 18253 7361 18265 7395
rect 18299 7392 18311 7395
rect 18509 7395 18567 7401
rect 18299 7364 18460 7392
rect 18299 7361 18311 7364
rect 18253 7355 18311 7361
rect 12894 7324 12900 7336
rect 12855 7296 12900 7324
rect 12894 7284 12900 7296
rect 12952 7284 12958 7336
rect 12989 7327 13047 7333
rect 12989 7293 13001 7327
rect 13035 7293 13047 7327
rect 14182 7324 14188 7336
rect 14095 7296 14188 7324
rect 12989 7287 13047 7293
rect 4890 7216 4896 7268
rect 4948 7256 4954 7268
rect 6917 7259 6975 7265
rect 6917 7256 6929 7259
rect 4948 7228 6929 7256
rect 4948 7216 4954 7228
rect 6917 7225 6929 7228
rect 6963 7256 6975 7259
rect 7374 7256 7380 7268
rect 6963 7228 7380 7256
rect 6963 7225 6975 7228
rect 6917 7219 6975 7225
rect 7374 7216 7380 7228
rect 7432 7216 7438 7268
rect 11330 7216 11336 7268
rect 11388 7256 11394 7268
rect 13004 7256 13032 7287
rect 14182 7284 14188 7296
rect 14240 7324 14246 7336
rect 14826 7324 14832 7336
rect 14240 7296 14832 7324
rect 14240 7284 14246 7296
rect 14826 7284 14832 7296
rect 14884 7284 14890 7336
rect 18432 7324 18460 7364
rect 18509 7361 18521 7395
rect 18555 7361 18567 7395
rect 19150 7392 19156 7404
rect 19111 7364 19156 7392
rect 18509 7355 18567 7361
rect 19150 7352 19156 7364
rect 19208 7352 19214 7404
rect 19337 7327 19395 7333
rect 18432 7296 18552 7324
rect 18524 7268 18552 7296
rect 19337 7293 19349 7327
rect 19383 7293 19395 7327
rect 19337 7287 19395 7293
rect 20349 7327 20407 7333
rect 20349 7293 20361 7327
rect 20395 7293 20407 7327
rect 20349 7287 20407 7293
rect 14921 7259 14979 7265
rect 14921 7256 14933 7259
rect 11388 7228 13032 7256
rect 13280 7228 14933 7256
rect 11388 7216 11394 7228
rect 5258 7188 5264 7200
rect 5219 7160 5264 7188
rect 5258 7148 5264 7160
rect 5316 7148 5322 7200
rect 5350 7148 5356 7200
rect 5408 7188 5414 7200
rect 5537 7191 5595 7197
rect 5537 7188 5549 7191
rect 5408 7160 5549 7188
rect 5408 7148 5414 7160
rect 5537 7157 5549 7160
rect 5583 7157 5595 7191
rect 5902 7188 5908 7200
rect 5863 7160 5908 7188
rect 5537 7151 5595 7157
rect 5902 7148 5908 7160
rect 5960 7148 5966 7200
rect 7285 7191 7343 7197
rect 7285 7157 7297 7191
rect 7331 7188 7343 7191
rect 7558 7188 7564 7200
rect 7331 7160 7564 7188
rect 7331 7157 7343 7160
rect 7285 7151 7343 7157
rect 7558 7148 7564 7160
rect 7616 7188 7622 7200
rect 9674 7188 9680 7200
rect 7616 7160 9680 7188
rect 7616 7148 7622 7160
rect 9674 7148 9680 7160
rect 9732 7148 9738 7200
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 12342 7188 12348 7200
rect 11112 7160 12348 7188
rect 11112 7148 11118 7160
rect 12342 7148 12348 7160
rect 12400 7148 12406 7200
rect 12434 7148 12440 7200
rect 12492 7188 12498 7200
rect 12492 7160 12537 7188
rect 12492 7148 12498 7160
rect 12710 7148 12716 7200
rect 12768 7188 12774 7200
rect 13280 7188 13308 7228
rect 14921 7225 14933 7228
rect 14967 7225 14979 7259
rect 14921 7219 14979 7225
rect 12768 7160 13308 7188
rect 12768 7148 12774 7160
rect 13354 7148 13360 7200
rect 13412 7188 13418 7200
rect 13541 7191 13599 7197
rect 13541 7188 13553 7191
rect 13412 7160 13553 7188
rect 13412 7148 13418 7160
rect 13541 7157 13553 7160
rect 13587 7157 13599 7191
rect 14936 7188 14964 7219
rect 18506 7216 18512 7268
rect 18564 7256 18570 7268
rect 19352 7256 19380 7287
rect 20364 7256 20392 7287
rect 18564 7228 20392 7256
rect 21361 7259 21419 7265
rect 18564 7216 18570 7228
rect 21361 7225 21373 7259
rect 21407 7256 21419 7259
rect 21542 7256 21548 7268
rect 21407 7228 21548 7256
rect 21407 7225 21419 7228
rect 21361 7219 21419 7225
rect 21542 7216 21548 7228
rect 21600 7256 21606 7268
rect 22278 7256 22284 7268
rect 21600 7228 22284 7256
rect 21600 7216 21606 7228
rect 22278 7216 22284 7228
rect 22336 7216 22342 7268
rect 16574 7188 16580 7200
rect 14936 7160 16580 7188
rect 13541 7151 13599 7157
rect 16574 7148 16580 7160
rect 16632 7148 16638 7200
rect 16669 7191 16727 7197
rect 16669 7157 16681 7191
rect 16715 7188 16727 7191
rect 17586 7188 17592 7200
rect 16715 7160 17592 7188
rect 16715 7157 16727 7160
rect 16669 7151 16727 7157
rect 17586 7148 17592 7160
rect 17644 7148 17650 7200
rect 18322 7148 18328 7200
rect 18380 7188 18386 7200
rect 19797 7191 19855 7197
rect 19797 7188 19809 7191
rect 18380 7160 19809 7188
rect 18380 7148 18386 7160
rect 19797 7157 19809 7160
rect 19843 7157 19855 7191
rect 19797 7151 19855 7157
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 5169 6987 5227 6993
rect 5169 6953 5181 6987
rect 5215 6984 5227 6987
rect 12342 6984 12348 6996
rect 5215 6956 12348 6984
rect 5215 6953 5227 6956
rect 5169 6947 5227 6953
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 12989 6987 13047 6993
rect 12989 6984 13001 6987
rect 12952 6956 13001 6984
rect 12952 6944 12958 6956
rect 12989 6953 13001 6956
rect 13035 6953 13047 6987
rect 12989 6947 13047 6953
rect 14292 6956 14964 6984
rect 8570 6916 8576 6928
rect 8531 6888 8576 6916
rect 8570 6876 8576 6888
rect 8628 6876 8634 6928
rect 9033 6919 9091 6925
rect 9033 6885 9045 6919
rect 9079 6916 9091 6919
rect 10962 6916 10968 6928
rect 9079 6888 10968 6916
rect 9079 6885 9091 6888
rect 9033 6879 9091 6885
rect 10962 6876 10968 6888
rect 11020 6876 11026 6928
rect 11330 6916 11336 6928
rect 11291 6888 11336 6916
rect 11330 6876 11336 6888
rect 11388 6876 11394 6928
rect 14292 6916 14320 6956
rect 14108 6888 14320 6916
rect 14936 6916 14964 6956
rect 15102 6944 15108 6996
rect 15160 6984 15166 6996
rect 15565 6987 15623 6993
rect 15565 6984 15577 6987
rect 15160 6956 15577 6984
rect 15160 6944 15166 6956
rect 15565 6953 15577 6956
rect 15611 6953 15623 6987
rect 15565 6947 15623 6953
rect 14936 6888 16160 6916
rect 4798 6848 4804 6860
rect 2746 6820 4804 6848
rect 1946 6740 1952 6792
rect 2004 6780 2010 6792
rect 2746 6780 2774 6820
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 5537 6851 5595 6857
rect 5537 6848 5549 6851
rect 5040 6820 5549 6848
rect 5040 6808 5046 6820
rect 5537 6817 5549 6820
rect 5583 6848 5595 6851
rect 6730 6848 6736 6860
rect 5583 6820 6736 6848
rect 5583 6817 5595 6820
rect 5537 6811 5595 6817
rect 6730 6808 6736 6820
rect 6788 6808 6794 6860
rect 6914 6848 6920 6860
rect 6875 6820 6920 6848
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 8021 6851 8079 6857
rect 8021 6817 8033 6851
rect 8067 6848 8079 6851
rect 8386 6848 8392 6860
rect 8067 6820 8392 6848
rect 8067 6817 8079 6820
rect 8021 6811 8079 6817
rect 8386 6808 8392 6820
rect 8444 6848 8450 6860
rect 9122 6848 9128 6860
rect 8444 6820 9128 6848
rect 8444 6808 8450 6820
rect 9122 6808 9128 6820
rect 9180 6848 9186 6860
rect 9401 6851 9459 6857
rect 9401 6848 9413 6851
rect 9180 6820 9413 6848
rect 9180 6808 9186 6820
rect 9401 6817 9413 6820
rect 9447 6817 9459 6851
rect 9401 6811 9459 6817
rect 9674 6808 9680 6860
rect 9732 6848 9738 6860
rect 10873 6851 10931 6857
rect 10873 6848 10885 6851
rect 9732 6820 10885 6848
rect 9732 6808 9738 6820
rect 10873 6817 10885 6820
rect 10919 6817 10931 6851
rect 10873 6811 10931 6817
rect 13078 6808 13084 6860
rect 13136 6848 13142 6860
rect 13633 6851 13691 6857
rect 13633 6848 13645 6851
rect 13136 6820 13645 6848
rect 13136 6808 13142 6820
rect 13633 6817 13645 6820
rect 13679 6848 13691 6851
rect 14108 6848 14136 6888
rect 14642 6848 14648 6860
rect 13679 6820 14136 6848
rect 14209 6820 14648 6848
rect 13679 6817 13691 6820
rect 13633 6811 13691 6817
rect 2004 6752 2774 6780
rect 2004 6740 2010 6752
rect 3050 6740 3056 6792
rect 3108 6780 3114 6792
rect 6181 6783 6239 6789
rect 6181 6780 6193 6783
rect 3108 6752 6193 6780
rect 3108 6740 3114 6752
rect 6181 6749 6193 6752
rect 6227 6780 6239 6783
rect 7466 6780 7472 6792
rect 6227 6752 7472 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 7466 6740 7472 6752
rect 7524 6740 7530 6792
rect 7561 6783 7619 6789
rect 7561 6749 7573 6783
rect 7607 6780 7619 6783
rect 7607 6752 8524 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 5905 6715 5963 6721
rect 5905 6681 5917 6715
rect 5951 6712 5963 6715
rect 6546 6712 6552 6724
rect 5951 6684 6552 6712
rect 5951 6681 5963 6684
rect 5905 6675 5963 6681
rect 6546 6672 6552 6684
rect 6604 6672 6610 6724
rect 6914 6672 6920 6724
rect 6972 6712 6978 6724
rect 7282 6712 7288 6724
rect 6972 6684 7288 6712
rect 6972 6672 6978 6684
rect 7282 6672 7288 6684
rect 7340 6672 7346 6724
rect 1302 6604 1308 6656
rect 1360 6644 1366 6656
rect 1397 6647 1455 6653
rect 1397 6644 1409 6647
rect 1360 6616 1409 6644
rect 1360 6604 1366 6616
rect 1397 6613 1409 6616
rect 1443 6613 1455 6647
rect 4154 6644 4160 6656
rect 4115 6616 4160 6644
rect 1397 6607 1455 6613
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4246 6604 4252 6656
rect 4304 6644 4310 6656
rect 5258 6644 5264 6656
rect 4304 6616 5264 6644
rect 4304 6604 4310 6616
rect 5258 6604 5264 6616
rect 5316 6644 5322 6656
rect 5810 6644 5816 6656
rect 5316 6616 5816 6644
rect 5316 6604 5322 6616
rect 5810 6604 5816 6616
rect 5868 6644 5874 6656
rect 6641 6647 6699 6653
rect 6641 6644 6653 6647
rect 5868 6616 6653 6644
rect 5868 6604 5874 6616
rect 6641 6613 6653 6616
rect 6687 6644 6699 6647
rect 6730 6644 6736 6656
rect 6687 6616 6736 6644
rect 6687 6613 6699 6616
rect 6641 6607 6699 6613
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 8110 6644 8116 6656
rect 8071 6616 8116 6644
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 8202 6604 8208 6656
rect 8260 6644 8266 6656
rect 8496 6644 8524 6752
rect 8570 6740 8576 6792
rect 8628 6780 8634 6792
rect 10689 6783 10747 6789
rect 10689 6780 10701 6783
rect 8628 6752 10701 6780
rect 8628 6740 8634 6752
rect 10689 6749 10701 6752
rect 10735 6749 10747 6783
rect 12713 6783 12771 6789
rect 12713 6780 12725 6783
rect 10689 6743 10747 6749
rect 12360 6752 12725 6780
rect 12360 6724 12388 6752
rect 12713 6749 12725 6752
rect 12759 6749 12771 6783
rect 13354 6780 13360 6792
rect 13315 6752 13360 6780
rect 12713 6743 12771 6749
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 13449 6783 13507 6789
rect 13449 6749 13461 6783
rect 13495 6780 13507 6783
rect 14209 6780 14237 6820
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 14737 6851 14795 6857
rect 14737 6817 14749 6851
rect 14783 6848 14795 6851
rect 14826 6848 14832 6860
rect 14783 6820 14832 6848
rect 14783 6817 14795 6820
rect 14737 6811 14795 6817
rect 14826 6808 14832 6820
rect 14884 6848 14890 6860
rect 16132 6857 16160 6888
rect 16574 6876 16580 6928
rect 16632 6916 16638 6928
rect 17586 6916 17592 6928
rect 16632 6888 17172 6916
rect 17547 6888 17592 6916
rect 16632 6876 16638 6888
rect 16117 6851 16175 6857
rect 14884 6820 16068 6848
rect 14884 6808 14890 6820
rect 13495 6752 14237 6780
rect 14277 6783 14335 6789
rect 13495 6749 13507 6752
rect 13449 6743 13507 6749
rect 14277 6749 14289 6783
rect 14323 6780 14335 6783
rect 15933 6783 15991 6789
rect 15933 6780 15945 6783
rect 14323 6752 15945 6780
rect 14323 6749 14335 6752
rect 14277 6743 14335 6749
rect 15933 6749 15945 6752
rect 15979 6749 15991 6783
rect 16040 6780 16068 6820
rect 16117 6817 16129 6851
rect 16163 6817 16175 6851
rect 17034 6848 17040 6860
rect 16995 6820 17040 6848
rect 16117 6811 16175 6817
rect 17034 6808 17040 6820
rect 17092 6808 17098 6860
rect 17144 6857 17172 6888
rect 17586 6876 17592 6888
rect 17644 6876 17650 6928
rect 17696 6888 18184 6916
rect 17129 6851 17187 6857
rect 17129 6817 17141 6851
rect 17175 6817 17187 6851
rect 17129 6811 17187 6817
rect 17696 6780 17724 6888
rect 17954 6808 17960 6860
rect 18012 6808 18018 6860
rect 18156 6857 18184 6888
rect 18141 6851 18199 6857
rect 18141 6817 18153 6851
rect 18187 6817 18199 6851
rect 18141 6811 18199 6817
rect 18874 6808 18880 6860
rect 18932 6848 18938 6860
rect 18932 6820 19564 6848
rect 18932 6808 18938 6820
rect 16040 6752 17724 6780
rect 15933 6743 15991 6749
rect 9585 6715 9643 6721
rect 9585 6681 9597 6715
rect 9631 6712 9643 6715
rect 9950 6712 9956 6724
rect 9631 6684 9956 6712
rect 9631 6681 9643 6684
rect 9585 6675 9643 6681
rect 9950 6672 9956 6684
rect 10008 6672 10014 6724
rect 10781 6715 10839 6721
rect 10781 6712 10793 6715
rect 10060 6684 10793 6712
rect 8570 6644 8576 6656
rect 8260 6616 8305 6644
rect 8496 6616 8576 6644
rect 8260 6604 8266 6616
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 9674 6604 9680 6656
rect 9732 6644 9738 6656
rect 10060 6653 10088 6684
rect 10781 6681 10793 6684
rect 10827 6681 10839 6715
rect 10781 6675 10839 6681
rect 11974 6672 11980 6724
rect 12032 6712 12038 6724
rect 12250 6712 12256 6724
rect 12032 6684 12256 6712
rect 12032 6672 12038 6684
rect 12250 6672 12256 6684
rect 12308 6672 12314 6724
rect 12342 6672 12348 6724
rect 12400 6672 12406 6724
rect 12468 6715 12526 6721
rect 12468 6681 12480 6715
rect 12514 6712 12526 6715
rect 13078 6712 13084 6724
rect 12514 6684 13084 6712
rect 12514 6681 12526 6684
rect 12468 6675 12526 6681
rect 13078 6672 13084 6684
rect 13136 6672 13142 6724
rect 13170 6672 13176 6724
rect 13228 6712 13234 6724
rect 14921 6715 14979 6721
rect 14921 6712 14933 6715
rect 13228 6684 14933 6712
rect 13228 6672 13234 6684
rect 14921 6681 14933 6684
rect 14967 6712 14979 6715
rect 15194 6712 15200 6724
rect 14967 6684 15200 6712
rect 14967 6681 14979 6684
rect 14921 6675 14979 6681
rect 15194 6672 15200 6684
rect 15252 6672 15258 6724
rect 16025 6715 16083 6721
rect 16025 6712 16037 6715
rect 15304 6684 16037 6712
rect 10045 6647 10103 6653
rect 9732 6616 9777 6644
rect 9732 6604 9738 6616
rect 10045 6613 10057 6647
rect 10091 6613 10103 6647
rect 10318 6644 10324 6656
rect 10279 6616 10324 6644
rect 10045 6607 10103 6613
rect 10318 6604 10324 6616
rect 10376 6604 10382 6656
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 14734 6644 14740 6656
rect 11020 6616 14740 6644
rect 11020 6604 11026 6616
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 14829 6647 14887 6653
rect 14829 6613 14841 6647
rect 14875 6644 14887 6647
rect 15010 6644 15016 6656
rect 14875 6616 15016 6644
rect 14875 6613 14887 6616
rect 14829 6607 14887 6613
rect 15010 6604 15016 6616
rect 15068 6604 15074 6656
rect 15304 6653 15332 6684
rect 16025 6681 16037 6684
rect 16071 6681 16083 6715
rect 17218 6712 17224 6724
rect 16025 6675 16083 6681
rect 16592 6684 17224 6712
rect 16592 6653 16620 6684
rect 17218 6672 17224 6684
rect 17276 6672 17282 6724
rect 17972 6721 18000 6808
rect 18598 6780 18604 6792
rect 18559 6752 18604 6780
rect 18598 6740 18604 6752
rect 18656 6740 18662 6792
rect 19426 6780 19432 6792
rect 19387 6752 19432 6780
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 19536 6780 19564 6820
rect 21085 6783 21143 6789
rect 21085 6780 21097 6783
rect 19536 6752 21097 6780
rect 21085 6749 21097 6752
rect 21131 6749 21143 6783
rect 21085 6743 21143 6749
rect 17957 6715 18015 6721
rect 17957 6681 17969 6715
rect 18003 6681 18015 6715
rect 17957 6675 18015 6681
rect 18049 6715 18107 6721
rect 18049 6681 18061 6715
rect 18095 6681 18107 6715
rect 18049 6675 18107 6681
rect 19696 6715 19754 6721
rect 19696 6681 19708 6715
rect 19742 6712 19754 6715
rect 20162 6712 20168 6724
rect 19742 6684 20168 6712
rect 19742 6681 19754 6684
rect 19696 6675 19754 6681
rect 15289 6647 15347 6653
rect 15289 6613 15301 6647
rect 15335 6613 15347 6647
rect 15289 6607 15347 6613
rect 16577 6647 16635 6653
rect 16577 6613 16589 6647
rect 16623 6613 16635 6647
rect 16577 6607 16635 6613
rect 16945 6647 17003 6653
rect 16945 6613 16957 6647
rect 16991 6644 17003 6647
rect 17494 6644 17500 6656
rect 16991 6616 17500 6644
rect 16991 6613 17003 6616
rect 16945 6607 17003 6613
rect 17494 6604 17500 6616
rect 17552 6604 17558 6656
rect 17678 6604 17684 6656
rect 17736 6644 17742 6656
rect 18064 6644 18092 6675
rect 20162 6672 20168 6684
rect 20220 6672 20226 6724
rect 20272 6684 21312 6712
rect 17736 6616 18092 6644
rect 17736 6604 17742 6616
rect 18138 6604 18144 6656
rect 18196 6644 18202 6656
rect 18785 6647 18843 6653
rect 18785 6644 18797 6647
rect 18196 6616 18797 6644
rect 18196 6604 18202 6616
rect 18785 6613 18797 6616
rect 18831 6613 18843 6647
rect 18785 6607 18843 6613
rect 18966 6604 18972 6656
rect 19024 6644 19030 6656
rect 20272 6644 20300 6684
rect 19024 6616 20300 6644
rect 19024 6604 19030 6616
rect 20622 6604 20628 6656
rect 20680 6644 20686 6656
rect 21284 6653 21312 6684
rect 20809 6647 20867 6653
rect 20809 6644 20821 6647
rect 20680 6616 20821 6644
rect 20680 6604 20686 6616
rect 20809 6613 20821 6616
rect 20855 6613 20867 6647
rect 20809 6607 20867 6613
rect 21269 6647 21327 6653
rect 21269 6613 21281 6647
rect 21315 6613 21327 6647
rect 21269 6607 21327 6613
rect 1104 6554 21896 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21896 6554
rect 1104 6480 21896 6502
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 3142 6440 3148 6452
rect 2832 6412 3148 6440
rect 2832 6400 2838 6412
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 3878 6440 3884 6452
rect 3839 6412 3884 6440
rect 3878 6400 3884 6412
rect 3936 6400 3942 6452
rect 4525 6443 4583 6449
rect 4525 6409 4537 6443
rect 4571 6440 4583 6443
rect 5074 6440 5080 6452
rect 4571 6412 5080 6440
rect 4571 6409 4583 6412
rect 4525 6403 4583 6409
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 5997 6443 6055 6449
rect 5997 6409 6009 6443
rect 6043 6440 6055 6443
rect 6730 6440 6736 6452
rect 6043 6412 6736 6440
rect 6043 6409 6055 6412
rect 5997 6403 6055 6409
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 7009 6443 7067 6449
rect 7009 6409 7021 6443
rect 7055 6440 7067 6443
rect 8202 6440 8208 6452
rect 7055 6412 8208 6440
rect 7055 6409 7067 6412
rect 7009 6403 7067 6409
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 9122 6440 9128 6452
rect 9083 6412 9128 6440
rect 9122 6400 9128 6412
rect 9180 6400 9186 6452
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 10321 6443 10379 6449
rect 10321 6440 10333 6443
rect 9732 6412 10333 6440
rect 9732 6400 9738 6412
rect 10321 6409 10333 6412
rect 10367 6409 10379 6443
rect 10321 6403 10379 6409
rect 10410 6400 10416 6452
rect 10468 6440 10474 6452
rect 10689 6443 10747 6449
rect 10689 6440 10701 6443
rect 10468 6412 10701 6440
rect 10468 6400 10474 6412
rect 10689 6409 10701 6412
rect 10735 6409 10747 6443
rect 10689 6403 10747 6409
rect 11146 6400 11152 6452
rect 11204 6440 11210 6452
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 11204 6412 11529 6440
rect 11204 6400 11210 6412
rect 11517 6409 11529 6412
rect 11563 6409 11575 6443
rect 11882 6440 11888 6452
rect 11843 6412 11888 6440
rect 11517 6403 11575 6409
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 11977 6443 12035 6449
rect 11977 6409 11989 6443
rect 12023 6440 12035 6443
rect 12526 6440 12532 6452
rect 12023 6412 12532 6440
rect 12023 6409 12035 6412
rect 11977 6403 12035 6409
rect 12526 6400 12532 6412
rect 12584 6400 12590 6452
rect 13078 6440 13084 6452
rect 13039 6412 13084 6440
rect 13078 6400 13084 6412
rect 13136 6400 13142 6452
rect 13630 6400 13636 6452
rect 13688 6440 13694 6452
rect 14366 6440 14372 6452
rect 13688 6412 14372 6440
rect 13688 6400 13694 6412
rect 14366 6400 14372 6412
rect 14424 6400 14430 6452
rect 14734 6400 14740 6452
rect 14792 6440 14798 6452
rect 17954 6440 17960 6452
rect 14792 6412 17960 6440
rect 14792 6400 14798 6412
rect 17954 6400 17960 6412
rect 18012 6400 18018 6452
rect 20530 6440 20536 6452
rect 20491 6412 20536 6440
rect 20530 6400 20536 6412
rect 20588 6400 20594 6452
rect 20898 6440 20904 6452
rect 20859 6412 20904 6440
rect 20898 6400 20904 6412
rect 20956 6400 20962 6452
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 8018 6381 8024 6384
rect 8012 6372 8024 6381
rect 5592 6344 7512 6372
rect 7979 6344 8024 6372
rect 5592 6332 5598 6344
rect 1394 6304 1400 6316
rect 1355 6276 1400 6304
rect 1394 6264 1400 6276
rect 1452 6304 1458 6316
rect 1857 6307 1915 6313
rect 1857 6304 1869 6307
rect 1452 6276 1869 6304
rect 1452 6264 1458 6276
rect 1857 6273 1869 6276
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6304 5687 6307
rect 7282 6304 7288 6316
rect 5675 6276 7288 6304
rect 5675 6273 5687 6276
rect 5629 6267 5687 6273
rect 7282 6264 7288 6276
rect 7340 6264 7346 6316
rect 7484 6304 7512 6344
rect 8012 6335 8024 6344
rect 8018 6332 8024 6335
rect 8076 6332 8082 6384
rect 8570 6332 8576 6384
rect 8628 6372 8634 6384
rect 11054 6372 11060 6384
rect 8628 6344 11060 6372
rect 8628 6332 8634 6344
rect 11054 6332 11060 6344
rect 11112 6332 11118 6384
rect 13354 6332 13360 6384
rect 13412 6372 13418 6384
rect 14642 6372 14648 6384
rect 13412 6344 14648 6372
rect 13412 6332 13418 6344
rect 14642 6332 14648 6344
rect 14700 6332 14706 6384
rect 14826 6372 14832 6384
rect 14752 6344 14832 6372
rect 10045 6307 10103 6313
rect 7484 6276 9674 6304
rect 6546 6236 6552 6248
rect 6507 6208 6552 6236
rect 6546 6196 6552 6208
rect 6604 6196 6610 6248
rect 7745 6239 7803 6245
rect 7745 6205 7757 6239
rect 7791 6205 7803 6239
rect 9646 6236 9674 6276
rect 10045 6273 10057 6307
rect 10091 6304 10103 6307
rect 11238 6304 11244 6316
rect 10091 6276 11244 6304
rect 10091 6273 10103 6276
rect 10045 6267 10103 6273
rect 11238 6264 11244 6276
rect 11296 6264 11302 6316
rect 12529 6307 12587 6313
rect 12529 6273 12541 6307
rect 12575 6304 12587 6307
rect 12618 6304 12624 6316
rect 12575 6276 12624 6304
rect 12575 6273 12587 6276
rect 12529 6267 12587 6273
rect 12618 6264 12624 6276
rect 12676 6264 12682 6316
rect 14205 6307 14263 6313
rect 14205 6273 14217 6307
rect 14251 6304 14263 6307
rect 14752 6304 14780 6344
rect 14826 6332 14832 6344
rect 14884 6332 14890 6384
rect 19426 6372 19432 6384
rect 14936 6344 19432 6372
rect 14936 6316 14964 6344
rect 17144 6316 17172 6344
rect 14918 6304 14924 6316
rect 14251 6276 14780 6304
rect 14879 6276 14924 6304
rect 14251 6273 14263 6276
rect 14205 6267 14263 6273
rect 14918 6264 14924 6276
rect 14976 6264 14982 6316
rect 15194 6313 15200 6316
rect 15188 6267 15200 6313
rect 15252 6304 15258 6316
rect 16669 6307 16727 6313
rect 15252 6276 15288 6304
rect 15194 6264 15200 6267
rect 15252 6264 15258 6276
rect 16669 6273 16681 6307
rect 16715 6304 16727 6307
rect 16942 6304 16948 6316
rect 16715 6276 16948 6304
rect 16715 6273 16727 6276
rect 16669 6267 16727 6273
rect 16942 6264 16948 6276
rect 17000 6264 17006 6316
rect 17126 6264 17132 6316
rect 17184 6304 17190 6316
rect 17396 6307 17454 6313
rect 17184 6276 17277 6304
rect 17184 6264 17190 6276
rect 17396 6273 17408 6307
rect 17442 6304 17454 6307
rect 17770 6304 17776 6316
rect 17442 6276 17776 6304
rect 17442 6273 17454 6276
rect 17396 6267 17454 6273
rect 17770 6264 17776 6276
rect 17828 6264 17834 6316
rect 18800 6313 18828 6344
rect 19426 6332 19432 6344
rect 19484 6332 19490 6384
rect 19058 6313 19064 6316
rect 18785 6307 18843 6313
rect 18785 6273 18797 6307
rect 18831 6273 18843 6307
rect 19052 6304 19064 6313
rect 19019 6276 19064 6304
rect 18785 6267 18843 6273
rect 19052 6267 19064 6276
rect 19058 6264 19064 6267
rect 19116 6264 19122 6316
rect 10594 6236 10600 6248
rect 9646 6208 10600 6236
rect 7745 6199 7803 6205
rect 6730 6128 6736 6180
rect 6788 6168 6794 6180
rect 7760 6168 7788 6199
rect 10594 6196 10600 6208
rect 10652 6196 10658 6248
rect 10778 6236 10784 6248
rect 10739 6208 10784 6236
rect 10778 6196 10784 6208
rect 10836 6196 10842 6248
rect 10870 6196 10876 6248
rect 10928 6236 10934 6248
rect 10928 6208 10973 6236
rect 10928 6196 10934 6208
rect 11698 6196 11704 6248
rect 11756 6236 11762 6248
rect 12069 6239 12127 6245
rect 12069 6236 12081 6239
rect 11756 6208 12081 6236
rect 11756 6196 11762 6208
rect 12069 6205 12081 6208
rect 12115 6205 12127 6239
rect 14458 6236 14464 6248
rect 14419 6208 14464 6236
rect 12069 6199 12127 6205
rect 14458 6196 14464 6208
rect 14516 6196 14522 6248
rect 20622 6196 20628 6248
rect 20680 6236 20686 6248
rect 20993 6239 21051 6245
rect 20993 6236 21005 6239
rect 20680 6208 21005 6236
rect 20680 6196 20686 6208
rect 20993 6205 21005 6208
rect 21039 6205 21051 6239
rect 21174 6236 21180 6248
rect 21135 6208 21180 6236
rect 20993 6199 21051 6205
rect 21174 6196 21180 6208
rect 21232 6196 21238 6248
rect 6788 6140 7788 6168
rect 6788 6128 6794 6140
rect 1578 6100 1584 6112
rect 1539 6072 1584 6100
rect 1578 6060 1584 6072
rect 1636 6060 1642 6112
rect 1670 6060 1676 6112
rect 1728 6100 1734 6112
rect 2225 6103 2283 6109
rect 2225 6100 2237 6103
rect 1728 6072 2237 6100
rect 1728 6060 1734 6072
rect 2225 6069 2237 6072
rect 2271 6069 2283 6103
rect 3418 6100 3424 6112
rect 3379 6072 3424 6100
rect 2225 6063 2283 6069
rect 3418 6060 3424 6072
rect 3476 6060 3482 6112
rect 4890 6100 4896 6112
rect 4851 6072 4896 6100
rect 4890 6060 4896 6072
rect 4948 6060 4954 6112
rect 5261 6103 5319 6109
rect 5261 6069 5273 6103
rect 5307 6100 5319 6103
rect 6546 6100 6552 6112
rect 5307 6072 6552 6100
rect 5307 6069 5319 6072
rect 5261 6063 5319 6069
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 7466 6100 7472 6112
rect 7427 6072 7472 6100
rect 7466 6060 7472 6072
rect 7524 6060 7530 6112
rect 7760 6100 7788 6140
rect 10502 6128 10508 6180
rect 10560 6168 10566 6180
rect 16942 6168 16948 6180
rect 10560 6140 13584 6168
rect 10560 6128 10566 6140
rect 8662 6100 8668 6112
rect 7760 6072 8668 6100
rect 8662 6060 8668 6072
rect 8720 6060 8726 6112
rect 9401 6103 9459 6109
rect 9401 6069 9413 6103
rect 9447 6100 9459 6103
rect 10962 6100 10968 6112
rect 9447 6072 10968 6100
rect 9447 6069 9459 6072
rect 9401 6063 9459 6069
rect 10962 6060 10968 6072
rect 11020 6060 11026 6112
rect 12713 6103 12771 6109
rect 12713 6069 12725 6103
rect 12759 6100 12771 6103
rect 13446 6100 13452 6112
rect 12759 6072 13452 6100
rect 12759 6069 12771 6072
rect 12713 6063 12771 6069
rect 13446 6060 13452 6072
rect 13504 6060 13510 6112
rect 13556 6100 13584 6140
rect 16316 6140 16948 6168
rect 16316 6109 16344 6140
rect 16942 6128 16948 6140
rect 17000 6128 17006 6180
rect 18340 6140 18828 6168
rect 16301 6103 16359 6109
rect 16301 6100 16313 6103
rect 13556 6072 16313 6100
rect 16301 6069 16313 6072
rect 16347 6069 16359 6103
rect 16301 6063 16359 6069
rect 16853 6103 16911 6109
rect 16853 6069 16865 6103
rect 16899 6100 16911 6103
rect 18340 6100 18368 6140
rect 18506 6100 18512 6112
rect 16899 6072 18368 6100
rect 18467 6072 18512 6100
rect 16899 6069 16911 6072
rect 16853 6063 16911 6069
rect 18506 6060 18512 6072
rect 18564 6060 18570 6112
rect 18800 6100 18828 6140
rect 19518 6100 19524 6112
rect 18800 6072 19524 6100
rect 19518 6060 19524 6072
rect 19576 6060 19582 6112
rect 20162 6100 20168 6112
rect 20123 6072 20168 6100
rect 20162 6060 20168 6072
rect 20220 6060 20226 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 3421 5899 3479 5905
rect 3421 5865 3433 5899
rect 3467 5896 3479 5899
rect 4246 5896 4252 5908
rect 3467 5868 4252 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 6457 5899 6515 5905
rect 6457 5865 6469 5899
rect 6503 5896 6515 5899
rect 6638 5896 6644 5908
rect 6503 5868 6644 5896
rect 6503 5865 6515 5868
rect 6457 5859 6515 5865
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 7466 5856 7472 5908
rect 7524 5896 7530 5908
rect 7524 5868 8064 5896
rect 7524 5856 7530 5868
rect 2406 5788 2412 5840
rect 2464 5828 2470 5840
rect 5810 5828 5816 5840
rect 2464 5800 5816 5828
rect 2464 5788 2470 5800
rect 5810 5788 5816 5800
rect 5868 5828 5874 5840
rect 5905 5831 5963 5837
rect 5905 5828 5917 5831
rect 5868 5800 5917 5828
rect 5868 5788 5874 5800
rect 5905 5797 5917 5800
rect 5951 5797 5963 5831
rect 8036 5828 8064 5868
rect 8110 5856 8116 5908
rect 8168 5896 8174 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8168 5868 9045 5896
rect 8168 5856 8174 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 10594 5896 10600 5908
rect 9033 5859 9091 5865
rect 9646 5868 10600 5896
rect 8294 5828 8300 5840
rect 8036 5800 8300 5828
rect 5905 5791 5963 5797
rect 8294 5788 8300 5800
rect 8352 5788 8358 5840
rect 8662 5788 8668 5840
rect 8720 5828 8726 5840
rect 9646 5828 9674 5868
rect 10594 5856 10600 5868
rect 10652 5896 10658 5908
rect 10689 5899 10747 5905
rect 10689 5896 10701 5899
rect 10652 5868 10701 5896
rect 10652 5856 10658 5868
rect 10689 5865 10701 5868
rect 10735 5865 10747 5899
rect 10689 5859 10747 5865
rect 10778 5856 10784 5908
rect 10836 5896 10842 5908
rect 14274 5896 14280 5908
rect 10836 5868 14280 5896
rect 10836 5856 10842 5868
rect 14274 5856 14280 5868
rect 14332 5856 14338 5908
rect 14642 5856 14648 5908
rect 14700 5896 14706 5908
rect 15289 5899 15347 5905
rect 15289 5896 15301 5899
rect 14700 5868 15301 5896
rect 14700 5856 14706 5868
rect 15289 5865 15301 5868
rect 15335 5896 15347 5899
rect 15746 5896 15752 5908
rect 15335 5868 15752 5896
rect 15335 5865 15347 5868
rect 15289 5859 15347 5865
rect 15746 5856 15752 5868
rect 15804 5856 15810 5908
rect 17126 5896 17132 5908
rect 17087 5868 17132 5896
rect 17126 5856 17132 5868
rect 17184 5856 17190 5908
rect 17494 5856 17500 5908
rect 17552 5896 17558 5908
rect 17865 5899 17923 5905
rect 17865 5896 17877 5899
rect 17552 5868 17877 5896
rect 17552 5856 17558 5868
rect 17865 5865 17877 5868
rect 17911 5865 17923 5899
rect 19058 5896 19064 5908
rect 17865 5859 17923 5865
rect 17972 5868 19064 5896
rect 8720 5800 9674 5828
rect 8720 5788 8726 5800
rect 9766 5788 9772 5840
rect 9824 5828 9830 5840
rect 9824 5800 12848 5828
rect 9824 5788 9830 5800
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 6730 5760 6736 5772
rect 1636 5732 6408 5760
rect 6691 5732 6736 5760
rect 1636 5720 1642 5732
rect 4430 5692 4436 5704
rect 4391 5664 4436 5692
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 5534 5692 5540 5704
rect 5495 5664 5540 5692
rect 5534 5652 5540 5664
rect 5592 5652 5598 5704
rect 5902 5652 5908 5704
rect 5960 5692 5966 5704
rect 6273 5695 6331 5701
rect 6273 5692 6285 5695
rect 5960 5664 6285 5692
rect 5960 5652 5966 5664
rect 6273 5661 6285 5664
rect 6319 5661 6331 5695
rect 6380 5692 6408 5732
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 8018 5720 8024 5772
rect 8076 5760 8082 5772
rect 9677 5763 9735 5769
rect 9677 5760 9689 5763
rect 8076 5732 9689 5760
rect 8076 5720 8082 5732
rect 6989 5695 7047 5701
rect 6989 5692 7001 5695
rect 6380 5664 7001 5692
rect 6273 5655 6331 5661
rect 6989 5661 7001 5664
rect 7035 5661 7047 5695
rect 6989 5655 7047 5661
rect 3053 5627 3111 5633
rect 3053 5593 3065 5627
rect 3099 5624 3111 5627
rect 4338 5624 4344 5636
rect 3099 5596 4344 5624
rect 3099 5593 3111 5596
rect 3053 5587 3111 5593
rect 4338 5584 4344 5596
rect 4396 5584 4402 5636
rect 4893 5627 4951 5633
rect 4893 5593 4905 5627
rect 4939 5624 4951 5627
rect 6288 5624 6316 5655
rect 6454 5624 6460 5636
rect 4939 5596 6224 5624
rect 6288 5596 6460 5624
rect 4939 5593 4951 5596
rect 4893 5587 4951 5593
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 1946 5556 1952 5568
rect 1907 5528 1952 5556
rect 1946 5516 1952 5528
rect 2004 5516 2010 5568
rect 2317 5559 2375 5565
rect 2317 5525 2329 5559
rect 2363 5556 2375 5559
rect 2498 5556 2504 5568
rect 2363 5528 2504 5556
rect 2363 5525 2375 5528
rect 2317 5519 2375 5525
rect 2498 5516 2504 5528
rect 2556 5516 2562 5568
rect 2682 5556 2688 5568
rect 2643 5528 2688 5556
rect 2682 5516 2688 5528
rect 2740 5516 2746 5568
rect 4062 5516 4068 5568
rect 4120 5556 4126 5568
rect 4157 5559 4215 5565
rect 4157 5556 4169 5559
rect 4120 5528 4169 5556
rect 4120 5516 4126 5528
rect 4157 5525 4169 5528
rect 4203 5525 4215 5559
rect 4157 5519 4215 5525
rect 4246 5516 4252 5568
rect 4304 5556 4310 5568
rect 4982 5556 4988 5568
rect 4304 5528 4988 5556
rect 4304 5516 4310 5528
rect 4982 5516 4988 5528
rect 5040 5516 5046 5568
rect 5261 5559 5319 5565
rect 5261 5525 5273 5559
rect 5307 5556 5319 5559
rect 5994 5556 6000 5568
rect 5307 5528 6000 5556
rect 5307 5525 5319 5528
rect 5261 5519 5319 5525
rect 5994 5516 6000 5528
rect 6052 5516 6058 5568
rect 6196 5556 6224 5596
rect 6454 5584 6460 5596
rect 6512 5584 6518 5636
rect 7374 5556 7380 5568
rect 6196 5528 7380 5556
rect 7374 5516 7380 5528
rect 7432 5556 7438 5568
rect 7926 5556 7932 5568
rect 7432 5528 7932 5556
rect 7432 5516 7438 5528
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 8128 5565 8156 5732
rect 9677 5729 9689 5732
rect 9723 5760 9735 5763
rect 10870 5760 10876 5772
rect 9723 5732 10876 5760
rect 9723 5729 9735 5732
rect 9677 5723 9735 5729
rect 10870 5720 10876 5732
rect 10928 5720 10934 5772
rect 12710 5760 12716 5772
rect 11992 5732 12434 5760
rect 12671 5732 12716 5760
rect 8570 5652 8576 5704
rect 8628 5692 8634 5704
rect 8628 5664 10180 5692
rect 8628 5652 8634 5664
rect 9122 5584 9128 5636
rect 9180 5624 9186 5636
rect 9401 5627 9459 5633
rect 9401 5624 9413 5627
rect 9180 5596 9413 5624
rect 9180 5584 9186 5596
rect 9401 5593 9413 5596
rect 9447 5593 9459 5627
rect 9401 5587 9459 5593
rect 9490 5584 9496 5636
rect 9548 5624 9554 5636
rect 9548 5596 9593 5624
rect 9548 5584 9554 5596
rect 8113 5559 8171 5565
rect 8113 5525 8125 5559
rect 8159 5525 8171 5559
rect 8570 5556 8576 5568
rect 8531 5528 8576 5556
rect 8113 5519 8171 5525
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 10152 5565 10180 5664
rect 10318 5652 10324 5704
rect 10376 5692 10382 5704
rect 11992 5692 12020 5732
rect 12158 5692 12164 5704
rect 10376 5664 12020 5692
rect 12119 5664 12164 5692
rect 10376 5652 10382 5664
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 12406 5692 12434 5732
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 12820 5769 12848 5800
rect 13170 5788 13176 5840
rect 13228 5828 13234 5840
rect 17972 5828 18000 5868
rect 19058 5856 19064 5868
rect 19116 5896 19122 5908
rect 20625 5899 20683 5905
rect 20625 5896 20637 5899
rect 19116 5868 20637 5896
rect 19116 5856 19122 5868
rect 20625 5865 20637 5868
rect 20671 5865 20683 5899
rect 20625 5859 20683 5865
rect 13228 5800 18000 5828
rect 13228 5788 13234 5800
rect 12805 5763 12863 5769
rect 12805 5729 12817 5763
rect 12851 5760 12863 5763
rect 12986 5760 12992 5772
rect 12851 5732 12992 5760
rect 12851 5729 12863 5732
rect 12805 5723 12863 5729
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 14366 5760 14372 5772
rect 13464 5732 13860 5760
rect 14327 5732 14372 5760
rect 13464 5692 13492 5732
rect 13722 5692 13728 5704
rect 12406 5664 13492 5692
rect 13683 5664 13728 5692
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 13832 5692 13860 5732
rect 14366 5720 14372 5732
rect 14424 5720 14430 5772
rect 18322 5760 18328 5772
rect 18283 5732 18328 5760
rect 18322 5720 18328 5732
rect 18380 5720 18386 5772
rect 18414 5720 18420 5772
rect 18472 5760 18478 5772
rect 18472 5732 18517 5760
rect 18472 5720 18478 5732
rect 18874 5720 18880 5772
rect 18932 5760 18938 5772
rect 18932 5732 19380 5760
rect 18932 5720 18938 5732
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 13832 5664 14565 5692
rect 14553 5661 14565 5664
rect 14599 5661 14611 5695
rect 14553 5655 14611 5661
rect 17126 5652 17132 5704
rect 17184 5692 17190 5704
rect 18966 5692 18972 5704
rect 17184 5664 18972 5692
rect 17184 5652 17190 5664
rect 18966 5652 18972 5664
rect 19024 5692 19030 5704
rect 19245 5695 19303 5701
rect 19245 5692 19257 5695
rect 19024 5664 19257 5692
rect 19024 5652 19030 5664
rect 19245 5661 19257 5664
rect 19291 5661 19303 5695
rect 19352 5692 19380 5732
rect 20901 5695 20959 5701
rect 20901 5692 20913 5695
rect 19352 5664 20913 5692
rect 19245 5655 19303 5661
rect 20901 5661 20913 5664
rect 20947 5661 20959 5695
rect 20901 5655 20959 5661
rect 20990 5652 20996 5704
rect 21048 5692 21054 5704
rect 21085 5695 21143 5701
rect 21085 5692 21097 5695
rect 21048 5664 21097 5692
rect 21048 5652 21054 5664
rect 21085 5661 21097 5664
rect 21131 5692 21143 5695
rect 21818 5692 21824 5704
rect 21131 5664 21824 5692
rect 21131 5661 21143 5664
rect 21085 5655 21143 5661
rect 21818 5652 21824 5664
rect 21876 5652 21882 5704
rect 10594 5584 10600 5636
rect 10652 5624 10658 5636
rect 11238 5624 11244 5636
rect 10652 5596 11244 5624
rect 10652 5584 10658 5596
rect 11238 5584 11244 5596
rect 11296 5584 11302 5636
rect 12176 5624 12204 5652
rect 15654 5624 15660 5636
rect 12176 5596 15660 5624
rect 15654 5584 15660 5596
rect 15712 5584 15718 5636
rect 19334 5584 19340 5636
rect 19392 5624 19398 5636
rect 19490 5627 19548 5633
rect 19490 5624 19502 5627
rect 19392 5596 19502 5624
rect 19392 5584 19398 5596
rect 19490 5593 19502 5596
rect 19536 5593 19548 5627
rect 19490 5587 19548 5593
rect 10137 5559 10195 5565
rect 10137 5525 10149 5559
rect 10183 5556 10195 5559
rect 12250 5556 12256 5568
rect 10183 5528 12256 5556
rect 10183 5525 10195 5528
rect 10137 5519 10195 5525
rect 12250 5516 12256 5528
rect 12308 5516 12314 5568
rect 12802 5516 12808 5568
rect 12860 5556 12866 5568
rect 12897 5559 12955 5565
rect 12897 5556 12909 5559
rect 12860 5528 12909 5556
rect 12860 5516 12866 5528
rect 12897 5525 12909 5528
rect 12943 5525 12955 5559
rect 12897 5519 12955 5525
rect 12986 5516 12992 5568
rect 13044 5556 13050 5568
rect 13265 5559 13323 5565
rect 13265 5556 13277 5559
rect 13044 5528 13277 5556
rect 13044 5516 13050 5528
rect 13265 5525 13277 5528
rect 13311 5525 13323 5559
rect 13265 5519 13323 5525
rect 13541 5559 13599 5565
rect 13541 5525 13553 5559
rect 13587 5556 13599 5559
rect 14274 5556 14280 5568
rect 13587 5528 14280 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 14550 5516 14556 5568
rect 14608 5556 14614 5568
rect 14645 5559 14703 5565
rect 14645 5556 14657 5559
rect 14608 5528 14657 5556
rect 14608 5516 14614 5528
rect 14645 5525 14657 5528
rect 14691 5525 14703 5559
rect 15010 5556 15016 5568
rect 14971 5528 15016 5556
rect 14645 5519 14703 5525
rect 15010 5516 15016 5528
rect 15068 5516 15074 5568
rect 18230 5556 18236 5568
rect 18191 5528 18236 5556
rect 18230 5516 18236 5528
rect 18288 5516 18294 5568
rect 1104 5466 21896 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21896 5466
rect 1104 5392 21896 5414
rect 1854 5352 1860 5364
rect 1815 5324 1860 5352
rect 1854 5312 1860 5324
rect 1912 5312 1918 5364
rect 4065 5355 4123 5361
rect 4065 5321 4077 5355
rect 4111 5352 4123 5355
rect 7650 5352 7656 5364
rect 4111 5324 7052 5352
rect 7611 5324 7656 5352
rect 4111 5321 4123 5324
rect 4065 5315 4123 5321
rect 4433 5287 4491 5293
rect 4433 5253 4445 5287
rect 4479 5284 4491 5287
rect 5442 5284 5448 5296
rect 4479 5256 5448 5284
rect 4479 5253 4491 5256
rect 4433 5247 4491 5253
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 5537 5287 5595 5293
rect 5537 5253 5549 5287
rect 5583 5284 5595 5287
rect 6086 5284 6092 5296
rect 5583 5256 6092 5284
rect 5583 5253 5595 5256
rect 5537 5247 5595 5253
rect 6086 5244 6092 5256
rect 6144 5284 6150 5296
rect 6822 5284 6828 5296
rect 6144 5256 6828 5284
rect 6144 5244 6150 5256
rect 6822 5244 6828 5256
rect 6880 5244 6886 5296
rect 7024 5228 7052 5324
rect 7650 5312 7656 5324
rect 7708 5312 7714 5364
rect 8386 5352 8392 5364
rect 8347 5324 8392 5352
rect 8386 5312 8392 5324
rect 8444 5312 8450 5364
rect 14366 5352 14372 5364
rect 9048 5324 14372 5352
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5216 3019 5219
rect 4614 5216 4620 5228
rect 3007 5188 4620 5216
rect 3007 5185 3019 5188
rect 2961 5179 3019 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 4801 5219 4859 5225
rect 4801 5185 4813 5219
rect 4847 5216 4859 5219
rect 5718 5216 5724 5228
rect 4847 5188 5724 5216
rect 4847 5185 4859 5188
rect 4801 5179 4859 5185
rect 5718 5176 5724 5188
rect 5776 5176 5782 5228
rect 5997 5219 6055 5225
rect 5997 5185 6009 5219
rect 6043 5216 6055 5219
rect 6454 5216 6460 5228
rect 6043 5188 6460 5216
rect 6043 5185 6055 5188
rect 5997 5179 6055 5185
rect 6454 5176 6460 5188
rect 6512 5176 6518 5228
rect 6549 5219 6607 5225
rect 6549 5185 6561 5219
rect 6595 5216 6607 5219
rect 6638 5216 6644 5228
rect 6595 5188 6644 5216
rect 6595 5185 6607 5188
rect 6549 5179 6607 5185
rect 6638 5176 6644 5188
rect 6696 5176 6702 5228
rect 7006 5216 7012 5228
rect 6919 5188 7012 5216
rect 7006 5176 7012 5188
rect 7064 5176 7070 5228
rect 7374 5176 7380 5228
rect 7432 5216 7438 5228
rect 7469 5219 7527 5225
rect 7469 5216 7481 5219
rect 7432 5188 7481 5216
rect 7432 5176 7438 5188
rect 7469 5185 7481 5188
rect 7515 5185 7527 5219
rect 7469 5179 7527 5185
rect 7929 5220 7987 5225
rect 8018 5220 8024 5228
rect 7929 5219 8024 5220
rect 7929 5185 7941 5219
rect 7975 5192 8024 5219
rect 7975 5185 7987 5192
rect 7929 5179 7987 5185
rect 8018 5176 8024 5192
rect 8076 5176 8082 5228
rect 9048 5225 9076 5324
rect 14366 5312 14372 5324
rect 14424 5312 14430 5364
rect 14553 5355 14611 5361
rect 14553 5321 14565 5355
rect 14599 5352 14611 5355
rect 14599 5324 14872 5352
rect 14599 5321 14611 5324
rect 14553 5315 14611 5321
rect 9306 5284 9312 5296
rect 9267 5256 9312 5284
rect 9306 5244 9312 5256
rect 9364 5244 9370 5296
rect 10686 5284 10692 5296
rect 10647 5256 10692 5284
rect 10686 5244 10692 5256
rect 10744 5244 10750 5296
rect 12342 5284 12348 5296
rect 11532 5256 12348 5284
rect 9033 5219 9091 5225
rect 9033 5185 9045 5219
rect 9079 5185 9091 5219
rect 9033 5179 9091 5185
rect 9953 5219 10011 5225
rect 9953 5185 9965 5219
rect 9999 5216 10011 5219
rect 10502 5216 10508 5228
rect 9999 5188 10508 5216
rect 9999 5185 10011 5188
rect 9953 5179 10011 5185
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 10594 5176 10600 5228
rect 10652 5216 10658 5228
rect 10652 5188 10697 5216
rect 10652 5176 10658 5188
rect 11238 5176 11244 5228
rect 11296 5216 11302 5228
rect 11532 5225 11560 5256
rect 12342 5244 12348 5256
rect 12400 5244 12406 5296
rect 13630 5284 13636 5296
rect 13188 5256 13636 5284
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 11296 5188 11529 5216
rect 11296 5176 11302 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 11773 5219 11831 5225
rect 11773 5216 11785 5219
rect 11517 5179 11575 5185
rect 11624 5188 11785 5216
rect 1489 5151 1547 5157
rect 1489 5117 1501 5151
rect 1535 5148 1547 5151
rect 3234 5148 3240 5160
rect 1535 5120 3240 5148
rect 1535 5117 1547 5120
rect 1489 5111 1547 5117
rect 3234 5108 3240 5120
rect 3292 5108 3298 5160
rect 5810 5148 5816 5160
rect 3620 5120 5816 5148
rect 2593 5083 2651 5089
rect 2593 5049 2605 5083
rect 2639 5080 2651 5083
rect 3620 5080 3648 5120
rect 5810 5108 5816 5120
rect 5868 5108 5874 5160
rect 9766 5148 9772 5160
rect 6748 5120 9772 5148
rect 2639 5052 3648 5080
rect 3697 5083 3755 5089
rect 2639 5049 2651 5052
rect 2593 5043 2651 5049
rect 3697 5049 3709 5083
rect 3743 5080 3755 5083
rect 5994 5080 6000 5092
rect 3743 5052 6000 5080
rect 3743 5049 3755 5052
rect 3697 5043 3755 5049
rect 5994 5040 6000 5052
rect 6052 5040 6058 5092
rect 6748 5089 6776 5120
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 10870 5148 10876 5160
rect 10831 5120 10876 5148
rect 10870 5108 10876 5120
rect 10928 5108 10934 5160
rect 10962 5108 10968 5160
rect 11020 5148 11026 5160
rect 11624 5148 11652 5188
rect 11773 5185 11785 5188
rect 11819 5185 11831 5219
rect 12360 5216 12388 5244
rect 13188 5225 13216 5256
rect 13630 5244 13636 5256
rect 13688 5284 13694 5296
rect 14458 5284 14464 5296
rect 13688 5256 14464 5284
rect 13688 5244 13694 5256
rect 14458 5244 14464 5256
rect 14516 5244 14522 5296
rect 14844 5284 14872 5324
rect 15304 5324 18000 5352
rect 15074 5287 15132 5293
rect 15074 5284 15086 5287
rect 14844 5256 15086 5284
rect 15074 5253 15086 5256
rect 15120 5284 15132 5287
rect 15194 5284 15200 5296
rect 15120 5256 15200 5284
rect 15120 5253 15132 5256
rect 15074 5247 15132 5253
rect 15194 5244 15200 5256
rect 15252 5244 15258 5296
rect 13173 5219 13231 5225
rect 13173 5216 13185 5219
rect 12360 5188 13185 5216
rect 11773 5179 11831 5185
rect 13173 5185 13185 5188
rect 13219 5185 13231 5219
rect 13429 5219 13487 5225
rect 13429 5216 13441 5219
rect 13173 5179 13231 5185
rect 13280 5188 13441 5216
rect 13280 5148 13308 5188
rect 13429 5185 13441 5188
rect 13475 5185 13487 5219
rect 13429 5179 13487 5185
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 15304 5216 15332 5324
rect 16574 5244 16580 5296
rect 16632 5284 16638 5296
rect 17190 5287 17248 5293
rect 17190 5284 17202 5287
rect 16632 5256 17202 5284
rect 16632 5244 16638 5256
rect 17190 5253 17202 5256
rect 17236 5253 17248 5287
rect 17190 5247 17248 5253
rect 13780 5188 15332 5216
rect 16945 5219 17003 5225
rect 13780 5176 13786 5188
rect 16945 5185 16957 5219
rect 16991 5216 17003 5219
rect 17034 5216 17040 5228
rect 16991 5188 17040 5216
rect 16991 5185 17003 5188
rect 16945 5179 17003 5185
rect 17034 5176 17040 5188
rect 17092 5176 17098 5228
rect 11020 5120 11652 5148
rect 12820 5120 13308 5148
rect 11020 5108 11026 5120
rect 6733 5083 6791 5089
rect 6733 5049 6745 5083
rect 6779 5049 6791 5083
rect 6733 5043 6791 5049
rect 9950 5040 9956 5092
rect 10008 5080 10014 5092
rect 10229 5083 10287 5089
rect 10229 5080 10241 5083
rect 10008 5052 10241 5080
rect 10008 5040 10014 5052
rect 10229 5049 10241 5052
rect 10275 5049 10287 5083
rect 10229 5043 10287 5049
rect 2222 5012 2228 5024
rect 2183 4984 2228 5012
rect 2222 4972 2228 4984
rect 2280 4972 2286 5024
rect 3329 5015 3387 5021
rect 3329 4981 3341 5015
rect 3375 5012 3387 5015
rect 4706 5012 4712 5024
rect 3375 4984 4712 5012
rect 3375 4981 3387 4984
rect 3329 4975 3387 4981
rect 4706 4972 4712 4984
rect 4764 4972 4770 5024
rect 4890 4972 4896 5024
rect 4948 5012 4954 5024
rect 5077 5015 5135 5021
rect 5077 5012 5089 5015
rect 4948 4984 5089 5012
rect 4948 4972 4954 4984
rect 5077 4981 5089 4984
rect 5123 4981 5135 5015
rect 5077 4975 5135 4981
rect 5534 4972 5540 5024
rect 5592 5012 5598 5024
rect 5813 5015 5871 5021
rect 5813 5012 5825 5015
rect 5592 4984 5825 5012
rect 5592 4972 5598 4984
rect 5813 4981 5825 4984
rect 5859 4981 5871 5015
rect 5813 4975 5871 4981
rect 7193 5015 7251 5021
rect 7193 4981 7205 5015
rect 7239 5012 7251 5015
rect 7742 5012 7748 5024
rect 7239 4984 7748 5012
rect 7239 4981 7251 4984
rect 7193 4975 7251 4981
rect 7742 4972 7748 4984
rect 7800 4972 7806 5024
rect 8110 5012 8116 5024
rect 8071 4984 8116 5012
rect 8110 4972 8116 4984
rect 8168 4972 8174 5024
rect 9490 4972 9496 5024
rect 9548 5012 9554 5024
rect 12820 5012 12848 5120
rect 14458 5108 14464 5160
rect 14516 5148 14522 5160
rect 14829 5151 14887 5157
rect 14829 5148 14841 5151
rect 14516 5120 14841 5148
rect 14516 5108 14522 5120
rect 14829 5117 14841 5120
rect 14875 5117 14887 5151
rect 17972 5148 18000 5324
rect 18046 5312 18052 5364
rect 18104 5352 18110 5364
rect 19429 5355 19487 5361
rect 19429 5352 19441 5355
rect 18104 5324 19441 5352
rect 18104 5312 18110 5324
rect 19429 5321 19441 5324
rect 19475 5321 19487 5355
rect 19429 5315 19487 5321
rect 19610 5312 19616 5364
rect 19668 5352 19674 5364
rect 19797 5355 19855 5361
rect 19797 5352 19809 5355
rect 19668 5324 19809 5352
rect 19668 5312 19674 5324
rect 19797 5321 19809 5324
rect 19843 5321 19855 5355
rect 20622 5352 20628 5364
rect 20583 5324 20628 5352
rect 19797 5315 19855 5321
rect 20622 5312 20628 5324
rect 20680 5312 20686 5364
rect 18506 5244 18512 5296
rect 18564 5284 18570 5296
rect 18564 5256 20024 5284
rect 18564 5244 18570 5256
rect 18598 5216 18604 5228
rect 18559 5188 18604 5216
rect 18598 5176 18604 5188
rect 18656 5176 18662 5228
rect 19886 5148 19892 5160
rect 17972 5120 18920 5148
rect 19847 5120 19892 5148
rect 14829 5111 14887 5117
rect 16022 5040 16028 5092
rect 16080 5080 16086 5092
rect 18785 5083 18843 5089
rect 18785 5080 18797 5083
rect 16080 5052 16344 5080
rect 16080 5040 16086 5052
rect 9548 4984 12848 5012
rect 9548 4972 9554 4984
rect 12894 4972 12900 5024
rect 12952 5012 12958 5024
rect 12952 4984 12997 5012
rect 12952 4972 12958 4984
rect 14366 4972 14372 5024
rect 14424 5012 14430 5024
rect 15930 5012 15936 5024
rect 14424 4984 15936 5012
rect 14424 4972 14430 4984
rect 15930 4972 15936 4984
rect 15988 5012 15994 5024
rect 16209 5015 16267 5021
rect 16209 5012 16221 5015
rect 15988 4984 16221 5012
rect 15988 4972 15994 4984
rect 16209 4981 16221 4984
rect 16255 4981 16267 5015
rect 16316 5012 16344 5052
rect 17880 5052 18797 5080
rect 17880 5012 17908 5052
rect 18785 5049 18797 5052
rect 18831 5049 18843 5083
rect 18892 5080 18920 5120
rect 19886 5108 19892 5120
rect 19944 5108 19950 5160
rect 19996 5157 20024 5256
rect 20622 5176 20628 5228
rect 20680 5216 20686 5228
rect 20993 5219 21051 5225
rect 20993 5216 21005 5219
rect 20680 5188 21005 5216
rect 20680 5176 20686 5188
rect 20993 5185 21005 5188
rect 21039 5185 21051 5219
rect 20993 5179 21051 5185
rect 19981 5151 20039 5157
rect 19981 5117 19993 5151
rect 20027 5117 20039 5151
rect 19981 5111 20039 5117
rect 21085 5151 21143 5157
rect 21085 5117 21097 5151
rect 21131 5117 21143 5151
rect 21085 5111 21143 5117
rect 21269 5151 21327 5157
rect 21269 5117 21281 5151
rect 21315 5148 21327 5151
rect 21450 5148 21456 5160
rect 21315 5120 21456 5148
rect 21315 5117 21327 5120
rect 21269 5111 21327 5117
rect 21100 5080 21128 5111
rect 21450 5108 21456 5120
rect 21508 5108 21514 5160
rect 18892 5052 21128 5080
rect 18785 5043 18843 5049
rect 16316 4984 17908 5012
rect 18325 5015 18383 5021
rect 16209 4975 16267 4981
rect 18325 4981 18337 5015
rect 18371 5012 18383 5015
rect 18598 5012 18604 5024
rect 18371 4984 18604 5012
rect 18371 4981 18383 4984
rect 18325 4975 18383 4981
rect 18598 4972 18604 4984
rect 18656 4972 18662 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 4525 4811 4583 4817
rect 4525 4777 4537 4811
rect 4571 4808 4583 4811
rect 4706 4808 4712 4820
rect 4571 4780 4712 4808
rect 4571 4777 4583 4780
rect 4525 4771 4583 4777
rect 4706 4768 4712 4780
rect 4764 4768 4770 4820
rect 5353 4811 5411 4817
rect 5353 4777 5365 4811
rect 5399 4808 5411 4811
rect 5442 4808 5448 4820
rect 5399 4780 5448 4808
rect 5399 4777 5411 4780
rect 5353 4771 5411 4777
rect 5442 4768 5448 4780
rect 5500 4768 5506 4820
rect 5813 4811 5871 4817
rect 5813 4777 5825 4811
rect 5859 4808 5871 4811
rect 6362 4808 6368 4820
rect 5859 4780 6368 4808
rect 5859 4777 5871 4780
rect 5813 4771 5871 4777
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 6730 4808 6736 4820
rect 6691 4780 6736 4808
rect 6730 4768 6736 4780
rect 6788 4768 6794 4820
rect 7193 4811 7251 4817
rect 7193 4777 7205 4811
rect 7239 4808 7251 4811
rect 9122 4808 9128 4820
rect 7239 4780 9128 4808
rect 7239 4777 7251 4780
rect 7193 4771 7251 4777
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 10594 4808 10600 4820
rect 9324 4780 10600 4808
rect 3421 4743 3479 4749
rect 3421 4709 3433 4743
rect 3467 4740 3479 4743
rect 6086 4740 6092 4752
rect 3467 4712 6092 4740
rect 3467 4709 3479 4712
rect 3421 4703 3479 4709
rect 6086 4700 6092 4712
rect 6144 4700 6150 4752
rect 6273 4743 6331 4749
rect 6273 4709 6285 4743
rect 6319 4740 6331 4743
rect 9324 4740 9352 4780
rect 10594 4768 10600 4780
rect 10652 4808 10658 4820
rect 10652 4780 14228 4808
rect 10652 4768 10658 4780
rect 6319 4712 9352 4740
rect 6319 4709 6331 4712
rect 6273 4703 6331 4709
rect 13538 4700 13544 4752
rect 13596 4740 13602 4752
rect 13633 4743 13691 4749
rect 13633 4740 13645 4743
rect 13596 4712 13645 4740
rect 13596 4700 13602 4712
rect 13633 4709 13645 4712
rect 13679 4709 13691 4743
rect 13633 4703 13691 4709
rect 4157 4675 4215 4681
rect 4157 4641 4169 4675
rect 4203 4672 4215 4675
rect 7650 4672 7656 4684
rect 4203 4644 7512 4672
rect 7611 4644 7656 4672
rect 4203 4641 4215 4644
rect 4157 4635 4215 4641
rect 2685 4607 2743 4613
rect 2685 4573 2697 4607
rect 2731 4604 2743 4607
rect 5074 4604 5080 4616
rect 2731 4576 5080 4604
rect 2731 4573 2743 4576
rect 2685 4567 2743 4573
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4604 5227 4607
rect 5534 4604 5540 4616
rect 5215 4576 5540 4604
rect 5215 4573 5227 4576
rect 5169 4567 5227 4573
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4573 5687 4607
rect 5629 4567 5687 4573
rect 3694 4496 3700 4548
rect 3752 4536 3758 4548
rect 4062 4536 4068 4548
rect 3752 4508 4068 4536
rect 3752 4496 3758 4508
rect 4062 4496 4068 4508
rect 4120 4536 4126 4548
rect 5644 4536 5672 4567
rect 5994 4564 6000 4616
rect 6052 4604 6058 4616
rect 6089 4607 6147 4613
rect 6089 4604 6101 4607
rect 6052 4576 6101 4604
rect 6052 4564 6058 4576
rect 6089 4573 6101 4576
rect 6135 4573 6147 4607
rect 6546 4604 6552 4616
rect 6507 4576 6552 4604
rect 6089 4567 6147 4573
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 6822 4564 6828 4616
rect 6880 4604 6886 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6880 4576 7021 4604
rect 6880 4564 6886 4576
rect 7009 4573 7021 4576
rect 7055 4604 7067 4607
rect 7374 4604 7380 4616
rect 7055 4576 7380 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 7374 4564 7380 4576
rect 7432 4564 7438 4616
rect 7484 4604 7512 4644
rect 7650 4632 7656 4644
rect 7708 4632 7714 4684
rect 8662 4632 8668 4684
rect 8720 4672 8726 4684
rect 9309 4675 9367 4681
rect 9309 4672 9321 4675
rect 8720 4644 9321 4672
rect 8720 4632 8726 4644
rect 9309 4641 9321 4644
rect 9355 4641 9367 4675
rect 12342 4672 12348 4684
rect 12303 4644 12348 4672
rect 9309 4635 9367 4641
rect 12342 4632 12348 4644
rect 12400 4632 12406 4684
rect 13173 4675 13231 4681
rect 13173 4641 13185 4675
rect 13219 4641 13231 4675
rect 13173 4635 13231 4641
rect 8202 4604 8208 4616
rect 7484 4576 8208 4604
rect 8202 4564 8208 4576
rect 8260 4564 8266 4616
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4604 8631 4607
rect 9214 4604 9220 4616
rect 8619 4576 9220 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 9214 4564 9220 4576
rect 9272 4564 9278 4616
rect 10686 4564 10692 4616
rect 10744 4604 10750 4616
rect 12078 4607 12136 4613
rect 12078 4604 12090 4607
rect 10744 4576 12090 4604
rect 10744 4564 10750 4576
rect 12078 4573 12090 4576
rect 12124 4604 12136 4607
rect 12986 4604 12992 4616
rect 12124 4576 12296 4604
rect 12947 4576 12992 4604
rect 12124 4573 12136 4576
rect 12078 4567 12136 4573
rect 4120 4508 5672 4536
rect 4120 4496 4126 4508
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 1949 4471 2007 4477
rect 1949 4437 1961 4471
rect 1995 4468 2007 4471
rect 2130 4468 2136 4480
rect 1995 4440 2136 4468
rect 1995 4437 2007 4440
rect 1949 4431 2007 4437
rect 2130 4428 2136 4440
rect 2188 4428 2194 4480
rect 2314 4468 2320 4480
rect 2275 4440 2320 4468
rect 2314 4428 2320 4440
rect 2372 4428 2378 4480
rect 2866 4428 2872 4480
rect 2924 4468 2930 4480
rect 2961 4471 3019 4477
rect 2961 4468 2973 4471
rect 2924 4440 2973 4468
rect 2924 4428 2930 4440
rect 2961 4437 2973 4440
rect 3007 4437 3019 4471
rect 2961 4431 3019 4437
rect 4430 4428 4436 4480
rect 4488 4468 4494 4480
rect 4614 4468 4620 4480
rect 4488 4440 4620 4468
rect 4488 4428 4494 4440
rect 4614 4428 4620 4440
rect 4672 4468 4678 4480
rect 4893 4471 4951 4477
rect 4893 4468 4905 4471
rect 4672 4440 4905 4468
rect 4672 4428 4678 4440
rect 4893 4437 4905 4440
rect 4939 4468 4951 4471
rect 4982 4468 4988 4480
rect 4939 4440 4988 4468
rect 4939 4437 4951 4440
rect 4893 4431 4951 4437
rect 4982 4428 4988 4440
rect 5040 4428 5046 4480
rect 5644 4468 5672 4508
rect 6362 4496 6368 4548
rect 6420 4536 6426 4548
rect 7929 4539 7987 4545
rect 6420 4508 7880 4536
rect 6420 4496 6426 4508
rect 6546 4468 6552 4480
rect 5644 4440 6552 4468
rect 6546 4428 6552 4440
rect 6604 4428 6610 4480
rect 7852 4468 7880 4508
rect 7929 4505 7941 4539
rect 7975 4536 7987 4539
rect 9398 4536 9404 4548
rect 7975 4508 9404 4536
rect 7975 4505 7987 4508
rect 7929 4499 7987 4505
rect 9398 4496 9404 4508
rect 9456 4496 9462 4548
rect 9576 4539 9634 4545
rect 9576 4505 9588 4539
rect 9622 4536 9634 4539
rect 11882 4536 11888 4548
rect 9622 4508 11888 4536
rect 9622 4505 9634 4508
rect 9576 4499 9634 4505
rect 11882 4496 11888 4508
rect 11940 4496 11946 4548
rect 12268 4536 12296 4576
rect 12986 4564 12992 4576
rect 13044 4564 13050 4616
rect 13188 4536 13216 4635
rect 14090 4604 14096 4616
rect 14051 4576 14096 4604
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 14200 4604 14228 4780
rect 16206 4768 16212 4820
rect 16264 4808 16270 4820
rect 17862 4808 17868 4820
rect 16264 4780 16988 4808
rect 17823 4780 17868 4808
rect 16264 4768 16270 4780
rect 14277 4743 14335 4749
rect 14277 4709 14289 4743
rect 14323 4740 14335 4743
rect 15470 4740 15476 4752
rect 14323 4712 15476 4740
rect 14323 4709 14335 4712
rect 14277 4703 14335 4709
rect 15470 4700 15476 4712
rect 15528 4700 15534 4752
rect 16577 4743 16635 4749
rect 16577 4709 16589 4743
rect 16623 4709 16635 4743
rect 16850 4740 16856 4752
rect 16811 4712 16856 4740
rect 16577 4703 16635 4709
rect 15013 4675 15071 4681
rect 15013 4641 15025 4675
rect 15059 4672 15071 4675
rect 15194 4672 15200 4684
rect 15059 4644 15200 4672
rect 15059 4641 15071 4644
rect 15013 4635 15071 4641
rect 15194 4632 15200 4644
rect 15252 4632 15258 4684
rect 15930 4672 15936 4684
rect 15891 4644 15936 4672
rect 15930 4632 15936 4644
rect 15988 4632 15994 4684
rect 16592 4672 16620 4703
rect 16850 4700 16856 4712
rect 16908 4700 16914 4752
rect 16960 4740 16988 4780
rect 17862 4768 17868 4780
rect 17920 4768 17926 4820
rect 19058 4740 19064 4752
rect 16960 4712 19064 4740
rect 19058 4700 19064 4712
rect 19116 4700 19122 4752
rect 16592 4644 16896 4672
rect 15105 4607 15163 4613
rect 15105 4604 15117 4607
rect 14200 4576 15117 4604
rect 15105 4573 15117 4576
rect 15151 4573 15163 4607
rect 15105 4567 15163 4573
rect 15488 4576 16344 4604
rect 12268 4508 13216 4536
rect 13262 4496 13268 4548
rect 13320 4536 13326 4548
rect 14734 4536 14740 4548
rect 13320 4508 14740 4536
rect 13320 4496 13326 4508
rect 14734 4496 14740 4508
rect 14792 4496 14798 4548
rect 15010 4496 15016 4548
rect 15068 4536 15074 4548
rect 15488 4536 15516 4576
rect 16209 4539 16267 4545
rect 16209 4536 16221 4539
rect 15068 4508 15516 4536
rect 15580 4508 16221 4536
rect 15068 4496 15074 4508
rect 8478 4468 8484 4480
rect 7852 4440 8484 4468
rect 8478 4428 8484 4440
rect 8536 4428 8542 4480
rect 9033 4471 9091 4477
rect 9033 4437 9045 4471
rect 9079 4468 9091 4471
rect 9122 4468 9128 4480
rect 9079 4440 9128 4468
rect 9079 4437 9091 4440
rect 9033 4431 9091 4437
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 10226 4428 10232 4480
rect 10284 4468 10290 4480
rect 10686 4468 10692 4480
rect 10284 4440 10692 4468
rect 10284 4428 10290 4440
rect 10686 4428 10692 4440
rect 10744 4428 10750 4480
rect 10962 4468 10968 4480
rect 10923 4440 10968 4468
rect 10962 4428 10968 4440
rect 11020 4428 11026 4480
rect 11054 4428 11060 4480
rect 11112 4468 11118 4480
rect 12621 4471 12679 4477
rect 12621 4468 12633 4471
rect 11112 4440 12633 4468
rect 11112 4428 11118 4440
rect 12621 4437 12633 4440
rect 12667 4437 12679 4471
rect 13078 4468 13084 4480
rect 13039 4440 13084 4468
rect 12621 4431 12679 4437
rect 13078 4428 13084 4440
rect 13136 4428 13142 4480
rect 14274 4428 14280 4480
rect 14332 4468 14338 4480
rect 15580 4477 15608 4508
rect 16209 4505 16221 4508
rect 16255 4505 16267 4539
rect 16209 4499 16267 4505
rect 15197 4471 15255 4477
rect 15197 4468 15209 4471
rect 14332 4440 15209 4468
rect 14332 4428 14338 4440
rect 15197 4437 15209 4440
rect 15243 4437 15255 4471
rect 15197 4431 15255 4437
rect 15565 4471 15623 4477
rect 15565 4437 15577 4471
rect 15611 4437 15623 4471
rect 16114 4468 16120 4480
rect 16075 4440 16120 4468
rect 15565 4431 15623 4437
rect 16114 4428 16120 4440
rect 16172 4428 16178 4480
rect 16316 4468 16344 4576
rect 16868 4536 16896 4644
rect 16942 4632 16948 4684
rect 17000 4672 17006 4684
rect 17405 4675 17463 4681
rect 17405 4672 17417 4675
rect 17000 4644 17417 4672
rect 17000 4632 17006 4644
rect 17405 4641 17417 4644
rect 17451 4641 17463 4675
rect 17405 4635 17463 4641
rect 18509 4675 18567 4681
rect 18509 4641 18521 4675
rect 18555 4672 18567 4675
rect 18598 4672 18604 4684
rect 18555 4644 18604 4672
rect 18555 4641 18567 4644
rect 18509 4635 18567 4641
rect 18598 4632 18604 4644
rect 18656 4632 18662 4684
rect 18966 4632 18972 4684
rect 19024 4672 19030 4684
rect 19245 4675 19303 4681
rect 19245 4672 19257 4675
rect 19024 4644 19257 4672
rect 19024 4632 19030 4644
rect 19245 4641 19257 4644
rect 19291 4641 19303 4675
rect 19245 4635 19303 4641
rect 17678 4564 17684 4616
rect 17736 4604 17742 4616
rect 18414 4604 18420 4616
rect 17736 4576 18420 4604
rect 17736 4564 17742 4576
rect 18414 4564 18420 4576
rect 18472 4564 18478 4616
rect 20898 4604 20904 4616
rect 20859 4576 20904 4604
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 17313 4539 17371 4545
rect 17313 4536 17325 4539
rect 16868 4508 17325 4536
rect 17313 4505 17325 4508
rect 17359 4505 17371 4539
rect 17313 4499 17371 4505
rect 17862 4496 17868 4548
rect 17920 4536 17926 4548
rect 19512 4539 19570 4545
rect 17920 4508 19334 4536
rect 17920 4496 17926 4508
rect 17221 4471 17279 4477
rect 17221 4468 17233 4471
rect 16316 4440 17233 4468
rect 17221 4437 17233 4440
rect 17267 4437 17279 4471
rect 17221 4431 17279 4437
rect 17954 4428 17960 4480
rect 18012 4468 18018 4480
rect 18233 4471 18291 4477
rect 18233 4468 18245 4471
rect 18012 4440 18245 4468
rect 18012 4428 18018 4440
rect 18233 4437 18245 4440
rect 18279 4437 18291 4471
rect 18233 4431 18291 4437
rect 18322 4428 18328 4480
rect 18380 4468 18386 4480
rect 19306 4468 19334 4508
rect 19512 4505 19524 4539
rect 19558 4536 19570 4539
rect 19794 4536 19800 4548
rect 19558 4508 19800 4536
rect 19558 4505 19570 4508
rect 19512 4499 19570 4505
rect 19794 4496 19800 4508
rect 19852 4496 19858 4548
rect 20625 4471 20683 4477
rect 20625 4468 20637 4471
rect 18380 4440 18425 4468
rect 19306 4440 20637 4468
rect 18380 4428 18386 4440
rect 20625 4437 20637 4440
rect 20671 4437 20683 4471
rect 20625 4431 20683 4437
rect 20990 4428 20996 4480
rect 21048 4468 21054 4480
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 21048 4440 21097 4468
rect 21048 4428 21054 4440
rect 21085 4437 21097 4440
rect 21131 4437 21143 4471
rect 21085 4431 21143 4437
rect 1104 4378 21896 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21896 4378
rect 1104 4304 21896 4326
rect 2593 4267 2651 4273
rect 2593 4233 2605 4267
rect 2639 4264 2651 4267
rect 2639 4236 5672 4264
rect 2639 4233 2651 4236
rect 2593 4227 2651 4233
rect 3694 4196 3700 4208
rect 3655 4168 3700 4196
rect 3694 4156 3700 4168
rect 3752 4156 3758 4208
rect 4798 4156 4804 4208
rect 4856 4196 4862 4208
rect 5644 4196 5672 4236
rect 5718 4224 5724 4276
rect 5776 4264 5782 4276
rect 11977 4267 12035 4273
rect 5776 4236 9168 4264
rect 5776 4224 5782 4236
rect 5810 4196 5816 4208
rect 4856 4168 5396 4196
rect 5644 4168 5816 4196
rect 4856 4156 4862 4168
rect 1489 4131 1547 4137
rect 1489 4097 1501 4131
rect 1535 4128 1547 4131
rect 2038 4128 2044 4140
rect 1535 4100 2044 4128
rect 1535 4097 1547 4100
rect 1489 4091 1547 4097
rect 2038 4088 2044 4100
rect 2096 4088 2102 4140
rect 2225 4131 2283 4137
rect 2225 4097 2237 4131
rect 2271 4128 2283 4131
rect 2590 4128 2596 4140
rect 2271 4100 2596 4128
rect 2271 4097 2283 4100
rect 2225 4091 2283 4097
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 3878 4088 3884 4140
rect 3936 4128 3942 4140
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3936 4100 3985 4128
rect 3936 4088 3942 4100
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 4430 4128 4436 4140
rect 4391 4100 4436 4128
rect 3973 4091 4031 4097
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 5368 4137 5396 4168
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 6822 4196 6828 4208
rect 6783 4168 6828 4196
rect 6822 4156 6828 4168
rect 6880 4156 6886 4208
rect 7392 4168 8156 4196
rect 5069 4131 5127 4137
rect 5069 4097 5081 4131
rect 5115 4097 5127 4131
rect 5069 4091 5127 4097
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 3329 4063 3387 4069
rect 3329 4029 3341 4063
rect 3375 4060 3387 4063
rect 4062 4060 4068 4072
rect 3375 4032 4068 4060
rect 3375 4029 3387 4032
rect 3329 4023 3387 4029
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 1578 3952 1584 4004
rect 1636 3992 1642 4004
rect 4614 3992 4620 4004
rect 1636 3964 4016 3992
rect 4575 3964 4620 3992
rect 1636 3952 1642 3964
rect 3988 3936 4016 3964
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 5092 3936 5120 4091
rect 6362 4088 6368 4140
rect 6420 4128 6426 4140
rect 6914 4128 6920 4140
rect 6420 4100 6920 4128
rect 6420 4088 6426 4100
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7285 4131 7343 4137
rect 7285 4097 7297 4131
rect 7331 4128 7343 4131
rect 7392 4128 7420 4168
rect 7561 4131 7619 4137
rect 7561 4128 7573 4131
rect 7331 4100 7420 4128
rect 7484 4100 7573 4128
rect 7331 4097 7343 4100
rect 7285 4091 7343 4097
rect 5997 4063 6055 4069
rect 5997 4029 6009 4063
rect 6043 4060 6055 4063
rect 6546 4060 6552 4072
rect 6043 4032 6552 4060
rect 6043 4029 6055 4032
rect 5997 4023 6055 4029
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 7190 4020 7196 4072
rect 7248 4060 7254 4072
rect 7484 4060 7512 4100
rect 7561 4097 7573 4100
rect 7607 4097 7619 4131
rect 7561 4091 7619 4097
rect 8128 4060 8156 4168
rect 8754 4156 8760 4208
rect 8812 4196 8818 4208
rect 9140 4205 9168 4236
rect 11977 4233 11989 4267
rect 12023 4264 12035 4267
rect 12250 4264 12256 4276
rect 12023 4236 12256 4264
rect 12023 4233 12035 4236
rect 11977 4227 12035 4233
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 12621 4267 12679 4273
rect 12621 4233 12633 4267
rect 12667 4264 12679 4267
rect 13078 4264 13084 4276
rect 12667 4236 13084 4264
rect 12667 4233 12679 4236
rect 12621 4227 12679 4233
rect 13078 4224 13084 4236
rect 13136 4224 13142 4276
rect 14182 4264 14188 4276
rect 14143 4236 14188 4264
rect 14182 4224 14188 4236
rect 14240 4224 14246 4276
rect 15197 4267 15255 4273
rect 15197 4233 15209 4267
rect 15243 4264 15255 4267
rect 15286 4264 15292 4276
rect 15243 4236 15292 4264
rect 15243 4233 15255 4236
rect 15197 4227 15255 4233
rect 15286 4224 15292 4236
rect 15344 4224 15350 4276
rect 15565 4267 15623 4273
rect 15565 4233 15577 4267
rect 15611 4264 15623 4267
rect 16114 4264 16120 4276
rect 15611 4236 16120 4264
rect 15611 4233 15623 4236
rect 15565 4227 15623 4233
rect 16114 4224 16120 4236
rect 16172 4224 16178 4276
rect 17497 4267 17555 4273
rect 17497 4233 17509 4267
rect 17543 4264 17555 4267
rect 17678 4264 17684 4276
rect 17543 4236 17684 4264
rect 17543 4233 17555 4236
rect 17497 4227 17555 4233
rect 17678 4224 17684 4236
rect 17736 4224 17742 4276
rect 17957 4267 18015 4273
rect 17957 4233 17969 4267
rect 18003 4264 18015 4267
rect 18322 4264 18328 4276
rect 18003 4236 18328 4264
rect 18003 4233 18015 4236
rect 17957 4227 18015 4233
rect 18322 4224 18328 4236
rect 18380 4224 18386 4276
rect 18966 4224 18972 4276
rect 19024 4224 19030 4276
rect 8941 4199 8999 4205
rect 8941 4196 8953 4199
rect 8812 4168 8953 4196
rect 8812 4156 8818 4168
rect 8941 4165 8953 4168
rect 8987 4165 8999 4199
rect 8941 4159 8999 4165
rect 9125 4199 9183 4205
rect 9125 4165 9137 4199
rect 9171 4196 9183 4199
rect 10042 4196 10048 4208
rect 9171 4168 10048 4196
rect 9171 4165 9183 4168
rect 9125 4159 9183 4165
rect 10042 4156 10048 4168
rect 10100 4156 10106 4208
rect 10962 4196 10968 4208
rect 10152 4168 10968 4196
rect 8205 4131 8263 4137
rect 8205 4097 8217 4131
rect 8251 4128 8263 4131
rect 8386 4128 8392 4140
rect 8251 4100 8392 4128
rect 8251 4097 8263 4100
rect 8205 4091 8263 4097
rect 8386 4088 8392 4100
rect 8444 4088 8450 4140
rect 8481 4131 8539 4137
rect 8481 4097 8493 4131
rect 8527 4128 8539 4131
rect 8662 4128 8668 4140
rect 8527 4100 8668 4128
rect 8527 4097 8539 4100
rect 8481 4091 8539 4097
rect 8662 4088 8668 4100
rect 8720 4088 8726 4140
rect 9490 4128 9496 4140
rect 9451 4100 9496 4128
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 10152 4137 10180 4168
rect 10962 4156 10968 4168
rect 11020 4156 11026 4208
rect 12986 4196 12992 4208
rect 11992 4168 12434 4196
rect 12947 4168 12992 4196
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4097 10195 4131
rect 10778 4128 10784 4140
rect 10739 4100 10784 4128
rect 10137 4091 10195 4097
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 10873 4131 10931 4137
rect 10873 4097 10885 4131
rect 10919 4128 10931 4131
rect 11054 4128 11060 4140
rect 10919 4100 11060 4128
rect 10919 4097 10931 4100
rect 10873 4091 10931 4097
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 7248 4032 7512 4060
rect 7576 4032 7972 4060
rect 8128 4032 10456 4060
rect 7248 4020 7254 4032
rect 5442 3952 5448 4004
rect 5500 3992 5506 4004
rect 7576 3992 7604 4032
rect 5500 3964 7604 3992
rect 7944 3992 7972 4032
rect 9674 3992 9680 4004
rect 7944 3964 9680 3992
rect 5500 3952 5506 3964
rect 9674 3952 9680 3964
rect 9732 3952 9738 4004
rect 10428 4001 10456 4032
rect 10962 4020 10968 4072
rect 11020 4060 11026 4072
rect 11020 4032 11065 4060
rect 11020 4020 11026 4032
rect 11882 4020 11888 4072
rect 11940 4060 11946 4072
rect 11992 4060 12020 4168
rect 12066 4088 12072 4140
rect 12124 4128 12130 4140
rect 12406 4128 12434 4168
rect 12986 4156 12992 4168
rect 13044 4156 13050 4208
rect 13446 4156 13452 4208
rect 13504 4196 13510 4208
rect 15838 4196 15844 4208
rect 13504 4168 15844 4196
rect 13504 4156 13510 4168
rect 15838 4156 15844 4168
rect 15896 4156 15902 4208
rect 16025 4199 16083 4205
rect 16025 4165 16037 4199
rect 16071 4196 16083 4199
rect 17034 4196 17040 4208
rect 16071 4168 17040 4196
rect 16071 4165 16083 4168
rect 16025 4159 16083 4165
rect 17034 4156 17040 4168
rect 17092 4156 17098 4208
rect 17589 4199 17647 4205
rect 17589 4165 17601 4199
rect 17635 4196 17647 4199
rect 18046 4196 18052 4208
rect 17635 4168 18052 4196
rect 17635 4165 17647 4168
rect 17589 4159 17647 4165
rect 18046 4156 18052 4168
rect 18104 4156 18110 4208
rect 18984 4196 19012 4224
rect 18248 4168 19012 4196
rect 12894 4128 12900 4140
rect 12124 4100 12169 4128
rect 12406 4100 12900 4128
rect 12124 4088 12130 4100
rect 12894 4088 12900 4100
rect 12952 4128 12958 4140
rect 12952 4100 13216 4128
rect 12952 4088 12958 4100
rect 12161 4063 12219 4069
rect 12161 4060 12173 4063
rect 11940 4032 12173 4060
rect 11940 4020 11946 4032
rect 12161 4029 12173 4032
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 12250 4020 12256 4072
rect 12308 4060 12314 4072
rect 13188 4069 13216 4100
rect 13630 4088 13636 4140
rect 13688 4128 13694 4140
rect 15562 4128 15568 4140
rect 13688 4100 15568 4128
rect 13688 4088 13694 4100
rect 15562 4088 15568 4100
rect 15620 4088 15626 4140
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4128 16727 4131
rect 16942 4128 16948 4140
rect 16715 4100 16948 4128
rect 16715 4097 16727 4100
rect 16669 4091 16727 4097
rect 16942 4088 16948 4100
rect 17000 4088 17006 4140
rect 18248 4137 18276 4168
rect 19610 4156 19616 4208
rect 19668 4196 19674 4208
rect 19668 4168 20024 4196
rect 19668 4156 19674 4168
rect 18233 4131 18291 4137
rect 18233 4097 18245 4131
rect 18279 4097 18291 4131
rect 18233 4091 18291 4097
rect 18489 4131 18547 4137
rect 18489 4097 18501 4131
rect 18535 4128 18547 4131
rect 18966 4128 18972 4140
rect 18535 4100 18972 4128
rect 18535 4097 18547 4100
rect 18489 4091 18547 4097
rect 18966 4088 18972 4100
rect 19024 4088 19030 4140
rect 19886 4128 19892 4140
rect 19847 4100 19892 4128
rect 19886 4088 19892 4100
rect 19944 4088 19950 4140
rect 19996 4128 20024 4168
rect 20254 4156 20260 4208
rect 20312 4196 20318 4208
rect 20809 4199 20867 4205
rect 20809 4196 20821 4199
rect 20312 4168 20821 4196
rect 20312 4156 20318 4168
rect 20809 4165 20821 4168
rect 20855 4165 20867 4199
rect 20809 4159 20867 4165
rect 20070 4128 20076 4140
rect 19996 4100 20076 4128
rect 20070 4088 20076 4100
rect 20128 4088 20134 4140
rect 20346 4088 20352 4140
rect 20404 4128 20410 4140
rect 21266 4128 21272 4140
rect 20404 4100 21272 4128
rect 20404 4088 20410 4100
rect 21266 4088 21272 4100
rect 21324 4088 21330 4140
rect 13081 4063 13139 4069
rect 13081 4060 13093 4063
rect 12308 4032 13093 4060
rect 12308 4020 12314 4032
rect 13081 4029 13093 4032
rect 13127 4029 13139 4063
rect 13081 4023 13139 4029
rect 13173 4063 13231 4069
rect 13173 4029 13185 4063
rect 13219 4029 13231 4063
rect 14274 4060 14280 4072
rect 14235 4032 14280 4060
rect 13173 4023 13231 4029
rect 14274 4020 14280 4032
rect 14332 4020 14338 4072
rect 14461 4063 14519 4069
rect 14461 4029 14473 4063
rect 14507 4029 14519 4063
rect 14461 4023 14519 4029
rect 15013 4063 15071 4069
rect 15013 4029 15025 4063
rect 15059 4029 15071 4063
rect 15013 4023 15071 4029
rect 15105 4063 15163 4069
rect 15105 4029 15117 4063
rect 15151 4060 15163 4063
rect 15286 4060 15292 4072
rect 15151 4032 15292 4060
rect 15151 4029 15163 4032
rect 15105 4023 15163 4029
rect 10413 3995 10471 4001
rect 10413 3961 10425 3995
rect 10459 3961 10471 3995
rect 10413 3955 10471 3961
rect 11054 3952 11060 4004
rect 11112 3992 11118 4004
rect 14366 3992 14372 4004
rect 11112 3964 14372 3992
rect 11112 3952 11118 3964
rect 14366 3952 14372 3964
rect 14424 3992 14430 4004
rect 14476 3992 14504 4023
rect 14424 3964 14504 3992
rect 15028 3992 15056 4023
rect 15286 4020 15292 4032
rect 15344 4020 15350 4072
rect 15654 4020 15660 4072
rect 15712 4060 15718 4072
rect 15841 4063 15899 4069
rect 15841 4060 15853 4063
rect 15712 4032 15853 4060
rect 15712 4020 15718 4032
rect 15841 4029 15853 4032
rect 15887 4029 15899 4063
rect 15841 4023 15899 4029
rect 17313 4063 17371 4069
rect 17313 4029 17325 4063
rect 17359 4029 17371 4063
rect 20898 4060 20904 4072
rect 17313 4023 17371 4029
rect 19536 4032 20760 4060
rect 20859 4032 20904 4060
rect 15194 3992 15200 4004
rect 15028 3964 15200 3992
rect 14424 3952 14430 3964
rect 15194 3952 15200 3964
rect 15252 3952 15258 4004
rect 17328 3992 17356 4023
rect 17862 3992 17868 4004
rect 15304 3964 17868 3992
rect 1854 3924 1860 3936
rect 1815 3896 1860 3924
rect 1854 3884 1860 3896
rect 1912 3884 1918 3936
rect 2961 3927 3019 3933
rect 2961 3893 2973 3927
rect 3007 3924 3019 3927
rect 3142 3924 3148 3936
rect 3007 3896 3148 3924
rect 3007 3893 3019 3896
rect 2961 3887 3019 3893
rect 3142 3884 3148 3896
rect 3200 3884 3206 3936
rect 3970 3884 3976 3936
rect 4028 3884 4034 3936
rect 4157 3927 4215 3933
rect 4157 3893 4169 3927
rect 4203 3924 4215 3927
rect 4798 3924 4804 3936
rect 4203 3896 4804 3924
rect 4203 3893 4215 3896
rect 4157 3887 4215 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 4890 3884 4896 3936
rect 4948 3924 4954 3936
rect 4948 3896 4993 3924
rect 4948 3884 4954 3896
rect 5074 3884 5080 3936
rect 5132 3884 5138 3936
rect 5537 3927 5595 3933
rect 5537 3893 5549 3927
rect 5583 3924 5595 3927
rect 5718 3924 5724 3936
rect 5583 3896 5724 3924
rect 5583 3893 5595 3896
rect 5537 3887 5595 3893
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 7101 3927 7159 3933
rect 7101 3924 7113 3927
rect 6788 3896 7113 3924
rect 6788 3884 6794 3896
rect 7101 3893 7113 3896
rect 7147 3893 7159 3927
rect 7101 3887 7159 3893
rect 7650 3884 7656 3936
rect 7708 3924 7714 3936
rect 7745 3927 7803 3933
rect 7745 3924 7757 3927
rect 7708 3896 7757 3924
rect 7708 3884 7714 3896
rect 7745 3893 7757 3896
rect 7791 3893 7803 3927
rect 8018 3924 8024 3936
rect 7979 3896 8024 3924
rect 7745 3887 7803 3893
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 8665 3927 8723 3933
rect 8665 3893 8677 3927
rect 8711 3924 8723 3927
rect 9766 3924 9772 3936
rect 8711 3896 9772 3924
rect 8711 3893 8723 3896
rect 8665 3887 8723 3893
rect 9766 3884 9772 3896
rect 9824 3884 9830 3936
rect 10502 3884 10508 3936
rect 10560 3924 10566 3936
rect 11609 3927 11667 3933
rect 11609 3924 11621 3927
rect 10560 3896 11621 3924
rect 10560 3884 10566 3896
rect 11609 3893 11621 3896
rect 11655 3893 11667 3927
rect 11609 3887 11667 3893
rect 13817 3927 13875 3933
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 14458 3924 14464 3936
rect 13863 3896 14464 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 15102 3884 15108 3936
rect 15160 3924 15166 3936
rect 15304 3924 15332 3964
rect 17862 3952 17868 3964
rect 17920 3952 17926 4004
rect 15160 3896 15332 3924
rect 15160 3884 15166 3896
rect 15378 3884 15384 3936
rect 15436 3924 15442 3936
rect 16482 3924 16488 3936
rect 15436 3896 16488 3924
rect 15436 3884 15442 3896
rect 16482 3884 16488 3896
rect 16540 3884 16546 3936
rect 16853 3927 16911 3933
rect 16853 3893 16865 3927
rect 16899 3924 16911 3927
rect 19536 3924 19564 4032
rect 19702 3952 19708 4004
rect 19760 3992 19766 4004
rect 20441 3995 20499 4001
rect 20441 3992 20453 3995
rect 19760 3964 20453 3992
rect 19760 3952 19766 3964
rect 20441 3961 20453 3964
rect 20487 3961 20499 3995
rect 20732 3992 20760 4032
rect 20898 4020 20904 4032
rect 20956 4020 20962 4072
rect 21082 4060 21088 4072
rect 21043 4032 21088 4060
rect 21082 4020 21088 4032
rect 21140 4020 21146 4072
rect 21542 3992 21548 4004
rect 20732 3964 21548 3992
rect 20441 3955 20499 3961
rect 21542 3952 21548 3964
rect 21600 3952 21606 4004
rect 16899 3896 19564 3924
rect 19613 3927 19671 3933
rect 16899 3893 16911 3896
rect 16853 3887 16911 3893
rect 19613 3893 19625 3927
rect 19659 3924 19671 3927
rect 19794 3924 19800 3936
rect 19659 3896 19800 3924
rect 19659 3893 19671 3896
rect 19613 3887 19671 3893
rect 19794 3884 19800 3896
rect 19852 3884 19858 3936
rect 20070 3924 20076 3936
rect 20031 3896 20076 3924
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 6457 3723 6515 3729
rect 6457 3689 6469 3723
rect 6503 3720 6515 3723
rect 7190 3720 7196 3732
rect 6503 3692 7196 3720
rect 6503 3689 6515 3692
rect 6457 3683 6515 3689
rect 7190 3680 7196 3692
rect 7248 3680 7254 3732
rect 7650 3680 7656 3732
rect 7708 3680 7714 3732
rect 7837 3723 7895 3729
rect 7837 3689 7849 3723
rect 7883 3720 7895 3723
rect 8110 3720 8116 3732
rect 7883 3692 8116 3720
rect 7883 3689 7895 3692
rect 7837 3683 7895 3689
rect 8110 3680 8116 3692
rect 8168 3680 8174 3732
rect 9122 3680 9128 3732
rect 9180 3720 9186 3732
rect 9858 3720 9864 3732
rect 9180 3692 9864 3720
rect 9180 3680 9186 3692
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 10778 3720 10784 3732
rect 10739 3692 10784 3720
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 11072 3692 12434 3720
rect 2593 3655 2651 3661
rect 2593 3621 2605 3655
rect 2639 3652 2651 3655
rect 3050 3652 3056 3664
rect 2639 3624 3056 3652
rect 2639 3621 2651 3624
rect 2593 3615 2651 3621
rect 3050 3612 3056 3624
rect 3108 3612 3114 3664
rect 3421 3655 3479 3661
rect 3421 3621 3433 3655
rect 3467 3652 3479 3655
rect 5442 3652 5448 3664
rect 3467 3624 5448 3652
rect 3467 3621 3479 3624
rect 3421 3615 3479 3621
rect 5442 3612 5448 3624
rect 5500 3612 5506 3664
rect 5997 3655 6055 3661
rect 5997 3621 6009 3655
rect 6043 3652 6055 3655
rect 6362 3652 6368 3664
rect 6043 3624 6368 3652
rect 6043 3621 6055 3624
rect 5997 3615 6055 3621
rect 6362 3612 6368 3624
rect 6420 3612 6426 3664
rect 6917 3655 6975 3661
rect 6917 3621 6929 3655
rect 6963 3652 6975 3655
rect 7668 3652 7696 3680
rect 8481 3655 8539 3661
rect 6963 3624 7328 3652
rect 7668 3624 8441 3652
rect 6963 3621 6975 3624
rect 6917 3615 6975 3621
rect 4706 3584 4712 3596
rect 3252 3556 4712 3584
rect 1857 3519 1915 3525
rect 1857 3485 1869 3519
rect 1903 3516 1915 3519
rect 2314 3516 2320 3528
rect 1903 3488 2320 3516
rect 1903 3485 1915 3488
rect 1857 3479 1915 3485
rect 2314 3476 2320 3488
rect 2372 3476 2378 3528
rect 2682 3476 2688 3528
rect 2740 3516 2746 3528
rect 3252 3525 3280 3556
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 5258 3544 5264 3596
rect 5316 3544 5322 3596
rect 7300 3584 7328 3624
rect 8413 3584 8441 3624
rect 8481 3621 8493 3655
rect 8527 3652 8539 3655
rect 11072 3652 11100 3692
rect 8527 3624 11100 3652
rect 12406 3652 12434 3692
rect 12710 3680 12716 3732
rect 12768 3720 12774 3732
rect 13722 3720 13728 3732
rect 12768 3692 13728 3720
rect 12768 3680 12774 3692
rect 13722 3680 13728 3692
rect 13780 3680 13786 3732
rect 14366 3680 14372 3732
rect 14424 3720 14430 3732
rect 15473 3723 15531 3729
rect 15473 3720 15485 3723
rect 14424 3692 15485 3720
rect 14424 3680 14430 3692
rect 15473 3689 15485 3692
rect 15519 3689 15531 3723
rect 15473 3683 15531 3689
rect 15562 3680 15568 3732
rect 15620 3720 15626 3732
rect 18785 3723 18843 3729
rect 18785 3720 18797 3723
rect 15620 3692 18797 3720
rect 15620 3680 15626 3692
rect 18785 3689 18797 3692
rect 18831 3689 18843 3723
rect 18785 3683 18843 3689
rect 19886 3680 19892 3732
rect 19944 3720 19950 3732
rect 20806 3720 20812 3732
rect 19944 3692 20812 3720
rect 19944 3680 19950 3692
rect 20806 3680 20812 3692
rect 20864 3680 20870 3732
rect 20898 3680 20904 3732
rect 20956 3720 20962 3732
rect 21177 3723 21235 3729
rect 21177 3720 21189 3723
rect 20956 3692 21189 3720
rect 20956 3680 20962 3692
rect 21177 3689 21189 3692
rect 21223 3689 21235 3723
rect 21177 3683 21235 3689
rect 14090 3652 14096 3664
rect 12406 3624 14096 3652
rect 8527 3621 8539 3624
rect 8481 3615 8539 3621
rect 14090 3612 14096 3624
rect 14148 3612 14154 3664
rect 20070 3652 20076 3664
rect 17236 3624 20076 3652
rect 10226 3584 10232 3596
rect 7300 3556 8340 3584
rect 8413 3556 9674 3584
rect 10187 3556 10232 3584
rect 3237 3519 3295 3525
rect 3237 3516 3249 3519
rect 2740 3488 3249 3516
rect 2740 3476 2746 3488
rect 3237 3485 3249 3488
rect 3283 3485 3295 3519
rect 3970 3516 3976 3528
rect 3883 3488 3976 3516
rect 3237 3479 3295 3485
rect 3970 3476 3976 3488
rect 4028 3516 4034 3528
rect 4430 3516 4436 3528
rect 4028 3488 4436 3516
rect 4028 3476 4034 3488
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 4522 3476 4528 3528
rect 4580 3516 4586 3528
rect 4617 3519 4675 3525
rect 4617 3516 4629 3519
rect 4580 3488 4629 3516
rect 4580 3476 4586 3488
rect 4617 3485 4629 3488
rect 4663 3485 4675 3519
rect 4890 3516 4896 3528
rect 4851 3488 4896 3516
rect 4617 3479 4675 3485
rect 4890 3476 4896 3488
rect 4948 3476 4954 3528
rect 5276 3516 5304 3544
rect 5353 3519 5411 3525
rect 5353 3516 5365 3519
rect 5276 3488 5365 3516
rect 5353 3485 5365 3488
rect 5399 3485 5411 3519
rect 5353 3479 5411 3485
rect 5718 3476 5724 3528
rect 5776 3516 5782 3528
rect 5813 3519 5871 3525
rect 5813 3516 5825 3519
rect 5776 3488 5825 3516
rect 5776 3476 5782 3488
rect 5813 3485 5825 3488
rect 5859 3485 5871 3519
rect 6270 3516 6276 3528
rect 6231 3488 6276 3516
rect 5813 3479 5871 3485
rect 6270 3476 6276 3488
rect 6328 3476 6334 3528
rect 6730 3516 6736 3528
rect 6691 3488 6736 3516
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 8312 3525 8340 3556
rect 7193 3519 7251 3525
rect 7193 3485 7205 3519
rect 7239 3512 7251 3519
rect 8297 3519 8355 3525
rect 7300 3512 8055 3516
rect 7239 3488 8055 3512
rect 7239 3485 7328 3488
rect 7193 3484 7328 3485
rect 7193 3479 7251 3484
rect 2225 3451 2283 3457
rect 2225 3417 2237 3451
rect 2271 3448 2283 3451
rect 2961 3451 3019 3457
rect 2271 3420 2912 3448
rect 2271 3417 2283 3420
rect 2225 3411 2283 3417
rect 1489 3383 1547 3389
rect 1489 3349 1501 3383
rect 1535 3380 1547 3383
rect 2590 3380 2596 3392
rect 1535 3352 2596 3380
rect 1535 3349 1547 3352
rect 1489 3343 1547 3349
rect 2590 3340 2596 3352
rect 2648 3340 2654 3392
rect 2884 3380 2912 3420
rect 2961 3417 2973 3451
rect 3007 3448 3019 3451
rect 3694 3448 3700 3460
rect 3007 3420 3700 3448
rect 3007 3417 3019 3420
rect 2961 3411 3019 3417
rect 3694 3408 3700 3420
rect 3752 3408 3758 3460
rect 7745 3451 7803 3457
rect 7745 3448 7757 3451
rect 4080 3420 7757 3448
rect 4080 3380 4108 3420
rect 7576 3392 7604 3420
rect 7745 3417 7757 3420
rect 7791 3417 7803 3451
rect 8027 3448 8055 3488
rect 8297 3485 8309 3519
rect 8343 3485 8355 3519
rect 8297 3479 8355 3485
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 9214 3516 9220 3528
rect 8720 3488 9220 3516
rect 8720 3476 8726 3488
rect 9214 3476 9220 3488
rect 9272 3476 9278 3528
rect 8110 3448 8116 3460
rect 8027 3420 8116 3448
rect 7745 3411 7803 3417
rect 8110 3408 8116 3420
rect 8168 3408 8174 3460
rect 8386 3408 8392 3460
rect 8444 3448 8450 3460
rect 9306 3448 9312 3460
rect 8444 3420 9312 3448
rect 8444 3408 8450 3420
rect 9306 3408 9312 3420
rect 9364 3408 9370 3460
rect 2884 3352 4108 3380
rect 4157 3383 4215 3389
rect 4157 3349 4169 3383
rect 4203 3380 4215 3383
rect 4246 3380 4252 3392
rect 4203 3352 4252 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 4430 3380 4436 3392
rect 4391 3352 4436 3380
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 5077 3383 5135 3389
rect 5077 3349 5089 3383
rect 5123 3380 5135 3383
rect 5258 3380 5264 3392
rect 5123 3352 5264 3380
rect 5123 3349 5135 3352
rect 5077 3343 5135 3349
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5534 3380 5540 3392
rect 5495 3352 5540 3380
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 5718 3340 5724 3392
rect 5776 3380 5782 3392
rect 6730 3380 6736 3392
rect 5776 3352 6736 3380
rect 5776 3340 5782 3352
rect 6730 3340 6736 3352
rect 6788 3340 6794 3392
rect 7190 3340 7196 3392
rect 7248 3380 7254 3392
rect 7377 3383 7435 3389
rect 7377 3380 7389 3383
rect 7248 3352 7389 3380
rect 7248 3340 7254 3352
rect 7377 3349 7389 3352
rect 7423 3349 7435 3383
rect 7377 3343 7435 3349
rect 7558 3340 7564 3392
rect 7616 3340 7622 3392
rect 7650 3340 7656 3392
rect 7708 3380 7714 3392
rect 8938 3380 8944 3392
rect 7708 3352 8944 3380
rect 7708 3340 7714 3352
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 9122 3380 9128 3392
rect 9083 3352 9128 3380
rect 9122 3340 9128 3352
rect 9180 3340 9186 3392
rect 9646 3380 9674 3556
rect 10226 3544 10232 3556
rect 10284 3544 10290 3596
rect 10321 3587 10379 3593
rect 10321 3553 10333 3587
rect 10367 3584 10379 3587
rect 10502 3584 10508 3596
rect 10367 3556 10508 3584
rect 10367 3553 10379 3556
rect 10321 3547 10379 3553
rect 10502 3544 10508 3556
rect 10560 3544 10566 3596
rect 12894 3544 12900 3596
rect 12952 3584 12958 3596
rect 13081 3587 13139 3593
rect 13081 3584 13093 3587
rect 12952 3556 13093 3584
rect 12952 3544 12958 3556
rect 13081 3553 13093 3556
rect 13127 3584 13139 3587
rect 13170 3584 13176 3596
rect 13127 3556 13176 3584
rect 13127 3553 13139 3556
rect 13081 3547 13139 3553
rect 13170 3544 13176 3556
rect 13228 3544 13234 3596
rect 9766 3516 9772 3528
rect 9727 3488 9772 3516
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 10134 3476 10140 3528
rect 10192 3516 10198 3528
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 10192 3488 10425 3516
rect 10192 3476 10198 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 11057 3519 11115 3525
rect 11057 3485 11069 3519
rect 11103 3516 11115 3519
rect 11146 3516 11152 3528
rect 11103 3488 11152 3516
rect 11103 3485 11115 3488
rect 11057 3479 11115 3485
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 11324 3519 11382 3525
rect 11324 3485 11336 3519
rect 11370 3516 11382 3519
rect 11606 3516 11612 3528
rect 11370 3488 11612 3516
rect 11370 3485 11382 3488
rect 11324 3479 11382 3485
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 13354 3516 13360 3528
rect 13315 3488 13360 3516
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 13596 3488 14105 3516
rect 13596 3476 13602 3488
rect 14093 3485 14105 3488
rect 14139 3516 14151 3519
rect 14642 3516 14648 3528
rect 14139 3488 14648 3516
rect 14139 3485 14151 3488
rect 14093 3479 14151 3485
rect 14642 3476 14648 3488
rect 14700 3476 14706 3528
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 15838 3516 15844 3528
rect 14792 3488 15844 3516
rect 14792 3476 14798 3488
rect 15838 3476 15844 3488
rect 15896 3476 15902 3528
rect 15933 3519 15991 3525
rect 15933 3485 15945 3519
rect 15979 3516 15991 3519
rect 17126 3516 17132 3528
rect 15979 3488 17132 3516
rect 15979 3485 15991 3488
rect 15933 3479 15991 3485
rect 11698 3408 11704 3460
rect 11756 3448 11762 3460
rect 14338 3451 14396 3457
rect 14338 3448 14350 3451
rect 11756 3420 14350 3448
rect 11756 3408 11762 3420
rect 14338 3417 14350 3420
rect 14384 3417 14396 3451
rect 14338 3411 14396 3417
rect 15562 3408 15568 3460
rect 15620 3448 15626 3460
rect 15948 3448 15976 3479
rect 17126 3476 17132 3488
rect 17184 3476 17190 3528
rect 16206 3457 16212 3460
rect 16200 3448 16212 3457
rect 15620 3420 15976 3448
rect 16167 3420 16212 3448
rect 15620 3408 15626 3420
rect 16200 3411 16212 3420
rect 16206 3408 16212 3411
rect 16264 3408 16270 3460
rect 16482 3408 16488 3460
rect 16540 3448 16546 3460
rect 17236 3448 17264 3624
rect 20070 3612 20076 3624
rect 20128 3612 20134 3664
rect 18141 3587 18199 3593
rect 18141 3584 18153 3587
rect 16540 3420 17264 3448
rect 17328 3556 18153 3584
rect 16540 3408 16546 3420
rect 12250 3380 12256 3392
rect 9646 3352 12256 3380
rect 12250 3340 12256 3352
rect 12308 3340 12314 3392
rect 12437 3383 12495 3389
rect 12437 3349 12449 3383
rect 12483 3380 12495 3383
rect 12526 3380 12532 3392
rect 12483 3352 12532 3380
rect 12483 3349 12495 3352
rect 12437 3343 12495 3349
rect 12526 3340 12532 3352
rect 12584 3340 12590 3392
rect 12802 3340 12808 3392
rect 12860 3380 12866 3392
rect 13265 3383 13323 3389
rect 13265 3380 13277 3383
rect 12860 3352 13277 3380
rect 12860 3340 12866 3352
rect 13265 3349 13277 3352
rect 13311 3349 13323 3383
rect 13722 3380 13728 3392
rect 13683 3352 13728 3380
rect 13265 3343 13323 3349
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 15654 3340 15660 3392
rect 15712 3380 15718 3392
rect 17328 3389 17356 3556
rect 18141 3553 18153 3556
rect 18187 3553 18199 3587
rect 18141 3547 18199 3553
rect 18414 3544 18420 3596
rect 18472 3584 18478 3596
rect 19150 3584 19156 3596
rect 18472 3556 19156 3584
rect 18472 3544 18478 3556
rect 19150 3544 19156 3556
rect 19208 3544 19214 3596
rect 19610 3544 19616 3596
rect 19668 3584 19674 3596
rect 19981 3587 20039 3593
rect 19668 3556 19932 3584
rect 19668 3544 19674 3556
rect 17957 3519 18015 3525
rect 17957 3485 17969 3519
rect 18003 3516 18015 3519
rect 18046 3516 18052 3528
rect 18003 3488 18052 3516
rect 18003 3485 18015 3488
rect 17957 3479 18015 3485
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 18506 3476 18512 3528
rect 18564 3516 18570 3528
rect 18601 3519 18659 3525
rect 18601 3516 18613 3519
rect 18564 3488 18613 3516
rect 18564 3476 18570 3488
rect 18601 3485 18613 3488
rect 18647 3485 18659 3519
rect 19797 3519 19855 3525
rect 19797 3516 19809 3519
rect 18601 3479 18659 3485
rect 18708 3488 19809 3516
rect 17494 3408 17500 3460
rect 17552 3448 17558 3460
rect 17552 3420 18276 3448
rect 17552 3408 17558 3420
rect 17313 3383 17371 3389
rect 17313 3380 17325 3383
rect 15712 3352 17325 3380
rect 15712 3340 15718 3352
rect 17313 3349 17325 3352
rect 17359 3349 17371 3383
rect 17586 3380 17592 3392
rect 17547 3352 17592 3380
rect 17313 3343 17371 3349
rect 17586 3340 17592 3352
rect 17644 3340 17650 3392
rect 18046 3340 18052 3392
rect 18104 3380 18110 3392
rect 18248 3380 18276 3420
rect 18414 3408 18420 3460
rect 18472 3448 18478 3460
rect 18708 3448 18736 3488
rect 19797 3485 19809 3488
rect 19843 3485 19855 3519
rect 19904 3516 19932 3556
rect 19981 3553 19993 3587
rect 20027 3584 20039 3587
rect 20530 3584 20536 3596
rect 20027 3556 20536 3584
rect 20027 3553 20039 3556
rect 19981 3547 20039 3553
rect 20530 3544 20536 3556
rect 20588 3544 20594 3596
rect 20625 3587 20683 3593
rect 20625 3553 20637 3587
rect 20671 3584 20683 3587
rect 20714 3584 20720 3596
rect 20671 3556 20720 3584
rect 20671 3553 20683 3556
rect 20625 3547 20683 3553
rect 20714 3544 20720 3556
rect 20772 3544 20778 3596
rect 20070 3516 20076 3528
rect 19904 3488 20076 3516
rect 19797 3479 19855 3485
rect 20070 3476 20076 3488
rect 20128 3476 20134 3528
rect 20809 3519 20867 3525
rect 20809 3485 20821 3519
rect 20855 3516 20867 3519
rect 21358 3516 21364 3528
rect 20855 3488 21364 3516
rect 20855 3485 20867 3488
rect 20809 3479 20867 3485
rect 21358 3476 21364 3488
rect 21416 3476 21422 3528
rect 18472 3420 18736 3448
rect 18472 3408 18478 3420
rect 19518 3408 19524 3460
rect 19576 3448 19582 3460
rect 19889 3451 19947 3457
rect 19889 3448 19901 3451
rect 19576 3420 19901 3448
rect 19576 3408 19582 3420
rect 19889 3417 19901 3420
rect 19935 3417 19947 3451
rect 19889 3411 19947 3417
rect 20717 3451 20775 3457
rect 20717 3417 20729 3451
rect 20763 3448 20775 3451
rect 22094 3448 22100 3460
rect 20763 3420 22100 3448
rect 20763 3417 20775 3420
rect 20717 3411 20775 3417
rect 22094 3408 22100 3420
rect 22152 3408 22158 3460
rect 19058 3380 19064 3392
rect 18104 3352 18149 3380
rect 18248 3352 19064 3380
rect 18104 3340 18110 3352
rect 19058 3340 19064 3352
rect 19116 3340 19122 3392
rect 19429 3383 19487 3389
rect 19429 3349 19441 3383
rect 19475 3380 19487 3383
rect 19610 3380 19616 3392
rect 19475 3352 19616 3380
rect 19475 3349 19487 3352
rect 19429 3343 19487 3349
rect 19610 3340 19616 3352
rect 19668 3340 19674 3392
rect 1104 3290 21896 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21896 3290
rect 1104 3216 21896 3238
rect 1762 3136 1768 3188
rect 1820 3176 1826 3188
rect 3421 3179 3479 3185
rect 1820 3148 3280 3176
rect 1820 3136 1826 3148
rect 1394 3040 1400 3052
rect 1307 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3040 1458 3052
rect 1670 3040 1676 3052
rect 1452 3012 1676 3040
rect 1452 3000 1458 3012
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 1857 3043 1915 3049
rect 1857 3009 1869 3043
rect 1903 3009 1915 3043
rect 1857 3003 1915 3009
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3040 2375 3043
rect 2498 3040 2504 3052
rect 2363 3012 2504 3040
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 842 2932 848 2984
rect 900 2972 906 2984
rect 1486 2972 1492 2984
rect 900 2944 1492 2972
rect 900 2932 906 2944
rect 1486 2932 1492 2944
rect 1544 2972 1550 2984
rect 1872 2972 1900 3003
rect 2498 3000 2504 3012
rect 2556 3000 2562 3052
rect 2774 3000 2780 3052
rect 2832 3040 2838 3052
rect 3252 3049 3280 3148
rect 3421 3145 3433 3179
rect 3467 3176 3479 3179
rect 3878 3176 3884 3188
rect 3467 3148 3884 3176
rect 3467 3145 3479 3148
rect 3421 3139 3479 3145
rect 3878 3136 3884 3148
rect 3936 3136 3942 3188
rect 4890 3176 4896 3188
rect 4448 3148 4896 3176
rect 3602 3068 3608 3120
rect 3660 3108 3666 3120
rect 3789 3111 3847 3117
rect 3789 3108 3801 3111
rect 3660 3080 3801 3108
rect 3660 3068 3666 3080
rect 3789 3077 3801 3080
rect 3835 3077 3847 3111
rect 3789 3071 3847 3077
rect 3237 3043 3295 3049
rect 2832 3012 2877 3040
rect 2832 3000 2838 3012
rect 3237 3009 3249 3043
rect 3283 3009 3295 3043
rect 3237 3003 3295 3009
rect 3878 3000 3884 3052
rect 3936 3040 3942 3052
rect 3973 3043 4031 3049
rect 3973 3040 3985 3043
rect 3936 3012 3985 3040
rect 3936 3000 3942 3012
rect 3973 3009 3985 3012
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 4338 3000 4344 3052
rect 4396 3040 4402 3052
rect 4448 3049 4476 3148
rect 4890 3136 4896 3148
rect 4948 3136 4954 3188
rect 5077 3179 5135 3185
rect 5077 3145 5089 3179
rect 5123 3176 5135 3179
rect 5166 3176 5172 3188
rect 5123 3148 5172 3176
rect 5123 3145 5135 3148
rect 5077 3139 5135 3145
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 8018 3176 8024 3188
rect 7668 3148 8024 3176
rect 4614 3068 4620 3120
rect 4672 3108 4678 3120
rect 4982 3108 4988 3120
rect 4672 3080 4988 3108
rect 4672 3068 4678 3080
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 7668 3108 7696 3148
rect 8018 3136 8024 3148
rect 8076 3136 8082 3188
rect 8297 3179 8355 3185
rect 8297 3145 8309 3179
rect 8343 3176 8355 3179
rect 8343 3148 8984 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 8662 3108 8668 3120
rect 5920 3080 6776 3108
rect 4433 3043 4491 3049
rect 4433 3040 4445 3043
rect 4396 3012 4445 3040
rect 4396 3000 4402 3012
rect 4433 3009 4445 3012
rect 4479 3009 4491 3043
rect 4433 3003 4491 3009
rect 4893 3043 4951 3049
rect 4893 3009 4905 3043
rect 4939 3009 4951 3043
rect 4893 3003 4951 3009
rect 1544 2944 1900 2972
rect 1544 2932 1550 2944
rect 2130 2932 2136 2984
rect 2188 2972 2194 2984
rect 4908 2972 4936 3003
rect 5166 3000 5172 3052
rect 5224 3040 5230 3052
rect 5353 3043 5411 3049
rect 5353 3040 5365 3043
rect 5224 3012 5365 3040
rect 5224 3000 5230 3012
rect 5353 3009 5365 3012
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 5813 3043 5871 3049
rect 5813 3009 5825 3043
rect 5859 3040 5871 3043
rect 5920 3040 5948 3080
rect 6641 3043 6699 3049
rect 6641 3040 6653 3043
rect 5859 3012 5948 3040
rect 6012 3012 6653 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 5718 2972 5724 2984
rect 2188 2944 5724 2972
rect 2188 2932 2194 2944
rect 5718 2932 5724 2944
rect 5776 2932 5782 2984
rect 6012 2972 6040 3012
rect 6641 3009 6653 3012
rect 6687 3009 6699 3043
rect 6748 3040 6776 3080
rect 7004 3080 7696 3108
rect 7944 3080 8668 3108
rect 7004 3040 7032 3080
rect 7282 3040 7288 3052
rect 6748 3012 7032 3040
rect 7243 3012 7288 3040
rect 6641 3003 6699 3009
rect 7282 3000 7288 3012
rect 7340 3000 7346 3052
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 7745 3044 7803 3049
rect 7745 3043 7880 3044
rect 7745 3009 7757 3043
rect 7791 3040 7880 3043
rect 7944 3040 7972 3080
rect 8662 3068 8668 3080
rect 8720 3068 8726 3120
rect 7791 3016 7972 3040
rect 7791 3009 7803 3016
rect 7852 3012 7972 3016
rect 7745 3003 7803 3009
rect 5920 2944 6040 2972
rect 5920 2916 5948 2944
rect 6822 2932 6828 2984
rect 6880 2972 6886 2984
rect 7576 2972 7604 3003
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 8113 3043 8171 3049
rect 8113 3040 8125 3043
rect 8076 3012 8125 3040
rect 8076 3000 8082 3012
rect 8113 3009 8125 3012
rect 8159 3009 8171 3043
rect 8113 3003 8171 3009
rect 7650 2972 7656 2984
rect 6880 2944 6925 2972
rect 7576 2944 7656 2972
rect 6880 2932 6886 2944
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 8956 2972 8984 3148
rect 9398 3136 9404 3188
rect 9456 3176 9462 3188
rect 11238 3176 11244 3188
rect 9456 3148 11244 3176
rect 9456 3136 9462 3148
rect 11238 3136 11244 3148
rect 11296 3136 11302 3188
rect 11609 3179 11667 3185
rect 11609 3145 11621 3179
rect 11655 3176 11667 3179
rect 11698 3176 11704 3188
rect 11655 3148 11704 3176
rect 11655 3145 11667 3148
rect 11609 3139 11667 3145
rect 11698 3136 11704 3148
rect 11756 3136 11762 3188
rect 14274 3176 14280 3188
rect 11808 3148 13676 3176
rect 14235 3148 14280 3176
rect 9030 3068 9036 3120
rect 9088 3108 9094 3120
rect 9950 3108 9956 3120
rect 9088 3080 9956 3108
rect 9088 3068 9094 3080
rect 9950 3068 9956 3080
rect 10008 3068 10014 3120
rect 10505 3111 10563 3117
rect 10505 3077 10517 3111
rect 10551 3108 10563 3111
rect 11808 3108 11836 3148
rect 10551 3080 11836 3108
rect 10551 3077 10563 3080
rect 10505 3071 10563 3077
rect 12710 3068 12716 3120
rect 12768 3068 12774 3120
rect 12897 3111 12955 3117
rect 12897 3077 12909 3111
rect 12943 3108 12955 3111
rect 13078 3108 13084 3120
rect 12943 3080 13084 3108
rect 12943 3077 12955 3080
rect 12897 3071 12955 3077
rect 13078 3068 13084 3080
rect 13136 3068 13142 3120
rect 13648 3108 13676 3148
rect 14274 3136 14280 3148
rect 14332 3136 14338 3188
rect 15746 3136 15752 3188
rect 15804 3176 15810 3188
rect 15804 3148 18736 3176
rect 15804 3136 15810 3148
rect 14890 3111 14948 3117
rect 14890 3108 14902 3111
rect 13648 3080 14902 3108
rect 14890 3077 14902 3080
rect 14936 3077 14948 3111
rect 14890 3071 14948 3077
rect 15010 3068 15016 3120
rect 15068 3108 15074 3120
rect 17282 3111 17340 3117
rect 17282 3108 17294 3111
rect 15068 3080 17294 3108
rect 15068 3068 15074 3080
rect 17282 3077 17294 3080
rect 17328 3077 17340 3111
rect 17282 3071 17340 3077
rect 17402 3068 17408 3120
rect 17460 3068 17466 3120
rect 9309 3043 9367 3049
rect 9309 3009 9321 3043
rect 9355 3040 9367 3043
rect 9398 3040 9404 3052
rect 9355 3012 9404 3040
rect 9355 3009 9367 3012
rect 9309 3003 9367 3009
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 9582 3000 9588 3052
rect 9640 3040 9646 3052
rect 10226 3040 10232 3052
rect 9640 3012 9685 3040
rect 10187 3012 10232 3040
rect 9640 3000 9646 3012
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11149 3043 11207 3049
rect 11149 3040 11161 3043
rect 11112 3012 11161 3040
rect 11112 3000 11118 3012
rect 11149 3009 11161 3012
rect 11195 3009 11207 3043
rect 11149 3003 11207 3009
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 11882 3040 11888 3052
rect 11296 3012 11888 3040
rect 11296 3000 11302 3012
rect 11882 3000 11888 3012
rect 11940 3000 11946 3052
rect 12253 3043 12311 3049
rect 12253 3009 12265 3043
rect 12299 3040 12311 3043
rect 12526 3040 12532 3052
rect 12299 3012 12532 3040
rect 12299 3009 12311 3012
rect 12253 3003 12311 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 12728 3040 12756 3068
rect 12805 3043 12863 3049
rect 12805 3040 12817 3043
rect 12728 3012 12817 3040
rect 12805 3009 12817 3012
rect 12851 3009 12863 3043
rect 13906 3040 13912 3052
rect 13867 3012 13912 3040
rect 12805 3003 12863 3009
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 14642 3040 14648 3052
rect 14603 3012 14648 3040
rect 14642 3000 14648 3012
rect 14700 3000 14706 3052
rect 15654 3000 15660 3052
rect 15712 3040 15718 3052
rect 17037 3043 17095 3049
rect 17037 3040 17049 3043
rect 15712 3012 17049 3040
rect 15712 3000 15718 3012
rect 17037 3009 17049 3012
rect 17083 3009 17095 3043
rect 17420 3040 17448 3068
rect 18708 3049 18736 3148
rect 19150 3136 19156 3188
rect 19208 3176 19214 3188
rect 20254 3176 20260 3188
rect 19208 3148 20024 3176
rect 20215 3148 20260 3176
rect 19208 3136 19214 3148
rect 17037 3003 17095 3009
rect 17144 3012 17448 3040
rect 18693 3043 18751 3049
rect 12434 2972 12440 2984
rect 8956 2944 12440 2972
rect 12434 2932 12440 2944
rect 12492 2932 12498 2984
rect 2590 2864 2596 2916
rect 2648 2904 2654 2916
rect 5902 2904 5908 2916
rect 2648 2876 5908 2904
rect 2648 2864 2654 2876
rect 5902 2864 5908 2876
rect 5960 2864 5966 2916
rect 5997 2907 6055 2913
rect 5997 2873 6009 2907
rect 6043 2904 6055 2907
rect 6914 2904 6920 2916
rect 6043 2876 6920 2904
rect 6043 2873 6055 2876
rect 5997 2867 6055 2873
rect 6914 2864 6920 2876
rect 6972 2864 6978 2916
rect 9030 2904 9036 2916
rect 7024 2876 9036 2904
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 2038 2836 2044 2848
rect 1999 2808 2044 2836
rect 2038 2796 2044 2808
rect 2096 2796 2102 2848
rect 2501 2839 2559 2845
rect 2501 2805 2513 2839
rect 2547 2836 2559 2839
rect 2682 2836 2688 2848
rect 2547 2808 2688 2836
rect 2547 2805 2559 2808
rect 2501 2799 2559 2805
rect 2682 2796 2688 2808
rect 2740 2796 2746 2848
rect 2958 2836 2964 2848
rect 2919 2808 2964 2836
rect 2958 2796 2964 2808
rect 3016 2796 3022 2848
rect 3878 2796 3884 2848
rect 3936 2836 3942 2848
rect 4062 2836 4068 2848
rect 3936 2808 4068 2836
rect 3936 2796 3942 2808
rect 4062 2796 4068 2808
rect 4120 2796 4126 2848
rect 4614 2836 4620 2848
rect 4575 2808 4620 2836
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 5537 2839 5595 2845
rect 5537 2805 5549 2839
rect 5583 2836 5595 2839
rect 5626 2836 5632 2848
rect 5583 2808 5632 2836
rect 5583 2805 5595 2808
rect 5537 2799 5595 2805
rect 5626 2796 5632 2808
rect 5684 2796 5690 2848
rect 5718 2796 5724 2848
rect 5776 2836 5782 2848
rect 7024 2836 7052 2876
rect 9030 2864 9036 2876
rect 9088 2864 9094 2916
rect 10226 2864 10232 2916
rect 10284 2904 10290 2916
rect 12342 2904 12348 2916
rect 10284 2876 12348 2904
rect 10284 2864 10290 2876
rect 12342 2864 12348 2876
rect 12400 2864 12406 2916
rect 5776 2808 7052 2836
rect 7101 2839 7159 2845
rect 5776 2796 5782 2808
rect 7101 2805 7113 2839
rect 7147 2836 7159 2839
rect 8110 2836 8116 2848
rect 7147 2808 8116 2836
rect 7147 2805 7159 2808
rect 7101 2799 7159 2805
rect 8110 2796 8116 2808
rect 8168 2796 8174 2848
rect 8665 2839 8723 2845
rect 8665 2805 8677 2839
rect 8711 2836 8723 2839
rect 11790 2836 11796 2848
rect 8711 2808 11796 2836
rect 8711 2805 8723 2808
rect 8665 2799 8723 2805
rect 11790 2796 11796 2808
rect 11848 2796 11854 2848
rect 12544 2836 12572 3000
rect 12621 2975 12679 2981
rect 12621 2941 12633 2975
rect 12667 2941 12679 2975
rect 13633 2975 13691 2981
rect 13633 2972 13645 2975
rect 12621 2935 12679 2941
rect 13004 2944 13645 2972
rect 12636 2904 12664 2935
rect 12894 2904 12900 2916
rect 12636 2876 12900 2904
rect 12894 2864 12900 2876
rect 12952 2864 12958 2916
rect 13004 2836 13032 2944
rect 13633 2941 13645 2944
rect 13679 2941 13691 2975
rect 13633 2935 13691 2941
rect 13817 2975 13875 2981
rect 13817 2941 13829 2975
rect 13863 2972 13875 2975
rect 14458 2972 14464 2984
rect 13863 2944 14464 2972
rect 13863 2941 13875 2944
rect 13817 2935 13875 2941
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 16761 2975 16819 2981
rect 16761 2941 16773 2975
rect 16807 2972 16819 2975
rect 17144 2972 17172 3012
rect 18693 3009 18705 3043
rect 18739 3009 18751 3043
rect 18693 3003 18751 3009
rect 19426 3000 19432 3052
rect 19484 3040 19490 3052
rect 19889 3043 19947 3049
rect 19889 3040 19901 3043
rect 19484 3012 19901 3040
rect 19484 3000 19490 3012
rect 19889 3009 19901 3012
rect 19935 3009 19947 3043
rect 19996 3040 20024 3148
rect 20254 3136 20260 3148
rect 20312 3136 20318 3188
rect 20809 3043 20867 3049
rect 20809 3040 20821 3043
rect 19996 3012 20821 3040
rect 19889 3003 19947 3009
rect 20809 3009 20821 3012
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 16807 2944 17172 2972
rect 16807 2941 16819 2944
rect 16761 2935 16819 2941
rect 18322 2932 18328 2984
rect 18380 2972 18386 2984
rect 18380 2944 19012 2972
rect 18380 2932 18386 2944
rect 16022 2904 16028 2916
rect 15983 2876 16028 2904
rect 16022 2864 16028 2876
rect 16080 2864 16086 2916
rect 18877 2907 18935 2913
rect 18877 2904 18889 2907
rect 16132 2876 17080 2904
rect 13262 2836 13268 2848
rect 12544 2808 13032 2836
rect 13223 2808 13268 2836
rect 13262 2796 13268 2808
rect 13320 2796 13326 2848
rect 14918 2796 14924 2848
rect 14976 2836 14982 2848
rect 16132 2836 16160 2876
rect 14976 2808 16160 2836
rect 17052 2836 17080 2876
rect 17972 2876 18889 2904
rect 17972 2836 18000 2876
rect 18877 2873 18889 2876
rect 18923 2873 18935 2907
rect 18877 2867 18935 2873
rect 17052 2808 18000 2836
rect 18417 2839 18475 2845
rect 14976 2796 14982 2808
rect 18417 2805 18429 2839
rect 18463 2836 18475 2839
rect 18690 2836 18696 2848
rect 18463 2808 18696 2836
rect 18463 2805 18475 2808
rect 18417 2799 18475 2805
rect 18690 2796 18696 2808
rect 18748 2796 18754 2848
rect 18984 2836 19012 2944
rect 19334 2932 19340 2984
rect 19392 2972 19398 2984
rect 19613 2975 19671 2981
rect 19613 2972 19625 2975
rect 19392 2944 19625 2972
rect 19392 2932 19398 2944
rect 19613 2941 19625 2944
rect 19659 2941 19671 2975
rect 19613 2935 19671 2941
rect 19797 2975 19855 2981
rect 19797 2941 19809 2975
rect 19843 2972 19855 2975
rect 20070 2972 20076 2984
rect 19843 2944 20076 2972
rect 19843 2941 19855 2944
rect 19797 2935 19855 2941
rect 20070 2932 20076 2944
rect 20128 2932 20134 2984
rect 20533 2975 20591 2981
rect 20533 2941 20545 2975
rect 20579 2972 20591 2975
rect 20622 2972 20628 2984
rect 20579 2944 20628 2972
rect 20579 2941 20591 2944
rect 20533 2935 20591 2941
rect 19058 2864 19064 2916
rect 19116 2904 19122 2916
rect 20548 2904 20576 2935
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 22646 2904 22652 2916
rect 19116 2876 20576 2904
rect 20640 2876 22652 2904
rect 19116 2864 19122 2876
rect 20640 2836 20668 2876
rect 22646 2864 22652 2876
rect 22704 2864 22710 2916
rect 18984 2808 20668 2836
rect 20714 2796 20720 2848
rect 20772 2836 20778 2848
rect 22094 2836 22100 2848
rect 20772 2808 22100 2836
rect 20772 2796 20778 2808
rect 22094 2796 22100 2808
rect 22152 2796 22158 2848
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 3326 2632 3332 2644
rect 3287 2604 3332 2632
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 3970 2592 3976 2644
rect 4028 2632 4034 2644
rect 4801 2635 4859 2641
rect 4801 2632 4813 2635
rect 4028 2604 4813 2632
rect 4028 2592 4034 2604
rect 4801 2601 4813 2604
rect 4847 2632 4859 2635
rect 5258 2632 5264 2644
rect 4847 2604 5264 2632
rect 4847 2601 4859 2604
rect 4801 2595 4859 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 5902 2632 5908 2644
rect 5863 2604 5908 2632
rect 5902 2592 5908 2604
rect 5960 2592 5966 2644
rect 7282 2632 7288 2644
rect 6012 2604 6776 2632
rect 7243 2604 7288 2632
rect 2777 2567 2835 2573
rect 2777 2533 2789 2567
rect 2823 2564 2835 2567
rect 3050 2564 3056 2576
rect 2823 2536 3056 2564
rect 2823 2533 2835 2536
rect 2777 2527 2835 2533
rect 3050 2524 3056 2536
rect 3108 2524 3114 2576
rect 3142 2524 3148 2576
rect 3200 2564 3206 2576
rect 3878 2564 3884 2576
rect 3200 2536 3884 2564
rect 3200 2524 3206 2536
rect 3878 2524 3884 2536
rect 3936 2524 3942 2576
rect 4525 2567 4583 2573
rect 4525 2533 4537 2567
rect 4571 2564 4583 2567
rect 5534 2564 5540 2576
rect 4571 2536 5540 2564
rect 4571 2533 4583 2536
rect 4525 2527 4583 2533
rect 5534 2524 5540 2536
rect 5592 2524 5598 2576
rect 290 2456 296 2508
rect 348 2496 354 2508
rect 1302 2496 1308 2508
rect 348 2468 1308 2496
rect 348 2456 354 2468
rect 1302 2456 1308 2468
rect 1360 2496 1366 2508
rect 1397 2499 1455 2505
rect 1397 2496 1409 2499
rect 1360 2468 1409 2496
rect 1360 2456 1366 2468
rect 1397 2465 1409 2468
rect 1443 2465 1455 2499
rect 1397 2459 1455 2465
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 2406 2496 2412 2508
rect 1719 2468 2412 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 2406 2456 2412 2468
rect 2464 2456 2470 2508
rect 4614 2456 4620 2508
rect 4672 2496 4678 2508
rect 6012 2496 6040 2604
rect 6641 2567 6699 2573
rect 6641 2533 6653 2567
rect 6687 2533 6699 2567
rect 6748 2564 6776 2604
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 8294 2632 8300 2644
rect 7392 2604 8300 2632
rect 7392 2564 7420 2604
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 9398 2632 9404 2644
rect 9359 2604 9404 2632
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 11790 2592 11796 2644
rect 11848 2632 11854 2644
rect 15194 2632 15200 2644
rect 11848 2604 15200 2632
rect 11848 2592 11854 2604
rect 15194 2592 15200 2604
rect 15252 2592 15258 2644
rect 15562 2632 15568 2644
rect 15523 2604 15568 2632
rect 15562 2592 15568 2604
rect 15620 2592 15626 2644
rect 17405 2635 17463 2641
rect 17405 2601 17417 2635
rect 17451 2632 17463 2635
rect 18046 2632 18052 2644
rect 17451 2604 18052 2632
rect 17451 2601 17463 2604
rect 17405 2595 17463 2601
rect 18046 2592 18052 2604
rect 18104 2592 18110 2644
rect 6748 2536 7420 2564
rect 8481 2567 8539 2573
rect 6641 2527 6699 2533
rect 8481 2533 8493 2567
rect 8527 2564 8539 2567
rect 11698 2564 11704 2576
rect 8527 2536 11560 2564
rect 11659 2536 11704 2564
rect 8527 2533 8539 2536
rect 8481 2527 8539 2533
rect 4672 2468 6040 2496
rect 6656 2496 6684 2527
rect 6730 2496 6736 2508
rect 6656 2468 6736 2496
rect 4672 2456 4678 2468
rect 6730 2456 6736 2468
rect 6788 2456 6794 2508
rect 6914 2456 6920 2508
rect 6972 2496 6978 2508
rect 10137 2499 10195 2505
rect 6972 2468 8340 2496
rect 6972 2456 6978 2468
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2593 2431 2651 2437
rect 2593 2428 2605 2431
rect 2004 2400 2605 2428
rect 2004 2388 2010 2400
rect 2593 2397 2605 2400
rect 2639 2397 2651 2431
rect 3234 2428 3240 2440
rect 3195 2400 3240 2428
rect 2593 2391 2651 2397
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 3789 2431 3847 2437
rect 3789 2397 3801 2431
rect 3835 2428 3847 2431
rect 4430 2428 4436 2440
rect 3835 2400 4436 2428
rect 3835 2397 3847 2400
rect 3789 2391 3847 2397
rect 4430 2388 4436 2400
rect 4488 2388 4494 2440
rect 5626 2388 5632 2440
rect 5684 2428 5690 2440
rect 8312 2437 8340 2468
rect 10137 2465 10149 2499
rect 10183 2496 10195 2499
rect 10410 2496 10416 2508
rect 10183 2468 10416 2496
rect 10183 2465 10195 2468
rect 10137 2459 10195 2465
rect 10410 2456 10416 2468
rect 10468 2456 10474 2508
rect 11532 2496 11560 2536
rect 11698 2524 11704 2536
rect 11756 2524 11762 2576
rect 12526 2564 12532 2576
rect 12406 2536 12532 2564
rect 12406 2496 12434 2536
rect 12526 2524 12532 2536
rect 12584 2524 12590 2576
rect 16022 2524 16028 2576
rect 16080 2564 16086 2576
rect 19659 2567 19717 2573
rect 19659 2564 19671 2567
rect 16080 2536 16804 2564
rect 16080 2524 16086 2536
rect 11532 2468 12434 2496
rect 13081 2499 13139 2505
rect 13081 2465 13093 2499
rect 13127 2496 13139 2499
rect 14734 2496 14740 2508
rect 13127 2468 14740 2496
rect 13127 2465 13139 2468
rect 13081 2459 13139 2465
rect 14734 2456 14740 2468
rect 14792 2456 14798 2508
rect 16776 2505 16804 2536
rect 16960 2536 19671 2564
rect 16960 2505 16988 2536
rect 19659 2533 19671 2536
rect 19705 2564 19717 2567
rect 20530 2564 20536 2576
rect 19705 2536 20536 2564
rect 19705 2533 19717 2536
rect 19659 2527 19717 2533
rect 20530 2524 20536 2536
rect 20588 2524 20594 2576
rect 16209 2499 16267 2505
rect 16209 2465 16221 2499
rect 16255 2465 16267 2499
rect 16209 2459 16267 2465
rect 16761 2499 16819 2505
rect 16761 2465 16773 2499
rect 16807 2465 16819 2499
rect 16761 2459 16819 2465
rect 16945 2499 17003 2505
rect 16945 2465 16957 2499
rect 16991 2465 17003 2499
rect 16945 2459 17003 2465
rect 17865 2499 17923 2505
rect 17865 2465 17877 2499
rect 17911 2496 17923 2499
rect 18230 2496 18236 2508
rect 17911 2468 18236 2496
rect 17911 2465 17923 2468
rect 17865 2459 17923 2465
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 5684 2400 7757 2428
rect 5684 2388 5690 2400
rect 7745 2397 7757 2400
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2397 8355 2431
rect 9674 2428 9680 2440
rect 8297 2391 8355 2397
rect 8404 2400 9680 2428
rect 4154 2320 4160 2372
rect 4212 2360 4218 2372
rect 4341 2363 4399 2369
rect 4341 2360 4353 2363
rect 4212 2332 4353 2360
rect 4212 2320 4218 2332
rect 4341 2329 4353 2332
rect 4387 2329 4399 2363
rect 5350 2360 5356 2372
rect 5311 2332 5356 2360
rect 4341 2323 4399 2329
rect 5350 2320 5356 2332
rect 5408 2320 5414 2372
rect 5810 2360 5816 2372
rect 5723 2332 5816 2360
rect 5810 2320 5816 2332
rect 5868 2360 5874 2372
rect 6086 2360 6092 2372
rect 5868 2332 6092 2360
rect 5868 2320 5874 2332
rect 6086 2320 6092 2332
rect 6144 2320 6150 2372
rect 6730 2320 6736 2372
rect 6788 2360 6794 2372
rect 6825 2363 6883 2369
rect 6825 2360 6837 2363
rect 6788 2332 6837 2360
rect 6788 2320 6794 2332
rect 6825 2329 6837 2332
rect 6871 2329 6883 2363
rect 6825 2323 6883 2329
rect 7098 2320 7104 2372
rect 7156 2360 7162 2372
rect 7377 2363 7435 2369
rect 7377 2360 7389 2363
rect 7156 2332 7389 2360
rect 7156 2320 7162 2332
rect 7377 2329 7389 2332
rect 7423 2360 7435 2363
rect 8404 2360 8432 2400
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 9766 2388 9772 2440
rect 9824 2428 9830 2440
rect 9861 2431 9919 2437
rect 9861 2428 9873 2431
rect 9824 2400 9873 2428
rect 9824 2388 9830 2400
rect 9861 2397 9873 2400
rect 9907 2397 9919 2431
rect 11146 2428 11152 2440
rect 11107 2400 11152 2428
rect 9861 2391 9919 2397
rect 11146 2388 11152 2400
rect 11204 2388 11210 2440
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 12710 2428 12716 2440
rect 12671 2400 12716 2428
rect 11517 2391 11575 2397
rect 7423 2332 8432 2360
rect 7423 2329 7435 2332
rect 7377 2323 7435 2329
rect 8478 2320 8484 2372
rect 8536 2360 8542 2372
rect 8536 2332 9076 2360
rect 8536 2320 8542 2332
rect 3970 2292 3976 2304
rect 3931 2264 3976 2292
rect 3970 2252 3976 2264
rect 4028 2252 4034 2304
rect 5261 2295 5319 2301
rect 5261 2261 5273 2295
rect 5307 2292 5319 2295
rect 7190 2292 7196 2304
rect 5307 2264 7196 2292
rect 5307 2261 5319 2264
rect 5261 2255 5319 2261
rect 7190 2252 7196 2264
rect 7248 2252 7254 2304
rect 7929 2295 7987 2301
rect 7929 2261 7941 2295
rect 7975 2292 7987 2295
rect 8202 2292 8208 2304
rect 7975 2264 8208 2292
rect 7975 2261 7987 2264
rect 7929 2255 7987 2261
rect 8202 2252 8208 2264
rect 8260 2252 8266 2304
rect 8938 2292 8944 2304
rect 8899 2264 8944 2292
rect 8938 2252 8944 2264
rect 8996 2252 9002 2304
rect 9048 2292 9076 2332
rect 9398 2320 9404 2372
rect 9456 2360 9462 2372
rect 9493 2363 9551 2369
rect 9493 2360 9505 2363
rect 9456 2332 9505 2360
rect 9456 2320 9462 2332
rect 9493 2329 9505 2332
rect 9539 2329 9551 2363
rect 11532 2360 11560 2391
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 13262 2388 13268 2440
rect 13320 2388 13326 2440
rect 13722 2388 13728 2440
rect 13780 2428 13786 2440
rect 14829 2431 14887 2437
rect 14829 2428 14841 2431
rect 13780 2400 14841 2428
rect 13780 2388 13786 2400
rect 14829 2397 14841 2400
rect 14875 2397 14887 2431
rect 16224 2428 16252 2459
rect 18230 2456 18236 2468
rect 18288 2456 18294 2508
rect 18690 2496 18696 2508
rect 18651 2468 18696 2496
rect 18690 2456 18696 2468
rect 18748 2456 18754 2508
rect 19794 2496 19800 2508
rect 18800 2468 19800 2496
rect 18800 2428 18828 2468
rect 19794 2456 19800 2468
rect 19852 2456 19858 2508
rect 16224 2400 18828 2428
rect 14829 2391 14887 2397
rect 19242 2388 19248 2440
rect 19300 2428 19306 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 19300 2400 19441 2428
rect 19300 2388 19306 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 21082 2428 21088 2440
rect 21043 2400 21088 2428
rect 19429 2391 19487 2397
rect 21082 2388 21088 2400
rect 21140 2388 21146 2440
rect 21358 2428 21364 2440
rect 21319 2400 21364 2428
rect 21358 2388 21364 2400
rect 21416 2388 21422 2440
rect 9493 2323 9551 2329
rect 10428 2332 11560 2360
rect 13280 2360 13308 2388
rect 14921 2363 14979 2369
rect 14921 2360 14933 2363
rect 13280 2332 14933 2360
rect 10428 2292 10456 2332
rect 14921 2329 14933 2332
rect 14967 2329 14979 2363
rect 14921 2323 14979 2329
rect 15010 2320 15016 2372
rect 15068 2360 15074 2372
rect 15933 2363 15991 2369
rect 15933 2360 15945 2363
rect 15068 2332 15945 2360
rect 15068 2320 15074 2332
rect 15933 2329 15945 2332
rect 15979 2329 15991 2363
rect 15933 2323 15991 2329
rect 16025 2363 16083 2369
rect 16025 2329 16037 2363
rect 16071 2360 16083 2363
rect 16071 2332 18184 2360
rect 16071 2329 16083 2332
rect 16025 2323 16083 2329
rect 10962 2292 10968 2304
rect 9048 2264 10456 2292
rect 10923 2264 10968 2292
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 12066 2292 12072 2304
rect 12027 2264 12072 2292
rect 12066 2252 12072 2264
rect 12124 2252 12130 2304
rect 13170 2252 13176 2304
rect 13228 2292 13234 2304
rect 13265 2295 13323 2301
rect 13265 2292 13277 2295
rect 13228 2264 13277 2292
rect 13228 2252 13234 2264
rect 13265 2261 13277 2264
rect 13311 2261 13323 2295
rect 13265 2255 13323 2261
rect 13354 2252 13360 2304
rect 13412 2292 13418 2304
rect 13722 2292 13728 2304
rect 13412 2264 13457 2292
rect 13683 2264 13728 2292
rect 13412 2252 13418 2264
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 14274 2292 14280 2304
rect 14235 2264 14280 2292
rect 14274 2252 14280 2264
rect 14332 2252 14338 2304
rect 15286 2292 15292 2304
rect 15247 2264 15292 2292
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 17034 2252 17040 2304
rect 17092 2292 17098 2304
rect 18156 2301 18184 2332
rect 18322 2320 18328 2372
rect 18380 2360 18386 2372
rect 18601 2363 18659 2369
rect 18601 2360 18613 2363
rect 18380 2332 18613 2360
rect 18380 2320 18386 2332
rect 18601 2329 18613 2332
rect 18647 2360 18659 2363
rect 22278 2360 22284 2372
rect 18647 2332 22284 2360
rect 18647 2329 18659 2332
rect 18601 2323 18659 2329
rect 22278 2320 22284 2332
rect 22336 2320 22342 2372
rect 18141 2295 18199 2301
rect 17092 2264 17137 2292
rect 17092 2252 17098 2264
rect 18141 2261 18153 2295
rect 18187 2261 18199 2295
rect 18506 2292 18512 2304
rect 18467 2264 18512 2292
rect 18141 2255 18199 2261
rect 18506 2252 18512 2264
rect 18564 2252 18570 2304
rect 1104 2202 21896 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21896 2202
rect 1104 2128 21896 2150
rect 2866 2048 2872 2100
rect 2924 2088 2930 2100
rect 7098 2088 7104 2100
rect 2924 2060 7104 2088
rect 2924 2048 2930 2060
rect 7098 2048 7104 2060
rect 7156 2048 7162 2100
rect 8570 2048 8576 2100
rect 8628 2088 8634 2100
rect 13354 2088 13360 2100
rect 8628 2060 13360 2088
rect 8628 2048 8634 2060
rect 13354 2048 13360 2060
rect 13412 2048 13418 2100
rect 14274 2048 14280 2100
rect 14332 2088 14338 2100
rect 17954 2088 17960 2100
rect 14332 2060 17960 2088
rect 14332 2048 14338 2060
rect 17954 2048 17960 2060
rect 18012 2048 18018 2100
rect 4982 1980 4988 2032
rect 5040 2020 5046 2032
rect 12158 2020 12164 2032
rect 5040 1992 12164 2020
rect 5040 1980 5046 1992
rect 12158 1980 12164 1992
rect 12216 1980 12222 2032
rect 12250 1980 12256 2032
rect 12308 2020 12314 2032
rect 12986 2020 12992 2032
rect 12308 1992 12992 2020
rect 12308 1980 12314 1992
rect 12986 1980 12992 1992
rect 13044 1980 13050 2032
rect 13722 1980 13728 2032
rect 13780 2020 13786 2032
rect 18414 2020 18420 2032
rect 13780 1992 18420 2020
rect 13780 1980 13786 1992
rect 18414 1980 18420 1992
rect 18472 1980 18478 2032
rect 5166 1912 5172 1964
rect 5224 1952 5230 1964
rect 10962 1952 10968 1964
rect 5224 1924 10968 1952
rect 5224 1912 5230 1924
rect 10962 1912 10968 1924
rect 11020 1912 11026 1964
rect 12710 1912 12716 1964
rect 12768 1952 12774 1964
rect 18598 1952 18604 1964
rect 12768 1924 18604 1952
rect 12768 1912 12774 1924
rect 18598 1912 18604 1924
rect 18656 1912 18662 1964
rect 2314 1844 2320 1896
rect 2372 1884 2378 1896
rect 6730 1884 6736 1896
rect 2372 1856 6736 1884
rect 2372 1844 2378 1856
rect 6730 1844 6736 1856
rect 6788 1884 6794 1896
rect 8110 1884 8116 1896
rect 6788 1856 8116 1884
rect 6788 1844 6794 1856
rect 8110 1844 8116 1856
rect 8168 1844 8174 1896
rect 8386 1844 8392 1896
rect 8444 1884 8450 1896
rect 13078 1884 13084 1896
rect 8444 1856 13084 1884
rect 8444 1844 8450 1856
rect 13078 1844 13084 1856
rect 13136 1844 13142 1896
rect 15286 1844 15292 1896
rect 15344 1884 15350 1896
rect 19518 1884 19524 1896
rect 15344 1856 19524 1884
rect 15344 1844 15350 1856
rect 19518 1844 19524 1856
rect 19576 1844 19582 1896
rect 7006 1776 7012 1828
rect 7064 1816 7070 1828
rect 16114 1816 16120 1828
rect 7064 1788 16120 1816
rect 7064 1776 7070 1788
rect 16114 1776 16120 1788
rect 16172 1776 16178 1828
rect 9674 1708 9680 1760
rect 9732 1748 9738 1760
rect 10870 1748 10876 1760
rect 9732 1720 10876 1748
rect 9732 1708 9738 1720
rect 10870 1708 10876 1720
rect 10928 1708 10934 1760
rect 11146 1708 11152 1760
rect 11204 1748 11210 1760
rect 11204 1720 14688 1748
rect 11204 1708 11210 1720
rect 8938 1640 8944 1692
rect 8996 1680 9002 1692
rect 12250 1680 12256 1692
rect 8996 1652 12256 1680
rect 8996 1640 9002 1652
rect 12250 1640 12256 1652
rect 12308 1640 12314 1692
rect 14660 1680 14688 1720
rect 14734 1708 14740 1760
rect 14792 1748 14798 1760
rect 20254 1748 20260 1760
rect 14792 1720 20260 1748
rect 14792 1708 14798 1720
rect 20254 1708 20260 1720
rect 20312 1708 20318 1760
rect 17218 1680 17224 1692
rect 14660 1652 17224 1680
rect 17218 1640 17224 1652
rect 17276 1640 17282 1692
rect 3878 1572 3884 1624
rect 3936 1612 3942 1624
rect 9398 1612 9404 1624
rect 3936 1584 9404 1612
rect 3936 1572 3942 1584
rect 9398 1572 9404 1584
rect 9456 1572 9462 1624
rect 9490 1572 9496 1624
rect 9548 1612 9554 1624
rect 15102 1612 15108 1624
rect 9548 1584 15108 1612
rect 9548 1572 9554 1584
rect 15102 1572 15108 1584
rect 15160 1572 15166 1624
rect 9950 1504 9956 1556
rect 10008 1544 10014 1556
rect 11422 1544 11428 1556
rect 10008 1516 11428 1544
rect 10008 1504 10014 1516
rect 11422 1504 11428 1516
rect 11480 1504 11486 1556
rect 12434 1504 12440 1556
rect 12492 1544 12498 1556
rect 14826 1544 14832 1556
rect 12492 1516 14832 1544
rect 12492 1504 12498 1516
rect 14826 1504 14832 1516
rect 14884 1504 14890 1556
rect 8202 1436 8208 1488
rect 8260 1476 8266 1488
rect 12066 1476 12072 1488
rect 8260 1448 12072 1476
rect 8260 1436 8266 1448
rect 12066 1436 12072 1448
rect 12124 1436 12130 1488
rect 13170 1436 13176 1488
rect 13228 1476 13234 1488
rect 14918 1476 14924 1488
rect 13228 1448 14924 1476
rect 13228 1436 13234 1448
rect 14918 1436 14924 1448
rect 14976 1436 14982 1488
rect 19334 1368 19340 1420
rect 19392 1408 19398 1420
rect 20162 1408 20168 1420
rect 19392 1380 20168 1408
rect 19392 1368 19398 1380
rect 20162 1368 20168 1380
rect 20220 1368 20226 1420
rect 9122 1300 9128 1352
rect 9180 1340 9186 1352
rect 16206 1340 16212 1352
rect 9180 1312 16212 1340
rect 9180 1300 9186 1312
rect 16206 1300 16212 1312
rect 16264 1300 16270 1352
rect 17126 1300 17132 1352
rect 17184 1340 17190 1352
rect 19242 1340 19248 1352
rect 17184 1312 19248 1340
rect 17184 1300 17190 1312
rect 19242 1300 19248 1312
rect 19300 1300 19306 1352
rect 7374 1232 7380 1284
rect 7432 1272 7438 1284
rect 15746 1272 15752 1284
rect 7432 1244 15752 1272
rect 7432 1232 7438 1244
rect 15746 1232 15752 1244
rect 15804 1232 15810 1284
rect 11882 1164 11888 1216
rect 11940 1204 11946 1216
rect 18690 1204 18696 1216
rect 11940 1176 18696 1204
rect 11940 1164 11946 1176
rect 18690 1164 18696 1176
rect 18748 1164 18754 1216
rect 6822 1096 6828 1148
rect 6880 1136 6886 1148
rect 18874 1136 18880 1148
rect 6880 1108 18880 1136
rect 6880 1096 6886 1108
rect 18874 1096 18880 1108
rect 18932 1096 18938 1148
rect 6638 1028 6644 1080
rect 6696 1068 6702 1080
rect 17494 1068 17500 1080
rect 6696 1040 17500 1068
rect 6696 1028 6702 1040
rect 17494 1028 17500 1040
rect 17552 1028 17558 1080
rect 9306 960 9312 1012
rect 9364 1000 9370 1012
rect 17862 1000 17868 1012
rect 9364 972 17868 1000
rect 9364 960 9370 972
rect 17862 960 17868 972
rect 17920 960 17926 1012
rect 5902 892 5908 944
rect 5960 932 5966 944
rect 8662 932 8668 944
rect 5960 904 8668 932
rect 5960 892 5966 904
rect 8662 892 8668 904
rect 8720 892 8726 944
rect 9398 892 9404 944
rect 9456 932 9462 944
rect 17954 932 17960 944
rect 9456 904 17960 932
rect 9456 892 9462 904
rect 17954 892 17960 904
rect 18012 892 18018 944
rect 4522 824 4528 876
rect 4580 864 4586 876
rect 19610 864 19616 876
rect 4580 836 19616 864
rect 4580 824 4586 836
rect 19610 824 19616 836
rect 19668 824 19674 876
rect 2958 756 2964 808
rect 3016 796 3022 808
rect 16942 796 16948 808
rect 3016 768 16948 796
rect 3016 756 3022 768
rect 16942 756 16948 768
rect 17000 756 17006 808
rect 5074 688 5080 740
rect 5132 728 5138 740
rect 18966 728 18972 740
rect 5132 700 18972 728
rect 5132 688 5138 700
rect 18966 688 18972 700
rect 19024 688 19030 740
rect 7926 620 7932 672
rect 7984 660 7990 672
rect 17586 660 17592 672
rect 7984 632 17592 660
rect 7984 620 7990 632
rect 17586 620 17592 632
rect 17644 620 17650 672
rect 4062 552 4068 604
rect 4120 592 4126 604
rect 14458 592 14464 604
rect 4120 564 14464 592
rect 4120 552 4126 564
rect 14458 552 14464 564
rect 14516 592 14522 604
rect 21082 592 21088 604
rect 14516 564 21088 592
rect 14516 552 14522 564
rect 21082 552 21088 564
rect 21140 552 21146 604
<< via1 >>
rect 6000 21292 6052 21344
rect 14648 21292 14700 21344
rect 8208 21224 8260 21276
rect 12348 21224 12400 21276
rect 4896 21156 4948 21208
rect 18420 21156 18472 21208
rect 4804 21088 4856 21140
rect 20352 21088 20404 21140
rect 9312 21020 9364 21072
rect 17592 21020 17644 21072
rect 7472 20952 7524 21004
rect 17132 20952 17184 21004
rect 7104 20884 7156 20936
rect 17224 20884 17276 20936
rect 7656 20816 7708 20868
rect 11428 20816 11480 20868
rect 7380 20748 7432 20800
rect 16212 20748 16264 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 7196 20544 7248 20596
rect 1952 20476 2004 20528
rect 3056 20476 3108 20528
rect 3608 20476 3660 20528
rect 4160 20476 4212 20528
rect 2504 20408 2556 20460
rect 3424 20408 3476 20460
rect 7012 20476 7064 20528
rect 9404 20476 9456 20528
rect 9956 20519 10008 20528
rect 9956 20485 9965 20519
rect 9965 20485 9999 20519
rect 9999 20485 10008 20519
rect 9956 20476 10008 20485
rect 11060 20476 11112 20528
rect 12624 20544 12676 20596
rect 14464 20544 14516 20596
rect 5172 20340 5224 20392
rect 5632 20408 5684 20460
rect 5816 20451 5868 20460
rect 5816 20417 5825 20451
rect 5825 20417 5859 20451
rect 5859 20417 5868 20451
rect 5816 20408 5868 20417
rect 6644 20451 6696 20460
rect 6644 20417 6653 20451
rect 6653 20417 6687 20451
rect 6687 20417 6696 20451
rect 6644 20408 6696 20417
rect 6828 20451 6880 20460
rect 6828 20417 6837 20451
rect 6837 20417 6871 20451
rect 6871 20417 6880 20451
rect 6828 20408 6880 20417
rect 5356 20340 5408 20392
rect 7288 20408 7340 20460
rect 7564 20408 7616 20460
rect 7932 20408 7984 20460
rect 8116 20408 8168 20460
rect 8668 20408 8720 20460
rect 9680 20408 9732 20460
rect 10324 20408 10376 20460
rect 11152 20451 11204 20460
rect 11152 20417 11161 20451
rect 11161 20417 11195 20451
rect 11195 20417 11204 20451
rect 11152 20408 11204 20417
rect 12256 20408 12308 20460
rect 13360 20408 13412 20460
rect 14372 20476 14424 20528
rect 7840 20340 7892 20392
rect 8024 20340 8076 20392
rect 2320 20315 2372 20324
rect 2320 20281 2329 20315
rect 2329 20281 2363 20315
rect 2363 20281 2372 20315
rect 2320 20272 2372 20281
rect 4528 20315 4580 20324
rect 4528 20281 4537 20315
rect 4537 20281 4571 20315
rect 4571 20281 4580 20315
rect 4528 20272 4580 20281
rect 6828 20272 6880 20324
rect 8300 20272 8352 20324
rect 11980 20340 12032 20392
rect 13176 20272 13228 20324
rect 15384 20544 15436 20596
rect 16396 20544 16448 20596
rect 15292 20476 15344 20528
rect 15752 20451 15804 20460
rect 15752 20417 15761 20451
rect 15761 20417 15795 20451
rect 15795 20417 15804 20451
rect 15752 20408 15804 20417
rect 16948 20408 17000 20460
rect 17224 20451 17276 20460
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 17684 20476 17736 20528
rect 21548 20544 21600 20596
rect 18052 20408 18104 20460
rect 18880 20408 18932 20460
rect 19800 20451 19852 20460
rect 19800 20417 19809 20451
rect 19809 20417 19843 20451
rect 19843 20417 19852 20451
rect 19800 20408 19852 20417
rect 20352 20451 20404 20460
rect 20352 20417 20361 20451
rect 20361 20417 20395 20451
rect 20395 20417 20404 20451
rect 20352 20408 20404 20417
rect 21088 20451 21140 20460
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 15292 20340 15344 20392
rect 2964 20204 3016 20256
rect 3332 20247 3384 20256
rect 3332 20213 3341 20247
rect 3341 20213 3375 20247
rect 3375 20213 3384 20247
rect 3332 20204 3384 20213
rect 5448 20204 5500 20256
rect 6276 20204 6328 20256
rect 7748 20204 7800 20256
rect 9496 20204 9548 20256
rect 10048 20247 10100 20256
rect 10048 20213 10057 20247
rect 10057 20213 10091 20247
rect 10091 20213 10100 20247
rect 10048 20204 10100 20213
rect 10876 20204 10928 20256
rect 13268 20247 13320 20256
rect 13268 20213 13277 20247
rect 13277 20213 13311 20247
rect 13311 20213 13320 20247
rect 13268 20204 13320 20213
rect 13452 20204 13504 20256
rect 13820 20204 13872 20256
rect 17040 20272 17092 20324
rect 22100 20272 22152 20324
rect 18972 20204 19024 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 4344 20043 4396 20052
rect 4344 20009 4353 20043
rect 4353 20009 4387 20043
rect 4387 20009 4396 20043
rect 4344 20000 4396 20009
rect 4804 20043 4856 20052
rect 4804 20009 4813 20043
rect 4813 20009 4847 20043
rect 4847 20009 4856 20043
rect 4804 20000 4856 20009
rect 1400 19932 1452 19984
rect 1676 19932 1728 19984
rect 3332 19932 3384 19984
rect 5540 19932 5592 19984
rect 2044 19864 2096 19916
rect 6920 20000 6972 20052
rect 5724 19975 5776 19984
rect 5724 19941 5733 19975
rect 5733 19941 5767 19975
rect 5767 19941 5776 19975
rect 5724 19932 5776 19941
rect 6736 19932 6788 19984
rect 296 19796 348 19848
rect 1400 19796 1452 19848
rect 848 19728 900 19780
rect 3148 19796 3200 19848
rect 3976 19796 4028 19848
rect 4436 19796 4488 19848
rect 4804 19796 4856 19848
rect 2780 19728 2832 19780
rect 1768 19703 1820 19712
rect 1768 19669 1777 19703
rect 1777 19669 1811 19703
rect 1811 19669 1820 19703
rect 1768 19660 1820 19669
rect 2228 19660 2280 19712
rect 3240 19660 3292 19712
rect 3792 19660 3844 19712
rect 4252 19728 4304 19780
rect 5724 19796 5776 19848
rect 6276 19864 6328 19916
rect 6000 19839 6052 19848
rect 6000 19805 6009 19839
rect 6009 19805 6043 19839
rect 6043 19805 6052 19839
rect 6000 19796 6052 19805
rect 6092 19796 6144 19848
rect 6736 19796 6788 19848
rect 7748 19864 7800 19916
rect 10140 19907 10192 19916
rect 10140 19873 10149 19907
rect 10149 19873 10183 19907
rect 10183 19873 10192 19907
rect 10140 19864 10192 19873
rect 7656 19796 7708 19848
rect 8208 19796 8260 19848
rect 8392 19796 8444 19848
rect 7656 19660 7708 19712
rect 8024 19703 8076 19712
rect 8024 19669 8033 19703
rect 8033 19669 8067 19703
rect 8067 19669 8076 19703
rect 8024 19660 8076 19669
rect 8116 19660 8168 19712
rect 10968 19839 11020 19848
rect 10968 19805 10977 19839
rect 10977 19805 11011 19839
rect 11011 19805 11020 19839
rect 10968 19796 11020 19805
rect 11244 19839 11296 19848
rect 11244 19805 11278 19839
rect 11278 19805 11296 19839
rect 11244 19796 11296 19805
rect 12164 20000 12216 20052
rect 15936 20000 15988 20052
rect 17868 20000 17920 20052
rect 18328 20043 18380 20052
rect 18328 20009 18337 20043
rect 18337 20009 18371 20043
rect 18371 20009 18380 20043
rect 18328 20000 18380 20009
rect 18880 20043 18932 20052
rect 18880 20009 18889 20043
rect 18889 20009 18923 20043
rect 18923 20009 18932 20043
rect 18880 20000 18932 20009
rect 12072 19932 12124 19984
rect 12992 19907 13044 19916
rect 12992 19873 13001 19907
rect 13001 19873 13035 19907
rect 13035 19873 13044 19907
rect 12992 19864 13044 19873
rect 18236 19932 18288 19984
rect 14832 19907 14884 19916
rect 14832 19873 14841 19907
rect 14841 19873 14875 19907
rect 14875 19873 14884 19907
rect 14832 19864 14884 19873
rect 17500 19864 17552 19916
rect 20536 19864 20588 19916
rect 15016 19839 15068 19848
rect 15016 19805 15025 19839
rect 15025 19805 15059 19839
rect 15059 19805 15068 19839
rect 15016 19796 15068 19805
rect 15108 19796 15160 19848
rect 16120 19839 16172 19848
rect 16120 19805 16129 19839
rect 16129 19805 16163 19839
rect 16163 19805 16172 19839
rect 16120 19796 16172 19805
rect 16212 19796 16264 19848
rect 17592 19839 17644 19848
rect 17592 19805 17601 19839
rect 17601 19805 17635 19839
rect 17635 19805 17644 19839
rect 17592 19796 17644 19805
rect 18144 19839 18196 19848
rect 18144 19805 18153 19839
rect 18153 19805 18187 19839
rect 18187 19805 18196 19839
rect 18144 19796 18196 19805
rect 18604 19796 18656 19848
rect 20812 19839 20864 19848
rect 8484 19703 8536 19712
rect 8484 19669 8493 19703
rect 8493 19669 8527 19703
rect 8527 19669 8536 19703
rect 9128 19703 9180 19712
rect 8484 19660 8536 19669
rect 9128 19669 9137 19703
rect 9137 19669 9171 19703
rect 9171 19669 9180 19703
rect 9128 19660 9180 19669
rect 9588 19703 9640 19712
rect 9588 19669 9597 19703
rect 9597 19669 9631 19703
rect 9631 19669 9640 19703
rect 9588 19660 9640 19669
rect 10232 19703 10284 19712
rect 10232 19669 10241 19703
rect 10241 19669 10275 19703
rect 10275 19669 10284 19703
rect 10232 19660 10284 19669
rect 10692 19703 10744 19712
rect 10692 19669 10701 19703
rect 10701 19669 10735 19703
rect 10735 19669 10744 19703
rect 10692 19660 10744 19669
rect 11888 19728 11940 19780
rect 16948 19728 17000 19780
rect 20812 19805 20821 19839
rect 20821 19805 20855 19839
rect 20855 19805 20864 19839
rect 20812 19796 20864 19805
rect 20168 19771 20220 19780
rect 20168 19737 20177 19771
rect 20177 19737 20211 19771
rect 20211 19737 20220 19771
rect 20168 19728 20220 19737
rect 21272 19771 21324 19780
rect 21272 19737 21281 19771
rect 21281 19737 21315 19771
rect 21315 19737 21324 19771
rect 21272 19728 21324 19737
rect 12072 19660 12124 19712
rect 12256 19660 12308 19712
rect 13084 19703 13136 19712
rect 13084 19669 13093 19703
rect 13093 19669 13127 19703
rect 13127 19669 13136 19703
rect 13084 19660 13136 19669
rect 13728 19660 13780 19712
rect 13820 19660 13872 19712
rect 15292 19660 15344 19712
rect 15752 19660 15804 19712
rect 18604 19660 18656 19712
rect 18788 19660 18840 19712
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 3884 19456 3936 19508
rect 4528 19456 4580 19508
rect 4712 19456 4764 19508
rect 7104 19499 7156 19508
rect 7104 19465 7113 19499
rect 7113 19465 7147 19499
rect 7147 19465 7156 19499
rect 7104 19456 7156 19465
rect 8392 19456 8444 19508
rect 4620 19388 4672 19440
rect 7012 19388 7064 19440
rect 16120 19499 16172 19508
rect 4344 19320 4396 19372
rect 4988 19320 5040 19372
rect 5172 19320 5224 19372
rect 5356 19320 5408 19372
rect 5816 19320 5868 19372
rect 6092 19320 6144 19372
rect 6920 19363 6972 19372
rect 6920 19329 6929 19363
rect 6929 19329 6963 19363
rect 6963 19329 6972 19363
rect 6920 19320 6972 19329
rect 7104 19320 7156 19372
rect 7288 19320 7340 19372
rect 7564 19320 7616 19372
rect 8300 19363 8352 19372
rect 8300 19329 8309 19363
rect 8309 19329 8343 19363
rect 8343 19329 8352 19363
rect 8300 19320 8352 19329
rect 8760 19363 8812 19372
rect 8760 19329 8769 19363
rect 8769 19329 8803 19363
rect 8803 19329 8812 19363
rect 8760 19320 8812 19329
rect 9220 19320 9272 19372
rect 9772 19363 9824 19372
rect 9772 19329 9781 19363
rect 9781 19329 9815 19363
rect 9815 19329 9824 19363
rect 9772 19320 9824 19329
rect 10508 19320 10560 19372
rect 11888 19363 11940 19372
rect 11888 19329 11897 19363
rect 11897 19329 11931 19363
rect 11931 19329 11940 19363
rect 11888 19320 11940 19329
rect 12164 19320 12216 19372
rect 14464 19388 14516 19440
rect 13636 19320 13688 19372
rect 15384 19388 15436 19440
rect 16120 19465 16129 19499
rect 16129 19465 16163 19499
rect 16163 19465 16172 19499
rect 16120 19456 16172 19465
rect 17316 19456 17368 19508
rect 18052 19456 18104 19508
rect 18512 19499 18564 19508
rect 18512 19465 18521 19499
rect 18521 19465 18555 19499
rect 18555 19465 18564 19499
rect 18512 19456 18564 19465
rect 19248 19456 19300 19508
rect 21272 19499 21324 19508
rect 17960 19388 18012 19440
rect 18788 19388 18840 19440
rect 21272 19465 21281 19499
rect 21281 19465 21315 19499
rect 21315 19465 21324 19499
rect 21272 19456 21324 19465
rect 14832 19320 14884 19372
rect 17040 19320 17092 19372
rect 17132 19320 17184 19372
rect 17776 19363 17828 19372
rect 17776 19329 17785 19363
rect 17785 19329 17819 19363
rect 17819 19329 17828 19363
rect 17776 19320 17828 19329
rect 17868 19320 17920 19372
rect 18880 19363 18932 19372
rect 18880 19329 18889 19363
rect 18889 19329 18923 19363
rect 18923 19329 18932 19363
rect 18880 19320 18932 19329
rect 19432 19363 19484 19372
rect 19432 19329 19441 19363
rect 19441 19329 19475 19363
rect 19475 19329 19484 19363
rect 19432 19320 19484 19329
rect 19616 19320 19668 19372
rect 20536 19363 20588 19372
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 21180 19320 21232 19372
rect 9036 19252 9088 19304
rect 2688 19184 2740 19236
rect 5080 19227 5132 19236
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 1860 19159 1912 19168
rect 1860 19125 1869 19159
rect 1869 19125 1903 19159
rect 1903 19125 1912 19159
rect 1860 19116 1912 19125
rect 2596 19159 2648 19168
rect 2596 19125 2605 19159
rect 2605 19125 2639 19159
rect 2639 19125 2648 19159
rect 2596 19116 2648 19125
rect 4804 19116 4856 19168
rect 5080 19193 5089 19227
rect 5089 19193 5123 19227
rect 5123 19193 5132 19227
rect 5080 19184 5132 19193
rect 5356 19159 5408 19168
rect 5356 19125 5365 19159
rect 5365 19125 5399 19159
rect 5399 19125 5408 19159
rect 5356 19116 5408 19125
rect 8116 19184 8168 19236
rect 9680 19252 9732 19304
rect 11244 19252 11296 19304
rect 12072 19295 12124 19304
rect 12072 19261 12081 19295
rect 12081 19261 12115 19295
rect 12115 19261 12124 19295
rect 13084 19295 13136 19304
rect 12072 19252 12124 19261
rect 13084 19261 13093 19295
rect 13093 19261 13127 19295
rect 13127 19261 13136 19295
rect 13084 19252 13136 19261
rect 9588 19184 9640 19236
rect 9312 19159 9364 19168
rect 9312 19125 9321 19159
rect 9321 19125 9355 19159
rect 9355 19125 9364 19159
rect 9312 19116 9364 19125
rect 11060 19116 11112 19168
rect 11244 19116 11296 19168
rect 14372 19116 14424 19168
rect 14556 19116 14608 19168
rect 19340 19252 19392 19304
rect 19524 19252 19576 19304
rect 22652 19252 22704 19304
rect 20996 19184 21048 19236
rect 19524 19116 19576 19168
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 1584 18955 1636 18964
rect 1584 18921 1593 18955
rect 1593 18921 1627 18955
rect 1627 18921 1636 18955
rect 1584 18912 1636 18921
rect 2412 18912 2464 18964
rect 4068 18912 4120 18964
rect 4804 18912 4856 18964
rect 5080 18912 5132 18964
rect 5356 18955 5408 18964
rect 5356 18921 5365 18955
rect 5365 18921 5399 18955
rect 5399 18921 5408 18955
rect 5356 18912 5408 18921
rect 5816 18955 5868 18964
rect 5816 18921 5825 18955
rect 5825 18921 5859 18955
rect 5859 18921 5868 18955
rect 5816 18912 5868 18921
rect 6552 18912 6604 18964
rect 6644 18844 6696 18896
rect 4068 18819 4120 18828
rect 4068 18785 4077 18819
rect 4077 18785 4111 18819
rect 4111 18785 4120 18819
rect 4068 18776 4120 18785
rect 4896 18776 4948 18828
rect 7104 18912 7156 18964
rect 7472 18912 7524 18964
rect 8208 18912 8260 18964
rect 8576 18912 8628 18964
rect 6828 18844 6880 18896
rect 8484 18844 8536 18896
rect 10232 18912 10284 18964
rect 10600 18955 10652 18964
rect 10600 18921 10609 18955
rect 10609 18921 10643 18955
rect 10643 18921 10652 18955
rect 10600 18912 10652 18921
rect 10416 18844 10468 18896
rect 4712 18751 4764 18760
rect 4712 18717 4721 18751
rect 4721 18717 4755 18751
rect 4755 18717 4764 18751
rect 4712 18708 4764 18717
rect 5172 18751 5224 18760
rect 5172 18717 5181 18751
rect 5181 18717 5215 18751
rect 5215 18717 5224 18751
rect 5172 18708 5224 18717
rect 5356 18708 5408 18760
rect 1860 18640 1912 18692
rect 4804 18640 4856 18692
rect 4896 18640 4948 18692
rect 6460 18708 6512 18760
rect 6644 18708 6696 18760
rect 8576 18751 8628 18760
rect 8300 18640 8352 18692
rect 2412 18572 2464 18624
rect 4712 18572 4764 18624
rect 7380 18572 7432 18624
rect 7656 18615 7708 18624
rect 7656 18581 7665 18615
rect 7665 18581 7699 18615
rect 7699 18581 7708 18615
rect 7656 18572 7708 18581
rect 8576 18717 8585 18751
rect 8585 18717 8619 18751
rect 8619 18717 8628 18751
rect 8576 18708 8628 18717
rect 9772 18708 9824 18760
rect 9956 18708 10008 18760
rect 11060 18776 11112 18828
rect 12256 18912 12308 18964
rect 12992 18912 13044 18964
rect 16948 18912 17000 18964
rect 18696 18912 18748 18964
rect 12900 18844 12952 18896
rect 14556 18844 14608 18896
rect 14372 18819 14424 18828
rect 14372 18785 14381 18819
rect 14381 18785 14415 18819
rect 14415 18785 14424 18819
rect 14372 18776 14424 18785
rect 10968 18708 11020 18760
rect 11888 18751 11940 18760
rect 11888 18717 11897 18751
rect 11897 18717 11931 18751
rect 11931 18717 11940 18751
rect 11888 18708 11940 18717
rect 13084 18708 13136 18760
rect 13544 18751 13596 18760
rect 13544 18717 13553 18751
rect 13553 18717 13587 18751
rect 13587 18717 13596 18751
rect 13544 18708 13596 18717
rect 13728 18708 13780 18760
rect 15384 18751 15436 18760
rect 15384 18717 15393 18751
rect 15393 18717 15427 18751
rect 15427 18717 15436 18751
rect 15384 18708 15436 18717
rect 16120 18708 16172 18760
rect 10784 18640 10836 18692
rect 11244 18683 11296 18692
rect 11244 18649 11253 18683
rect 11253 18649 11287 18683
rect 11287 18649 11296 18683
rect 11244 18640 11296 18649
rect 13268 18640 13320 18692
rect 10876 18615 10928 18624
rect 10876 18581 10885 18615
rect 10885 18581 10919 18615
rect 10919 18581 10928 18615
rect 10876 18572 10928 18581
rect 11704 18572 11756 18624
rect 11796 18572 11848 18624
rect 15476 18640 15528 18692
rect 15752 18640 15804 18692
rect 17224 18751 17276 18760
rect 17224 18717 17233 18751
rect 17233 18717 17267 18751
rect 17267 18717 17276 18751
rect 17224 18708 17276 18717
rect 18052 18708 18104 18760
rect 18420 18708 18472 18760
rect 19524 18708 19576 18760
rect 20904 18708 20956 18760
rect 14464 18572 14516 18624
rect 14924 18615 14976 18624
rect 14924 18581 14933 18615
rect 14933 18581 14967 18615
rect 14967 18581 14976 18615
rect 14924 18572 14976 18581
rect 15016 18572 15068 18624
rect 16488 18640 16540 18692
rect 18696 18640 18748 18692
rect 19708 18640 19760 18692
rect 16396 18572 16448 18624
rect 16948 18572 17000 18624
rect 17316 18572 17368 18624
rect 18972 18572 19024 18624
rect 20260 18615 20312 18624
rect 20260 18581 20269 18615
rect 20269 18581 20303 18615
rect 20303 18581 20312 18615
rect 20260 18572 20312 18581
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 2136 18411 2188 18420
rect 2136 18377 2145 18411
rect 2145 18377 2179 18411
rect 2179 18377 2188 18411
rect 2136 18368 2188 18377
rect 2872 18411 2924 18420
rect 2872 18377 2881 18411
rect 2881 18377 2915 18411
rect 2915 18377 2924 18411
rect 2872 18368 2924 18377
rect 4068 18368 4120 18420
rect 4160 18300 4212 18352
rect 5356 18300 5408 18352
rect 5908 18368 5960 18420
rect 6552 18368 6604 18420
rect 7288 18411 7340 18420
rect 7288 18377 7297 18411
rect 7297 18377 7331 18411
rect 7331 18377 7340 18411
rect 7288 18368 7340 18377
rect 9036 18368 9088 18420
rect 9312 18368 9364 18420
rect 10232 18368 10284 18420
rect 10508 18411 10560 18420
rect 10508 18377 10517 18411
rect 10517 18377 10551 18411
rect 10551 18377 10560 18411
rect 10508 18368 10560 18377
rect 10784 18368 10836 18420
rect 5632 18232 5684 18284
rect 3240 18207 3292 18216
rect 3240 18173 3249 18207
rect 3249 18173 3283 18207
rect 3283 18173 3292 18207
rect 3240 18164 3292 18173
rect 7012 18300 7064 18352
rect 7196 18300 7248 18352
rect 8208 18300 8260 18352
rect 8668 18300 8720 18352
rect 6736 18232 6788 18284
rect 9036 18232 9088 18284
rect 9496 18232 9548 18284
rect 9680 18300 9732 18352
rect 10600 18300 10652 18352
rect 11704 18368 11756 18420
rect 11888 18368 11940 18420
rect 12256 18368 12308 18420
rect 12900 18411 12952 18420
rect 12900 18377 12909 18411
rect 12909 18377 12943 18411
rect 12943 18377 12952 18411
rect 12900 18368 12952 18377
rect 13636 18368 13688 18420
rect 14924 18368 14976 18420
rect 15476 18368 15528 18420
rect 17408 18368 17460 18420
rect 18604 18368 18656 18420
rect 18696 18368 18748 18420
rect 20812 18368 20864 18420
rect 10876 18232 10928 18284
rect 15292 18300 15344 18352
rect 11888 18275 11940 18284
rect 11888 18241 11897 18275
rect 11897 18241 11931 18275
rect 11931 18241 11940 18275
rect 11888 18232 11940 18241
rect 12716 18275 12768 18284
rect 12716 18241 12725 18275
rect 12725 18241 12759 18275
rect 12759 18241 12768 18275
rect 12716 18232 12768 18241
rect 12992 18232 13044 18284
rect 14280 18232 14332 18284
rect 14924 18232 14976 18284
rect 16304 18300 16356 18352
rect 16396 18300 16448 18352
rect 16028 18275 16080 18284
rect 16028 18241 16037 18275
rect 16037 18241 16071 18275
rect 16071 18241 16080 18275
rect 16028 18232 16080 18241
rect 7104 18164 7156 18216
rect 7288 18164 7340 18216
rect 8668 18164 8720 18216
rect 9404 18164 9456 18216
rect 2688 18096 2740 18148
rect 2780 18096 2832 18148
rect 6828 18139 6880 18148
rect 4804 18028 4856 18080
rect 5080 18071 5132 18080
rect 5080 18037 5089 18071
rect 5089 18037 5123 18071
rect 5123 18037 5132 18071
rect 5080 18028 5132 18037
rect 6828 18105 6837 18139
rect 6837 18105 6871 18139
rect 6871 18105 6880 18139
rect 6828 18096 6880 18105
rect 7012 18096 7064 18148
rect 7196 18096 7248 18148
rect 10600 18164 10652 18216
rect 10692 18164 10744 18216
rect 12072 18207 12124 18216
rect 12072 18173 12081 18207
rect 12081 18173 12115 18207
rect 12115 18173 12124 18207
rect 12072 18164 12124 18173
rect 9772 18096 9824 18148
rect 10508 18096 10560 18148
rect 14372 18164 14424 18216
rect 15108 18164 15160 18216
rect 12348 18096 12400 18148
rect 16764 18164 16816 18216
rect 19800 18300 19852 18352
rect 19984 18343 20036 18352
rect 19984 18309 19993 18343
rect 19993 18309 20027 18343
rect 20027 18309 20036 18343
rect 19984 18300 20036 18309
rect 18236 18275 18288 18284
rect 18236 18241 18270 18275
rect 18270 18241 18288 18275
rect 18236 18232 18288 18241
rect 17040 18207 17092 18216
rect 17040 18173 17049 18207
rect 17049 18173 17083 18207
rect 17083 18173 17092 18207
rect 17040 18164 17092 18173
rect 17960 18207 18012 18216
rect 17960 18173 17969 18207
rect 17969 18173 18003 18207
rect 18003 18173 18012 18207
rect 17960 18164 18012 18173
rect 20812 18232 20864 18284
rect 17868 18096 17920 18148
rect 7932 18028 7984 18080
rect 8392 18028 8444 18080
rect 8668 18071 8720 18080
rect 8668 18037 8677 18071
rect 8677 18037 8711 18071
rect 8711 18037 8720 18071
rect 8668 18028 8720 18037
rect 9588 18028 9640 18080
rect 10140 18071 10192 18080
rect 10140 18037 10149 18071
rect 10149 18037 10183 18071
rect 10183 18037 10192 18071
rect 10140 18028 10192 18037
rect 10232 18028 10284 18080
rect 12072 18028 12124 18080
rect 17408 18028 17460 18080
rect 18144 18028 18196 18080
rect 19524 18028 19576 18080
rect 20352 18071 20404 18080
rect 20352 18037 20361 18071
rect 20361 18037 20395 18071
rect 20395 18037 20404 18071
rect 20352 18028 20404 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 5172 17867 5224 17876
rect 5172 17833 5181 17867
rect 5181 17833 5215 17867
rect 5215 17833 5224 17867
rect 5172 17824 5224 17833
rect 6920 17824 6972 17876
rect 7012 17824 7064 17876
rect 7288 17824 7340 17876
rect 10600 17867 10652 17876
rect 10600 17833 10609 17867
rect 10609 17833 10643 17867
rect 10643 17833 10652 17867
rect 10600 17824 10652 17833
rect 11060 17824 11112 17876
rect 12716 17867 12768 17876
rect 12716 17833 12725 17867
rect 12725 17833 12759 17867
rect 12759 17833 12768 17867
rect 12716 17824 12768 17833
rect 13360 17824 13412 17876
rect 10968 17756 11020 17808
rect 11244 17756 11296 17808
rect 4344 17688 4396 17740
rect 5172 17688 5224 17740
rect 3516 17620 3568 17672
rect 3976 17620 4028 17672
rect 5632 17620 5684 17672
rect 6920 17620 6972 17672
rect 10232 17688 10284 17740
rect 13176 17731 13228 17740
rect 13176 17697 13185 17731
rect 13185 17697 13219 17731
rect 13219 17697 13228 17731
rect 13176 17688 13228 17697
rect 13544 17756 13596 17808
rect 15108 17756 15160 17808
rect 14280 17731 14332 17740
rect 14280 17697 14289 17731
rect 14289 17697 14323 17731
rect 14323 17697 14332 17731
rect 14280 17688 14332 17697
rect 19892 17756 19944 17808
rect 19984 17799 20036 17808
rect 19984 17765 19993 17799
rect 19993 17765 20027 17799
rect 20027 17765 20036 17799
rect 19984 17756 20036 17765
rect 18052 17688 18104 17740
rect 18236 17688 18288 17740
rect 19524 17688 19576 17740
rect 8392 17620 8444 17672
rect 9956 17620 10008 17672
rect 10324 17620 10376 17672
rect 11704 17620 11756 17672
rect 13820 17620 13872 17672
rect 14556 17620 14608 17672
rect 16120 17663 16172 17672
rect 16120 17629 16129 17663
rect 16129 17629 16163 17663
rect 16163 17629 16172 17663
rect 16120 17620 16172 17629
rect 16396 17663 16448 17672
rect 16396 17629 16430 17663
rect 16430 17629 16448 17663
rect 16396 17620 16448 17629
rect 18144 17663 18196 17672
rect 18144 17629 18153 17663
rect 18153 17629 18187 17663
rect 18187 17629 18196 17663
rect 18144 17620 18196 17629
rect 20352 17620 20404 17672
rect 6736 17552 6788 17604
rect 7012 17552 7064 17604
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 1952 17527 2004 17536
rect 1952 17493 1961 17527
rect 1961 17493 1995 17527
rect 1995 17493 2004 17527
rect 1952 17484 2004 17493
rect 2688 17527 2740 17536
rect 2688 17493 2697 17527
rect 2697 17493 2731 17527
rect 2731 17493 2740 17527
rect 2688 17484 2740 17493
rect 4252 17484 4304 17536
rect 4712 17527 4764 17536
rect 4712 17493 4721 17527
rect 4721 17493 4755 17527
rect 4755 17493 4764 17527
rect 4712 17484 4764 17493
rect 8116 17484 8168 17536
rect 9496 17552 9548 17604
rect 11336 17552 11388 17604
rect 13636 17552 13688 17604
rect 16304 17552 16356 17604
rect 19524 17595 19576 17604
rect 19524 17561 19533 17595
rect 19533 17561 19567 17595
rect 19567 17561 19576 17595
rect 19524 17552 19576 17561
rect 19984 17552 20036 17604
rect 10232 17484 10284 17536
rect 10324 17527 10376 17536
rect 10324 17493 10333 17527
rect 10333 17493 10367 17527
rect 10367 17493 10376 17527
rect 10968 17527 11020 17536
rect 10324 17484 10376 17493
rect 10968 17493 10977 17527
rect 10977 17493 11011 17527
rect 11011 17493 11020 17527
rect 10968 17484 11020 17493
rect 13544 17484 13596 17536
rect 14464 17527 14516 17536
rect 14464 17493 14473 17527
rect 14473 17493 14507 17527
rect 14507 17493 14516 17527
rect 14832 17527 14884 17536
rect 14464 17484 14516 17493
rect 14832 17493 14841 17527
rect 14841 17493 14875 17527
rect 14875 17493 14884 17527
rect 14832 17484 14884 17493
rect 18052 17527 18104 17536
rect 18052 17493 18061 17527
rect 18061 17493 18095 17527
rect 18095 17493 18104 17527
rect 18052 17484 18104 17493
rect 18144 17484 18196 17536
rect 21548 17552 21600 17604
rect 21456 17484 21508 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 1400 17323 1452 17332
rect 1400 17289 1409 17323
rect 1409 17289 1443 17323
rect 1443 17289 1452 17323
rect 1400 17280 1452 17289
rect 2044 17280 2096 17332
rect 2228 17323 2280 17332
rect 2228 17289 2237 17323
rect 2237 17289 2271 17323
rect 2271 17289 2280 17323
rect 2228 17280 2280 17289
rect 3056 17323 3108 17332
rect 3056 17289 3065 17323
rect 3065 17289 3099 17323
rect 3099 17289 3108 17323
rect 3056 17280 3108 17289
rect 3424 17323 3476 17332
rect 3424 17289 3433 17323
rect 3433 17289 3467 17323
rect 3467 17289 3476 17323
rect 3424 17280 3476 17289
rect 5264 17280 5316 17332
rect 3148 17212 3200 17264
rect 1584 17076 1636 17128
rect 5908 17212 5960 17264
rect 6552 17280 6604 17332
rect 7656 17280 7708 17332
rect 6092 17212 6144 17264
rect 4896 17187 4948 17196
rect 4896 17153 4905 17187
rect 4905 17153 4939 17187
rect 4939 17153 4948 17187
rect 4896 17144 4948 17153
rect 5356 17076 5408 17128
rect 6736 17144 6788 17196
rect 6920 17187 6972 17196
rect 6920 17153 6929 17187
rect 6929 17153 6963 17187
rect 6963 17153 6972 17187
rect 6920 17144 6972 17153
rect 7932 17144 7984 17196
rect 8116 17255 8168 17264
rect 8116 17221 8150 17255
rect 8150 17221 8168 17255
rect 8116 17212 8168 17221
rect 9680 17280 9732 17332
rect 9772 17280 9824 17332
rect 9128 17212 9180 17264
rect 10968 17280 11020 17332
rect 14556 17323 14608 17332
rect 10876 17212 10928 17264
rect 12440 17212 12492 17264
rect 7104 17076 7156 17128
rect 11520 17144 11572 17196
rect 14556 17289 14565 17323
rect 14565 17289 14599 17323
rect 14599 17289 14608 17323
rect 14556 17280 14608 17289
rect 17500 17280 17552 17332
rect 17684 17280 17736 17332
rect 18144 17280 18196 17332
rect 18236 17280 18288 17332
rect 15108 17212 15160 17264
rect 16304 17212 16356 17264
rect 13176 17187 13228 17196
rect 13176 17153 13210 17187
rect 13210 17153 13228 17187
rect 13176 17144 13228 17153
rect 14280 17144 14332 17196
rect 16764 17144 16816 17196
rect 9312 17076 9364 17128
rect 10232 17119 10284 17128
rect 10232 17085 10241 17119
rect 10241 17085 10275 17119
rect 10275 17085 10284 17119
rect 10232 17076 10284 17085
rect 1676 17008 1728 17060
rect 4252 16940 4304 16992
rect 6092 16940 6144 16992
rect 6828 16940 6880 16992
rect 7564 16983 7616 16992
rect 7564 16949 7573 16983
rect 7573 16949 7607 16983
rect 7607 16949 7616 16983
rect 7564 16940 7616 16949
rect 9496 16940 9548 16992
rect 9680 16940 9732 16992
rect 11704 17076 11756 17128
rect 12256 17076 12308 17128
rect 10876 17008 10928 17060
rect 12808 17008 12860 17060
rect 16120 17076 16172 17128
rect 16304 17076 16356 17128
rect 17960 17212 18012 17264
rect 18972 17255 19024 17264
rect 17316 17187 17368 17196
rect 17316 17153 17350 17187
rect 17350 17153 17368 17187
rect 17316 17144 17368 17153
rect 18972 17221 19006 17255
rect 19006 17221 19024 17255
rect 18972 17212 19024 17221
rect 18144 17076 18196 17128
rect 20628 17144 20680 17196
rect 20996 17187 21048 17196
rect 20996 17153 21005 17187
rect 21005 17153 21039 17187
rect 21039 17153 21048 17187
rect 20996 17144 21048 17153
rect 10784 16940 10836 16992
rect 11888 16940 11940 16992
rect 12164 16940 12216 16992
rect 13820 16940 13872 16992
rect 15660 16940 15712 16992
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 19984 16940 20036 16992
rect 20444 16940 20496 16992
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 1860 16779 1912 16788
rect 1860 16745 1869 16779
rect 1869 16745 1903 16779
rect 1903 16745 1912 16779
rect 1860 16736 1912 16745
rect 2504 16779 2556 16788
rect 2504 16745 2513 16779
rect 2513 16745 2547 16779
rect 2547 16745 2556 16779
rect 2504 16736 2556 16745
rect 4620 16736 4672 16788
rect 4988 16779 5040 16788
rect 4988 16745 4997 16779
rect 4997 16745 5031 16779
rect 5031 16745 5040 16779
rect 4988 16736 5040 16745
rect 5356 16779 5408 16788
rect 5356 16745 5365 16779
rect 5365 16745 5399 16779
rect 5399 16745 5408 16779
rect 5356 16736 5408 16745
rect 5540 16736 5592 16788
rect 6920 16779 6972 16788
rect 6920 16745 6929 16779
rect 6929 16745 6963 16779
rect 6963 16745 6972 16779
rect 6920 16736 6972 16745
rect 7932 16736 7984 16788
rect 6000 16668 6052 16720
rect 8392 16736 8444 16788
rect 9680 16736 9732 16788
rect 9956 16736 10008 16788
rect 5356 16600 5408 16652
rect 5632 16600 5684 16652
rect 9312 16643 9364 16652
rect 9312 16609 9321 16643
rect 9321 16609 9355 16643
rect 9355 16609 9364 16643
rect 9312 16600 9364 16609
rect 9496 16643 9548 16652
rect 9496 16609 9505 16643
rect 9505 16609 9539 16643
rect 9539 16609 9548 16643
rect 9496 16600 9548 16609
rect 9588 16600 9640 16652
rect 11152 16736 11204 16788
rect 12256 16736 12308 16788
rect 12808 16736 12860 16788
rect 15200 16736 15252 16788
rect 15936 16779 15988 16788
rect 15936 16745 15945 16779
rect 15945 16745 15979 16779
rect 15979 16745 15988 16779
rect 15936 16736 15988 16745
rect 18052 16736 18104 16788
rect 20628 16736 20680 16788
rect 13176 16668 13228 16720
rect 9956 16532 10008 16584
rect 12164 16575 12216 16584
rect 10232 16464 10284 16516
rect 10692 16464 10744 16516
rect 11520 16464 11572 16516
rect 12164 16541 12198 16575
rect 12198 16541 12216 16575
rect 12164 16532 12216 16541
rect 14556 16668 14608 16720
rect 15844 16668 15896 16720
rect 20168 16668 20220 16720
rect 14832 16600 14884 16652
rect 14740 16532 14792 16584
rect 16764 16643 16816 16652
rect 15568 16575 15620 16584
rect 15568 16541 15577 16575
rect 15577 16541 15611 16575
rect 15611 16541 15620 16575
rect 15568 16532 15620 16541
rect 16764 16609 16773 16643
rect 16773 16609 16807 16643
rect 16807 16609 16816 16643
rect 16764 16600 16816 16609
rect 19248 16600 19300 16652
rect 17684 16575 17736 16584
rect 17684 16541 17693 16575
rect 17693 16541 17727 16575
rect 17727 16541 17736 16575
rect 18880 16575 18932 16584
rect 17684 16532 17736 16541
rect 18880 16541 18889 16575
rect 18889 16541 18923 16575
rect 18923 16541 18932 16575
rect 18880 16532 18932 16541
rect 2688 16396 2740 16448
rect 6552 16396 6604 16448
rect 9312 16396 9364 16448
rect 9588 16439 9640 16448
rect 9588 16405 9597 16439
rect 9597 16405 9631 16439
rect 9631 16405 9640 16439
rect 9588 16396 9640 16405
rect 9680 16396 9732 16448
rect 13544 16396 13596 16448
rect 13912 16396 13964 16448
rect 14372 16396 14424 16448
rect 14556 16396 14608 16448
rect 15016 16396 15068 16448
rect 15568 16396 15620 16448
rect 15936 16464 15988 16516
rect 16948 16464 17000 16516
rect 19616 16532 19668 16584
rect 19800 16643 19852 16652
rect 19800 16609 19809 16643
rect 19809 16609 19843 16643
rect 19843 16609 19852 16643
rect 19800 16600 19852 16609
rect 20996 16600 21048 16652
rect 19524 16464 19576 16516
rect 20076 16464 20128 16516
rect 17592 16439 17644 16448
rect 17592 16405 17601 16439
rect 17601 16405 17635 16439
rect 17635 16405 17644 16439
rect 17592 16396 17644 16405
rect 17776 16396 17828 16448
rect 19800 16396 19852 16448
rect 20260 16439 20312 16448
rect 20260 16405 20269 16439
rect 20269 16405 20303 16439
rect 20303 16405 20312 16439
rect 20260 16396 20312 16405
rect 20352 16396 20404 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 4528 16192 4580 16244
rect 9680 16235 9732 16244
rect 5816 16124 5868 16176
rect 4620 15920 4672 15972
rect 5448 16056 5500 16108
rect 7932 16124 7984 16176
rect 9680 16201 9689 16235
rect 9689 16201 9723 16235
rect 9723 16201 9732 16235
rect 9680 16192 9732 16201
rect 11704 16235 11756 16244
rect 7564 16056 7616 16108
rect 5264 15988 5316 16040
rect 5632 16031 5684 16040
rect 5632 15997 5641 16031
rect 5641 15997 5675 16031
rect 5675 15997 5684 16031
rect 5632 15988 5684 15997
rect 9772 15988 9824 16040
rect 10692 16124 10744 16176
rect 10784 16099 10836 16108
rect 10784 16065 10793 16099
rect 10793 16065 10827 16099
rect 10827 16065 10836 16099
rect 10784 16056 10836 16065
rect 10876 16031 10928 16040
rect 10876 15997 10885 16031
rect 10885 15997 10919 16031
rect 10919 15997 10928 16031
rect 10876 15988 10928 15997
rect 10968 16031 11020 16040
rect 10968 15997 10977 16031
rect 10977 15997 11011 16031
rect 11011 15997 11020 16031
rect 11704 16201 11713 16235
rect 11713 16201 11747 16235
rect 11747 16201 11756 16235
rect 11704 16192 11756 16201
rect 13728 16192 13780 16244
rect 17684 16124 17736 16176
rect 19248 16192 19300 16244
rect 20076 16235 20128 16244
rect 20076 16201 20085 16235
rect 20085 16201 20119 16235
rect 20119 16201 20128 16235
rect 20076 16192 20128 16201
rect 20352 16235 20404 16244
rect 20352 16201 20361 16235
rect 20361 16201 20395 16235
rect 20395 16201 20404 16235
rect 20352 16192 20404 16201
rect 12440 16056 12492 16108
rect 10968 15988 11020 15997
rect 13544 16031 13596 16040
rect 13544 15997 13553 16031
rect 13553 15997 13587 16031
rect 13587 15997 13596 16031
rect 13544 15988 13596 15997
rect 6920 15920 6972 15972
rect 4988 15852 5040 15904
rect 7288 15920 7340 15972
rect 14372 16056 14424 16108
rect 16212 16056 16264 16108
rect 17408 16099 17460 16108
rect 17408 16065 17417 16099
rect 17417 16065 17451 16099
rect 17451 16065 17460 16099
rect 17408 16056 17460 16065
rect 19984 16124 20036 16176
rect 16304 16031 16356 16040
rect 16304 15997 16313 16031
rect 16313 15997 16347 16031
rect 16347 15997 16356 16031
rect 16304 15988 16356 15997
rect 13912 15920 13964 15972
rect 8116 15852 8168 15904
rect 9128 15852 9180 15904
rect 9404 15852 9456 15904
rect 10968 15852 11020 15904
rect 12532 15852 12584 15904
rect 14280 15852 14332 15904
rect 14924 15895 14976 15904
rect 14924 15861 14933 15895
rect 14933 15861 14967 15895
rect 14967 15861 14976 15895
rect 14924 15852 14976 15861
rect 16948 15920 17000 15972
rect 18972 15920 19024 15972
rect 20720 16099 20772 16108
rect 20720 16065 20729 16099
rect 20729 16065 20763 16099
rect 20763 16065 20772 16099
rect 20720 16056 20772 16065
rect 18420 15852 18472 15904
rect 18604 15852 18656 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 7012 15648 7064 15700
rect 5540 15580 5592 15632
rect 6736 15580 6788 15632
rect 9588 15648 9640 15700
rect 9956 15691 10008 15700
rect 9956 15657 9965 15691
rect 9965 15657 9999 15691
rect 9999 15657 10008 15691
rect 9956 15648 10008 15657
rect 11152 15648 11204 15700
rect 12440 15691 12492 15700
rect 12440 15657 12449 15691
rect 12449 15657 12483 15691
rect 12483 15657 12492 15691
rect 12440 15648 12492 15657
rect 14464 15648 14516 15700
rect 16028 15648 16080 15700
rect 17684 15691 17736 15700
rect 17684 15657 17693 15691
rect 17693 15657 17727 15691
rect 17727 15657 17736 15691
rect 17684 15648 17736 15657
rect 10232 15580 10284 15632
rect 13636 15580 13688 15632
rect 14004 15580 14056 15632
rect 16304 15580 16356 15632
rect 17408 15580 17460 15632
rect 20260 15648 20312 15700
rect 18696 15623 18748 15632
rect 18696 15589 18705 15623
rect 18705 15589 18739 15623
rect 18739 15589 18748 15623
rect 18696 15580 18748 15589
rect 8116 15555 8168 15564
rect 8116 15521 8125 15555
rect 8125 15521 8159 15555
rect 8159 15521 8168 15555
rect 8116 15512 8168 15521
rect 9128 15555 9180 15564
rect 9128 15521 9137 15555
rect 9137 15521 9171 15555
rect 9171 15521 9180 15555
rect 9128 15512 9180 15521
rect 10968 15512 11020 15564
rect 6460 15487 6512 15496
rect 6460 15453 6469 15487
rect 6469 15453 6503 15487
rect 6503 15453 6512 15487
rect 6460 15444 6512 15453
rect 7748 15444 7800 15496
rect 9312 15487 9364 15496
rect 9312 15453 9321 15487
rect 9321 15453 9355 15487
rect 9355 15453 9364 15487
rect 9312 15444 9364 15453
rect 10140 15487 10192 15496
rect 10140 15453 10149 15487
rect 10149 15453 10183 15487
rect 10183 15453 10192 15487
rect 10140 15444 10192 15453
rect 13820 15512 13872 15564
rect 14464 15512 14516 15564
rect 14740 15555 14792 15564
rect 14740 15521 14749 15555
rect 14749 15521 14783 15555
rect 14783 15521 14792 15555
rect 14740 15512 14792 15521
rect 14924 15512 14976 15564
rect 6184 15419 6236 15428
rect 6184 15385 6193 15419
rect 6193 15385 6227 15419
rect 6227 15385 6236 15419
rect 6184 15376 6236 15385
rect 5816 15308 5868 15360
rect 6920 15376 6972 15428
rect 7288 15376 7340 15428
rect 8208 15419 8260 15428
rect 8208 15385 8217 15419
rect 8217 15385 8251 15419
rect 8251 15385 8260 15419
rect 8208 15376 8260 15385
rect 10876 15376 10928 15428
rect 12164 15419 12216 15428
rect 12164 15385 12173 15419
rect 12173 15385 12207 15419
rect 12207 15385 12216 15419
rect 12164 15376 12216 15385
rect 13544 15376 13596 15428
rect 18052 15444 18104 15496
rect 20628 15487 20680 15496
rect 15660 15419 15712 15428
rect 15660 15385 15669 15419
rect 15669 15385 15703 15419
rect 15703 15385 15712 15419
rect 15660 15376 15712 15385
rect 6644 15351 6696 15360
rect 6644 15317 6653 15351
rect 6653 15317 6687 15351
rect 6687 15317 6696 15351
rect 6644 15308 6696 15317
rect 8668 15308 8720 15360
rect 8760 15308 8812 15360
rect 9588 15308 9640 15360
rect 9864 15308 9916 15360
rect 12256 15308 12308 15360
rect 13820 15308 13872 15360
rect 14556 15351 14608 15360
rect 14556 15317 14565 15351
rect 14565 15317 14599 15351
rect 14599 15317 14608 15351
rect 14556 15308 14608 15317
rect 15108 15308 15160 15360
rect 18236 15376 18288 15428
rect 18972 15376 19024 15428
rect 19800 15376 19852 15428
rect 20628 15453 20637 15487
rect 20637 15453 20671 15487
rect 20671 15453 20680 15487
rect 20628 15444 20680 15453
rect 20444 15376 20496 15428
rect 19248 15351 19300 15360
rect 19248 15317 19257 15351
rect 19257 15317 19291 15351
rect 19291 15317 19300 15351
rect 19248 15308 19300 15317
rect 20076 15308 20128 15360
rect 21364 15308 21416 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 7196 15104 7248 15156
rect 8760 15104 8812 15156
rect 8116 14968 8168 15020
rect 9128 15104 9180 15156
rect 9772 15147 9824 15156
rect 9772 15113 9781 15147
rect 9781 15113 9815 15147
rect 9815 15113 9824 15147
rect 9772 15104 9824 15113
rect 11244 15104 11296 15156
rect 11704 15104 11756 15156
rect 12072 15104 12124 15156
rect 12256 15104 12308 15156
rect 10876 15011 10928 15020
rect 10876 14977 10894 15011
rect 10894 14977 10928 15011
rect 11796 15036 11848 15088
rect 12440 15036 12492 15088
rect 14280 15079 14332 15088
rect 14280 15045 14314 15079
rect 14314 15045 14332 15079
rect 14280 15036 14332 15045
rect 16212 15104 16264 15156
rect 18328 15104 18380 15156
rect 17040 15036 17092 15088
rect 17592 15036 17644 15088
rect 18512 15104 18564 15156
rect 19432 15104 19484 15156
rect 20628 15104 20680 15156
rect 20812 15147 20864 15156
rect 20812 15113 20821 15147
rect 20821 15113 20855 15147
rect 20855 15113 20864 15147
rect 20812 15104 20864 15113
rect 11152 15011 11204 15020
rect 10876 14968 10928 14977
rect 11152 14977 11161 15011
rect 11161 14977 11195 15011
rect 11195 14977 11204 15011
rect 11152 14968 11204 14977
rect 12532 15011 12584 15020
rect 12532 14977 12541 15011
rect 12541 14977 12575 15011
rect 12575 14977 12584 15011
rect 12532 14968 12584 14977
rect 14004 15011 14056 15020
rect 14004 14977 14013 15011
rect 14013 14977 14047 15011
rect 14047 14977 14056 15011
rect 14004 14968 14056 14977
rect 14556 14968 14608 15020
rect 14740 14968 14792 15020
rect 9864 14900 9916 14952
rect 11980 14943 12032 14952
rect 11980 14909 11989 14943
rect 11989 14909 12023 14943
rect 12023 14909 12032 14943
rect 11980 14900 12032 14909
rect 13268 14943 13320 14952
rect 6828 14832 6880 14884
rect 6460 14807 6512 14816
rect 6460 14773 6469 14807
rect 6469 14773 6503 14807
rect 6503 14773 6512 14807
rect 6460 14764 6512 14773
rect 7012 14807 7064 14816
rect 7012 14773 7021 14807
rect 7021 14773 7055 14807
rect 7055 14773 7064 14807
rect 7012 14764 7064 14773
rect 7748 14807 7800 14816
rect 7748 14773 7757 14807
rect 7757 14773 7791 14807
rect 7791 14773 7800 14807
rect 7748 14764 7800 14773
rect 11152 14832 11204 14884
rect 13268 14909 13277 14943
rect 13277 14909 13311 14943
rect 13311 14909 13320 14943
rect 13268 14900 13320 14909
rect 13820 14832 13872 14884
rect 11244 14764 11296 14816
rect 13636 14764 13688 14816
rect 14372 14764 14424 14816
rect 14648 14764 14700 14816
rect 16948 14968 17000 15020
rect 17868 15011 17920 15020
rect 17868 14977 17877 15011
rect 17877 14977 17911 15011
rect 17911 14977 17920 15011
rect 17868 14968 17920 14977
rect 15476 14900 15528 14952
rect 17592 14900 17644 14952
rect 19248 15036 19300 15088
rect 20996 15036 21048 15088
rect 19432 15011 19484 15020
rect 19432 14977 19441 15011
rect 19441 14977 19475 15011
rect 19475 14977 19484 15011
rect 19432 14968 19484 14977
rect 18696 14943 18748 14952
rect 18696 14909 18705 14943
rect 18705 14909 18739 14943
rect 18739 14909 18748 14943
rect 18696 14900 18748 14909
rect 20720 14968 20772 15020
rect 21088 15011 21140 15020
rect 21088 14977 21097 15011
rect 21097 14977 21131 15011
rect 21131 14977 21140 15011
rect 21088 14968 21140 14977
rect 15568 14832 15620 14884
rect 17316 14807 17368 14816
rect 17316 14773 17325 14807
rect 17325 14773 17359 14807
rect 17359 14773 17368 14807
rect 17316 14764 17368 14773
rect 20444 14764 20496 14816
rect 21272 14807 21324 14816
rect 21272 14773 21281 14807
rect 21281 14773 21315 14807
rect 21315 14773 21324 14807
rect 21272 14764 21324 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 6552 14560 6604 14612
rect 7012 14560 7064 14612
rect 4436 14492 4488 14544
rect 7748 14492 7800 14544
rect 11888 14535 11940 14544
rect 7012 14424 7064 14476
rect 7196 14467 7248 14476
rect 7196 14433 7205 14467
rect 7205 14433 7239 14467
rect 7239 14433 7248 14467
rect 7196 14424 7248 14433
rect 5540 14356 5592 14408
rect 6000 14356 6052 14408
rect 9128 14424 9180 14476
rect 11888 14501 11897 14535
rect 11897 14501 11931 14535
rect 11931 14501 11940 14535
rect 11888 14492 11940 14501
rect 11244 14424 11296 14476
rect 14004 14492 14056 14544
rect 14188 14467 14240 14476
rect 9588 14399 9640 14408
rect 9312 14288 9364 14340
rect 9588 14365 9597 14399
rect 9597 14365 9631 14399
rect 9631 14365 9640 14399
rect 9588 14356 9640 14365
rect 10876 14356 10928 14408
rect 12348 14399 12400 14408
rect 10048 14288 10100 14340
rect 10968 14288 11020 14340
rect 12348 14365 12357 14399
rect 12357 14365 12391 14399
rect 12391 14365 12400 14399
rect 12348 14356 12400 14365
rect 14188 14433 14197 14467
rect 14197 14433 14231 14467
rect 14231 14433 14240 14467
rect 14188 14424 14240 14433
rect 14372 14467 14424 14476
rect 14372 14433 14381 14467
rect 14381 14433 14415 14467
rect 14415 14433 14424 14467
rect 14372 14424 14424 14433
rect 15568 14467 15620 14476
rect 15568 14433 15577 14467
rect 15577 14433 15611 14467
rect 15611 14433 15620 14467
rect 15568 14424 15620 14433
rect 12256 14288 12308 14340
rect 13820 14288 13872 14340
rect 14096 14288 14148 14340
rect 17868 14560 17920 14612
rect 18788 14603 18840 14612
rect 18788 14569 18797 14603
rect 18797 14569 18831 14603
rect 18831 14569 18840 14603
rect 18788 14560 18840 14569
rect 19616 14603 19668 14612
rect 19616 14569 19625 14603
rect 19625 14569 19659 14603
rect 19659 14569 19668 14603
rect 19616 14560 19668 14569
rect 19524 14424 19576 14476
rect 20444 14467 20496 14476
rect 20444 14433 20453 14467
rect 20453 14433 20487 14467
rect 20487 14433 20496 14467
rect 20444 14424 20496 14433
rect 20812 14424 20864 14476
rect 19432 14399 19484 14408
rect 19432 14365 19441 14399
rect 19441 14365 19475 14399
rect 19475 14365 19484 14399
rect 19432 14356 19484 14365
rect 17776 14288 17828 14340
rect 18236 14288 18288 14340
rect 7748 14220 7800 14272
rect 8300 14220 8352 14272
rect 11704 14220 11756 14272
rect 11888 14220 11940 14272
rect 14004 14220 14056 14272
rect 14464 14263 14516 14272
rect 14464 14229 14473 14263
rect 14473 14229 14507 14263
rect 14507 14229 14516 14263
rect 14832 14263 14884 14272
rect 14464 14220 14516 14229
rect 14832 14229 14841 14263
rect 14841 14229 14875 14263
rect 14875 14229 14884 14263
rect 14832 14220 14884 14229
rect 14924 14220 14976 14272
rect 15476 14263 15528 14272
rect 15476 14229 15485 14263
rect 15485 14229 15519 14263
rect 15519 14229 15528 14263
rect 15476 14220 15528 14229
rect 16212 14220 16264 14272
rect 17224 14220 17276 14272
rect 20352 14263 20404 14272
rect 20352 14229 20361 14263
rect 20361 14229 20395 14263
rect 20395 14229 20404 14263
rect 20352 14220 20404 14229
rect 21180 14263 21232 14272
rect 21180 14229 21189 14263
rect 21189 14229 21223 14263
rect 21223 14229 21232 14263
rect 21180 14220 21232 14229
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 8116 14059 8168 14068
rect 8116 14025 8125 14059
rect 8125 14025 8159 14059
rect 8159 14025 8168 14059
rect 8116 14016 8168 14025
rect 9312 14016 9364 14068
rect 11152 14016 11204 14068
rect 8208 13948 8260 14000
rect 3884 13880 3936 13932
rect 8300 13923 8352 13932
rect 7104 13812 7156 13864
rect 8300 13889 8309 13923
rect 8309 13889 8343 13923
rect 8343 13889 8352 13923
rect 8300 13880 8352 13889
rect 9864 13948 9916 14000
rect 12992 14016 13044 14068
rect 14280 14016 14332 14068
rect 14464 14016 14516 14068
rect 14924 14016 14976 14068
rect 15568 14016 15620 14068
rect 19616 14016 19668 14068
rect 19800 14016 19852 14068
rect 20352 14059 20404 14068
rect 20352 14025 20361 14059
rect 20361 14025 20395 14059
rect 20395 14025 20404 14059
rect 20352 14016 20404 14025
rect 12348 13948 12400 14000
rect 10324 13880 10376 13932
rect 10876 13923 10928 13932
rect 10876 13889 10885 13923
rect 10885 13889 10919 13923
rect 10919 13889 10928 13923
rect 12624 13923 12676 13932
rect 15476 13948 15528 14000
rect 10876 13880 10928 13889
rect 12624 13889 12642 13923
rect 12642 13889 12676 13923
rect 12624 13880 12676 13889
rect 9864 13812 9916 13864
rect 13728 13812 13780 13864
rect 14096 13855 14148 13864
rect 14096 13821 14105 13855
rect 14105 13821 14139 13855
rect 14139 13821 14148 13855
rect 14096 13812 14148 13821
rect 14740 13880 14792 13932
rect 17224 13880 17276 13932
rect 15108 13812 15160 13864
rect 15476 13855 15528 13864
rect 15476 13821 15485 13855
rect 15485 13821 15519 13855
rect 15519 13821 15528 13855
rect 15476 13812 15528 13821
rect 8208 13744 8260 13796
rect 9496 13744 9548 13796
rect 14188 13744 14240 13796
rect 16120 13812 16172 13864
rect 19984 13948 20036 14000
rect 20168 13948 20220 14000
rect 17868 13880 17920 13932
rect 20352 13880 20404 13932
rect 9312 13676 9364 13728
rect 12716 13676 12768 13728
rect 12900 13676 12952 13728
rect 15016 13719 15068 13728
rect 15016 13685 15025 13719
rect 15025 13685 15059 13719
rect 15059 13685 15068 13719
rect 15016 13676 15068 13685
rect 18236 13812 18288 13864
rect 18328 13812 18380 13864
rect 18880 13855 18932 13864
rect 18880 13821 18889 13855
rect 18889 13821 18923 13855
rect 18923 13821 18932 13855
rect 19892 13855 19944 13864
rect 18880 13812 18932 13821
rect 17408 13676 17460 13728
rect 17776 13676 17828 13728
rect 19892 13821 19901 13855
rect 19901 13821 19935 13855
rect 19935 13821 19944 13855
rect 19892 13812 19944 13821
rect 20996 13855 21048 13864
rect 20996 13821 21005 13855
rect 21005 13821 21039 13855
rect 21039 13821 21048 13855
rect 20996 13812 21048 13821
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 5448 13472 5500 13524
rect 9680 13472 9732 13524
rect 10876 13515 10928 13524
rect 10876 13481 10885 13515
rect 10885 13481 10919 13515
rect 10919 13481 10928 13515
rect 10876 13472 10928 13481
rect 12440 13515 12492 13524
rect 12440 13481 12449 13515
rect 12449 13481 12483 13515
rect 12483 13481 12492 13515
rect 12440 13472 12492 13481
rect 12716 13472 12768 13524
rect 17960 13472 18012 13524
rect 20720 13472 20772 13524
rect 5172 13404 5224 13456
rect 8208 13336 8260 13388
rect 9220 13379 9272 13388
rect 9220 13345 9229 13379
rect 9229 13345 9263 13379
rect 9263 13345 9272 13379
rect 9220 13336 9272 13345
rect 10784 13404 10836 13456
rect 11796 13404 11848 13456
rect 14280 13404 14332 13456
rect 12900 13379 12952 13388
rect 12900 13345 12909 13379
rect 12909 13345 12943 13379
rect 12943 13345 12952 13379
rect 12900 13336 12952 13345
rect 12992 13379 13044 13388
rect 12992 13345 13001 13379
rect 13001 13345 13035 13379
rect 13035 13345 13044 13379
rect 14648 13379 14700 13388
rect 12992 13336 13044 13345
rect 14648 13345 14657 13379
rect 14657 13345 14691 13379
rect 14691 13345 14700 13379
rect 14648 13336 14700 13345
rect 14832 13379 14884 13388
rect 14832 13345 14841 13379
rect 14841 13345 14875 13379
rect 14875 13345 14884 13379
rect 14832 13336 14884 13345
rect 18052 13404 18104 13456
rect 21088 13404 21140 13456
rect 2320 13268 2372 13320
rect 5448 13268 5500 13320
rect 8576 13311 8628 13320
rect 8576 13277 8585 13311
rect 8585 13277 8619 13311
rect 8619 13277 8628 13311
rect 8576 13268 8628 13277
rect 9404 13311 9456 13320
rect 9404 13277 9413 13311
rect 9413 13277 9447 13311
rect 9447 13277 9456 13311
rect 9404 13268 9456 13277
rect 12164 13311 12216 13320
rect 12164 13277 12173 13311
rect 12173 13277 12207 13311
rect 12207 13277 12216 13311
rect 13636 13311 13688 13320
rect 12164 13268 12216 13277
rect 6920 13200 6972 13252
rect 7196 13132 7248 13184
rect 8208 13132 8260 13184
rect 11244 13200 11296 13252
rect 13636 13277 13645 13311
rect 13645 13277 13679 13311
rect 13679 13277 13688 13311
rect 13636 13268 13688 13277
rect 14556 13268 14608 13320
rect 15016 13268 15068 13320
rect 16304 13268 16356 13320
rect 15660 13243 15712 13252
rect 15660 13209 15669 13243
rect 15669 13209 15703 13243
rect 15703 13209 15712 13243
rect 15660 13200 15712 13209
rect 17408 13243 17460 13252
rect 17408 13209 17417 13243
rect 17417 13209 17451 13243
rect 17451 13209 17460 13243
rect 17408 13200 17460 13209
rect 18696 13336 18748 13388
rect 19892 13379 19944 13388
rect 19892 13345 19901 13379
rect 19901 13345 19935 13379
rect 19935 13345 19944 13379
rect 19892 13336 19944 13345
rect 20720 13336 20772 13388
rect 18604 13311 18656 13320
rect 18604 13277 18613 13311
rect 18613 13277 18647 13311
rect 18647 13277 18656 13311
rect 18604 13268 18656 13277
rect 19064 13268 19116 13320
rect 20536 13311 20588 13320
rect 20536 13277 20545 13311
rect 20545 13277 20579 13311
rect 20579 13277 20588 13311
rect 20536 13268 20588 13277
rect 21456 13268 21508 13320
rect 12348 13132 12400 13184
rect 12808 13175 12860 13184
rect 12808 13141 12817 13175
rect 12817 13141 12851 13175
rect 12851 13141 12860 13175
rect 12808 13132 12860 13141
rect 14464 13132 14516 13184
rect 14648 13132 14700 13184
rect 14924 13132 14976 13184
rect 15936 13132 15988 13184
rect 18880 13132 18932 13184
rect 19984 13132 20036 13184
rect 20260 13132 20312 13184
rect 20628 13175 20680 13184
rect 20628 13141 20637 13175
rect 20637 13141 20671 13175
rect 20671 13141 20680 13175
rect 20996 13175 21048 13184
rect 20628 13132 20680 13141
rect 20996 13141 21005 13175
rect 21005 13141 21039 13175
rect 21039 13141 21048 13175
rect 20996 13132 21048 13141
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 7472 12928 7524 12980
rect 8116 12928 8168 12980
rect 9404 12928 9456 12980
rect 10324 12971 10376 12980
rect 10324 12937 10333 12971
rect 10333 12937 10367 12971
rect 10367 12937 10376 12971
rect 10324 12928 10376 12937
rect 12808 12928 12860 12980
rect 14556 12971 14608 12980
rect 14556 12937 14565 12971
rect 14565 12937 14599 12971
rect 14599 12937 14608 12971
rect 14556 12928 14608 12937
rect 15200 12928 15252 12980
rect 15476 12928 15528 12980
rect 15752 12928 15804 12980
rect 18696 12928 18748 12980
rect 20260 12971 20312 12980
rect 20260 12937 20269 12971
rect 20269 12937 20303 12971
rect 20303 12937 20312 12971
rect 20260 12928 20312 12937
rect 20996 12928 21048 12980
rect 21548 12928 21600 12980
rect 4988 12860 5040 12912
rect 10416 12860 10468 12912
rect 12532 12860 12584 12912
rect 12624 12860 12676 12912
rect 15108 12860 15160 12912
rect 17408 12860 17460 12912
rect 7748 12792 7800 12844
rect 8852 12792 8904 12844
rect 10232 12792 10284 12844
rect 12348 12792 12400 12844
rect 12072 12724 12124 12776
rect 12992 12767 13044 12776
rect 12992 12733 13001 12767
rect 13001 12733 13035 12767
rect 13035 12733 13044 12767
rect 12992 12724 13044 12733
rect 11980 12656 12032 12708
rect 13360 12835 13412 12844
rect 13360 12801 13369 12835
rect 13369 12801 13403 12835
rect 13403 12801 13412 12835
rect 13360 12792 13412 12801
rect 13544 12724 13596 12776
rect 14740 12724 14792 12776
rect 15016 12767 15068 12776
rect 15016 12733 15025 12767
rect 15025 12733 15059 12767
rect 15059 12733 15068 12767
rect 15016 12724 15068 12733
rect 16948 12792 17000 12844
rect 19524 12860 19576 12912
rect 16212 12767 16264 12776
rect 14556 12656 14608 12708
rect 14832 12656 14884 12708
rect 16212 12733 16221 12767
rect 16221 12733 16255 12767
rect 16255 12733 16264 12767
rect 16212 12724 16264 12733
rect 19708 12835 19760 12844
rect 19708 12801 19726 12835
rect 19726 12801 19760 12835
rect 19708 12792 19760 12801
rect 8116 12588 8168 12640
rect 11704 12588 11756 12640
rect 13360 12588 13412 12640
rect 13820 12588 13872 12640
rect 16672 12631 16724 12640
rect 16672 12597 16681 12631
rect 16681 12597 16715 12631
rect 16715 12597 16724 12631
rect 16672 12588 16724 12597
rect 18788 12724 18840 12776
rect 20536 12724 20588 12776
rect 20904 12767 20956 12776
rect 20904 12733 20913 12767
rect 20913 12733 20947 12767
rect 20947 12733 20956 12767
rect 20904 12724 20956 12733
rect 18512 12656 18564 12708
rect 18696 12656 18748 12708
rect 20628 12588 20680 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 7656 12359 7708 12368
rect 7656 12325 7665 12359
rect 7665 12325 7699 12359
rect 7699 12325 7708 12359
rect 7656 12316 7708 12325
rect 8760 12316 8812 12368
rect 9220 12384 9272 12436
rect 8392 12248 8444 12300
rect 12072 12427 12124 12436
rect 12072 12393 12081 12427
rect 12081 12393 12115 12427
rect 12115 12393 12124 12427
rect 12072 12384 12124 12393
rect 15108 12384 15160 12436
rect 17684 12427 17736 12436
rect 17684 12393 17693 12427
rect 17693 12393 17727 12427
rect 17727 12393 17736 12427
rect 17684 12384 17736 12393
rect 18604 12384 18656 12436
rect 20904 12384 20956 12436
rect 8116 12180 8168 12232
rect 8944 12180 8996 12232
rect 9036 12180 9088 12232
rect 10876 12248 10928 12300
rect 11704 12248 11756 12300
rect 10784 12223 10836 12232
rect 10784 12189 10793 12223
rect 10793 12189 10827 12223
rect 10827 12189 10836 12223
rect 10784 12180 10836 12189
rect 11796 12180 11848 12232
rect 15476 12316 15528 12368
rect 17776 12316 17828 12368
rect 16304 12291 16356 12300
rect 15200 12223 15252 12232
rect 15200 12189 15218 12223
rect 15218 12189 15252 12223
rect 15200 12180 15252 12189
rect 9864 12112 9916 12164
rect 11612 12155 11664 12164
rect 11612 12121 11621 12155
rect 11621 12121 11655 12155
rect 11655 12121 11664 12155
rect 11612 12112 11664 12121
rect 12164 12112 12216 12164
rect 12440 12112 12492 12164
rect 10508 12044 10560 12096
rect 11152 12044 11204 12096
rect 14280 12112 14332 12164
rect 13912 12044 13964 12096
rect 16304 12257 16313 12291
rect 16313 12257 16347 12291
rect 16347 12257 16356 12291
rect 16304 12248 16356 12257
rect 16672 12248 16724 12300
rect 17224 12248 17276 12300
rect 17684 12248 17736 12300
rect 18788 12248 18840 12300
rect 19524 12248 19576 12300
rect 17408 12180 17460 12232
rect 18236 12180 18288 12232
rect 19708 12180 19760 12232
rect 16120 12155 16172 12164
rect 16120 12121 16129 12155
rect 16129 12121 16163 12155
rect 16163 12121 16172 12155
rect 16120 12112 16172 12121
rect 16212 12087 16264 12096
rect 16212 12053 16221 12087
rect 16221 12053 16255 12087
rect 16255 12053 16264 12087
rect 16212 12044 16264 12053
rect 17868 12044 17920 12096
rect 20720 12112 20772 12164
rect 18144 12044 18196 12096
rect 18512 12044 18564 12096
rect 19892 12044 19944 12096
rect 20444 12044 20496 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 4896 11840 4948 11892
rect 6920 11883 6972 11892
rect 6920 11849 6929 11883
rect 6929 11849 6963 11883
rect 6963 11849 6972 11883
rect 6920 11840 6972 11849
rect 7196 11840 7248 11892
rect 8484 11840 8536 11892
rect 8944 11840 8996 11892
rect 9680 11840 9732 11892
rect 9496 11772 9548 11824
rect 11152 11772 11204 11824
rect 8024 11704 8076 11756
rect 8760 11747 8812 11756
rect 8760 11713 8769 11747
rect 8769 11713 8803 11747
rect 8803 11713 8812 11747
rect 8760 11704 8812 11713
rect 9036 11747 9088 11756
rect 9036 11713 9045 11747
rect 9045 11713 9079 11747
rect 9079 11713 9088 11747
rect 9036 11704 9088 11713
rect 11796 11840 11848 11892
rect 13820 11883 13872 11892
rect 13820 11849 13829 11883
rect 13829 11849 13863 11883
rect 13863 11849 13872 11883
rect 13820 11840 13872 11849
rect 6552 11636 6604 11688
rect 10048 11636 10100 11688
rect 14740 11772 14792 11824
rect 15844 11815 15896 11824
rect 15844 11781 15853 11815
rect 15853 11781 15887 11815
rect 15887 11781 15896 11815
rect 15844 11772 15896 11781
rect 18052 11840 18104 11892
rect 18328 11883 18380 11892
rect 18328 11849 18337 11883
rect 18337 11849 18371 11883
rect 18371 11849 18380 11883
rect 18328 11840 18380 11849
rect 18880 11840 18932 11892
rect 11980 11747 12032 11756
rect 11980 11713 12014 11747
rect 12014 11713 12032 11747
rect 17316 11772 17368 11824
rect 19616 11772 19668 11824
rect 11980 11704 12032 11713
rect 15108 11636 15160 11688
rect 18604 11704 18656 11756
rect 18972 11704 19024 11756
rect 20720 11747 20772 11756
rect 20720 11713 20729 11747
rect 20729 11713 20763 11747
rect 20763 11713 20772 11747
rect 20720 11704 20772 11713
rect 16672 11679 16724 11688
rect 16672 11645 16681 11679
rect 16681 11645 16715 11679
rect 16715 11645 16724 11679
rect 16672 11636 16724 11645
rect 17684 11636 17736 11688
rect 19800 11679 19852 11688
rect 19800 11645 19809 11679
rect 19809 11645 19843 11679
rect 19843 11645 19852 11679
rect 19800 11636 19852 11645
rect 19984 11679 20036 11688
rect 19984 11645 19993 11679
rect 19993 11645 20027 11679
rect 20027 11645 20036 11679
rect 19984 11636 20036 11645
rect 5080 11568 5132 11620
rect 7656 11568 7708 11620
rect 10324 11568 10376 11620
rect 11336 11568 11388 11620
rect 7472 11500 7524 11552
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 15660 11500 15712 11552
rect 16304 11543 16356 11552
rect 16304 11509 16313 11543
rect 16313 11509 16347 11543
rect 16347 11509 16356 11543
rect 16304 11500 16356 11509
rect 20628 11568 20680 11620
rect 16856 11500 16908 11552
rect 18052 11543 18104 11552
rect 18052 11509 18061 11543
rect 18061 11509 18095 11543
rect 18095 11509 18104 11543
rect 18052 11500 18104 11509
rect 18236 11500 18288 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 7748 11296 7800 11348
rect 8576 11339 8628 11348
rect 8576 11305 8585 11339
rect 8585 11305 8619 11339
rect 8619 11305 8628 11339
rect 8576 11296 8628 11305
rect 9220 11296 9272 11348
rect 9496 11296 9548 11348
rect 10784 11296 10836 11348
rect 1768 11228 1820 11280
rect 5724 11228 5776 11280
rect 11244 11296 11296 11348
rect 13636 11296 13688 11348
rect 14832 11339 14884 11348
rect 14832 11305 14841 11339
rect 14841 11305 14875 11339
rect 14875 11305 14884 11339
rect 14832 11296 14884 11305
rect 14924 11296 14976 11348
rect 16580 11296 16632 11348
rect 17132 11296 17184 11348
rect 18696 11296 18748 11348
rect 5540 11160 5592 11212
rect 8208 11160 8260 11212
rect 11336 11160 11388 11212
rect 13084 11160 13136 11212
rect 16304 11228 16356 11280
rect 17684 11228 17736 11280
rect 17868 11228 17920 11280
rect 17040 11203 17092 11212
rect 7656 11092 7708 11144
rect 3148 11024 3200 11076
rect 5816 11024 5868 11076
rect 9220 11024 9272 11076
rect 9404 11024 9456 11076
rect 9772 10999 9824 11008
rect 9772 10965 9781 10999
rect 9781 10965 9815 10999
rect 9815 10965 9824 10999
rect 9772 10956 9824 10965
rect 10508 11024 10560 11076
rect 11796 11092 11848 11144
rect 13728 11092 13780 11144
rect 14280 11092 14332 11144
rect 15108 11092 15160 11144
rect 17040 11169 17049 11203
rect 17049 11169 17083 11203
rect 17083 11169 17092 11203
rect 20996 11228 21048 11280
rect 21456 11228 21508 11280
rect 17040 11160 17092 11169
rect 15476 11092 15528 11144
rect 15936 11135 15988 11144
rect 15936 11101 15954 11135
rect 15954 11101 15988 11135
rect 15936 11092 15988 11101
rect 16672 11092 16724 11144
rect 18144 11092 18196 11144
rect 19248 11092 19300 11144
rect 16580 11024 16632 11076
rect 12716 10999 12768 11008
rect 12716 10965 12725 10999
rect 12725 10965 12759 10999
rect 12759 10965 12768 10999
rect 12716 10956 12768 10965
rect 12808 10999 12860 11008
rect 12808 10965 12817 10999
rect 12817 10965 12851 10999
rect 12851 10965 12860 10999
rect 12808 10956 12860 10965
rect 16396 10956 16448 11008
rect 17132 11024 17184 11076
rect 18236 11024 18288 11076
rect 18420 11024 18472 11076
rect 21640 11024 21692 11076
rect 17224 10956 17276 11008
rect 17500 10999 17552 11008
rect 17500 10965 17509 10999
rect 17509 10965 17543 10999
rect 17543 10965 17552 10999
rect 17500 10956 17552 10965
rect 17684 10956 17736 11008
rect 17960 10999 18012 11008
rect 17960 10965 17969 10999
rect 17969 10965 18003 10999
rect 18003 10965 18012 10999
rect 17960 10956 18012 10965
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 8116 10752 8168 10804
rect 9312 10684 9364 10736
rect 10048 10752 10100 10804
rect 10232 10752 10284 10804
rect 10784 10795 10836 10804
rect 10784 10761 10793 10795
rect 10793 10761 10827 10795
rect 10827 10761 10836 10795
rect 10784 10752 10836 10761
rect 12808 10752 12860 10804
rect 11796 10684 11848 10736
rect 12072 10684 12124 10736
rect 12256 10684 12308 10736
rect 15016 10752 15068 10804
rect 15292 10752 15344 10804
rect 16212 10752 16264 10804
rect 19984 10752 20036 10804
rect 14924 10684 14976 10736
rect 9312 10548 9364 10600
rect 9496 10548 9548 10600
rect 9772 10616 9824 10668
rect 11152 10616 11204 10668
rect 12348 10616 12400 10668
rect 17500 10684 17552 10736
rect 15292 10659 15344 10668
rect 15292 10625 15301 10659
rect 15301 10625 15335 10659
rect 15335 10625 15344 10659
rect 15936 10659 15988 10668
rect 15292 10616 15344 10625
rect 15936 10625 15945 10659
rect 15945 10625 15979 10659
rect 15979 10625 15988 10659
rect 17960 10684 18012 10736
rect 18052 10684 18104 10736
rect 19248 10684 19300 10736
rect 15936 10616 15988 10625
rect 18236 10616 18288 10668
rect 20260 10727 20312 10736
rect 20260 10693 20294 10727
rect 20294 10693 20312 10727
rect 20260 10684 20312 10693
rect 10140 10548 10192 10600
rect 5632 10480 5684 10532
rect 7748 10523 7800 10532
rect 7748 10489 7757 10523
rect 7757 10489 7791 10523
rect 7791 10489 7800 10523
rect 7748 10480 7800 10489
rect 8392 10480 8444 10532
rect 9128 10480 9180 10532
rect 6644 10412 6696 10464
rect 6828 10412 6880 10464
rect 10232 10412 10284 10464
rect 11060 10548 11112 10600
rect 13268 10548 13320 10600
rect 13820 10548 13872 10600
rect 15200 10548 15252 10600
rect 17040 10548 17092 10600
rect 18144 10548 18196 10600
rect 11244 10412 11296 10464
rect 12808 10480 12860 10532
rect 15568 10480 15620 10532
rect 13820 10412 13872 10464
rect 14280 10412 14332 10464
rect 16212 10412 16264 10464
rect 16672 10455 16724 10464
rect 16672 10421 16681 10455
rect 16681 10421 16715 10455
rect 16715 10421 16724 10455
rect 16672 10412 16724 10421
rect 18052 10412 18104 10464
rect 20628 10412 20680 10464
rect 20904 10412 20956 10464
rect 21180 10412 21232 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 4252 10208 4304 10260
rect 7656 10208 7708 10260
rect 7932 10208 7984 10260
rect 8392 10140 8444 10192
rect 7288 10072 7340 10124
rect 5816 10004 5868 10056
rect 6736 10004 6788 10056
rect 7472 10047 7524 10056
rect 7472 10013 7481 10047
rect 7481 10013 7515 10047
rect 7515 10013 7524 10047
rect 7472 10004 7524 10013
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 9496 10115 9548 10124
rect 9496 10081 9505 10115
rect 9505 10081 9539 10115
rect 9539 10081 9548 10115
rect 10232 10208 10284 10260
rect 10140 10183 10192 10192
rect 10140 10149 10149 10183
rect 10149 10149 10183 10183
rect 10183 10149 10192 10183
rect 10140 10140 10192 10149
rect 12072 10140 12124 10192
rect 12716 10208 12768 10260
rect 13820 10208 13872 10260
rect 15568 10208 15620 10260
rect 15936 10140 15988 10192
rect 16120 10208 16172 10260
rect 20352 10208 20404 10260
rect 20628 10251 20680 10260
rect 20628 10217 20637 10251
rect 20637 10217 20671 10251
rect 20671 10217 20680 10251
rect 20628 10208 20680 10217
rect 9496 10072 9548 10081
rect 10416 10004 10468 10056
rect 12256 10072 12308 10124
rect 13544 10072 13596 10124
rect 14556 10072 14608 10124
rect 14004 10004 14056 10056
rect 14740 10004 14792 10056
rect 17224 10072 17276 10124
rect 6644 9936 6696 9988
rect 7932 9979 7984 9988
rect 5908 9868 5960 9920
rect 6552 9868 6604 9920
rect 7656 9911 7708 9920
rect 7656 9877 7665 9911
rect 7665 9877 7699 9911
rect 7699 9877 7708 9911
rect 7656 9868 7708 9877
rect 7932 9945 7941 9979
rect 7941 9945 7975 9979
rect 7975 9945 7984 9979
rect 7932 9936 7984 9945
rect 8392 9936 8444 9988
rect 10324 9936 10376 9988
rect 11060 9936 11112 9988
rect 11704 9936 11756 9988
rect 12164 9936 12216 9988
rect 12992 9911 13044 9920
rect 12992 9877 13001 9911
rect 13001 9877 13035 9911
rect 13035 9877 13044 9911
rect 12992 9868 13044 9877
rect 14280 9868 14332 9920
rect 14464 9911 14516 9920
rect 14464 9877 14473 9911
rect 14473 9877 14507 9911
rect 14507 9877 14516 9911
rect 14464 9868 14516 9877
rect 14556 9911 14608 9920
rect 14556 9877 14565 9911
rect 14565 9877 14599 9911
rect 14599 9877 14608 9911
rect 14556 9868 14608 9877
rect 15200 9868 15252 9920
rect 16672 10004 16724 10056
rect 17684 10004 17736 10056
rect 18144 10004 18196 10056
rect 18604 10047 18656 10056
rect 18604 10013 18613 10047
rect 18613 10013 18647 10047
rect 18647 10013 18656 10047
rect 18604 10004 18656 10013
rect 19340 10004 19392 10056
rect 20720 10004 20772 10056
rect 20168 9936 20220 9988
rect 15844 9868 15896 9920
rect 17868 9868 17920 9920
rect 19892 9868 19944 9920
rect 20812 9868 20864 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 7472 9707 7524 9716
rect 7472 9673 7481 9707
rect 7481 9673 7515 9707
rect 7515 9673 7524 9707
rect 7472 9664 7524 9673
rect 7656 9664 7708 9716
rect 12072 9664 12124 9716
rect 12992 9664 13044 9716
rect 14556 9664 14608 9716
rect 15108 9664 15160 9716
rect 1860 9596 1912 9648
rect 6828 9596 6880 9648
rect 7288 9596 7340 9648
rect 8300 9596 8352 9648
rect 8668 9639 8720 9648
rect 8668 9605 8677 9639
rect 8677 9605 8711 9639
rect 8711 9605 8720 9639
rect 8668 9596 8720 9605
rect 9128 9596 9180 9648
rect 7104 9571 7156 9580
rect 7104 9537 7113 9571
rect 7113 9537 7147 9571
rect 7147 9537 7156 9571
rect 7104 9528 7156 9537
rect 8392 9571 8444 9580
rect 8392 9537 8401 9571
rect 8401 9537 8435 9571
rect 8435 9537 8444 9571
rect 8392 9528 8444 9537
rect 9496 9596 9548 9648
rect 11704 9596 11756 9648
rect 11980 9596 12032 9648
rect 12440 9639 12492 9648
rect 12440 9605 12449 9639
rect 12449 9605 12483 9639
rect 12483 9605 12492 9639
rect 12440 9596 12492 9605
rect 14372 9596 14424 9648
rect 15844 9664 15896 9716
rect 16212 9664 16264 9716
rect 20904 9664 20956 9716
rect 16120 9596 16172 9648
rect 5724 9324 5776 9376
rect 6828 9324 6880 9376
rect 9864 9528 9916 9580
rect 11244 9528 11296 9580
rect 12256 9528 12308 9580
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 11060 9460 11112 9512
rect 11612 9460 11664 9512
rect 14280 9528 14332 9580
rect 15936 9528 15988 9580
rect 13636 9460 13688 9512
rect 14004 9503 14056 9512
rect 14004 9469 14013 9503
rect 14013 9469 14047 9503
rect 14047 9469 14056 9503
rect 14004 9460 14056 9469
rect 14832 9503 14884 9512
rect 14832 9469 14841 9503
rect 14841 9469 14875 9503
rect 14875 9469 14884 9503
rect 14832 9460 14884 9469
rect 9588 9367 9640 9376
rect 9588 9333 9597 9367
rect 9597 9333 9631 9367
rect 9631 9333 9640 9367
rect 9588 9324 9640 9333
rect 10232 9324 10284 9376
rect 13544 9392 13596 9444
rect 15292 9460 15344 9512
rect 15752 9460 15804 9512
rect 16120 9503 16172 9512
rect 16120 9469 16129 9503
rect 16129 9469 16163 9503
rect 16163 9469 16172 9503
rect 16120 9460 16172 9469
rect 16396 9528 16448 9580
rect 16856 9596 16908 9648
rect 17960 9596 18012 9648
rect 16948 9528 17000 9580
rect 17040 9528 17092 9580
rect 18696 9528 18748 9580
rect 20168 9571 20220 9580
rect 20168 9537 20177 9571
rect 20177 9537 20211 9571
rect 20211 9537 20220 9571
rect 20168 9528 20220 9537
rect 21088 9571 21140 9580
rect 21088 9537 21097 9571
rect 21097 9537 21131 9571
rect 21131 9537 21140 9571
rect 21088 9528 21140 9537
rect 18144 9503 18196 9512
rect 13452 9324 13504 9376
rect 13820 9324 13872 9376
rect 14740 9324 14792 9376
rect 15292 9324 15344 9376
rect 15844 9324 15896 9376
rect 16580 9324 16632 9376
rect 16672 9324 16724 9376
rect 16948 9324 17000 9376
rect 18144 9469 18153 9503
rect 18153 9469 18187 9503
rect 18187 9469 18196 9503
rect 18144 9460 18196 9469
rect 20260 9503 20312 9512
rect 20260 9469 20269 9503
rect 20269 9469 20303 9503
rect 20303 9469 20312 9503
rect 20260 9460 20312 9469
rect 20352 9460 20404 9512
rect 20628 9460 20680 9512
rect 19524 9435 19576 9444
rect 19524 9401 19533 9435
rect 19533 9401 19567 9435
rect 19567 9401 19576 9435
rect 19524 9392 19576 9401
rect 19800 9435 19852 9444
rect 19800 9401 19809 9435
rect 19809 9401 19843 9435
rect 19843 9401 19852 9435
rect 19800 9392 19852 9401
rect 17408 9324 17460 9376
rect 20352 9324 20404 9376
rect 20628 9324 20680 9376
rect 21272 9367 21324 9376
rect 21272 9333 21281 9367
rect 21281 9333 21315 9367
rect 21315 9333 21324 9367
rect 21272 9324 21324 9333
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 10232 9120 10284 9172
rect 10416 9163 10468 9172
rect 10416 9129 10425 9163
rect 10425 9129 10459 9163
rect 10459 9129 10468 9163
rect 10416 9120 10468 9129
rect 14372 9120 14424 9172
rect 7288 9095 7340 9104
rect 7288 9061 7297 9095
rect 7297 9061 7331 9095
rect 7331 9061 7340 9095
rect 7288 9052 7340 9061
rect 11612 9052 11664 9104
rect 13544 9052 13596 9104
rect 14464 9052 14516 9104
rect 6920 9027 6972 9036
rect 6920 8993 6929 9027
rect 6929 8993 6963 9027
rect 6963 8993 6972 9027
rect 6920 8984 6972 8993
rect 7104 8984 7156 9036
rect 6828 8916 6880 8968
rect 8484 8984 8536 9036
rect 9496 9027 9548 9036
rect 9496 8993 9505 9027
rect 9505 8993 9539 9027
rect 9539 8993 9548 9027
rect 9496 8984 9548 8993
rect 9588 8984 9640 9036
rect 11060 8984 11112 9036
rect 12164 9027 12216 9036
rect 12164 8993 12173 9027
rect 12173 8993 12207 9027
rect 12207 8993 12216 9027
rect 12164 8984 12216 8993
rect 13728 8984 13780 9036
rect 15384 9120 15436 9172
rect 15936 9120 15988 9172
rect 16580 9120 16632 9172
rect 17224 9120 17276 9172
rect 17408 9120 17460 9172
rect 17132 9052 17184 9104
rect 16304 8984 16356 9036
rect 16580 9027 16632 9036
rect 16580 8993 16589 9027
rect 16589 8993 16623 9027
rect 16623 8993 16632 9027
rect 16580 8984 16632 8993
rect 17500 8984 17552 9036
rect 8024 8916 8076 8968
rect 6552 8891 6604 8900
rect 6552 8857 6561 8891
rect 6561 8857 6595 8891
rect 6595 8857 6604 8891
rect 6552 8848 6604 8857
rect 10692 8916 10744 8968
rect 14280 8916 14332 8968
rect 7564 8823 7616 8832
rect 7564 8789 7573 8823
rect 7573 8789 7607 8823
rect 7607 8789 7616 8823
rect 7564 8780 7616 8789
rect 8576 8823 8628 8832
rect 8576 8789 8585 8823
rect 8585 8789 8619 8823
rect 8619 8789 8628 8823
rect 8576 8780 8628 8789
rect 13084 8848 13136 8900
rect 11152 8780 11204 8832
rect 12348 8780 12400 8832
rect 13452 8780 13504 8832
rect 14372 8823 14424 8832
rect 14372 8789 14381 8823
rect 14381 8789 14415 8823
rect 14415 8789 14424 8823
rect 14372 8780 14424 8789
rect 14464 8780 14516 8832
rect 15936 8916 15988 8968
rect 16120 8916 16172 8968
rect 16672 8916 16724 8968
rect 16948 8916 17000 8968
rect 17316 8916 17368 8968
rect 15844 8780 15896 8832
rect 16028 8780 16080 8832
rect 16856 8848 16908 8900
rect 17224 8848 17276 8900
rect 18052 9120 18104 9172
rect 18512 9120 18564 9172
rect 20260 9163 20312 9172
rect 20260 9129 20269 9163
rect 20269 9129 20303 9163
rect 20303 9129 20312 9163
rect 20260 9120 20312 9129
rect 20352 9120 20404 9172
rect 19156 9052 19208 9104
rect 19432 9052 19484 9104
rect 19524 9052 19576 9104
rect 18236 9027 18288 9036
rect 18236 8993 18245 9027
rect 18245 8993 18279 9027
rect 18279 8993 18288 9027
rect 18236 8984 18288 8993
rect 17868 8916 17920 8968
rect 19432 8916 19484 8968
rect 20168 8916 20220 8968
rect 18328 8891 18380 8900
rect 18328 8857 18337 8891
rect 18337 8857 18371 8891
rect 18371 8857 18380 8891
rect 18328 8848 18380 8857
rect 18696 8848 18748 8900
rect 18972 8848 19024 8900
rect 21364 8848 21416 8900
rect 18788 8823 18840 8832
rect 18788 8789 18797 8823
rect 18797 8789 18831 8823
rect 18831 8789 18840 8823
rect 18788 8780 18840 8789
rect 18880 8780 18932 8832
rect 19616 8823 19668 8832
rect 19616 8789 19625 8823
rect 19625 8789 19659 8823
rect 19659 8789 19668 8823
rect 19616 8780 19668 8789
rect 19800 8780 19852 8832
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 8024 8576 8076 8628
rect 8116 8483 8168 8492
rect 8116 8449 8125 8483
rect 8125 8449 8159 8483
rect 8159 8449 8168 8483
rect 8116 8440 8168 8449
rect 3332 8372 3384 8424
rect 7748 8415 7800 8424
rect 7748 8381 7757 8415
rect 7757 8381 7791 8415
rect 7791 8381 7800 8415
rect 7748 8372 7800 8381
rect 16028 8576 16080 8628
rect 17040 8619 17092 8628
rect 17040 8585 17049 8619
rect 17049 8585 17083 8619
rect 17083 8585 17092 8619
rect 17040 8576 17092 8585
rect 17224 8576 17276 8628
rect 18788 8576 18840 8628
rect 21088 8576 21140 8628
rect 8576 8508 8628 8560
rect 18144 8508 18196 8560
rect 10324 8440 10376 8492
rect 10600 8483 10652 8492
rect 10600 8449 10618 8483
rect 10618 8449 10652 8483
rect 10600 8440 10652 8449
rect 9864 8372 9916 8424
rect 11060 8372 11112 8424
rect 7840 8304 7892 8356
rect 9496 8347 9548 8356
rect 9496 8313 9505 8347
rect 9505 8313 9539 8347
rect 9539 8313 9548 8347
rect 9496 8304 9548 8313
rect 10968 8304 11020 8356
rect 11980 8440 12032 8492
rect 12164 8440 12216 8492
rect 12624 8440 12676 8492
rect 13544 8440 13596 8492
rect 14372 8483 14424 8492
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 12072 8372 12124 8424
rect 15936 8440 15988 8492
rect 16672 8440 16724 8492
rect 17132 8440 17184 8492
rect 14924 8415 14976 8424
rect 11888 8304 11940 8356
rect 14924 8381 14933 8415
rect 14933 8381 14967 8415
rect 14967 8381 14976 8415
rect 14924 8372 14976 8381
rect 16120 8372 16172 8424
rect 18880 8440 18932 8492
rect 18972 8440 19024 8492
rect 20720 8508 20772 8560
rect 7288 8236 7340 8288
rect 9588 8236 9640 8288
rect 13728 8304 13780 8356
rect 14004 8304 14056 8356
rect 15936 8304 15988 8356
rect 17500 8304 17552 8356
rect 17684 8304 17736 8356
rect 16120 8236 16172 8288
rect 19156 8304 19208 8356
rect 18420 8236 18472 8288
rect 18880 8236 18932 8288
rect 18972 8236 19024 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 7012 8032 7064 8084
rect 9588 8032 9640 8084
rect 9772 8032 9824 8084
rect 13636 8075 13688 8084
rect 9956 7964 10008 8016
rect 10508 7964 10560 8016
rect 10600 7964 10652 8016
rect 13636 8041 13645 8075
rect 13645 8041 13679 8075
rect 13679 8041 13688 8075
rect 13636 8032 13688 8041
rect 14832 8075 14884 8084
rect 14832 8041 14841 8075
rect 14841 8041 14875 8075
rect 14875 8041 14884 8075
rect 14832 8032 14884 8041
rect 15384 8032 15436 8084
rect 16120 8032 16172 8084
rect 16672 8032 16724 8084
rect 18144 8032 18196 8084
rect 19984 8032 20036 8084
rect 20628 8032 20680 8084
rect 8484 7896 8536 7948
rect 14740 7964 14792 8016
rect 18512 7964 18564 8016
rect 18972 7964 19024 8016
rect 19524 7964 19576 8016
rect 6552 7871 6604 7880
rect 6552 7837 6561 7871
rect 6561 7837 6595 7871
rect 6595 7837 6604 7871
rect 6552 7828 6604 7837
rect 7564 7871 7616 7880
rect 7564 7837 7573 7871
rect 7573 7837 7607 7871
rect 7607 7837 7616 7871
rect 7564 7828 7616 7837
rect 12716 7828 12768 7880
rect 13084 7896 13136 7948
rect 14464 7896 14516 7948
rect 17960 7896 18012 7948
rect 18420 7896 18472 7948
rect 15108 7871 15160 7880
rect 15108 7837 15117 7871
rect 15117 7837 15151 7871
rect 15151 7837 15160 7871
rect 15108 7828 15160 7837
rect 15292 7828 15344 7880
rect 7840 7760 7892 7812
rect 8944 7760 8996 7812
rect 11060 7760 11112 7812
rect 12164 7803 12216 7812
rect 12164 7769 12173 7803
rect 12173 7769 12207 7803
rect 12207 7769 12216 7803
rect 12164 7760 12216 7769
rect 12808 7803 12860 7812
rect 12808 7769 12817 7803
rect 12817 7769 12851 7803
rect 12851 7769 12860 7803
rect 12808 7760 12860 7769
rect 13728 7760 13780 7812
rect 14188 7760 14240 7812
rect 15200 7760 15252 7812
rect 15660 7803 15712 7812
rect 15660 7769 15669 7803
rect 15669 7769 15703 7803
rect 15703 7769 15712 7803
rect 15660 7760 15712 7769
rect 17776 7828 17828 7880
rect 19524 7828 19576 7880
rect 19708 7828 19760 7880
rect 20168 7760 20220 7812
rect 7104 7692 7156 7744
rect 8208 7735 8260 7744
rect 8208 7701 8217 7735
rect 8217 7701 8251 7735
rect 8251 7701 8260 7735
rect 8208 7692 8260 7701
rect 10140 7692 10192 7744
rect 12532 7692 12584 7744
rect 12992 7692 13044 7744
rect 16396 7692 16448 7744
rect 17040 7692 17092 7744
rect 18052 7735 18104 7744
rect 18052 7701 18061 7735
rect 18061 7701 18095 7735
rect 18095 7701 18104 7735
rect 18052 7692 18104 7701
rect 18788 7692 18840 7744
rect 20720 7692 20772 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 5448 7488 5500 7540
rect 7748 7488 7800 7540
rect 8208 7420 8260 7472
rect 10600 7488 10652 7540
rect 10692 7531 10744 7540
rect 10692 7497 10701 7531
rect 10701 7497 10735 7531
rect 10735 7497 10744 7531
rect 10692 7488 10744 7497
rect 11244 7488 11296 7540
rect 12624 7488 12676 7540
rect 13636 7488 13688 7540
rect 15016 7488 15068 7540
rect 16212 7488 16264 7540
rect 18420 7488 18472 7540
rect 18788 7531 18840 7540
rect 18788 7497 18797 7531
rect 18797 7497 18831 7531
rect 18831 7497 18840 7531
rect 18788 7488 18840 7497
rect 19064 7488 19116 7540
rect 20168 7531 20220 7540
rect 20168 7497 20177 7531
rect 20177 7497 20211 7531
rect 20211 7497 20220 7531
rect 20168 7488 20220 7497
rect 14648 7420 14700 7472
rect 14924 7420 14976 7472
rect 8392 7395 8444 7404
rect 8392 7361 8410 7395
rect 8410 7361 8444 7395
rect 8392 7352 8444 7361
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 12348 7352 12400 7404
rect 15108 7352 15160 7404
rect 16212 7352 16264 7404
rect 16948 7352 17000 7404
rect 18696 7420 18748 7472
rect 20996 7420 21048 7472
rect 22008 7420 22060 7472
rect 12900 7327 12952 7336
rect 12900 7293 12909 7327
rect 12909 7293 12943 7327
rect 12943 7293 12952 7327
rect 12900 7284 12952 7293
rect 14188 7327 14240 7336
rect 4896 7216 4948 7268
rect 7380 7216 7432 7268
rect 11336 7216 11388 7268
rect 14188 7293 14197 7327
rect 14197 7293 14231 7327
rect 14231 7293 14240 7327
rect 14188 7284 14240 7293
rect 14832 7284 14884 7336
rect 19156 7395 19208 7404
rect 19156 7361 19165 7395
rect 19165 7361 19199 7395
rect 19199 7361 19208 7395
rect 19156 7352 19208 7361
rect 5264 7191 5316 7200
rect 5264 7157 5273 7191
rect 5273 7157 5307 7191
rect 5307 7157 5316 7191
rect 5264 7148 5316 7157
rect 5356 7148 5408 7200
rect 5908 7191 5960 7200
rect 5908 7157 5917 7191
rect 5917 7157 5951 7191
rect 5951 7157 5960 7191
rect 5908 7148 5960 7157
rect 7564 7148 7616 7200
rect 9680 7148 9732 7200
rect 11060 7148 11112 7200
rect 12348 7148 12400 7200
rect 12440 7191 12492 7200
rect 12440 7157 12449 7191
rect 12449 7157 12483 7191
rect 12483 7157 12492 7191
rect 12440 7148 12492 7157
rect 12716 7148 12768 7200
rect 13360 7148 13412 7200
rect 18512 7216 18564 7268
rect 21548 7216 21600 7268
rect 22284 7216 22336 7268
rect 16580 7148 16632 7200
rect 17592 7148 17644 7200
rect 18328 7148 18380 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 12348 6944 12400 6996
rect 12900 6944 12952 6996
rect 8576 6919 8628 6928
rect 8576 6885 8585 6919
rect 8585 6885 8619 6919
rect 8619 6885 8628 6919
rect 8576 6876 8628 6885
rect 10968 6876 11020 6928
rect 11336 6919 11388 6928
rect 11336 6885 11345 6919
rect 11345 6885 11379 6919
rect 11379 6885 11388 6919
rect 11336 6876 11388 6885
rect 15108 6944 15160 6996
rect 4804 6851 4856 6860
rect 1952 6740 2004 6792
rect 4804 6817 4813 6851
rect 4813 6817 4847 6851
rect 4847 6817 4856 6851
rect 4804 6808 4856 6817
rect 4988 6808 5040 6860
rect 6736 6808 6788 6860
rect 6920 6851 6972 6860
rect 6920 6817 6929 6851
rect 6929 6817 6963 6851
rect 6963 6817 6972 6851
rect 6920 6808 6972 6817
rect 8392 6808 8444 6860
rect 9128 6808 9180 6860
rect 9680 6808 9732 6860
rect 13084 6808 13136 6860
rect 3056 6740 3108 6792
rect 7472 6740 7524 6792
rect 6552 6672 6604 6724
rect 6920 6672 6972 6724
rect 7288 6672 7340 6724
rect 1308 6604 1360 6656
rect 4160 6647 4212 6656
rect 4160 6613 4169 6647
rect 4169 6613 4203 6647
rect 4203 6613 4212 6647
rect 4160 6604 4212 6613
rect 4252 6604 4304 6656
rect 5264 6604 5316 6656
rect 5816 6604 5868 6656
rect 6736 6604 6788 6656
rect 8116 6647 8168 6656
rect 8116 6613 8125 6647
rect 8125 6613 8159 6647
rect 8159 6613 8168 6647
rect 8116 6604 8168 6613
rect 8208 6647 8260 6656
rect 8208 6613 8217 6647
rect 8217 6613 8251 6647
rect 8251 6613 8260 6647
rect 8576 6740 8628 6792
rect 13360 6783 13412 6792
rect 13360 6749 13369 6783
rect 13369 6749 13403 6783
rect 13403 6749 13412 6783
rect 13360 6740 13412 6749
rect 14648 6808 14700 6860
rect 14832 6808 14884 6860
rect 16580 6876 16632 6928
rect 17592 6919 17644 6928
rect 17040 6851 17092 6860
rect 17040 6817 17049 6851
rect 17049 6817 17083 6851
rect 17083 6817 17092 6851
rect 17040 6808 17092 6817
rect 17592 6885 17601 6919
rect 17601 6885 17635 6919
rect 17635 6885 17644 6919
rect 17592 6876 17644 6885
rect 17960 6808 18012 6860
rect 18880 6808 18932 6860
rect 9956 6672 10008 6724
rect 8208 6604 8260 6613
rect 8576 6604 8628 6656
rect 9680 6647 9732 6656
rect 9680 6613 9689 6647
rect 9689 6613 9723 6647
rect 9723 6613 9732 6647
rect 11980 6672 12032 6724
rect 12256 6672 12308 6724
rect 12348 6672 12400 6724
rect 13084 6672 13136 6724
rect 13176 6672 13228 6724
rect 15200 6672 15252 6724
rect 9680 6604 9732 6613
rect 10324 6647 10376 6656
rect 10324 6613 10333 6647
rect 10333 6613 10367 6647
rect 10367 6613 10376 6647
rect 10324 6604 10376 6613
rect 10968 6604 11020 6656
rect 14740 6604 14792 6656
rect 15016 6604 15068 6656
rect 17224 6672 17276 6724
rect 18604 6783 18656 6792
rect 18604 6749 18613 6783
rect 18613 6749 18647 6783
rect 18647 6749 18656 6783
rect 18604 6740 18656 6749
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 17500 6604 17552 6656
rect 17684 6604 17736 6656
rect 20168 6672 20220 6724
rect 18144 6604 18196 6656
rect 18972 6604 19024 6656
rect 20628 6604 20680 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 2780 6400 2832 6452
rect 3148 6443 3200 6452
rect 3148 6409 3157 6443
rect 3157 6409 3191 6443
rect 3191 6409 3200 6443
rect 3148 6400 3200 6409
rect 3884 6443 3936 6452
rect 3884 6409 3893 6443
rect 3893 6409 3927 6443
rect 3927 6409 3936 6443
rect 3884 6400 3936 6409
rect 5080 6400 5132 6452
rect 6736 6400 6788 6452
rect 8208 6400 8260 6452
rect 9128 6443 9180 6452
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 9680 6400 9732 6452
rect 10416 6400 10468 6452
rect 11152 6400 11204 6452
rect 11888 6443 11940 6452
rect 11888 6409 11897 6443
rect 11897 6409 11931 6443
rect 11931 6409 11940 6443
rect 11888 6400 11940 6409
rect 12532 6400 12584 6452
rect 13084 6443 13136 6452
rect 13084 6409 13093 6443
rect 13093 6409 13127 6443
rect 13127 6409 13136 6443
rect 13084 6400 13136 6409
rect 13636 6400 13688 6452
rect 14372 6400 14424 6452
rect 14740 6400 14792 6452
rect 17960 6400 18012 6452
rect 20536 6443 20588 6452
rect 20536 6409 20545 6443
rect 20545 6409 20579 6443
rect 20579 6409 20588 6443
rect 20536 6400 20588 6409
rect 20904 6443 20956 6452
rect 20904 6409 20913 6443
rect 20913 6409 20947 6443
rect 20947 6409 20956 6443
rect 20904 6400 20956 6409
rect 5540 6332 5592 6384
rect 8024 6375 8076 6384
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 8024 6341 8058 6375
rect 8058 6341 8076 6375
rect 8024 6332 8076 6341
rect 8576 6332 8628 6384
rect 11060 6332 11112 6384
rect 13360 6332 13412 6384
rect 14648 6332 14700 6384
rect 6552 6239 6604 6248
rect 6552 6205 6561 6239
rect 6561 6205 6595 6239
rect 6595 6205 6604 6239
rect 6552 6196 6604 6205
rect 11244 6264 11296 6316
rect 12624 6264 12676 6316
rect 14832 6332 14884 6384
rect 14924 6307 14976 6316
rect 14924 6273 14933 6307
rect 14933 6273 14967 6307
rect 14967 6273 14976 6307
rect 14924 6264 14976 6273
rect 15200 6307 15252 6316
rect 15200 6273 15234 6307
rect 15234 6273 15252 6307
rect 15200 6264 15252 6273
rect 16948 6264 17000 6316
rect 17132 6307 17184 6316
rect 17132 6273 17141 6307
rect 17141 6273 17175 6307
rect 17175 6273 17184 6307
rect 17132 6264 17184 6273
rect 17776 6264 17828 6316
rect 19432 6332 19484 6384
rect 19064 6307 19116 6316
rect 19064 6273 19098 6307
rect 19098 6273 19116 6307
rect 19064 6264 19116 6273
rect 6736 6128 6788 6180
rect 10600 6196 10652 6248
rect 10784 6239 10836 6248
rect 10784 6205 10793 6239
rect 10793 6205 10827 6239
rect 10827 6205 10836 6239
rect 10784 6196 10836 6205
rect 10876 6239 10928 6248
rect 10876 6205 10885 6239
rect 10885 6205 10919 6239
rect 10919 6205 10928 6239
rect 10876 6196 10928 6205
rect 11704 6196 11756 6248
rect 14464 6239 14516 6248
rect 14464 6205 14473 6239
rect 14473 6205 14507 6239
rect 14507 6205 14516 6239
rect 14464 6196 14516 6205
rect 20628 6196 20680 6248
rect 21180 6239 21232 6248
rect 21180 6205 21189 6239
rect 21189 6205 21223 6239
rect 21223 6205 21232 6239
rect 21180 6196 21232 6205
rect 1584 6103 1636 6112
rect 1584 6069 1593 6103
rect 1593 6069 1627 6103
rect 1627 6069 1636 6103
rect 1584 6060 1636 6069
rect 1676 6060 1728 6112
rect 3424 6103 3476 6112
rect 3424 6069 3433 6103
rect 3433 6069 3467 6103
rect 3467 6069 3476 6103
rect 3424 6060 3476 6069
rect 4896 6103 4948 6112
rect 4896 6069 4905 6103
rect 4905 6069 4939 6103
rect 4939 6069 4948 6103
rect 4896 6060 4948 6069
rect 6552 6060 6604 6112
rect 7472 6103 7524 6112
rect 7472 6069 7481 6103
rect 7481 6069 7515 6103
rect 7515 6069 7524 6103
rect 7472 6060 7524 6069
rect 10508 6128 10560 6180
rect 8668 6060 8720 6112
rect 10968 6060 11020 6112
rect 13452 6060 13504 6112
rect 16948 6128 17000 6180
rect 18512 6103 18564 6112
rect 18512 6069 18521 6103
rect 18521 6069 18555 6103
rect 18555 6069 18564 6103
rect 18512 6060 18564 6069
rect 19524 6060 19576 6112
rect 20168 6103 20220 6112
rect 20168 6069 20177 6103
rect 20177 6069 20211 6103
rect 20211 6069 20220 6103
rect 20168 6060 20220 6069
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 4252 5856 4304 5908
rect 6644 5856 6696 5908
rect 7472 5856 7524 5908
rect 2412 5788 2464 5840
rect 5816 5788 5868 5840
rect 8116 5856 8168 5908
rect 8300 5788 8352 5840
rect 8668 5788 8720 5840
rect 10600 5856 10652 5908
rect 10784 5856 10836 5908
rect 14280 5856 14332 5908
rect 14648 5856 14700 5908
rect 15752 5856 15804 5908
rect 17132 5899 17184 5908
rect 17132 5865 17141 5899
rect 17141 5865 17175 5899
rect 17175 5865 17184 5899
rect 17132 5856 17184 5865
rect 17500 5856 17552 5908
rect 9772 5788 9824 5840
rect 1584 5720 1636 5772
rect 6736 5763 6788 5772
rect 4436 5695 4488 5704
rect 4436 5661 4445 5695
rect 4445 5661 4479 5695
rect 4479 5661 4488 5695
rect 4436 5652 4488 5661
rect 5540 5695 5592 5704
rect 5540 5661 5549 5695
rect 5549 5661 5583 5695
rect 5583 5661 5592 5695
rect 5540 5652 5592 5661
rect 5908 5652 5960 5704
rect 6736 5729 6745 5763
rect 6745 5729 6779 5763
rect 6779 5729 6788 5763
rect 6736 5720 6788 5729
rect 8024 5720 8076 5772
rect 4344 5584 4396 5636
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 1952 5559 2004 5568
rect 1952 5525 1961 5559
rect 1961 5525 1995 5559
rect 1995 5525 2004 5559
rect 1952 5516 2004 5525
rect 2504 5516 2556 5568
rect 2688 5559 2740 5568
rect 2688 5525 2697 5559
rect 2697 5525 2731 5559
rect 2731 5525 2740 5559
rect 2688 5516 2740 5525
rect 4068 5516 4120 5568
rect 4252 5516 4304 5568
rect 4988 5516 5040 5568
rect 6000 5516 6052 5568
rect 6460 5584 6512 5636
rect 7380 5516 7432 5568
rect 7932 5516 7984 5568
rect 10876 5720 10928 5772
rect 12716 5763 12768 5772
rect 8576 5652 8628 5704
rect 9128 5584 9180 5636
rect 9496 5627 9548 5636
rect 9496 5593 9505 5627
rect 9505 5593 9539 5627
rect 9539 5593 9548 5627
rect 9496 5584 9548 5593
rect 8576 5559 8628 5568
rect 8576 5525 8585 5559
rect 8585 5525 8619 5559
rect 8619 5525 8628 5559
rect 8576 5516 8628 5525
rect 10324 5652 10376 5704
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 12716 5729 12725 5763
rect 12725 5729 12759 5763
rect 12759 5729 12768 5763
rect 12716 5720 12768 5729
rect 13176 5788 13228 5840
rect 19064 5856 19116 5908
rect 12992 5720 13044 5772
rect 14372 5763 14424 5772
rect 13728 5695 13780 5704
rect 13728 5661 13737 5695
rect 13737 5661 13771 5695
rect 13771 5661 13780 5695
rect 13728 5652 13780 5661
rect 14372 5729 14381 5763
rect 14381 5729 14415 5763
rect 14415 5729 14424 5763
rect 14372 5720 14424 5729
rect 18328 5763 18380 5772
rect 18328 5729 18337 5763
rect 18337 5729 18371 5763
rect 18371 5729 18380 5763
rect 18328 5720 18380 5729
rect 18420 5763 18472 5772
rect 18420 5729 18429 5763
rect 18429 5729 18463 5763
rect 18463 5729 18472 5763
rect 18420 5720 18472 5729
rect 18880 5720 18932 5772
rect 17132 5652 17184 5704
rect 18972 5652 19024 5704
rect 20996 5652 21048 5704
rect 21824 5652 21876 5704
rect 10600 5584 10652 5636
rect 11244 5584 11296 5636
rect 15660 5627 15712 5636
rect 15660 5593 15669 5627
rect 15669 5593 15703 5627
rect 15703 5593 15712 5627
rect 15660 5584 15712 5593
rect 19340 5584 19392 5636
rect 12256 5516 12308 5568
rect 12808 5516 12860 5568
rect 12992 5516 13044 5568
rect 14280 5516 14332 5568
rect 14556 5516 14608 5568
rect 15016 5559 15068 5568
rect 15016 5525 15025 5559
rect 15025 5525 15059 5559
rect 15059 5525 15068 5559
rect 15016 5516 15068 5525
rect 18236 5559 18288 5568
rect 18236 5525 18245 5559
rect 18245 5525 18279 5559
rect 18279 5525 18288 5559
rect 18236 5516 18288 5525
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 1860 5355 1912 5364
rect 1860 5321 1869 5355
rect 1869 5321 1903 5355
rect 1903 5321 1912 5355
rect 1860 5312 1912 5321
rect 7656 5355 7708 5364
rect 5448 5244 5500 5296
rect 6092 5244 6144 5296
rect 6828 5244 6880 5296
rect 7656 5321 7665 5355
rect 7665 5321 7699 5355
rect 7699 5321 7708 5355
rect 7656 5312 7708 5321
rect 8392 5355 8444 5364
rect 8392 5321 8401 5355
rect 8401 5321 8435 5355
rect 8435 5321 8444 5355
rect 8392 5312 8444 5321
rect 4620 5176 4672 5228
rect 5724 5176 5776 5228
rect 6460 5176 6512 5228
rect 6644 5176 6696 5228
rect 7012 5219 7064 5228
rect 7012 5185 7021 5219
rect 7021 5185 7055 5219
rect 7055 5185 7064 5219
rect 7012 5176 7064 5185
rect 7380 5176 7432 5228
rect 8024 5176 8076 5228
rect 14372 5312 14424 5364
rect 9312 5287 9364 5296
rect 9312 5253 9321 5287
rect 9321 5253 9355 5287
rect 9355 5253 9364 5287
rect 9312 5244 9364 5253
rect 10692 5287 10744 5296
rect 10692 5253 10701 5287
rect 10701 5253 10735 5287
rect 10735 5253 10744 5287
rect 10692 5244 10744 5253
rect 10508 5176 10560 5228
rect 10600 5219 10652 5228
rect 10600 5185 10609 5219
rect 10609 5185 10643 5219
rect 10643 5185 10652 5219
rect 10600 5176 10652 5185
rect 11244 5176 11296 5228
rect 12348 5244 12400 5296
rect 3240 5108 3292 5160
rect 5816 5108 5868 5160
rect 6000 5040 6052 5092
rect 9772 5108 9824 5160
rect 10876 5151 10928 5160
rect 10876 5117 10885 5151
rect 10885 5117 10919 5151
rect 10919 5117 10928 5151
rect 10876 5108 10928 5117
rect 10968 5108 11020 5160
rect 13636 5244 13688 5296
rect 14464 5244 14516 5296
rect 15200 5244 15252 5296
rect 13728 5176 13780 5228
rect 16580 5244 16632 5296
rect 17040 5176 17092 5228
rect 9956 5040 10008 5092
rect 2228 5015 2280 5024
rect 2228 4981 2237 5015
rect 2237 4981 2271 5015
rect 2271 4981 2280 5015
rect 2228 4972 2280 4981
rect 4712 4972 4764 5024
rect 4896 4972 4948 5024
rect 5540 4972 5592 5024
rect 7748 4972 7800 5024
rect 8116 5015 8168 5024
rect 8116 4981 8125 5015
rect 8125 4981 8159 5015
rect 8159 4981 8168 5015
rect 8116 4972 8168 4981
rect 9496 4972 9548 5024
rect 14464 5108 14516 5160
rect 18052 5312 18104 5364
rect 19616 5312 19668 5364
rect 20628 5355 20680 5364
rect 20628 5321 20637 5355
rect 20637 5321 20671 5355
rect 20671 5321 20680 5355
rect 20628 5312 20680 5321
rect 18512 5244 18564 5296
rect 18604 5219 18656 5228
rect 18604 5185 18613 5219
rect 18613 5185 18647 5219
rect 18647 5185 18656 5219
rect 18604 5176 18656 5185
rect 19892 5151 19944 5160
rect 16028 5040 16080 5092
rect 12900 5015 12952 5024
rect 12900 4981 12909 5015
rect 12909 4981 12943 5015
rect 12943 4981 12952 5015
rect 12900 4972 12952 4981
rect 14372 4972 14424 5024
rect 15936 4972 15988 5024
rect 19892 5117 19901 5151
rect 19901 5117 19935 5151
rect 19935 5117 19944 5151
rect 19892 5108 19944 5117
rect 20628 5176 20680 5228
rect 21456 5108 21508 5160
rect 18604 4972 18656 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 4712 4768 4764 4820
rect 5448 4768 5500 4820
rect 6368 4768 6420 4820
rect 6736 4811 6788 4820
rect 6736 4777 6745 4811
rect 6745 4777 6779 4811
rect 6779 4777 6788 4811
rect 6736 4768 6788 4777
rect 9128 4768 9180 4820
rect 6092 4700 6144 4752
rect 10600 4768 10652 4820
rect 13544 4700 13596 4752
rect 7656 4675 7708 4684
rect 5080 4564 5132 4616
rect 5540 4564 5592 4616
rect 3700 4496 3752 4548
rect 4068 4496 4120 4548
rect 6000 4564 6052 4616
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 6828 4564 6880 4616
rect 7380 4564 7432 4616
rect 7656 4641 7665 4675
rect 7665 4641 7699 4675
rect 7699 4641 7708 4675
rect 7656 4632 7708 4641
rect 8668 4632 8720 4684
rect 12348 4675 12400 4684
rect 12348 4641 12357 4675
rect 12357 4641 12391 4675
rect 12391 4641 12400 4675
rect 12348 4632 12400 4641
rect 8208 4564 8260 4616
rect 9220 4564 9272 4616
rect 10692 4564 10744 4616
rect 12992 4607 13044 4616
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 2136 4428 2188 4480
rect 2320 4471 2372 4480
rect 2320 4437 2329 4471
rect 2329 4437 2363 4471
rect 2363 4437 2372 4471
rect 2320 4428 2372 4437
rect 2872 4428 2924 4480
rect 4436 4428 4488 4480
rect 4620 4428 4672 4480
rect 4988 4428 5040 4480
rect 6368 4496 6420 4548
rect 6552 4428 6604 4480
rect 9404 4496 9456 4548
rect 11888 4496 11940 4548
rect 12992 4573 13001 4607
rect 13001 4573 13035 4607
rect 13035 4573 13044 4607
rect 12992 4564 13044 4573
rect 14096 4607 14148 4616
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 16212 4768 16264 4820
rect 17868 4811 17920 4820
rect 15476 4700 15528 4752
rect 16856 4743 16908 4752
rect 15200 4632 15252 4684
rect 15936 4675 15988 4684
rect 15936 4641 15945 4675
rect 15945 4641 15979 4675
rect 15979 4641 15988 4675
rect 15936 4632 15988 4641
rect 16856 4709 16865 4743
rect 16865 4709 16899 4743
rect 16899 4709 16908 4743
rect 16856 4700 16908 4709
rect 17868 4777 17877 4811
rect 17877 4777 17911 4811
rect 17911 4777 17920 4811
rect 17868 4768 17920 4777
rect 19064 4700 19116 4752
rect 13268 4496 13320 4548
rect 14740 4496 14792 4548
rect 15016 4496 15068 4548
rect 8484 4428 8536 4480
rect 9128 4428 9180 4480
rect 10232 4428 10284 4480
rect 10692 4471 10744 4480
rect 10692 4437 10701 4471
rect 10701 4437 10735 4471
rect 10735 4437 10744 4471
rect 10692 4428 10744 4437
rect 10968 4471 11020 4480
rect 10968 4437 10977 4471
rect 10977 4437 11011 4471
rect 11011 4437 11020 4471
rect 10968 4428 11020 4437
rect 11060 4428 11112 4480
rect 13084 4471 13136 4480
rect 13084 4437 13093 4471
rect 13093 4437 13127 4471
rect 13127 4437 13136 4471
rect 13084 4428 13136 4437
rect 14280 4428 14332 4480
rect 16120 4471 16172 4480
rect 16120 4437 16129 4471
rect 16129 4437 16163 4471
rect 16163 4437 16172 4471
rect 16120 4428 16172 4437
rect 16948 4632 17000 4684
rect 18604 4632 18656 4684
rect 18972 4632 19024 4684
rect 17684 4564 17736 4616
rect 18420 4564 18472 4616
rect 20904 4607 20956 4616
rect 20904 4573 20913 4607
rect 20913 4573 20947 4607
rect 20947 4573 20956 4607
rect 20904 4564 20956 4573
rect 17868 4496 17920 4548
rect 17960 4428 18012 4480
rect 18328 4471 18380 4480
rect 18328 4437 18337 4471
rect 18337 4437 18371 4471
rect 18371 4437 18380 4471
rect 19800 4496 19852 4548
rect 18328 4428 18380 4437
rect 20996 4428 21048 4480
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 3700 4199 3752 4208
rect 3700 4165 3709 4199
rect 3709 4165 3743 4199
rect 3743 4165 3752 4199
rect 3700 4156 3752 4165
rect 4804 4156 4856 4208
rect 5724 4224 5776 4276
rect 2044 4088 2096 4140
rect 2596 4088 2648 4140
rect 3884 4088 3936 4140
rect 4436 4131 4488 4140
rect 4436 4097 4445 4131
rect 4445 4097 4479 4131
rect 4479 4097 4488 4131
rect 4436 4088 4488 4097
rect 5816 4156 5868 4208
rect 6828 4199 6880 4208
rect 6828 4165 6837 4199
rect 6837 4165 6871 4199
rect 6871 4165 6880 4199
rect 6828 4156 6880 4165
rect 4068 4020 4120 4072
rect 1584 3952 1636 4004
rect 4620 3995 4672 4004
rect 4620 3961 4629 3995
rect 4629 3961 4663 3995
rect 4663 3961 4672 3995
rect 4620 3952 4672 3961
rect 6368 4088 6420 4140
rect 6920 4088 6972 4140
rect 6552 4020 6604 4072
rect 7196 4020 7248 4072
rect 8760 4156 8812 4208
rect 12256 4224 12308 4276
rect 13084 4224 13136 4276
rect 14188 4267 14240 4276
rect 14188 4233 14197 4267
rect 14197 4233 14231 4267
rect 14231 4233 14240 4267
rect 14188 4224 14240 4233
rect 15292 4224 15344 4276
rect 16120 4224 16172 4276
rect 17684 4224 17736 4276
rect 18328 4224 18380 4276
rect 18972 4224 19024 4276
rect 10048 4156 10100 4208
rect 8392 4088 8444 4140
rect 8668 4088 8720 4140
rect 9496 4131 9548 4140
rect 9496 4097 9505 4131
rect 9505 4097 9539 4131
rect 9539 4097 9548 4131
rect 9496 4088 9548 4097
rect 10968 4156 11020 4208
rect 12992 4199 13044 4208
rect 10784 4131 10836 4140
rect 10784 4097 10793 4131
rect 10793 4097 10827 4131
rect 10827 4097 10836 4131
rect 10784 4088 10836 4097
rect 11060 4088 11112 4140
rect 5448 3952 5500 4004
rect 9680 3952 9732 4004
rect 10968 4063 11020 4072
rect 10968 4029 10977 4063
rect 10977 4029 11011 4063
rect 11011 4029 11020 4063
rect 10968 4020 11020 4029
rect 11888 4020 11940 4072
rect 12072 4131 12124 4140
rect 12072 4097 12081 4131
rect 12081 4097 12115 4131
rect 12115 4097 12124 4131
rect 12992 4165 13001 4199
rect 13001 4165 13035 4199
rect 13035 4165 13044 4199
rect 12992 4156 13044 4165
rect 13452 4156 13504 4208
rect 15844 4156 15896 4208
rect 17040 4156 17092 4208
rect 18052 4156 18104 4208
rect 12072 4088 12124 4097
rect 12900 4088 12952 4140
rect 12256 4020 12308 4072
rect 13636 4088 13688 4140
rect 15568 4088 15620 4140
rect 16948 4088 17000 4140
rect 19616 4156 19668 4208
rect 18972 4088 19024 4140
rect 19892 4131 19944 4140
rect 19892 4097 19901 4131
rect 19901 4097 19935 4131
rect 19935 4097 19944 4131
rect 19892 4088 19944 4097
rect 20260 4156 20312 4208
rect 20076 4088 20128 4140
rect 20352 4088 20404 4140
rect 21272 4088 21324 4140
rect 14280 4063 14332 4072
rect 14280 4029 14289 4063
rect 14289 4029 14323 4063
rect 14323 4029 14332 4063
rect 14280 4020 14332 4029
rect 11060 3952 11112 4004
rect 14372 3952 14424 4004
rect 15292 4020 15344 4072
rect 15660 4020 15712 4072
rect 20904 4063 20956 4072
rect 15200 3952 15252 4004
rect 1860 3927 1912 3936
rect 1860 3893 1869 3927
rect 1869 3893 1903 3927
rect 1903 3893 1912 3927
rect 1860 3884 1912 3893
rect 3148 3884 3200 3936
rect 3976 3884 4028 3936
rect 4804 3884 4856 3936
rect 4896 3927 4948 3936
rect 4896 3893 4905 3927
rect 4905 3893 4939 3927
rect 4939 3893 4948 3927
rect 4896 3884 4948 3893
rect 5080 3884 5132 3936
rect 5724 3884 5776 3936
rect 6736 3884 6788 3936
rect 7656 3884 7708 3936
rect 8024 3927 8076 3936
rect 8024 3893 8033 3927
rect 8033 3893 8067 3927
rect 8067 3893 8076 3927
rect 8024 3884 8076 3893
rect 9772 3884 9824 3936
rect 10508 3884 10560 3936
rect 14464 3884 14516 3936
rect 15108 3884 15160 3936
rect 17868 3952 17920 4004
rect 15384 3884 15436 3936
rect 16488 3884 16540 3936
rect 19708 3952 19760 4004
rect 20904 4029 20913 4063
rect 20913 4029 20947 4063
rect 20947 4029 20956 4063
rect 20904 4020 20956 4029
rect 21088 4063 21140 4072
rect 21088 4029 21097 4063
rect 21097 4029 21131 4063
rect 21131 4029 21140 4063
rect 21088 4020 21140 4029
rect 21548 3952 21600 4004
rect 19800 3884 19852 3936
rect 20076 3927 20128 3936
rect 20076 3893 20085 3927
rect 20085 3893 20119 3927
rect 20119 3893 20128 3927
rect 20076 3884 20128 3893
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 7196 3680 7248 3732
rect 7656 3680 7708 3732
rect 8116 3680 8168 3732
rect 9128 3680 9180 3732
rect 9864 3680 9916 3732
rect 10784 3723 10836 3732
rect 10784 3689 10793 3723
rect 10793 3689 10827 3723
rect 10827 3689 10836 3723
rect 10784 3680 10836 3689
rect 3056 3612 3108 3664
rect 5448 3612 5500 3664
rect 6368 3612 6420 3664
rect 2320 3476 2372 3528
rect 2688 3476 2740 3528
rect 4712 3544 4764 3596
rect 5264 3544 5316 3596
rect 12716 3680 12768 3732
rect 13728 3680 13780 3732
rect 14372 3680 14424 3732
rect 15568 3680 15620 3732
rect 19892 3680 19944 3732
rect 20812 3680 20864 3732
rect 20904 3680 20956 3732
rect 14096 3612 14148 3664
rect 10232 3587 10284 3596
rect 3976 3519 4028 3528
rect 3976 3485 3985 3519
rect 3985 3485 4019 3519
rect 4019 3485 4028 3519
rect 3976 3476 4028 3485
rect 4436 3476 4488 3528
rect 4528 3476 4580 3528
rect 4896 3519 4948 3528
rect 4896 3485 4905 3519
rect 4905 3485 4939 3519
rect 4939 3485 4948 3519
rect 4896 3476 4948 3485
rect 5724 3476 5776 3528
rect 6276 3519 6328 3528
rect 6276 3485 6285 3519
rect 6285 3485 6319 3519
rect 6319 3485 6328 3519
rect 6276 3476 6328 3485
rect 6736 3519 6788 3528
rect 6736 3485 6745 3519
rect 6745 3485 6779 3519
rect 6779 3485 6788 3519
rect 6736 3476 6788 3485
rect 2596 3340 2648 3392
rect 3700 3408 3752 3460
rect 8668 3476 8720 3528
rect 9220 3476 9272 3528
rect 8116 3408 8168 3460
rect 8392 3408 8444 3460
rect 9312 3408 9364 3460
rect 4252 3340 4304 3392
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 4436 3340 4488 3349
rect 5264 3340 5316 3392
rect 5540 3383 5592 3392
rect 5540 3349 5549 3383
rect 5549 3349 5583 3383
rect 5583 3349 5592 3383
rect 5540 3340 5592 3349
rect 5724 3340 5776 3392
rect 6736 3340 6788 3392
rect 7196 3340 7248 3392
rect 7564 3340 7616 3392
rect 7656 3340 7708 3392
rect 8944 3340 8996 3392
rect 9128 3383 9180 3392
rect 9128 3349 9137 3383
rect 9137 3349 9171 3383
rect 9171 3349 9180 3383
rect 9128 3340 9180 3349
rect 10232 3553 10241 3587
rect 10241 3553 10275 3587
rect 10275 3553 10284 3587
rect 10232 3544 10284 3553
rect 10508 3544 10560 3596
rect 12900 3544 12952 3596
rect 13176 3544 13228 3596
rect 9772 3519 9824 3528
rect 9772 3485 9781 3519
rect 9781 3485 9815 3519
rect 9815 3485 9824 3519
rect 9772 3476 9824 3485
rect 10140 3476 10192 3528
rect 11152 3476 11204 3528
rect 11612 3476 11664 3528
rect 13360 3519 13412 3528
rect 13360 3485 13369 3519
rect 13369 3485 13403 3519
rect 13403 3485 13412 3519
rect 13360 3476 13412 3485
rect 13544 3476 13596 3528
rect 14648 3476 14700 3528
rect 14740 3476 14792 3528
rect 15844 3476 15896 3528
rect 11704 3408 11756 3460
rect 15568 3408 15620 3460
rect 17132 3476 17184 3528
rect 16212 3451 16264 3460
rect 16212 3417 16246 3451
rect 16246 3417 16264 3451
rect 16212 3408 16264 3417
rect 16488 3408 16540 3460
rect 20076 3612 20128 3664
rect 12256 3340 12308 3392
rect 12532 3340 12584 3392
rect 12808 3340 12860 3392
rect 13728 3383 13780 3392
rect 13728 3349 13737 3383
rect 13737 3349 13771 3383
rect 13771 3349 13780 3383
rect 13728 3340 13780 3349
rect 15660 3340 15712 3392
rect 18420 3544 18472 3596
rect 19156 3544 19208 3596
rect 19616 3544 19668 3596
rect 18052 3476 18104 3528
rect 18512 3476 18564 3528
rect 17500 3408 17552 3460
rect 17592 3383 17644 3392
rect 17592 3349 17601 3383
rect 17601 3349 17635 3383
rect 17635 3349 17644 3383
rect 17592 3340 17644 3349
rect 18052 3383 18104 3392
rect 18052 3349 18061 3383
rect 18061 3349 18095 3383
rect 18095 3349 18104 3383
rect 18420 3408 18472 3460
rect 20536 3544 20588 3596
rect 20720 3544 20772 3596
rect 20076 3476 20128 3528
rect 21364 3476 21416 3528
rect 19524 3408 19576 3460
rect 22100 3408 22152 3460
rect 18052 3340 18104 3349
rect 19064 3340 19116 3392
rect 19616 3340 19668 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 1768 3136 1820 3188
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 1676 3000 1728 3052
rect 848 2932 900 2984
rect 1492 2932 1544 2984
rect 2504 3000 2556 3052
rect 2780 3043 2832 3052
rect 2780 3009 2789 3043
rect 2789 3009 2823 3043
rect 2823 3009 2832 3043
rect 3884 3136 3936 3188
rect 3608 3068 3660 3120
rect 2780 3000 2832 3009
rect 3884 3000 3936 3052
rect 4344 3000 4396 3052
rect 4896 3136 4948 3188
rect 5172 3136 5224 3188
rect 4620 3068 4672 3120
rect 4988 3068 5040 3120
rect 8024 3136 8076 3188
rect 2136 2932 2188 2984
rect 5172 3000 5224 3052
rect 5724 2932 5776 2984
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 8668 3068 8720 3120
rect 6828 2975 6880 2984
rect 6828 2941 6837 2975
rect 6837 2941 6871 2975
rect 6871 2941 6880 2975
rect 8024 3000 8076 3052
rect 6828 2932 6880 2941
rect 7656 2932 7708 2984
rect 9404 3136 9456 3188
rect 11244 3136 11296 3188
rect 11704 3136 11756 3188
rect 14280 3179 14332 3188
rect 9036 3068 9088 3120
rect 9956 3068 10008 3120
rect 12716 3068 12768 3120
rect 13084 3068 13136 3120
rect 14280 3145 14289 3179
rect 14289 3145 14323 3179
rect 14323 3145 14332 3179
rect 14280 3136 14332 3145
rect 15752 3136 15804 3188
rect 15016 3068 15068 3120
rect 17408 3068 17460 3120
rect 9404 3000 9456 3052
rect 9588 3043 9640 3052
rect 9588 3009 9597 3043
rect 9597 3009 9631 3043
rect 9631 3009 9640 3043
rect 10232 3043 10284 3052
rect 9588 3000 9640 3009
rect 10232 3009 10241 3043
rect 10241 3009 10275 3043
rect 10275 3009 10284 3043
rect 10232 3000 10284 3009
rect 11060 3000 11112 3052
rect 11244 3000 11296 3052
rect 11888 3000 11940 3052
rect 12532 3000 12584 3052
rect 13912 3043 13964 3052
rect 13912 3009 13921 3043
rect 13921 3009 13955 3043
rect 13955 3009 13964 3043
rect 13912 3000 13964 3009
rect 14648 3043 14700 3052
rect 14648 3009 14657 3043
rect 14657 3009 14691 3043
rect 14691 3009 14700 3043
rect 14648 3000 14700 3009
rect 15660 3000 15712 3052
rect 19156 3136 19208 3188
rect 20260 3179 20312 3188
rect 12440 2932 12492 2984
rect 2596 2864 2648 2916
rect 5908 2864 5960 2916
rect 6920 2864 6972 2916
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 2044 2839 2096 2848
rect 2044 2805 2053 2839
rect 2053 2805 2087 2839
rect 2087 2805 2096 2839
rect 2044 2796 2096 2805
rect 2688 2796 2740 2848
rect 2964 2839 3016 2848
rect 2964 2805 2973 2839
rect 2973 2805 3007 2839
rect 3007 2805 3016 2839
rect 2964 2796 3016 2805
rect 3884 2796 3936 2848
rect 4068 2796 4120 2848
rect 4620 2839 4672 2848
rect 4620 2805 4629 2839
rect 4629 2805 4663 2839
rect 4663 2805 4672 2839
rect 4620 2796 4672 2805
rect 5632 2796 5684 2848
rect 5724 2796 5776 2848
rect 9036 2864 9088 2916
rect 10232 2864 10284 2916
rect 12348 2864 12400 2916
rect 8116 2796 8168 2848
rect 11796 2796 11848 2848
rect 12900 2864 12952 2916
rect 14464 2932 14516 2984
rect 19432 3000 19484 3052
rect 20260 3145 20269 3179
rect 20269 3145 20303 3179
rect 20303 3145 20312 3179
rect 20260 3136 20312 3145
rect 18328 2932 18380 2984
rect 16028 2907 16080 2916
rect 16028 2873 16037 2907
rect 16037 2873 16071 2907
rect 16071 2873 16080 2907
rect 16028 2864 16080 2873
rect 13268 2839 13320 2848
rect 13268 2805 13277 2839
rect 13277 2805 13311 2839
rect 13311 2805 13320 2839
rect 13268 2796 13320 2805
rect 14924 2796 14976 2848
rect 18696 2796 18748 2848
rect 19340 2932 19392 2984
rect 20076 2932 20128 2984
rect 19064 2864 19116 2916
rect 20628 2932 20680 2984
rect 22652 2864 22704 2916
rect 20720 2796 20772 2848
rect 22100 2796 22152 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 3332 2635 3384 2644
rect 3332 2601 3341 2635
rect 3341 2601 3375 2635
rect 3375 2601 3384 2635
rect 3332 2592 3384 2601
rect 3976 2592 4028 2644
rect 5264 2592 5316 2644
rect 5908 2635 5960 2644
rect 5908 2601 5917 2635
rect 5917 2601 5951 2635
rect 5951 2601 5960 2635
rect 5908 2592 5960 2601
rect 7288 2635 7340 2644
rect 3056 2524 3108 2576
rect 3148 2524 3200 2576
rect 3884 2524 3936 2576
rect 5540 2524 5592 2576
rect 296 2456 348 2508
rect 1308 2456 1360 2508
rect 2412 2456 2464 2508
rect 4620 2456 4672 2508
rect 7288 2601 7297 2635
rect 7297 2601 7331 2635
rect 7331 2601 7340 2635
rect 7288 2592 7340 2601
rect 8300 2592 8352 2644
rect 9404 2635 9456 2644
rect 9404 2601 9413 2635
rect 9413 2601 9447 2635
rect 9447 2601 9456 2635
rect 9404 2592 9456 2601
rect 11796 2592 11848 2644
rect 15200 2592 15252 2644
rect 15568 2635 15620 2644
rect 15568 2601 15577 2635
rect 15577 2601 15611 2635
rect 15611 2601 15620 2635
rect 15568 2592 15620 2601
rect 18052 2592 18104 2644
rect 11704 2567 11756 2576
rect 6736 2456 6788 2508
rect 6920 2456 6972 2508
rect 1952 2388 2004 2440
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 4436 2388 4488 2440
rect 5632 2388 5684 2440
rect 10416 2456 10468 2508
rect 11704 2533 11713 2567
rect 11713 2533 11747 2567
rect 11747 2533 11756 2567
rect 11704 2524 11756 2533
rect 12532 2524 12584 2576
rect 16028 2524 16080 2576
rect 14740 2499 14792 2508
rect 14740 2465 14749 2499
rect 14749 2465 14783 2499
rect 14783 2465 14792 2499
rect 14740 2456 14792 2465
rect 20536 2524 20588 2576
rect 4160 2320 4212 2372
rect 5356 2363 5408 2372
rect 5356 2329 5365 2363
rect 5365 2329 5399 2363
rect 5399 2329 5408 2363
rect 5356 2320 5408 2329
rect 5816 2363 5868 2372
rect 5816 2329 5825 2363
rect 5825 2329 5859 2363
rect 5859 2329 5868 2363
rect 5816 2320 5868 2329
rect 6092 2320 6144 2372
rect 6736 2320 6788 2372
rect 7104 2320 7156 2372
rect 9680 2388 9732 2440
rect 9772 2388 9824 2440
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 12716 2431 12768 2440
rect 8484 2320 8536 2372
rect 3976 2295 4028 2304
rect 3976 2261 3985 2295
rect 3985 2261 4019 2295
rect 4019 2261 4028 2295
rect 3976 2252 4028 2261
rect 7196 2252 7248 2304
rect 8208 2252 8260 2304
rect 8944 2295 8996 2304
rect 8944 2261 8953 2295
rect 8953 2261 8987 2295
rect 8987 2261 8996 2295
rect 8944 2252 8996 2261
rect 9404 2320 9456 2372
rect 12716 2397 12725 2431
rect 12725 2397 12759 2431
rect 12759 2397 12768 2431
rect 12716 2388 12768 2397
rect 13268 2388 13320 2440
rect 13728 2388 13780 2440
rect 18236 2456 18288 2508
rect 18696 2499 18748 2508
rect 18696 2465 18705 2499
rect 18705 2465 18739 2499
rect 18739 2465 18748 2499
rect 18696 2456 18748 2465
rect 19800 2456 19852 2508
rect 19248 2388 19300 2440
rect 21088 2431 21140 2440
rect 21088 2397 21097 2431
rect 21097 2397 21131 2431
rect 21131 2397 21140 2431
rect 21088 2388 21140 2397
rect 21364 2431 21416 2440
rect 21364 2397 21373 2431
rect 21373 2397 21407 2431
rect 21407 2397 21416 2431
rect 21364 2388 21416 2397
rect 15016 2320 15068 2372
rect 10968 2295 11020 2304
rect 10968 2261 10977 2295
rect 10977 2261 11011 2295
rect 11011 2261 11020 2295
rect 10968 2252 11020 2261
rect 12072 2295 12124 2304
rect 12072 2261 12081 2295
rect 12081 2261 12115 2295
rect 12115 2261 12124 2295
rect 12072 2252 12124 2261
rect 13176 2252 13228 2304
rect 13360 2295 13412 2304
rect 13360 2261 13369 2295
rect 13369 2261 13403 2295
rect 13403 2261 13412 2295
rect 13728 2295 13780 2304
rect 13360 2252 13412 2261
rect 13728 2261 13737 2295
rect 13737 2261 13771 2295
rect 13771 2261 13780 2295
rect 13728 2252 13780 2261
rect 14280 2295 14332 2304
rect 14280 2261 14289 2295
rect 14289 2261 14323 2295
rect 14323 2261 14332 2295
rect 14280 2252 14332 2261
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 15292 2252 15344 2261
rect 17040 2295 17092 2304
rect 17040 2261 17049 2295
rect 17049 2261 17083 2295
rect 17083 2261 17092 2295
rect 18328 2320 18380 2372
rect 22284 2320 22336 2372
rect 17040 2252 17092 2261
rect 18512 2295 18564 2304
rect 18512 2261 18521 2295
rect 18521 2261 18555 2295
rect 18555 2261 18564 2295
rect 18512 2252 18564 2261
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 2872 2048 2924 2100
rect 7104 2048 7156 2100
rect 8576 2048 8628 2100
rect 13360 2048 13412 2100
rect 14280 2048 14332 2100
rect 17960 2048 18012 2100
rect 4988 1980 5040 2032
rect 12164 1980 12216 2032
rect 12256 1980 12308 2032
rect 12992 1980 13044 2032
rect 13728 1980 13780 2032
rect 18420 1980 18472 2032
rect 5172 1912 5224 1964
rect 10968 1912 11020 1964
rect 12716 1912 12768 1964
rect 18604 1912 18656 1964
rect 2320 1844 2372 1896
rect 6736 1844 6788 1896
rect 8116 1844 8168 1896
rect 8392 1844 8444 1896
rect 13084 1844 13136 1896
rect 15292 1844 15344 1896
rect 19524 1844 19576 1896
rect 7012 1776 7064 1828
rect 16120 1776 16172 1828
rect 9680 1708 9732 1760
rect 10876 1708 10928 1760
rect 11152 1708 11204 1760
rect 8944 1640 8996 1692
rect 12256 1640 12308 1692
rect 14740 1708 14792 1760
rect 20260 1708 20312 1760
rect 17224 1640 17276 1692
rect 3884 1572 3936 1624
rect 9404 1572 9456 1624
rect 9496 1572 9548 1624
rect 15108 1572 15160 1624
rect 9956 1504 10008 1556
rect 11428 1504 11480 1556
rect 12440 1504 12492 1556
rect 14832 1504 14884 1556
rect 8208 1436 8260 1488
rect 12072 1436 12124 1488
rect 13176 1436 13228 1488
rect 14924 1436 14976 1488
rect 19340 1368 19392 1420
rect 20168 1368 20220 1420
rect 9128 1300 9180 1352
rect 16212 1300 16264 1352
rect 17132 1300 17184 1352
rect 19248 1300 19300 1352
rect 7380 1232 7432 1284
rect 15752 1232 15804 1284
rect 11888 1164 11940 1216
rect 18696 1164 18748 1216
rect 6828 1096 6880 1148
rect 18880 1096 18932 1148
rect 6644 1028 6696 1080
rect 17500 1028 17552 1080
rect 9312 960 9364 1012
rect 17868 960 17920 1012
rect 5908 892 5960 944
rect 8668 892 8720 944
rect 9404 892 9456 944
rect 17960 892 18012 944
rect 4528 824 4580 876
rect 19616 824 19668 876
rect 2964 756 3016 808
rect 16948 756 17000 808
rect 5080 688 5132 740
rect 18972 688 19024 740
rect 7932 620 7984 672
rect 17592 620 17644 672
rect 4068 552 4120 604
rect 14464 552 14516 604
rect 21088 552 21140 604
<< metal2 >>
rect 294 22200 350 23000
rect 846 22200 902 23000
rect 1398 22200 1454 23000
rect 1950 22200 2006 23000
rect 2502 22200 2558 23000
rect 3054 22200 3110 23000
rect 3606 22200 3662 23000
rect 4158 22200 4214 23000
rect 4710 22200 4766 23000
rect 5262 22200 5318 23000
rect 5814 22200 5870 23000
rect 6458 22200 6514 23000
rect 7010 22200 7066 23000
rect 7562 22200 7618 23000
rect 8114 22200 8170 23000
rect 8666 22200 8722 23000
rect 9218 22200 9274 23000
rect 9770 22200 9826 23000
rect 10322 22200 10378 23000
rect 10874 22200 10930 23000
rect 11426 22200 11482 23000
rect 12070 22200 12126 23000
rect 12622 22200 12678 23000
rect 13174 22200 13230 23000
rect 13726 22200 13782 23000
rect 14278 22200 14334 23000
rect 14830 22200 14886 23000
rect 14936 22222 15148 22250
rect 308 19854 336 22200
rect 296 19848 348 19854
rect 296 19790 348 19796
rect 860 19786 888 22200
rect 1412 19990 1440 22200
rect 1964 20534 1992 22200
rect 1952 20528 2004 20534
rect 1952 20470 2004 20476
rect 1400 19984 1452 19990
rect 1400 19926 1452 19932
rect 1676 19984 1728 19990
rect 1676 19926 1728 19932
rect 1400 19848 1452 19854
rect 1400 19790 1452 19796
rect 1582 19816 1638 19825
rect 848 19780 900 19786
rect 848 19722 900 19728
rect 1412 17338 1440 19790
rect 1582 19751 1638 19760
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1504 17626 1532 19110
rect 1596 18970 1624 19751
rect 1584 18964 1636 18970
rect 1584 18906 1636 18912
rect 1504 17598 1624 17626
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1504 17241 1532 17478
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1596 17134 1624 17598
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1688 17066 1716 19926
rect 1768 19712 1820 19718
rect 1768 19654 1820 19660
rect 1676 17060 1728 17066
rect 1676 17002 1728 17008
rect 1780 11286 1808 19654
rect 1860 19168 1912 19174
rect 1860 19110 1912 19116
rect 1872 18698 1900 19110
rect 1860 18692 1912 18698
rect 1860 18634 1912 18640
rect 1964 17864 1992 20470
rect 2516 20466 2544 22200
rect 3068 20618 3096 22200
rect 3068 20590 3188 20618
rect 3056 20528 3108 20534
rect 3056 20470 3108 20476
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2320 20324 2372 20330
rect 2320 20266 2372 20272
rect 2044 19916 2096 19922
rect 2044 19858 2096 19864
rect 1872 17836 1992 17864
rect 1872 16794 1900 17836
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 1768 11280 1820 11286
rect 1768 11222 1820 11228
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 1308 6656 1360 6662
rect 1308 6598 1360 6604
rect 848 2984 900 2990
rect 848 2926 900 2932
rect 296 2508 348 2514
rect 296 2450 348 2456
rect 308 800 336 2450
rect 860 800 888 2926
rect 1320 2514 1348 6598
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1412 5817 1440 6258
rect 1584 6112 1636 6118
rect 1584 6054 1636 6060
rect 1676 6112 1728 6118
rect 1676 6054 1728 6060
rect 1398 5808 1454 5817
rect 1596 5778 1624 6054
rect 1398 5743 1454 5752
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1492 5568 1544 5574
rect 1492 5510 1544 5516
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1308 2508 1360 2514
rect 1308 2450 1360 2456
rect 1412 800 1440 2994
rect 1504 2990 1532 5510
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1596 4010 1624 4422
rect 1584 4004 1636 4010
rect 1584 3946 1636 3952
rect 1688 3058 1716 6054
rect 1872 5370 1900 9590
rect 1964 6798 1992 17478
rect 2056 17338 2084 19858
rect 2228 19712 2280 19718
rect 2228 19654 2280 19660
rect 2134 18456 2190 18465
rect 2134 18391 2136 18400
rect 2188 18391 2190 18400
rect 2136 18362 2188 18368
rect 2240 17338 2268 19654
rect 2044 17332 2096 17338
rect 2044 17274 2096 17280
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2332 13326 2360 20266
rect 2410 19272 2466 19281
rect 2410 19207 2466 19216
rect 2424 18970 2452 19207
rect 2412 18964 2464 18970
rect 2412 18906 2464 18912
rect 2412 18624 2464 18630
rect 2410 18592 2412 18601
rect 2464 18592 2466 18601
rect 2410 18527 2466 18536
rect 2516 16794 2544 20402
rect 2964 20256 3016 20262
rect 2964 20198 3016 20204
rect 2870 19816 2926 19825
rect 2780 19780 2832 19786
rect 2870 19751 2926 19760
rect 2780 19722 2832 19728
rect 2688 19236 2740 19242
rect 2688 19178 2740 19184
rect 2596 19168 2648 19174
rect 2596 19110 2648 19116
rect 2608 18465 2636 19110
rect 2594 18456 2650 18465
rect 2594 18391 2650 18400
rect 2700 18154 2728 19178
rect 2792 18154 2820 19722
rect 2884 18426 2912 19751
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2688 18148 2740 18154
rect 2688 18090 2740 18096
rect 2780 18148 2832 18154
rect 2780 18090 2832 18096
rect 2976 17785 3004 20198
rect 2962 17776 3018 17785
rect 2962 17711 3018 17720
rect 2688 17536 2740 17542
rect 2688 17478 2740 17484
rect 2504 16788 2556 16794
rect 2504 16730 2556 16736
rect 2700 16454 2728 17478
rect 3068 17338 3096 20470
rect 3160 19854 3188 20590
rect 3620 20534 3648 22200
rect 4172 20534 4200 22200
rect 4342 21448 4398 21457
rect 4342 21383 4398 21392
rect 3608 20528 3660 20534
rect 4160 20528 4212 20534
rect 3608 20470 3660 20476
rect 3882 20496 3938 20505
rect 3424 20460 3476 20466
rect 4160 20470 4212 20476
rect 3882 20431 3938 20440
rect 3424 20402 3476 20408
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 3344 19990 3372 20198
rect 3332 19984 3384 19990
rect 3332 19926 3384 19932
rect 3148 19848 3200 19854
rect 3148 19790 3200 19796
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3160 17270 3188 19790
rect 3240 19712 3292 19718
rect 3240 19654 3292 19660
rect 3252 19530 3280 19654
rect 3252 19502 3372 19530
rect 3238 19408 3294 19417
rect 3238 19343 3294 19352
rect 3252 18222 3280 19343
rect 3240 18216 3292 18222
rect 3240 18158 3292 18164
rect 3148 17264 3200 17270
rect 3148 17206 3200 17212
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 3344 15065 3372 19502
rect 3436 17338 3464 20402
rect 3549 20156 3857 20176
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20080 3857 20100
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 3804 19156 3832 19654
rect 3896 19514 3924 20431
rect 3976 19848 4028 19854
rect 3976 19790 4028 19796
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 3804 19128 3924 19156
rect 3549 19068 3857 19088
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 18992 3857 19012
rect 3549 17980 3857 18000
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17904 3857 17924
rect 3516 17672 3568 17678
rect 3514 17640 3516 17649
rect 3568 17640 3570 17649
rect 3514 17575 3570 17584
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 3549 16892 3857 16912
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16816 3857 16836
rect 3549 15804 3857 15824
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15728 3857 15748
rect 3330 15056 3386 15065
rect 3330 14991 3386 15000
rect 3549 14716 3857 14736
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14640 3857 14660
rect 3896 13938 3924 19128
rect 3988 17678 4016 19790
rect 4066 19136 4122 19145
rect 4066 19071 4122 19080
rect 4080 18970 4108 19071
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 4066 18864 4122 18873
rect 4066 18799 4068 18808
rect 4120 18799 4122 18808
rect 4068 18770 4120 18776
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 3976 17672 4028 17678
rect 3976 17614 4028 17620
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 3238 13832 3294 13841
rect 3238 13767 3294 13776
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 3056 6792 3108 6798
rect 3056 6734 3108 6740
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2412 5840 2464 5846
rect 2412 5782 2464 5788
rect 2042 5672 2098 5681
rect 2042 5607 2098 5616
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1860 5364 1912 5370
rect 1780 5324 1860 5352
rect 1780 3194 1808 5324
rect 1860 5306 1912 5312
rect 1860 3936 1912 3942
rect 1860 3878 1912 3884
rect 1768 3188 1820 3194
rect 1768 3130 1820 3136
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1492 2984 1544 2990
rect 1492 2926 1544 2932
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1596 921 1624 2790
rect 1872 2417 1900 3878
rect 1964 2446 1992 5510
rect 2056 4146 2084 5607
rect 2228 5024 2280 5030
rect 2228 4966 2280 4972
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2148 2990 2176 4422
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 2044 2848 2096 2854
rect 2044 2790 2096 2796
rect 1952 2440 2004 2446
rect 1858 2408 1914 2417
rect 1952 2382 2004 2388
rect 1858 2343 1914 2352
rect 1582 912 1638 921
rect 1582 847 1638 856
rect 1964 800 1992 2382
rect 294 0 350 800
rect 846 0 902 800
rect 1398 0 1454 800
rect 1950 0 2006 800
rect 2056 649 2084 2790
rect 2240 2009 2268 4966
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2332 4185 2360 4422
rect 2318 4176 2374 4185
rect 2318 4111 2374 4120
rect 2320 3528 2372 3534
rect 2320 3470 2372 3476
rect 2226 2000 2282 2009
rect 2226 1935 2282 1944
rect 2332 1902 2360 3470
rect 2424 2514 2452 5782
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2516 3058 2544 5510
rect 2594 4176 2650 4185
rect 2594 4111 2596 4120
rect 2648 4111 2650 4120
rect 2596 4082 2648 4088
rect 2700 3534 2728 5510
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 2412 2508 2464 2514
rect 2412 2450 2464 2456
rect 2320 1896 2372 1902
rect 2320 1838 2372 1844
rect 2516 800 2544 2994
rect 2608 2922 2636 3334
rect 2792 3058 2820 6394
rect 3068 5522 3096 6734
rect 3160 6458 3188 11018
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3252 5681 3280 13767
rect 3549 13628 3857 13648
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13552 3857 13572
rect 3549 12540 3857 12560
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12464 3857 12484
rect 3549 11452 3857 11472
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11376 3857 11396
rect 3549 10364 3857 10384
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10288 3857 10308
rect 3549 9276 3857 9296
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9200 3857 9220
rect 3332 8424 3384 8430
rect 3332 8366 3384 8372
rect 3238 5672 3294 5681
rect 3238 5607 3294 5616
rect 2976 5494 3096 5522
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2596 2916 2648 2922
rect 2596 2858 2648 2864
rect 2688 2848 2740 2854
rect 2688 2790 2740 2796
rect 2700 1873 2728 2790
rect 2686 1864 2742 1873
rect 2686 1799 2742 1808
rect 2792 1601 2820 2994
rect 2884 2106 2912 4422
rect 2976 3482 3004 5494
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3054 4040 3110 4049
rect 3054 3975 3110 3984
rect 3068 3670 3096 3975
rect 3148 3936 3200 3942
rect 3148 3878 3200 3884
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 2976 3454 3096 3482
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 2778 1592 2834 1601
rect 2778 1527 2834 1536
rect 2976 814 3004 2790
rect 3068 2582 3096 3454
rect 3160 2582 3188 3878
rect 3056 2576 3108 2582
rect 3056 2518 3108 2524
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 3252 2446 3280 5102
rect 3344 2650 3372 8366
rect 3549 8188 3857 8208
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8112 3857 8132
rect 3549 7100 3857 7120
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7024 3857 7044
rect 3896 6458 3924 13874
rect 4080 12434 4108 18362
rect 4172 18358 4200 20470
rect 4356 20058 4384 21383
rect 4528 20324 4580 20330
rect 4528 20266 4580 20272
rect 4540 20097 4568 20266
rect 4526 20088 4582 20097
rect 4344 20052 4396 20058
rect 4526 20023 4582 20032
rect 4344 19994 4396 20000
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4252 19780 4304 19786
rect 4252 19722 4304 19728
rect 4160 18352 4212 18358
rect 4160 18294 4212 18300
rect 4264 17542 4292 19722
rect 4344 19372 4396 19378
rect 4344 19314 4396 19320
rect 4356 17746 4384 19314
rect 4344 17740 4396 17746
rect 4344 17682 4396 17688
rect 4252 17536 4304 17542
rect 4252 17478 4304 17484
rect 4264 16998 4292 17478
rect 4252 16992 4304 16998
rect 4252 16934 4304 16940
rect 4158 14376 4214 14385
rect 4158 14311 4214 14320
rect 3988 12406 4108 12434
rect 3988 11801 4016 12406
rect 3974 11792 4030 11801
rect 3974 11727 4030 11736
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3436 2938 3464 6054
rect 3549 6012 3857 6032
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5936 3857 5956
rect 3549 4924 3857 4944
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4848 3857 4868
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3712 4214 3740 4490
rect 3700 4208 3752 4214
rect 3700 4150 3752 4156
rect 3896 4146 3924 6394
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3988 4026 4016 11727
rect 4172 6746 4200 14311
rect 4264 10266 4292 16934
rect 4448 14550 4476 19790
rect 4724 19666 4752 22200
rect 4896 21208 4948 21214
rect 4896 21150 4948 21156
rect 4804 21140 4856 21146
rect 4804 21082 4856 21088
rect 4816 20058 4844 21082
rect 4804 20052 4856 20058
rect 4804 19994 4856 20000
rect 4802 19952 4858 19961
rect 4802 19887 4858 19896
rect 4816 19854 4844 19887
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4816 19689 4844 19790
rect 4632 19638 4752 19666
rect 4802 19680 4858 19689
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4540 16250 4568 19450
rect 4632 19446 4660 19638
rect 4802 19615 4858 19624
rect 4712 19508 4764 19514
rect 4712 19450 4764 19456
rect 4620 19440 4672 19446
rect 4620 19382 4672 19388
rect 4632 16794 4660 19382
rect 4724 18766 4752 19450
rect 4908 19394 4936 21150
rect 5170 21040 5226 21049
rect 5170 20975 5226 20984
rect 5184 20398 5212 20975
rect 5172 20392 5224 20398
rect 5078 20360 5134 20369
rect 5172 20334 5224 20340
rect 5276 20380 5304 22200
rect 5722 21176 5778 21185
rect 5722 21111 5778 21120
rect 5632 20460 5684 20466
rect 5632 20402 5684 20408
rect 5356 20392 5408 20398
rect 5276 20352 5356 20380
rect 5078 20295 5134 20304
rect 4816 19366 4936 19394
rect 4988 19372 5040 19378
rect 4816 19174 4844 19366
rect 4988 19314 5040 19320
rect 4894 19272 4950 19281
rect 4894 19207 4950 19216
rect 4804 19168 4856 19174
rect 4804 19110 4856 19116
rect 4804 18964 4856 18970
rect 4908 18952 4936 19207
rect 4856 18924 4936 18952
rect 4804 18906 4856 18912
rect 4896 18828 4948 18834
rect 4816 18788 4896 18816
rect 4712 18760 4764 18766
rect 4712 18702 4764 18708
rect 4816 18698 4844 18788
rect 4896 18770 4948 18776
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 4896 18692 4948 18698
rect 4896 18634 4948 18640
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 4724 18068 4752 18566
rect 4804 18080 4856 18086
rect 4724 18040 4804 18068
rect 4804 18022 4856 18028
rect 4712 17536 4764 17542
rect 4712 17478 4764 17484
rect 4620 16788 4672 16794
rect 4620 16730 4672 16736
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4724 16130 4752 17478
rect 4816 17241 4844 18022
rect 4802 17232 4858 17241
rect 4908 17202 4936 18634
rect 5000 17649 5028 19314
rect 5092 19242 5120 20295
rect 5172 19372 5224 19378
rect 5172 19314 5224 19320
rect 5080 19236 5132 19242
rect 5080 19178 5132 19184
rect 5078 19000 5134 19009
rect 5078 18935 5080 18944
rect 5132 18935 5134 18944
rect 5080 18906 5132 18912
rect 5184 18766 5212 19314
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5080 18080 5132 18086
rect 5080 18022 5132 18028
rect 4986 17640 5042 17649
rect 4986 17575 5042 17584
rect 4802 17167 4858 17176
rect 4896 17196 4948 17202
rect 4896 17138 4948 17144
rect 4540 16102 4752 16130
rect 4436 14544 4488 14550
rect 4436 14486 4488 14492
rect 4252 10260 4304 10266
rect 4252 10202 4304 10208
rect 4080 6718 4200 6746
rect 4080 5574 4108 6718
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4068 5568 4120 5574
rect 4068 5510 4120 5516
rect 4080 4554 4108 5510
rect 4068 4548 4120 4554
rect 4068 4490 4120 4496
rect 3896 3998 4016 4026
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3549 3836 3857 3856
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3760 3857 3780
rect 3896 3720 3924 3998
rect 3976 3936 4028 3942
rect 4080 3913 4108 4014
rect 3976 3878 4028 3884
rect 4066 3904 4122 3913
rect 3804 3692 3924 3720
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3608 3120 3660 3126
rect 3608 3062 3660 3068
rect 3620 2938 3648 3062
rect 3436 2910 3648 2938
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3240 2440 3292 2446
rect 3068 2400 3240 2428
rect 2964 808 3016 814
rect 2042 640 2098 649
rect 2042 575 2098 584
rect 2502 0 2558 800
rect 3068 800 3096 2400
rect 3240 2382 3292 2388
rect 3252 2317 3280 2382
rect 3436 1442 3464 2910
rect 3712 2836 3740 3402
rect 3804 3040 3832 3692
rect 3882 3632 3938 3641
rect 3882 3567 3938 3576
rect 3896 3194 3924 3567
rect 3988 3534 4016 3878
rect 4066 3839 4122 3848
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3884 3052 3936 3058
rect 3804 3012 3884 3040
rect 3884 2994 3936 3000
rect 3884 2848 3936 2854
rect 3712 2808 3884 2836
rect 3884 2790 3936 2796
rect 3549 2748 3857 2768
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2672 3857 2692
rect 3988 2650 4016 3470
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 3896 1630 3924 2518
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3884 1624 3936 1630
rect 3884 1566 3936 1572
rect 3988 1465 4016 2246
rect 3974 1456 4030 1465
rect 3436 1414 3648 1442
rect 3620 800 3648 1414
rect 3974 1391 4030 1400
rect 2964 750 3016 756
rect 3054 0 3110 800
rect 3606 0 3662 800
rect 4080 610 4108 2790
rect 4172 2378 4200 6598
rect 4264 5914 4292 6598
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4436 5704 4488 5710
rect 4434 5672 4436 5681
rect 4488 5672 4490 5681
rect 4344 5636 4396 5642
rect 4434 5607 4490 5616
rect 4344 5578 4396 5584
rect 4252 5568 4304 5574
rect 4252 5510 4304 5516
rect 4264 3398 4292 5510
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4356 3058 4384 5578
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4448 4146 4476 4422
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4540 3618 4568 16102
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 4632 12434 4660 15914
rect 4632 12406 4752 12434
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4632 4486 4660 5170
rect 4724 5030 4752 12406
rect 4908 11898 4936 17138
rect 4986 16824 5042 16833
rect 4986 16759 4988 16768
rect 5040 16759 5042 16768
rect 4988 16730 5040 16736
rect 5092 16697 5120 18022
rect 5170 17912 5226 17921
rect 5170 17847 5172 17856
rect 5224 17847 5226 17856
rect 5172 17818 5224 17824
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 5184 17218 5212 17682
rect 5276 17338 5304 20352
rect 5356 20334 5408 20340
rect 5448 20256 5500 20262
rect 5448 20198 5500 20204
rect 5356 19372 5408 19378
rect 5356 19314 5408 19320
rect 5368 19174 5396 19314
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 5354 19000 5410 19009
rect 5354 18935 5356 18944
rect 5408 18935 5410 18944
rect 5356 18906 5408 18912
rect 5356 18760 5408 18766
rect 5354 18728 5356 18737
rect 5408 18728 5410 18737
rect 5354 18663 5410 18672
rect 5356 18352 5408 18358
rect 5356 18294 5408 18300
rect 5368 18057 5396 18294
rect 5354 18048 5410 18057
rect 5354 17983 5410 17992
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5184 17190 5304 17218
rect 5078 16688 5134 16697
rect 5078 16623 5134 16632
rect 4986 16552 5042 16561
rect 4986 16487 5042 16496
rect 5000 15910 5028 16487
rect 5276 16046 5304 17190
rect 5368 17134 5396 17165
rect 5356 17128 5408 17134
rect 5354 17096 5356 17105
rect 5408 17096 5410 17105
rect 5354 17031 5410 17040
rect 5368 16794 5396 17031
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5264 16040 5316 16046
rect 5264 15982 5316 15988
rect 4988 15904 5040 15910
rect 4988 15846 5040 15852
rect 5000 12918 5028 15846
rect 5368 15688 5396 16594
rect 5460 16114 5488 20198
rect 5540 19984 5592 19990
rect 5540 19926 5592 19932
rect 5552 16794 5580 19926
rect 5644 18290 5672 20402
rect 5736 19990 5764 21111
rect 5828 20466 5856 22200
rect 6000 21344 6052 21350
rect 6000 21286 6052 21292
rect 5816 20460 5868 20466
rect 5816 20402 5868 20408
rect 5724 19984 5776 19990
rect 5724 19926 5776 19932
rect 6012 19854 6040 21286
rect 6472 20890 6500 22200
rect 6734 21312 6790 21321
rect 6734 21247 6790 21256
rect 6472 20862 6592 20890
rect 6148 20700 6456 20720
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20624 6456 20644
rect 6564 20448 6592 20862
rect 6644 20460 6696 20466
rect 6564 20420 6644 20448
rect 6644 20402 6696 20408
rect 6276 20256 6328 20262
rect 6276 20198 6328 20204
rect 6288 19922 6316 20198
rect 6276 19916 6328 19922
rect 6276 19858 6328 19864
rect 5724 19848 5776 19854
rect 5724 19790 5776 19796
rect 6000 19848 6052 19854
rect 6092 19848 6144 19854
rect 6000 19790 6052 19796
rect 6090 19816 6092 19825
rect 6144 19816 6146 19825
rect 5632 18284 5684 18290
rect 5632 18226 5684 18232
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5368 15660 5488 15688
rect 5460 15450 5488 15660
rect 5552 15638 5580 16730
rect 5644 16658 5672 17614
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5632 16040 5684 16046
rect 5630 16008 5632 16017
rect 5684 16008 5686 16017
rect 5630 15943 5686 15952
rect 5630 15872 5686 15881
rect 5630 15807 5686 15816
rect 5540 15632 5592 15638
rect 5540 15574 5592 15580
rect 5460 15422 5580 15450
rect 5552 14414 5580 15422
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5448 13524 5500 13530
rect 5448 13466 5500 13472
rect 5172 13456 5224 13462
rect 5172 13398 5224 13404
rect 4988 12912 5040 12918
rect 4988 12854 5040 12860
rect 4896 11892 4948 11898
rect 4896 11834 4948 11840
rect 5080 11620 5132 11626
rect 5080 11562 5132 11568
rect 4896 7268 4948 7274
rect 4896 7210 4948 7216
rect 4802 6896 4858 6905
rect 4802 6831 4804 6840
rect 4856 6831 4858 6840
rect 4804 6802 4856 6808
rect 4908 6746 4936 7210
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4816 6718 4936 6746
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4724 4826 4752 4966
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4448 3590 4568 3618
rect 4448 3534 4476 3590
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4344 3052 4396 3058
rect 4344 2994 4396 3000
rect 4448 2446 4476 3334
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 4160 2372 4212 2378
rect 4160 2314 4212 2320
rect 4172 800 4200 2314
rect 4540 882 4568 3470
rect 4632 3126 4660 3946
rect 4724 3777 4752 4762
rect 4816 4214 4844 6718
rect 4896 6112 4948 6118
rect 4896 6054 4948 6060
rect 4908 5030 4936 6054
rect 5000 5574 5028 6802
rect 5092 6458 5120 11562
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 4896 5024 4948 5030
rect 4896 4966 4948 4972
rect 4804 4208 4856 4214
rect 4802 4176 4804 4185
rect 4856 4176 4858 4185
rect 4802 4111 4858 4120
rect 4908 3942 4936 4966
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4710 3768 4766 3777
rect 4710 3703 4766 3712
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4620 3120 4672 3126
rect 4620 3062 4672 3068
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4632 2514 4660 2790
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4528 876 4580 882
rect 4528 818 4580 824
rect 4724 800 4752 3538
rect 4816 2825 4844 3878
rect 4908 3641 4936 3878
rect 4894 3632 4950 3641
rect 4894 3567 4950 3576
rect 4896 3528 4948 3534
rect 4894 3496 4896 3505
rect 4948 3496 4950 3505
rect 4894 3431 4950 3440
rect 5000 3369 5028 4422
rect 5092 3942 5120 4558
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 4986 3360 5042 3369
rect 4986 3295 5042 3304
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 4802 2816 4858 2825
rect 4802 2751 4858 2760
rect 4908 2553 4936 3130
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 4894 2544 4950 2553
rect 4894 2479 4950 2488
rect 5000 2038 5028 3062
rect 4988 2032 5040 2038
rect 4988 1974 5040 1980
rect 4068 604 4120 610
rect 4068 546 4120 552
rect 4158 0 4214 800
rect 4710 0 4766 800
rect 5092 746 5120 3878
rect 5184 3194 5212 13398
rect 5460 13326 5488 13466
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 7546 5488 13262
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5264 7200 5316 7206
rect 5264 7142 5316 7148
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5276 7041 5304 7142
rect 5262 7032 5318 7041
rect 5262 6967 5318 6976
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5276 3602 5304 6598
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5262 3496 5318 3505
rect 5262 3431 5318 3440
rect 5276 3398 5304 3431
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5184 1970 5212 2994
rect 5262 2952 5318 2961
rect 5262 2887 5318 2896
rect 5276 2650 5304 2887
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5368 2378 5396 7142
rect 5460 5302 5488 7482
rect 5552 6390 5580 11154
rect 5644 10538 5672 15807
rect 5736 11286 5764 19790
rect 6090 19751 6146 19760
rect 6550 19816 6606 19825
rect 6550 19751 6606 19760
rect 6148 19612 6456 19632
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19536 6456 19556
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 5828 19224 5856 19314
rect 5828 19196 6040 19224
rect 5816 18964 5868 18970
rect 5816 18906 5868 18912
rect 5828 16182 5856 18906
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5920 18329 5948 18362
rect 5906 18320 5962 18329
rect 5906 18255 5962 18264
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 5816 16176 5868 16182
rect 5816 16118 5868 16124
rect 5816 15360 5868 15366
rect 5816 15302 5868 15308
rect 5724 11280 5776 11286
rect 5724 11222 5776 11228
rect 5828 11082 5856 15302
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5632 10532 5684 10538
rect 5632 10474 5684 10480
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5552 5710 5580 6326
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5448 5296 5500 5302
rect 5446 5264 5448 5273
rect 5500 5264 5502 5273
rect 5446 5199 5502 5208
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5446 4856 5502 4865
rect 5446 4791 5448 4800
rect 5500 4791 5502 4800
rect 5448 4762 5500 4768
rect 5552 4622 5580 4966
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 5538 4176 5594 4185
rect 5538 4111 5594 4120
rect 5446 4040 5502 4049
rect 5446 3975 5448 3984
rect 5500 3975 5502 3984
rect 5448 3946 5500 3952
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5460 3097 5488 3606
rect 5552 3398 5580 4111
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5644 3210 5672 10474
rect 5920 10146 5948 17206
rect 6012 16726 6040 19196
rect 6104 19009 6132 19314
rect 6458 19136 6514 19145
rect 6458 19071 6514 19080
rect 6090 19000 6146 19009
rect 6090 18935 6146 18944
rect 6472 18766 6500 19071
rect 6564 18970 6592 19751
rect 6552 18964 6604 18970
rect 6552 18906 6604 18912
rect 6656 18902 6684 20402
rect 6748 19990 6776 21247
rect 6826 20632 6882 20641
rect 6826 20567 6882 20576
rect 6840 20466 6868 20567
rect 7024 20534 7052 22200
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7104 20936 7156 20942
rect 7104 20878 7156 20884
rect 7012 20528 7064 20534
rect 6918 20496 6974 20505
rect 6828 20460 6880 20466
rect 7012 20470 7064 20476
rect 6918 20431 6974 20440
rect 6828 20402 6880 20408
rect 6828 20324 6880 20330
rect 6828 20266 6880 20272
rect 6736 19984 6788 19990
rect 6736 19926 6788 19932
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6644 18896 6696 18902
rect 6644 18838 6696 18844
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6550 18592 6606 18601
rect 6148 18524 6456 18544
rect 6550 18527 6606 18536
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18448 6456 18468
rect 6564 18426 6592 18527
rect 6552 18420 6604 18426
rect 6552 18362 6604 18368
rect 6148 17436 6456 17456
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17360 6456 17380
rect 6550 17368 6606 17377
rect 6550 17303 6552 17312
rect 6604 17303 6606 17312
rect 6552 17274 6604 17280
rect 6092 17264 6144 17270
rect 6092 17206 6144 17212
rect 6104 16998 6132 17206
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6104 16436 6132 16934
rect 6550 16552 6606 16561
rect 6550 16487 6606 16496
rect 6564 16454 6592 16487
rect 6012 16408 6132 16436
rect 6552 16448 6604 16454
rect 6012 14498 6040 16408
rect 6552 16390 6604 16396
rect 6148 16348 6456 16368
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16272 6456 16292
rect 6656 16289 6684 18702
rect 6748 18290 6776 19790
rect 6840 19145 6868 20266
rect 6932 20058 6960 20431
rect 6920 20052 6972 20058
rect 6920 19994 6972 20000
rect 7010 19952 7066 19961
rect 7010 19887 7066 19896
rect 7024 19446 7052 19887
rect 7116 19514 7144 20878
rect 7380 20800 7432 20806
rect 7380 20742 7432 20748
rect 7196 20596 7248 20602
rect 7196 20538 7248 20544
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 7012 19440 7064 19446
rect 6918 19408 6974 19417
rect 7012 19382 7064 19388
rect 6918 19343 6920 19352
rect 6972 19343 6974 19352
rect 7104 19372 7156 19378
rect 6920 19314 6972 19320
rect 7104 19314 7156 19320
rect 6826 19136 6882 19145
rect 6826 19071 6882 19080
rect 7116 18970 7144 19314
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 6828 18896 6880 18902
rect 6828 18838 6880 18844
rect 6840 18737 6868 18838
rect 6826 18728 6882 18737
rect 6826 18663 6882 18672
rect 6918 18456 6974 18465
rect 6918 18391 6974 18400
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6748 17610 6776 18226
rect 6826 18184 6882 18193
rect 6826 18119 6828 18128
rect 6880 18119 6882 18128
rect 6828 18090 6880 18096
rect 6932 17882 6960 18391
rect 7208 18358 7236 20538
rect 7288 20460 7340 20466
rect 7288 20402 7340 20408
rect 7300 19378 7328 20402
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7286 18728 7342 18737
rect 7286 18663 7342 18672
rect 7300 18426 7328 18663
rect 7392 18630 7420 20742
rect 7484 18970 7512 20946
rect 7576 20466 7604 22200
rect 7656 20868 7708 20874
rect 7656 20810 7708 20816
rect 7564 20460 7616 20466
rect 7564 20402 7616 20408
rect 7668 19854 7696 20810
rect 8128 20466 8156 22200
rect 8482 21720 8538 21729
rect 8482 21655 8538 21664
rect 8208 21276 8260 21282
rect 8208 21218 8260 21224
rect 7932 20460 7984 20466
rect 7932 20402 7984 20408
rect 8116 20460 8168 20466
rect 8116 20402 8168 20408
rect 7840 20392 7892 20398
rect 7840 20334 7892 20340
rect 7748 20256 7800 20262
rect 7746 20224 7748 20233
rect 7800 20224 7802 20233
rect 7746 20159 7802 20168
rect 7748 19916 7800 19922
rect 7748 19858 7800 19864
rect 7656 19848 7708 19854
rect 7656 19790 7708 19796
rect 7668 19718 7696 19790
rect 7656 19712 7708 19718
rect 7656 19654 7708 19660
rect 7564 19372 7616 19378
rect 7564 19314 7616 19320
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7380 18624 7432 18630
rect 7380 18566 7432 18572
rect 7288 18420 7340 18426
rect 7288 18362 7340 18368
rect 7012 18352 7064 18358
rect 7012 18294 7064 18300
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7024 18154 7052 18294
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 7288 18216 7340 18222
rect 7288 18158 7340 18164
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 7024 17762 7052 17818
rect 6932 17734 7052 17762
rect 6932 17678 6960 17734
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6736 17604 6788 17610
rect 6736 17546 6788 17552
rect 7012 17604 7064 17610
rect 7012 17546 7064 17552
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6920 17196 6972 17202
rect 6920 17138 6972 17144
rect 6748 16425 6776 17138
rect 6828 16992 6880 16998
rect 6828 16934 6880 16940
rect 6734 16416 6790 16425
rect 6734 16351 6790 16360
rect 6642 16280 6698 16289
rect 6642 16215 6698 16224
rect 6458 16144 6514 16153
rect 6458 16079 6514 16088
rect 6472 15502 6500 16079
rect 6550 16008 6606 16017
rect 6550 15943 6606 15952
rect 6460 15496 6512 15502
rect 6182 15464 6238 15473
rect 6460 15438 6512 15444
rect 6182 15399 6184 15408
rect 6236 15399 6238 15408
rect 6184 15370 6236 15376
rect 6148 15260 6456 15280
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15184 6456 15204
rect 6460 14816 6512 14822
rect 6460 14758 6512 14764
rect 6472 14657 6500 14758
rect 6458 14648 6514 14657
rect 6564 14618 6592 15943
rect 6656 15881 6684 16215
rect 6642 15872 6698 15881
rect 6642 15807 6698 15816
rect 6736 15632 6788 15638
rect 6736 15574 6788 15580
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6458 14583 6514 14592
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 6656 14521 6684 15302
rect 6642 14512 6698 14521
rect 6012 14470 6592 14498
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 5736 10118 5948 10146
rect 5736 9382 5764 10118
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 5724 9376 5776 9382
rect 5724 9318 5776 9324
rect 5736 5545 5764 9318
rect 5828 6662 5856 9998
rect 5908 9920 5960 9926
rect 5906 9888 5908 9897
rect 5960 9888 5962 9897
rect 5906 9823 5962 9832
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5920 6440 5948 7142
rect 5828 6412 5948 6440
rect 5828 5953 5856 6412
rect 5814 5944 5870 5953
rect 5814 5879 5870 5888
rect 5828 5846 5856 5879
rect 5816 5840 5868 5846
rect 6012 5817 6040 14350
rect 6148 14172 6456 14192
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14096 6456 14116
rect 6148 13084 6456 13104
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13008 6456 13028
rect 6564 12434 6592 14470
rect 6642 14447 6698 14456
rect 6564 12406 6684 12434
rect 6148 11996 6456 12016
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11920 6456 11940
rect 6552 11688 6604 11694
rect 6552 11630 6604 11636
rect 6148 10908 6456 10928
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10832 6456 10852
rect 6564 9926 6592 11630
rect 6656 10470 6684 12406
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6748 10062 6776 15574
rect 6840 14890 6868 16934
rect 6932 16794 6960 17138
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6932 15978 6960 16730
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 7024 15706 7052 17546
rect 7116 17134 7144 18158
rect 7196 18148 7248 18154
rect 7196 18090 7248 18096
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6932 15337 6960 15370
rect 6918 15328 6974 15337
rect 6918 15263 6974 15272
rect 6828 14884 6880 14890
rect 6828 14826 6880 14832
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7024 14618 7052 14758
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7012 14476 7064 14482
rect 7012 14418 7064 14424
rect 6920 13252 6972 13258
rect 6920 13194 6972 13200
rect 6932 11898 6960 13194
rect 6920 11892 6972 11898
rect 6920 11834 6972 11840
rect 6826 11656 6882 11665
rect 6826 11591 6882 11600
rect 6840 11354 6868 11591
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 7024 10996 7052 14418
rect 7116 13870 7144 17070
rect 7208 15162 7236 18090
rect 7300 17882 7328 18158
rect 7470 18048 7526 18057
rect 7470 17983 7526 17992
rect 7288 17876 7340 17882
rect 7288 17818 7340 17824
rect 7288 15972 7340 15978
rect 7288 15914 7340 15920
rect 7300 15434 7328 15914
rect 7288 15428 7340 15434
rect 7288 15370 7340 15376
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7208 14482 7236 15098
rect 7196 14476 7248 14482
rect 7196 14418 7248 14424
rect 7104 13864 7156 13870
rect 7104 13806 7156 13812
rect 6932 10968 7052 10996
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6644 9988 6696 9994
rect 6644 9930 6696 9936
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6148 9820 6456 9840
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9744 6456 9764
rect 6550 8936 6606 8945
rect 6550 8871 6552 8880
rect 6604 8871 6606 8880
rect 6552 8842 6604 8848
rect 6148 8732 6456 8752
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8656 6456 8676
rect 6552 7880 6604 7886
rect 6550 7848 6552 7857
rect 6604 7848 6606 7857
rect 6550 7783 6606 7792
rect 6148 7644 6456 7664
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7568 6456 7588
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6148 6556 6456 6576
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6480 6456 6500
rect 6564 6440 6592 6666
rect 6472 6412 6592 6440
rect 5816 5782 5868 5788
rect 5998 5808 6054 5817
rect 5998 5743 6054 5752
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5722 5536 5778 5545
rect 5722 5471 5778 5480
rect 5920 5409 5948 5646
rect 6012 5574 6040 5743
rect 6472 5642 6500 6412
rect 6552 6248 6604 6254
rect 6550 6216 6552 6225
rect 6604 6216 6606 6225
rect 6550 6151 6606 6160
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6564 5794 6592 6054
rect 6656 5914 6684 9930
rect 6734 9888 6790 9897
rect 6734 9823 6790 9832
rect 6748 6866 6776 9823
rect 6840 9654 6868 10406
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6826 9480 6882 9489
rect 6826 9415 6882 9424
rect 6840 9382 6868 9415
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6932 9042 6960 10968
rect 7116 9738 7144 13806
rect 7194 13424 7250 13433
rect 7194 13359 7250 13368
rect 7208 13190 7236 13359
rect 7196 13184 7248 13190
rect 7194 13152 7196 13161
rect 7248 13152 7250 13161
rect 7194 13087 7250 13096
rect 7484 12986 7512 17983
rect 7576 17513 7604 19314
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7562 17504 7618 17513
rect 7562 17439 7618 17448
rect 7576 17241 7604 17439
rect 7668 17338 7696 18566
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7562 17232 7618 17241
rect 7562 17167 7618 17176
rect 7576 17082 7604 17167
rect 7576 17054 7696 17082
rect 7564 16992 7616 16998
rect 7564 16934 7616 16940
rect 7576 16114 7604 16934
rect 7564 16108 7616 16114
rect 7564 16050 7616 16056
rect 7668 15994 7696 17054
rect 7576 15966 7696 15994
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7286 12880 7342 12889
rect 7286 12815 7342 12824
rect 7196 11892 7248 11898
rect 7196 11834 7248 11840
rect 7024 9710 7144 9738
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6734 6760 6790 6769
rect 6734 6695 6790 6704
rect 6748 6662 6776 6695
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6734 6488 6790 6497
rect 6734 6423 6736 6432
rect 6788 6423 6790 6432
rect 6736 6394 6788 6400
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6564 5766 6684 5794
rect 6748 5778 6776 6122
rect 6550 5672 6606 5681
rect 6460 5636 6512 5642
rect 6550 5607 6606 5616
rect 6460 5578 6512 5584
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 6148 5468 6456 5488
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 5906 5400 5962 5409
rect 6148 5392 6456 5412
rect 5906 5335 5962 5344
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5736 4282 5764 5170
rect 5816 5160 5868 5166
rect 5868 5120 5948 5148
rect 5816 5102 5868 5108
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5722 4040 5778 4049
rect 5722 3975 5778 3984
rect 5736 3942 5764 3975
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5722 3768 5778 3777
rect 5722 3703 5778 3712
rect 5736 3534 5764 3703
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5736 3398 5764 3470
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5552 3182 5672 3210
rect 5446 3088 5502 3097
rect 5446 3023 5502 3032
rect 5552 2582 5580 3182
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5736 2854 5764 2926
rect 5632 2848 5684 2854
rect 5632 2790 5684 2796
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 5644 2446 5672 2790
rect 5828 2530 5856 4150
rect 5920 3040 5948 5120
rect 6000 5092 6052 5098
rect 6000 5034 6052 5040
rect 6012 4622 6040 5034
rect 6104 4758 6132 5238
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6092 4752 6144 4758
rect 6092 4694 6144 4700
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 6012 3176 6040 4558
rect 6380 4554 6408 4762
rect 6472 4593 6500 5170
rect 6564 4622 6592 5607
rect 6656 5234 6684 5766
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6840 5302 6868 8910
rect 7024 8090 7052 9710
rect 7102 9616 7158 9625
rect 7102 9551 7104 9560
rect 7156 9551 7158 9560
rect 7104 9522 7156 9528
rect 7104 9036 7156 9042
rect 7104 8978 7156 8984
rect 7012 8084 7064 8090
rect 7012 8026 7064 8032
rect 6918 7984 6974 7993
rect 7116 7970 7144 8978
rect 6918 7919 6974 7928
rect 7024 7942 7144 7970
rect 6932 6866 6960 7919
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6828 5296 6880 5302
rect 6828 5238 6880 5244
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6552 4616 6604 4622
rect 6458 4584 6514 4593
rect 6368 4548 6420 4554
rect 6552 4558 6604 4564
rect 6458 4519 6514 4528
rect 6368 4490 6420 4496
rect 6552 4480 6604 4486
rect 6550 4448 6552 4457
rect 6604 4448 6606 4457
rect 6148 4380 6456 4400
rect 6550 4383 6606 4392
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4304 6456 4324
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 6274 3768 6330 3777
rect 6274 3703 6330 3712
rect 6288 3534 6316 3703
rect 6380 3670 6408 4082
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6368 3664 6420 3670
rect 6368 3606 6420 3612
rect 6276 3528 6328 3534
rect 6276 3470 6328 3476
rect 6148 3292 6456 3312
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3216 6456 3236
rect 6012 3148 6316 3176
rect 5920 3012 6132 3040
rect 5908 2916 5960 2922
rect 5960 2876 6040 2904
rect 5908 2858 5960 2864
rect 5906 2680 5962 2689
rect 5906 2615 5908 2624
rect 5960 2615 5962 2624
rect 5908 2586 5960 2592
rect 5828 2502 5948 2530
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5356 2372 5408 2378
rect 5356 2314 5408 2320
rect 5816 2372 5868 2378
rect 5816 2314 5868 2320
rect 5172 1964 5224 1970
rect 5172 1906 5224 1912
rect 5368 1714 5396 2314
rect 5276 1686 5396 1714
rect 5276 800 5304 1686
rect 5828 800 5856 2314
rect 5920 950 5948 2502
rect 5908 944 5960 950
rect 5908 886 5960 892
rect 5080 740 5132 746
rect 5080 682 5132 688
rect 5262 0 5318 800
rect 5814 0 5870 800
rect 6012 762 6040 2876
rect 6104 2378 6132 3012
rect 6288 2689 6316 3148
rect 6274 2680 6330 2689
rect 6274 2615 6330 2624
rect 6092 2372 6144 2378
rect 6092 2314 6144 2320
rect 6148 2204 6456 2224
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2128 6456 2148
rect 6564 1737 6592 4014
rect 6550 1728 6606 1737
rect 6550 1663 6606 1672
rect 6656 1086 6684 5170
rect 6734 4992 6790 5001
rect 6734 4927 6790 4936
rect 6748 4826 6776 4927
rect 6736 4820 6788 4826
rect 6736 4762 6788 4768
rect 6840 4622 6868 5238
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6828 4208 6880 4214
rect 6826 4176 6828 4185
rect 6880 4176 6882 4185
rect 6932 4146 6960 6666
rect 7024 5522 7052 7942
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7116 7449 7144 7686
rect 7102 7440 7158 7449
rect 7102 7375 7158 7384
rect 7208 6089 7236 11834
rect 7300 10130 7328 12815
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7484 10062 7512 11494
rect 7472 10056 7524 10062
rect 7472 9998 7524 10004
rect 7484 9722 7512 9998
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7300 9217 7328 9590
rect 7286 9208 7342 9217
rect 7286 9143 7342 9152
rect 7300 9110 7328 9143
rect 7288 9104 7340 9110
rect 7288 9046 7340 9052
rect 7576 8838 7604 15966
rect 7760 15892 7788 19858
rect 7852 15994 7880 20334
rect 7944 18086 7972 20402
rect 8024 20392 8076 20398
rect 8024 20334 8076 20340
rect 8036 19718 8064 20334
rect 8220 19854 8248 21218
rect 8300 20324 8352 20330
rect 8300 20266 8352 20272
rect 8208 19848 8260 19854
rect 8208 19790 8260 19796
rect 8024 19712 8076 19718
rect 8024 19654 8076 19660
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8128 19242 8156 19654
rect 8206 19408 8262 19417
rect 8312 19378 8340 20266
rect 8392 19848 8444 19854
rect 8392 19790 8444 19796
rect 8404 19514 8432 19790
rect 8496 19718 8524 21655
rect 8680 20466 8708 22200
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 8574 20088 8630 20097
rect 8574 20023 8630 20032
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 8392 19508 8444 19514
rect 8392 19450 8444 19456
rect 8206 19343 8262 19352
rect 8300 19372 8352 19378
rect 8116 19236 8168 19242
rect 8116 19178 8168 19184
rect 8022 19136 8078 19145
rect 8022 19071 8078 19080
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 8036 17241 8064 19071
rect 8220 18970 8248 19343
rect 8588 19334 8616 20023
rect 8300 19314 8352 19320
rect 8404 19306 8616 19334
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 8208 18352 8260 18358
rect 8208 18294 8260 18300
rect 8220 18057 8248 18294
rect 8206 18048 8262 18057
rect 8206 17983 8262 17992
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8128 17270 8156 17478
rect 8116 17264 8168 17270
rect 8022 17232 8078 17241
rect 7932 17196 7984 17202
rect 8116 17206 8168 17212
rect 8022 17167 8078 17176
rect 7932 17138 7984 17144
rect 7944 16794 7972 17138
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7944 16182 7972 16730
rect 7932 16176 7984 16182
rect 7932 16118 7984 16124
rect 7852 15966 7972 15994
rect 7760 15864 7880 15892
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7760 14822 7788 15438
rect 7748 14816 7800 14822
rect 7748 14758 7800 14764
rect 7760 14550 7788 14758
rect 7748 14544 7800 14550
rect 7748 14486 7800 14492
rect 7748 14272 7800 14278
rect 7748 14214 7800 14220
rect 7760 12850 7788 14214
rect 7748 12844 7800 12850
rect 7748 12786 7800 12792
rect 7746 12744 7802 12753
rect 7746 12679 7802 12688
rect 7656 12368 7708 12374
rect 7654 12336 7656 12345
rect 7708 12336 7710 12345
rect 7654 12271 7710 12280
rect 7654 12200 7710 12209
rect 7654 12135 7710 12144
rect 7668 11626 7696 12135
rect 7656 11620 7708 11626
rect 7656 11562 7708 11568
rect 7668 11150 7696 11562
rect 7760 11354 7788 12679
rect 7748 11348 7800 11354
rect 7748 11290 7800 11296
rect 7656 11144 7708 11150
rect 7656 11086 7708 11092
rect 7654 10840 7710 10849
rect 7654 10775 7710 10784
rect 7668 10266 7696 10775
rect 7746 10568 7802 10577
rect 7746 10503 7748 10512
rect 7800 10503 7802 10512
rect 7748 10474 7800 10480
rect 7656 10260 7708 10266
rect 7708 10220 7788 10248
rect 7656 10202 7708 10208
rect 7656 9920 7708 9926
rect 7656 9862 7708 9868
rect 7668 9722 7696 9862
rect 7656 9716 7708 9722
rect 7656 9658 7708 9664
rect 7564 8832 7616 8838
rect 7562 8800 7564 8809
rect 7616 8800 7618 8809
rect 7562 8735 7618 8744
rect 7760 8616 7788 10220
rect 7668 8588 7788 8616
rect 7286 8392 7342 8401
rect 7286 8327 7342 8336
rect 7300 8294 7328 8327
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7300 6730 7328 8230
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7378 7576 7434 7585
rect 7378 7511 7434 7520
rect 7392 7274 7420 7511
rect 7470 7304 7526 7313
rect 7380 7268 7432 7274
rect 7470 7239 7526 7248
rect 7380 7210 7432 7216
rect 7484 6882 7512 7239
rect 7576 7206 7604 7822
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7668 7018 7696 8588
rect 7746 8528 7802 8537
rect 7746 8463 7802 8472
rect 7760 8430 7788 8463
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7852 8362 7880 15864
rect 7944 10266 7972 15966
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8128 15570 8156 15846
rect 8312 15586 8340 18634
rect 8404 18086 8432 19306
rect 8680 19258 8708 20402
rect 8747 20156 9055 20176
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20080 9055 20100
rect 9232 19802 9260 22200
rect 9586 21856 9642 21865
rect 9586 21791 9642 21800
rect 9312 21072 9364 21078
rect 9312 21014 9364 21020
rect 9048 19774 9260 19802
rect 8760 19372 8812 19378
rect 8760 19314 8812 19320
rect 8588 19230 8708 19258
rect 8588 19224 8616 19230
rect 8496 19196 8616 19224
rect 8496 18902 8524 19196
rect 8772 19156 8800 19314
rect 9048 19310 9076 19774
rect 9128 19712 9180 19718
rect 9128 19654 9180 19660
rect 9036 19304 9088 19310
rect 9036 19246 9088 19252
rect 8680 19128 8800 19156
rect 8576 18964 8628 18970
rect 8576 18906 8628 18912
rect 8484 18896 8536 18902
rect 8484 18838 8536 18844
rect 8588 18766 8616 18906
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8392 18080 8444 18086
rect 8588 18057 8616 18702
rect 8680 18358 8708 19128
rect 8747 19068 9055 19088
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 18992 9055 19012
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 8668 18352 8720 18358
rect 8668 18294 8720 18300
rect 9048 18290 9076 18362
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8680 18086 8708 18158
rect 8668 18080 8720 18086
rect 8392 18022 8444 18028
rect 8574 18048 8630 18057
rect 8668 18022 8720 18028
rect 8574 17983 8630 17992
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8404 16794 8432 17614
rect 8392 16788 8444 16794
rect 8392 16730 8444 16736
rect 8680 16266 8708 18022
rect 8747 17980 9055 18000
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17904 9055 17924
rect 9140 17270 9168 19654
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 8747 16892 9055 16912
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16816 9055 16836
rect 8588 16238 8708 16266
rect 8116 15564 8168 15570
rect 8312 15558 8432 15586
rect 8116 15506 8168 15512
rect 8208 15428 8260 15434
rect 8208 15370 8260 15376
rect 8116 15020 8168 15026
rect 8116 14962 8168 14968
rect 8022 14920 8078 14929
rect 8022 14855 8078 14864
rect 8036 11762 8064 14855
rect 8128 14074 8156 14962
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8220 14006 8248 15370
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8220 13802 8248 13942
rect 8312 13938 8340 14214
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8208 13796 8260 13802
rect 8208 13738 8260 13744
rect 8220 13394 8248 13738
rect 8208 13388 8260 13394
rect 8208 13330 8260 13336
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8114 13016 8170 13025
rect 8114 12951 8116 12960
rect 8168 12951 8170 12960
rect 8116 12922 8168 12928
rect 8116 12640 8168 12646
rect 8116 12582 8168 12588
rect 8128 12238 8156 12582
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8114 11792 8170 11801
rect 8024 11756 8076 11762
rect 8114 11727 8170 11736
rect 8024 11698 8076 11704
rect 8128 11370 8156 11727
rect 8036 11342 8156 11370
rect 7932 10260 7984 10266
rect 7932 10202 7984 10208
rect 7930 10024 7986 10033
rect 7930 9959 7932 9968
rect 7984 9959 7986 9968
rect 7932 9930 7984 9936
rect 8036 8974 8064 11342
rect 8114 11248 8170 11257
rect 8220 11218 8248 13126
rect 8404 12306 8432 15558
rect 8482 15056 8538 15065
rect 8482 14991 8538 15000
rect 8392 12300 8444 12306
rect 8392 12242 8444 12248
rect 8496 11898 8524 14991
rect 8588 14804 8616 16238
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 8747 15804 9055 15824
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15728 9055 15748
rect 9140 15570 9168 15846
rect 9232 15609 9260 19314
rect 9324 19174 9352 21014
rect 9404 20528 9456 20534
rect 9404 20470 9456 20476
rect 9312 19168 9364 19174
rect 9312 19110 9364 19116
rect 9416 18986 9444 20470
rect 9496 20256 9548 20262
rect 9496 20198 9548 20204
rect 9324 18958 9444 18986
rect 9324 18426 9352 18958
rect 9402 18864 9458 18873
rect 9402 18799 9458 18808
rect 9416 18601 9444 18799
rect 9402 18592 9458 18601
rect 9402 18527 9458 18536
rect 9508 18465 9536 20198
rect 9600 19718 9628 21791
rect 9784 21049 9812 22200
rect 9770 21040 9826 21049
rect 9770 20975 9826 20984
rect 9954 21040 10010 21049
rect 9954 20975 10010 20984
rect 9968 20534 9996 20975
rect 10230 20632 10286 20641
rect 10230 20567 10286 20576
rect 9956 20528 10008 20534
rect 9956 20470 10008 20476
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9692 19310 9720 20402
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 9772 19372 9824 19378
rect 9772 19314 9824 19320
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9588 19236 9640 19242
rect 9588 19178 9640 19184
rect 9600 19145 9628 19178
rect 9586 19136 9642 19145
rect 9586 19071 9642 19080
rect 9784 18766 9812 19314
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9956 18760 10008 18766
rect 9956 18702 10008 18708
rect 9494 18456 9550 18465
rect 9312 18420 9364 18426
rect 9494 18391 9550 18400
rect 9862 18456 9918 18465
rect 9862 18391 9918 18400
rect 9312 18362 9364 18368
rect 9324 17134 9352 18362
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 9496 18284 9548 18290
rect 9496 18226 9548 18232
rect 9404 18216 9456 18222
rect 9404 18158 9456 18164
rect 9416 18057 9444 18158
rect 9402 18048 9458 18057
rect 9402 17983 9458 17992
rect 9402 17912 9458 17921
rect 9402 17847 9458 17856
rect 9416 17513 9444 17847
rect 9508 17610 9536 18226
rect 9588 18080 9640 18086
rect 9588 18022 9640 18028
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9402 17504 9458 17513
rect 9402 17439 9458 17448
rect 9312 17128 9364 17134
rect 9312 17070 9364 17076
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 16658 9536 16934
rect 9600 16658 9628 18022
rect 9692 17338 9720 18294
rect 9772 18148 9824 18154
rect 9772 18090 9824 18096
rect 9784 17513 9812 18090
rect 9770 17504 9826 17513
rect 9770 17439 9826 17448
rect 9770 17368 9826 17377
rect 9680 17332 9732 17338
rect 9770 17303 9772 17312
rect 9680 17274 9732 17280
rect 9824 17303 9826 17312
rect 9772 17274 9824 17280
rect 9680 16992 9732 16998
rect 9680 16934 9732 16940
rect 9692 16794 9720 16934
rect 9680 16788 9732 16794
rect 9680 16730 9732 16736
rect 9312 16652 9364 16658
rect 9312 16594 9364 16600
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9324 16538 9352 16594
rect 9324 16510 9444 16538
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9218 15600 9274 15609
rect 9128 15564 9180 15570
rect 9218 15535 9274 15544
rect 9128 15506 9180 15512
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8760 15360 8812 15366
rect 8760 15302 8812 15308
rect 8680 14906 8708 15302
rect 8772 15162 8800 15302
rect 9140 15162 9168 15506
rect 9324 15502 9352 16390
rect 9416 15910 9444 16510
rect 9588 16448 9640 16454
rect 9588 16390 9640 16396
rect 9680 16448 9732 16454
rect 9680 16390 9732 16396
rect 9770 16416 9826 16425
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9600 15706 9628 16390
rect 9692 16250 9720 16390
rect 9770 16351 9826 16360
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9784 16153 9812 16351
rect 9770 16144 9826 16153
rect 9770 16079 9826 16088
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9588 15700 9640 15706
rect 9588 15642 9640 15648
rect 9312 15496 9364 15502
rect 9312 15438 9364 15444
rect 9588 15360 9640 15366
rect 9588 15302 9640 15308
rect 9402 15192 9458 15201
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 9128 15156 9180 15162
rect 9402 15127 9458 15136
rect 9128 15098 9180 15104
rect 9416 14929 9444 15127
rect 9402 14920 9458 14929
rect 8680 14878 9168 14906
rect 8588 14776 8708 14804
rect 8576 13320 8628 13326
rect 8574 13288 8576 13297
rect 8628 13288 8630 13297
rect 8574 13223 8630 13232
rect 8574 12336 8630 12345
rect 8574 12271 8630 12280
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8588 11354 8616 12271
rect 8576 11348 8628 11354
rect 8576 11290 8628 11296
rect 8680 11234 8708 14776
rect 8747 14716 9055 14736
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14640 9055 14660
rect 9140 14482 9168 14878
rect 9402 14855 9458 14864
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 9600 14414 9628 15302
rect 9784 15162 9812 15982
rect 9876 15450 9904 18391
rect 9968 17678 9996 18702
rect 9956 17672 10008 17678
rect 9956 17614 10008 17620
rect 9968 16794 9996 17614
rect 10060 16833 10088 20198
rect 10140 19916 10192 19922
rect 10140 19858 10192 19864
rect 10152 18952 10180 19858
rect 10244 19718 10272 20567
rect 10336 20466 10364 22200
rect 10414 21992 10470 22001
rect 10414 21927 10470 21936
rect 10428 21185 10456 21927
rect 10414 21176 10470 21185
rect 10414 21111 10470 21120
rect 10888 20618 10916 22200
rect 11440 20874 11468 22200
rect 11428 20868 11480 20874
rect 11428 20810 11480 20816
rect 11346 20700 11654 20720
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20624 11654 20644
rect 11794 20632 11850 20641
rect 10888 20590 11100 20618
rect 11072 20534 11100 20590
rect 11794 20567 11850 20576
rect 11060 20528 11112 20534
rect 11060 20470 11112 20476
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10876 20256 10928 20262
rect 10876 20198 10928 20204
rect 10782 20088 10838 20097
rect 10782 20023 10838 20032
rect 10232 19712 10284 19718
rect 10232 19654 10284 19660
rect 10692 19712 10744 19718
rect 10692 19654 10744 19660
rect 10244 19394 10272 19654
rect 10244 19366 10364 19394
rect 10232 18964 10284 18970
rect 10152 18924 10232 18952
rect 10232 18906 10284 18912
rect 10232 18420 10284 18426
rect 10232 18362 10284 18368
rect 10244 18086 10272 18362
rect 10336 18204 10364 19366
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 10416 18896 10468 18902
rect 10416 18838 10468 18844
rect 10428 18306 10456 18838
rect 10520 18426 10548 19314
rect 10600 18964 10652 18970
rect 10600 18906 10652 18912
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10612 18358 10640 18906
rect 10600 18352 10652 18358
rect 10428 18278 10548 18306
rect 10600 18294 10652 18300
rect 10336 18176 10456 18204
rect 10140 18080 10192 18086
rect 10140 18022 10192 18028
rect 10232 18080 10284 18086
rect 10232 18022 10284 18028
rect 10046 16824 10102 16833
rect 9956 16788 10008 16794
rect 10046 16759 10102 16768
rect 9956 16730 10008 16736
rect 9956 16584 10008 16590
rect 9956 16526 10008 16532
rect 9968 15706 9996 16526
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9876 15422 9996 15450
rect 9864 15360 9916 15366
rect 9864 15302 9916 15308
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 9876 14958 9904 15302
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 9324 14074 9352 14282
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9876 14006 9904 14894
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9496 13796 9548 13802
rect 9496 13738 9548 13744
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 8747 13628 9055 13648
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13552 9055 13572
rect 9220 13388 9272 13394
rect 9220 13330 9272 13336
rect 8864 12850 9168 12866
rect 8852 12844 9168 12850
rect 8904 12838 9168 12844
rect 8852 12786 8904 12792
rect 8747 12540 9055 12560
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12464 9055 12484
rect 9140 12434 9168 12838
rect 9232 12442 9260 13330
rect 9048 12406 9168 12434
rect 9220 12436 9272 12442
rect 8760 12368 8812 12374
rect 8760 12310 8812 12316
rect 8772 11762 8800 12310
rect 9048 12238 9076 12406
rect 9220 12378 9272 12384
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 9036 12232 9088 12238
rect 9036 12174 9088 12180
rect 8956 11898 8984 12174
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 9048 11762 9076 12174
rect 9126 11928 9182 11937
rect 9126 11863 9182 11872
rect 8760 11756 8812 11762
rect 8760 11698 8812 11704
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9140 11529 9168 11863
rect 9126 11520 9182 11529
rect 8747 11452 9055 11472
rect 9126 11455 9182 11464
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11376 9055 11396
rect 9220 11348 9272 11354
rect 9220 11290 9272 11296
rect 8114 11183 8170 11192
rect 8208 11212 8260 11218
rect 8128 10810 8156 11183
rect 8208 11154 8260 11160
rect 8496 11206 8708 11234
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8298 10704 8354 10713
rect 8298 10639 8354 10648
rect 8114 10160 8170 10169
rect 8114 10095 8170 10104
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 8036 8634 8064 8910
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 8128 8498 8156 10095
rect 8312 9654 8340 10639
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8404 10198 8432 10474
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8404 9994 8432 10134
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8300 9648 8352 9654
rect 8300 9590 8352 9596
rect 8390 9616 8446 9625
rect 8390 9551 8392 9560
rect 8444 9551 8446 9560
rect 8392 9522 8444 9528
rect 8496 9042 8524 11206
rect 8574 11112 8630 11121
rect 9232 11082 9260 11290
rect 8574 11047 8630 11056
rect 9220 11076 9272 11082
rect 8588 10062 8616 11047
rect 9220 11018 9272 11024
rect 9128 10532 9180 10538
rect 9128 10474 9180 10480
rect 9140 10441 9168 10474
rect 9126 10432 9182 10441
rect 8747 10364 9055 10384
rect 9126 10367 9182 10376
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10288 9055 10308
rect 9126 10296 9182 10305
rect 9126 10231 9182 10240
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 9140 9897 9168 10231
rect 9126 9888 9182 9897
rect 9126 9823 9182 9832
rect 8666 9752 8722 9761
rect 8666 9687 8722 9696
rect 8680 9654 8708 9687
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 8747 9276 9055 9296
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9200 9055 9220
rect 8666 9072 8722 9081
rect 8484 9036 8536 9042
rect 8666 9007 8722 9016
rect 8484 8978 8536 8984
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8588 8566 8616 8774
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 7840 8356 7892 8362
rect 7840 8298 7892 8304
rect 8680 8106 8708 9007
rect 8747 8188 9055 8208
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8112 9055 8132
rect 8496 8078 8708 8106
rect 8496 7954 8524 8078
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7392 6854 7512 6882
rect 7576 6990 7696 7018
rect 7288 6724 7340 6730
rect 7288 6666 7340 6672
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7194 6080 7250 6089
rect 7194 6015 7250 6024
rect 7300 5817 7328 6258
rect 7286 5808 7342 5817
rect 7286 5743 7342 5752
rect 7392 5658 7420 6854
rect 7472 6792 7524 6798
rect 7472 6734 7524 6740
rect 7484 6361 7512 6734
rect 7470 6352 7526 6361
rect 7470 6287 7526 6296
rect 7472 6112 7524 6118
rect 7472 6054 7524 6060
rect 7484 5914 7512 6054
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7392 5630 7512 5658
rect 7380 5568 7432 5574
rect 7024 5494 7236 5522
rect 7380 5510 7432 5516
rect 7012 5228 7064 5234
rect 7012 5170 7064 5176
rect 6826 4111 6882 4120
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6826 4040 6882 4049
rect 6826 3975 6882 3984
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 3534 6776 3878
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6736 3392 6788 3398
rect 6734 3360 6736 3369
rect 6788 3360 6790 3369
rect 6734 3295 6790 3304
rect 6734 3224 6790 3233
rect 6734 3159 6790 3168
rect 6748 2514 6776 3159
rect 6840 2990 6868 3975
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6920 2916 6972 2922
rect 6920 2858 6972 2864
rect 6826 2680 6882 2689
rect 6826 2615 6882 2624
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 6748 1902 6776 2314
rect 6736 1896 6788 1902
rect 6736 1838 6788 1844
rect 6840 1154 6868 2615
rect 6932 2514 6960 2858
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7024 1834 7052 5170
rect 7208 4468 7236 5494
rect 7392 5234 7420 5510
rect 7380 5228 7432 5234
rect 7380 5170 7432 5176
rect 7380 4616 7432 4622
rect 7380 4558 7432 4564
rect 7116 4440 7236 4468
rect 7116 2774 7144 4440
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7208 3738 7236 4014
rect 7392 3754 7420 4558
rect 7484 4264 7512 5630
rect 7576 4842 7604 6990
rect 7656 5364 7708 5370
rect 7656 5306 7708 5312
rect 7668 5273 7696 5306
rect 7654 5264 7710 5273
rect 7654 5199 7710 5208
rect 7760 5030 7788 7482
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7576 4814 7788 4842
rect 7654 4720 7710 4729
rect 7654 4655 7656 4664
rect 7708 4655 7710 4664
rect 7656 4626 7708 4632
rect 7484 4236 7696 4264
rect 7668 3942 7696 4236
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7392 3738 7696 3754
rect 7196 3732 7248 3738
rect 7392 3732 7708 3738
rect 7392 3726 7656 3732
rect 7196 3674 7248 3680
rect 7656 3674 7708 3680
rect 7484 3454 7696 3482
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7208 2836 7236 3334
rect 7484 3176 7512 3454
rect 7668 3398 7696 3454
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7300 3148 7512 3176
rect 7300 3058 7328 3148
rect 7288 3052 7340 3058
rect 7576 3040 7604 3334
rect 7288 2994 7340 3000
rect 7484 3012 7604 3040
rect 7208 2808 7420 2836
rect 7116 2746 7236 2774
rect 7104 2372 7156 2378
rect 7104 2314 7156 2320
rect 7116 2106 7144 2314
rect 7208 2310 7236 2746
rect 7286 2680 7342 2689
rect 7286 2615 7288 2624
rect 7340 2615 7342 2624
rect 7288 2586 7340 2592
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 7104 2100 7156 2106
rect 7104 2042 7156 2048
rect 7012 1828 7064 1834
rect 7012 1770 7064 1776
rect 7010 1320 7066 1329
rect 7392 1290 7420 2808
rect 7484 2292 7512 3012
rect 7656 2984 7708 2990
rect 7760 2972 7788 4814
rect 7708 2944 7788 2972
rect 7656 2926 7708 2932
rect 7484 2264 7604 2292
rect 7010 1255 7066 1264
rect 7380 1284 7432 1290
rect 6828 1148 6880 1154
rect 6828 1090 6880 1096
rect 6644 1080 6696 1086
rect 6644 1022 6696 1028
rect 6380 836 6500 864
rect 6380 762 6408 836
rect 6472 800 6500 836
rect 7024 800 7052 1255
rect 7380 1226 7432 1232
rect 7576 800 7604 2264
rect 6012 734 6408 762
rect 6458 0 6514 800
rect 7010 0 7066 800
rect 7562 0 7618 800
rect 7852 785 7880 7754
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 7478 8248 7686
rect 8208 7472 8260 7478
rect 8208 7414 8260 7420
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8404 6866 8432 7346
rect 8392 6860 8444 6866
rect 8392 6802 8444 6808
rect 8390 6760 8446 6769
rect 8390 6695 8446 6704
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8024 6384 8076 6390
rect 8024 6326 8076 6332
rect 8036 5778 8064 6326
rect 8128 5914 8156 6598
rect 8220 6458 8248 6598
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8300 5840 8352 5846
rect 8300 5782 8352 5788
rect 8024 5772 8076 5778
rect 8024 5714 8076 5720
rect 8206 5672 8262 5681
rect 8206 5607 8262 5616
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7838 776 7894 785
rect 7838 711 7894 720
rect 7944 678 7972 5510
rect 8022 5400 8078 5409
rect 8022 5335 8078 5344
rect 8036 5234 8064 5335
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8114 5128 8170 5137
rect 8114 5063 8170 5072
rect 8128 5030 8156 5063
rect 8116 5024 8168 5030
rect 8116 4966 8168 4972
rect 8220 4706 8248 5607
rect 8128 4678 8248 4706
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 8036 3194 8064 3878
rect 8128 3738 8156 4678
rect 8208 4616 8260 4622
rect 8208 4558 8260 4564
rect 8116 3732 8168 3738
rect 8116 3674 8168 3680
rect 8116 3460 8168 3466
rect 8116 3402 8168 3408
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 8036 2825 8064 2994
rect 8128 2854 8156 3402
rect 8116 2848 8168 2854
rect 8022 2816 8078 2825
rect 8116 2790 8168 2796
rect 8022 2751 8078 2760
rect 8220 2530 8248 4558
rect 8312 3346 8340 5782
rect 8404 5370 8432 6695
rect 8392 5364 8444 5370
rect 8392 5306 8444 5312
rect 8496 4593 8524 7890
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 8956 7410 8984 7754
rect 9140 7585 9168 9590
rect 9126 7576 9182 7585
rect 9126 7511 9182 7520
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 9140 7177 9168 7511
rect 9126 7168 9182 7177
rect 8747 7100 9055 7120
rect 9126 7103 9182 7112
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7024 9055 7044
rect 8576 6928 8628 6934
rect 8576 6870 8628 6876
rect 8588 6798 8616 6870
rect 9128 6860 9180 6866
rect 9128 6802 9180 6808
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8588 6390 8616 6598
rect 9140 6458 9168 6802
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 8668 6112 8720 6118
rect 9232 6089 9260 11018
rect 9324 10742 9352 13670
rect 9404 13320 9456 13326
rect 9404 13262 9456 13268
rect 9416 12986 9444 13262
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9402 12608 9458 12617
rect 9402 12543 9458 12552
rect 9416 11200 9444 12543
rect 9508 11830 9536 13738
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9692 13433 9720 13466
rect 9678 13424 9734 13433
rect 9678 13359 9734 13368
rect 9586 13016 9642 13025
rect 9586 12951 9642 12960
rect 9600 12617 9628 12951
rect 9586 12608 9642 12617
rect 9586 12543 9642 12552
rect 9876 12170 9904 13806
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9496 11824 9548 11830
rect 9496 11766 9548 11772
rect 9508 11354 9536 11766
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9416 11172 9536 11200
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9312 10736 9364 10742
rect 9312 10678 9364 10684
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 9324 6361 9352 10542
rect 9310 6352 9366 6361
rect 9310 6287 9366 6296
rect 8668 6054 8720 6060
rect 9218 6080 9274 6089
rect 8574 5944 8630 5953
rect 8574 5879 8630 5888
rect 8588 5710 8616 5879
rect 8680 5846 8708 6054
rect 8747 6012 9055 6032
rect 9218 6015 9274 6024
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5936 9055 5956
rect 9218 5944 9274 5953
rect 9218 5879 9274 5888
rect 8668 5840 8720 5846
rect 8668 5782 8720 5788
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8482 4584 8538 4593
rect 8482 4519 8538 4528
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8404 3466 8432 4082
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8312 3318 8432 3346
rect 8298 3224 8354 3233
rect 8298 3159 8354 3168
rect 8312 2650 8340 3159
rect 8300 2644 8352 2650
rect 8300 2586 8352 2592
rect 8220 2502 8340 2530
rect 8208 2304 8260 2310
rect 8208 2246 8260 2252
rect 8116 1896 8168 1902
rect 8116 1838 8168 1844
rect 8128 800 8156 1838
rect 8220 1494 8248 2246
rect 8208 1488 8260 1494
rect 8208 1430 8260 1436
rect 8312 1329 8340 2502
rect 8404 1902 8432 3318
rect 8496 2378 8524 4422
rect 8484 2372 8536 2378
rect 8484 2314 8536 2320
rect 8588 2106 8616 5510
rect 8680 4690 8708 5782
rect 9126 5672 9182 5681
rect 9126 5607 9128 5616
rect 9180 5607 9182 5616
rect 9128 5578 9180 5584
rect 9126 4992 9182 5001
rect 8747 4924 9055 4944
rect 9126 4927 9182 4936
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4848 9055 4868
rect 9140 4826 9168 4927
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9232 4706 9260 5879
rect 9310 5672 9366 5681
rect 9310 5607 9366 5616
rect 9324 5302 9352 5607
rect 9312 5296 9364 5302
rect 9312 5238 9364 5244
rect 9416 5114 9444 11018
rect 9508 10606 9536 11172
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9692 10248 9720 11834
rect 9772 11008 9824 11014
rect 9772 10950 9824 10956
rect 9784 10674 9812 10950
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9508 10220 9720 10248
rect 9508 10130 9536 10220
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9968 9738 9996 15422
rect 10060 15337 10088 16759
rect 10152 15502 10180 18022
rect 10232 17740 10284 17746
rect 10232 17682 10284 17688
rect 10244 17542 10272 17682
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10336 17542 10364 17614
rect 10232 17536 10284 17542
rect 10324 17536 10376 17542
rect 10232 17478 10284 17484
rect 10322 17504 10324 17513
rect 10376 17504 10378 17513
rect 10244 17134 10272 17478
rect 10322 17439 10378 17448
rect 10322 17232 10378 17241
rect 10322 17167 10378 17176
rect 10232 17128 10284 17134
rect 10232 17070 10284 17076
rect 10232 16516 10284 16522
rect 10232 16458 10284 16464
rect 10244 15638 10272 16458
rect 10336 16425 10364 17167
rect 10322 16416 10378 16425
rect 10322 16351 10378 16360
rect 10322 16280 10378 16289
rect 10322 16215 10378 16224
rect 10336 16017 10364 16215
rect 10322 16008 10378 16017
rect 10322 15943 10378 15952
rect 10232 15632 10284 15638
rect 10232 15574 10284 15580
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 10046 15328 10102 15337
rect 10046 15263 10102 15272
rect 10048 14340 10100 14346
rect 10048 14282 10100 14288
rect 10060 12889 10088 14282
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10336 12986 10364 13874
rect 10428 13841 10456 18176
rect 10520 18154 10548 18278
rect 10704 18222 10732 19654
rect 10796 19553 10824 20023
rect 10782 19544 10838 19553
rect 10782 19479 10838 19488
rect 10888 19145 10916 20198
rect 10968 19848 11020 19854
rect 10968 19790 11020 19796
rect 10874 19136 10930 19145
rect 10874 19071 10930 19080
rect 10980 18766 11008 19790
rect 11072 19174 11100 20470
rect 11152 20460 11204 20466
rect 11152 20402 11204 20408
rect 11060 19168 11112 19174
rect 11060 19110 11112 19116
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 10968 18760 11020 18766
rect 10968 18702 11020 18708
rect 10784 18692 10836 18698
rect 10784 18634 10836 18640
rect 10796 18426 10824 18634
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 10784 18420 10836 18426
rect 10784 18362 10836 18368
rect 10888 18290 10916 18566
rect 10966 18456 11022 18465
rect 10966 18391 11022 18400
rect 10876 18284 10928 18290
rect 10876 18226 10928 18232
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10692 18216 10744 18222
rect 10980 18170 11008 18391
rect 10692 18158 10744 18164
rect 10508 18148 10560 18154
rect 10508 18090 10560 18096
rect 10612 17882 10640 18158
rect 10888 18142 11008 18170
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10888 17354 10916 18142
rect 11072 17882 11100 18770
rect 11060 17876 11112 17882
rect 11060 17818 11112 17824
rect 10968 17808 11020 17814
rect 10968 17750 11020 17756
rect 10980 17542 11008 17750
rect 10968 17536 11020 17542
rect 10968 17478 11020 17484
rect 10888 17338 11008 17354
rect 10888 17332 11020 17338
rect 10888 17326 10968 17332
rect 10968 17274 11020 17280
rect 10876 17264 10928 17270
rect 10876 17206 10928 17212
rect 10888 17066 10916 17206
rect 10876 17060 10928 17066
rect 10876 17002 10928 17008
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 11164 16946 11192 20402
rect 11808 20369 11836 20567
rect 11980 20392 12032 20398
rect 11794 20360 11850 20369
rect 11980 20334 12032 20340
rect 11794 20295 11850 20304
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 11256 19310 11284 19790
rect 11888 19780 11940 19786
rect 11888 19722 11940 19728
rect 11346 19612 11654 19632
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19536 11654 19556
rect 11900 19378 11928 19722
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11244 19304 11296 19310
rect 11244 19246 11296 19252
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11256 18698 11284 19110
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11796 18624 11848 18630
rect 11796 18566 11848 18572
rect 11346 18524 11654 18544
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18448 11654 18468
rect 11716 18426 11744 18566
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11334 18048 11390 18057
rect 11334 17983 11390 17992
rect 11244 17808 11296 17814
rect 11242 17776 11244 17785
rect 11296 17776 11298 17785
rect 11242 17711 11298 17720
rect 11348 17610 11376 17983
rect 11704 17672 11756 17678
rect 11704 17614 11756 17620
rect 11336 17604 11388 17610
rect 11336 17546 11388 17552
rect 11346 17436 11654 17456
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17360 11654 17380
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 10796 16697 10824 16934
rect 11164 16918 11284 16946
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 10782 16688 10838 16697
rect 10782 16623 10838 16632
rect 10692 16516 10744 16522
rect 10692 16458 10744 16464
rect 10704 16182 10732 16458
rect 10692 16176 10744 16182
rect 10692 16118 10744 16124
rect 10796 16114 10824 16623
rect 10784 16108 10836 16114
rect 10784 16050 10836 16056
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10968 16040 11020 16046
rect 10968 15982 11020 15988
rect 10888 15434 10916 15982
rect 10980 15910 11008 15982
rect 10968 15904 11020 15910
rect 10968 15846 11020 15852
rect 10980 15570 11008 15846
rect 11164 15706 11192 16730
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 10968 15564 11020 15570
rect 10968 15506 11020 15512
rect 10876 15428 10928 15434
rect 10876 15370 10928 15376
rect 10876 15020 10928 15026
rect 10980 15008 11008 15506
rect 11164 15026 11192 15642
rect 11256 15162 11284 16918
rect 11532 16522 11560 17138
rect 11716 17134 11744 17614
rect 11704 17128 11756 17134
rect 11704 17070 11756 17076
rect 11702 16688 11758 16697
rect 11702 16623 11758 16632
rect 11520 16516 11572 16522
rect 11520 16458 11572 16464
rect 11346 16348 11654 16368
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16272 11654 16292
rect 11716 16250 11744 16623
rect 11704 16244 11756 16250
rect 11704 16186 11756 16192
rect 11346 15260 11654 15280
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15184 11654 15204
rect 11244 15156 11296 15162
rect 11244 15098 11296 15104
rect 11704 15156 11756 15162
rect 11704 15098 11756 15104
rect 10928 14980 11008 15008
rect 11152 15020 11204 15026
rect 10876 14962 10928 14968
rect 11152 14962 11204 14968
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 10782 14784 10838 14793
rect 10782 14719 10838 14728
rect 10796 14385 10824 14719
rect 10876 14408 10928 14414
rect 10782 14376 10838 14385
rect 10876 14350 10928 14356
rect 10966 14376 11022 14385
rect 10782 14311 10838 14320
rect 10888 13938 10916 14350
rect 10966 14311 10968 14320
rect 11020 14311 11022 14320
rect 10968 14282 11020 14288
rect 11164 14074 11192 14826
rect 11244 14816 11296 14822
rect 11244 14758 11296 14764
rect 11256 14482 11284 14758
rect 11244 14476 11296 14482
rect 11244 14418 11296 14424
rect 11716 14362 11744 15098
rect 11808 15094 11836 18566
rect 11900 18426 11928 18702
rect 11888 18420 11940 18426
rect 11888 18362 11940 18368
rect 11888 18284 11940 18290
rect 11888 18226 11940 18232
rect 11900 16998 11928 18226
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11886 15600 11942 15609
rect 11886 15535 11942 15544
rect 11796 15088 11848 15094
rect 11796 15030 11848 15036
rect 11900 14550 11928 15535
rect 11992 15042 12020 20334
rect 12084 20074 12112 22200
rect 12348 21276 12400 21282
rect 12348 21218 12400 21224
rect 12256 20460 12308 20466
rect 12256 20402 12308 20408
rect 12084 20058 12204 20074
rect 12084 20052 12216 20058
rect 12084 20046 12164 20052
rect 12164 19994 12216 20000
rect 12072 19984 12124 19990
rect 12072 19926 12124 19932
rect 12084 19718 12112 19926
rect 12268 19718 12296 20402
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 12256 19712 12308 19718
rect 12256 19654 12308 19660
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 12072 19304 12124 19310
rect 12176 19281 12204 19314
rect 12072 19246 12124 19252
rect 12162 19272 12218 19281
rect 12084 18222 12112 19246
rect 12162 19207 12218 19216
rect 12268 18970 12296 19654
rect 12256 18964 12308 18970
rect 12256 18906 12308 18912
rect 12360 18816 12388 21218
rect 12636 20602 12664 22200
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 13188 20330 13216 22200
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13176 20324 13228 20330
rect 13176 20266 13228 20272
rect 13268 20256 13320 20262
rect 13268 20198 13320 20204
rect 13082 20088 13138 20097
rect 13082 20023 13138 20032
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 13004 18970 13032 19858
rect 13096 19825 13124 20023
rect 13082 19816 13138 19825
rect 13082 19751 13138 19760
rect 13096 19718 13124 19751
rect 13084 19712 13136 19718
rect 13084 19654 13136 19660
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 12992 18964 13044 18970
rect 12992 18906 13044 18912
rect 12900 18896 12952 18902
rect 12900 18838 12952 18844
rect 12176 18788 12388 18816
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 12084 17377 12112 18022
rect 12070 17368 12126 17377
rect 12070 17303 12126 17312
rect 12176 17082 12204 18788
rect 12912 18426 12940 18838
rect 12256 18420 12308 18426
rect 12256 18362 12308 18368
rect 12900 18420 12952 18426
rect 12900 18362 12952 18368
rect 12268 17134 12296 18362
rect 13004 18290 13032 18906
rect 13096 18766 13124 19246
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 13280 18698 13308 20198
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 12348 18148 12400 18154
rect 12348 18090 12400 18096
rect 12084 17054 12204 17082
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 12084 15162 12112 17054
rect 12164 16992 12216 16998
rect 12164 16934 12216 16940
rect 12176 16590 12204 16934
rect 12268 16794 12296 17070
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12164 16584 12216 16590
rect 12164 16526 12216 16532
rect 12164 15428 12216 15434
rect 12164 15370 12216 15376
rect 12072 15156 12124 15162
rect 12072 15098 12124 15104
rect 11992 15014 12112 15042
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11716 14334 11836 14362
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11346 14172 11654 14192
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14096 11654 14116
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10414 13832 10470 13841
rect 10414 13767 10470 13776
rect 10888 13530 10916 13874
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 10784 13456 10836 13462
rect 10784 13398 10836 13404
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10046 12880 10102 12889
rect 10046 12815 10102 12824
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10048 11688 10100 11694
rect 10048 11630 10100 11636
rect 10060 10810 10088 11630
rect 10244 10810 10272 12786
rect 10336 11626 10364 12922
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10140 10600 10192 10606
rect 10140 10542 10192 10548
rect 10152 10198 10180 10542
rect 10232 10464 10284 10470
rect 10232 10406 10284 10412
rect 10244 10266 10272 10406
rect 10232 10260 10284 10266
rect 10232 10202 10284 10208
rect 10140 10192 10192 10198
rect 10428 10146 10456 12854
rect 10796 12238 10824 13398
rect 10888 12306 10916 13466
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 10876 12300 10928 12306
rect 10876 12242 10928 12248
rect 10784 12232 10836 12238
rect 10784 12174 10836 12180
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 10520 11082 10548 12038
rect 11164 11830 11192 12038
rect 11152 11824 11204 11830
rect 11152 11766 11204 11772
rect 11256 11354 11284 13194
rect 11346 13084 11654 13104
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13008 11654 13028
rect 11716 12646 11744 14214
rect 11808 13462 11836 14334
rect 11888 14272 11940 14278
rect 11888 14214 11940 14220
rect 11796 13456 11848 13462
rect 11796 13398 11848 13404
rect 11794 13152 11850 13161
rect 11794 13087 11850 13096
rect 11704 12640 11756 12646
rect 11808 12617 11836 13087
rect 11704 12582 11756 12588
rect 11794 12608 11850 12617
rect 11716 12306 11744 12582
rect 11794 12543 11850 12552
rect 11704 12300 11756 12306
rect 11704 12242 11756 12248
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11612 12164 11664 12170
rect 11664 12124 11744 12152
rect 11612 12106 11664 12112
rect 11346 11996 11654 12016
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11920 11654 11940
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10796 10810 10824 11290
rect 11348 11218 11376 11562
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11346 10908 11654 10928
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11150 10840 11206 10849
rect 10784 10804 10836 10810
rect 11346 10832 11654 10852
rect 11150 10775 11206 10784
rect 10784 10746 10836 10752
rect 11164 10674 11192 10775
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10140 10134 10192 10140
rect 9876 9710 9996 9738
rect 10244 10118 10456 10146
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9508 9042 9536 9590
rect 9876 9586 9904 9710
rect 10244 9674 10272 10118
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10324 9988 10376 9994
rect 10324 9930 10376 9936
rect 10336 9761 10364 9930
rect 10322 9752 10378 9761
rect 10322 9687 10378 9696
rect 9968 9646 10272 9674
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 9600 9042 9628 9318
rect 9496 9036 9548 9042
rect 9496 8978 9548 8984
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9508 8362 9536 8978
rect 9864 8424 9916 8430
rect 9864 8366 9916 8372
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9588 8288 9640 8294
rect 9588 8230 9640 8236
rect 9600 8090 9628 8230
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9680 7200 9732 7206
rect 9680 7142 9732 7148
rect 9692 6866 9720 7142
rect 9680 6860 9732 6866
rect 9680 6802 9732 6808
rect 9680 6656 9732 6662
rect 9680 6598 9732 6604
rect 9692 6458 9720 6598
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9494 6352 9550 6361
rect 9784 6338 9812 8026
rect 9876 7834 9904 8366
rect 9968 8022 9996 9646
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10244 9178 10272 9318
rect 10428 9178 10456 9998
rect 11072 9994 11100 10542
rect 11244 10464 11296 10470
rect 11244 10406 11296 10412
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11072 9518 11100 9930
rect 11256 9586 11284 10406
rect 11716 9994 11744 12124
rect 11808 11898 11836 12174
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11808 11150 11836 11834
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11346 9820 11654 9840
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9744 11654 9764
rect 11704 9648 11756 9654
rect 11704 9590 11756 9596
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11060 9512 11112 9518
rect 11060 9454 11112 9460
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 10782 9344 10838 9353
rect 10782 9279 10838 9288
rect 10232 9172 10284 9178
rect 10232 9114 10284 9120
rect 10416 9172 10468 9178
rect 10416 9114 10468 9120
rect 10692 8968 10744 8974
rect 10692 8910 10744 8916
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 9956 8016 10008 8022
rect 9956 7958 10008 7964
rect 9876 7806 10272 7834
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 9862 7032 9918 7041
rect 9862 6967 9918 6976
rect 9494 6287 9550 6296
rect 9692 6310 9812 6338
rect 9508 5642 9536 6287
rect 9496 5636 9548 5642
rect 9496 5578 9548 5584
rect 9416 5086 9628 5114
rect 9496 5024 9548 5030
rect 9496 4966 9548 4972
rect 9310 4856 9366 4865
rect 9310 4791 9366 4800
rect 8668 4684 8720 4690
rect 8668 4626 8720 4632
rect 9140 4678 9260 4706
rect 8758 4584 8814 4593
rect 8758 4519 8814 4528
rect 8772 4214 8800 4519
rect 9140 4486 9168 4678
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 8760 4208 8812 4214
rect 8760 4150 8812 4156
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 8680 4049 8708 4082
rect 8666 4040 8722 4049
rect 8666 3975 8722 3984
rect 8680 3534 8708 3975
rect 9232 3913 9260 4558
rect 9324 4321 9352 4791
rect 9402 4584 9458 4593
rect 9402 4519 9404 4528
rect 9456 4519 9458 4528
rect 9404 4490 9456 4496
rect 9310 4312 9366 4321
rect 9310 4247 9366 4256
rect 9508 4146 9536 4966
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9218 3904 9274 3913
rect 8747 3836 9055 3856
rect 9218 3839 9274 3848
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3760 9055 3780
rect 9128 3732 9180 3738
rect 8956 3692 9128 3720
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8956 3398 8984 3692
rect 9128 3674 9180 3680
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 9036 3120 9088 3126
rect 9036 3062 9088 3068
rect 8576 2100 8628 2106
rect 8576 2042 8628 2048
rect 8392 1896 8444 1902
rect 8392 1838 8444 1844
rect 8298 1320 8354 1329
rect 8298 1255 8354 1264
rect 8680 950 8708 3062
rect 9048 2922 9076 3062
rect 9036 2916 9088 2922
rect 9036 2858 9088 2864
rect 8747 2748 9055 2768
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2672 9055 2692
rect 8944 2304 8996 2310
rect 8944 2246 8996 2252
rect 8956 1698 8984 2246
rect 8944 1692 8996 1698
rect 8944 1634 8996 1640
rect 8956 1601 8984 1634
rect 8942 1592 8998 1601
rect 8942 1527 8998 1536
rect 9140 1358 9168 3334
rect 9232 2632 9260 3470
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 9324 2774 9352 3402
rect 9600 3233 9628 5086
rect 9692 5012 9720 6310
rect 9772 5840 9824 5846
rect 9772 5782 9824 5788
rect 9784 5166 9812 5782
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 9692 4984 9812 5012
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 9586 3224 9642 3233
rect 9404 3188 9456 3194
rect 9586 3159 9642 3168
rect 9404 3130 9456 3136
rect 9416 3058 9444 3130
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9600 2961 9628 2994
rect 9586 2952 9642 2961
rect 9586 2887 9642 2896
rect 9692 2774 9720 3946
rect 9784 3942 9812 4984
rect 9772 3936 9824 3942
rect 9772 3878 9824 3884
rect 9876 3738 9904 6967
rect 9956 6724 10008 6730
rect 9956 6666 10008 6672
rect 9968 5098 9996 6666
rect 9956 5092 10008 5098
rect 9956 5034 10008 5040
rect 10048 4208 10100 4214
rect 10048 4150 10100 4156
rect 9954 4040 10010 4049
rect 9954 3975 10010 3984
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9772 3528 9824 3534
rect 9770 3496 9772 3505
rect 9824 3496 9826 3505
rect 9770 3431 9826 3440
rect 9968 3369 9996 3975
rect 9954 3360 10010 3369
rect 9954 3295 10010 3304
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 9324 2746 9628 2774
rect 9692 2746 9812 2774
rect 9600 2689 9628 2746
rect 9402 2680 9458 2689
rect 9232 2604 9352 2632
rect 9402 2615 9404 2624
rect 9218 2544 9274 2553
rect 9218 2479 9274 2488
rect 9128 1352 9180 1358
rect 9128 1294 9180 1300
rect 8668 944 8720 950
rect 8668 886 8720 892
rect 8680 800 8708 886
rect 9232 800 9260 2479
rect 9324 1018 9352 2604
rect 9456 2615 9458 2624
rect 9586 2680 9642 2689
rect 9586 2615 9642 2624
rect 9404 2586 9456 2592
rect 9784 2446 9812 2746
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 9416 1630 9444 2314
rect 9494 2136 9550 2145
rect 9494 2071 9550 2080
rect 9508 1630 9536 2071
rect 9692 1766 9720 2382
rect 9680 1760 9732 1766
rect 9680 1702 9732 1708
rect 9404 1624 9456 1630
rect 9404 1566 9456 1572
rect 9496 1624 9548 1630
rect 9496 1566 9548 1572
rect 9312 1012 9364 1018
rect 9312 954 9364 960
rect 9416 950 9444 1566
rect 9404 944 9456 950
rect 9404 886 9456 892
rect 9784 800 9812 2382
rect 9968 1562 9996 3062
rect 9956 1556 10008 1562
rect 9956 1498 10008 1504
rect 7932 672 7984 678
rect 7932 614 7984 620
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9218 0 9274 800
rect 9770 0 9826 800
rect 10060 762 10088 4150
rect 10152 3534 10180 7686
rect 10244 6440 10272 7806
rect 10336 6662 10364 8434
rect 10612 8022 10640 8434
rect 10508 8016 10560 8022
rect 10508 7958 10560 7964
rect 10600 8016 10652 8022
rect 10600 7958 10652 7964
rect 10324 6656 10376 6662
rect 10324 6598 10376 6604
rect 10416 6452 10468 6458
rect 10244 6412 10416 6440
rect 10336 5710 10364 6412
rect 10416 6394 10468 6400
rect 10520 6338 10548 7958
rect 10612 7546 10640 7958
rect 10704 7546 10732 8910
rect 10600 7540 10652 7546
rect 10600 7482 10652 7488
rect 10692 7540 10744 7546
rect 10692 7482 10744 7488
rect 10598 7440 10654 7449
rect 10598 7375 10654 7384
rect 10612 6497 10640 7375
rect 10598 6488 10654 6497
rect 10598 6423 10654 6432
rect 10796 6338 10824 9279
rect 11072 9042 11100 9454
rect 11624 9110 11652 9454
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 10966 8528 11022 8537
rect 10966 8463 11022 8472
rect 10980 8362 11008 8463
rect 11072 8430 11100 8978
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 11072 7818 11100 8366
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 11058 7712 11114 7721
rect 11058 7647 11114 7656
rect 10968 7404 11020 7410
rect 10968 7346 11020 7352
rect 10980 6934 11008 7346
rect 11072 7206 11100 7647
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 10980 6662 11008 6870
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 11164 6458 11192 8774
rect 11346 8732 11654 8752
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8656 11654 8676
rect 11242 8528 11298 8537
rect 11242 8463 11298 8472
rect 11256 7546 11284 8463
rect 11346 7644 11654 7664
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7568 11654 7588
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11336 7268 11388 7274
rect 11336 7210 11388 7216
rect 11348 6934 11376 7210
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11348 6746 11376 6870
rect 11256 6718 11376 6746
rect 11152 6452 11204 6458
rect 11152 6394 11204 6400
rect 11060 6384 11112 6390
rect 10428 6310 10548 6338
rect 10612 6310 10824 6338
rect 11058 6352 11060 6361
rect 11112 6352 11114 6361
rect 10428 6089 10456 6310
rect 10612 6254 10640 6310
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10414 6080 10470 6089
rect 10414 6015 10470 6024
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10232 4480 10284 4486
rect 10232 4422 10284 4428
rect 10244 3602 10272 4422
rect 10232 3596 10284 3602
rect 10232 3538 10284 3544
rect 10140 3528 10192 3534
rect 10140 3470 10192 3476
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10244 2922 10272 2994
rect 10232 2916 10284 2922
rect 10232 2858 10284 2864
rect 10428 2514 10456 6015
rect 10520 5234 10548 6122
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10612 5642 10640 5850
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10704 5302 10732 6310
rect 11256 6322 11284 6718
rect 11346 6556 11654 6576
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6480 11654 6500
rect 11058 6287 11114 6296
rect 11244 6316 11296 6322
rect 11244 6258 11296 6264
rect 11716 6254 11744 9590
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10876 6248 10928 6254
rect 10876 6190 10928 6196
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 10796 5914 10824 6190
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10888 5778 10916 6190
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10876 5772 10928 5778
rect 10876 5714 10928 5720
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10600 5228 10652 5234
rect 10600 5170 10652 5176
rect 10612 4826 10640 5170
rect 10888 5166 10916 5714
rect 10980 5166 11008 6054
rect 11244 5636 11296 5642
rect 11244 5578 11296 5584
rect 11256 5234 11284 5578
rect 11808 5522 11836 10678
rect 11900 9330 11928 14214
rect 11992 12714 12020 14894
rect 12084 13172 12112 15014
rect 12176 13326 12204 15370
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12268 15162 12296 15302
rect 12256 15156 12308 15162
rect 12256 15098 12308 15104
rect 12360 14498 12388 18090
rect 12728 17882 12756 18226
rect 13372 17882 13400 20402
rect 13740 20346 13768 22200
rect 14186 21040 14242 21049
rect 14186 20975 14242 20984
rect 14200 20482 14228 20975
rect 14292 20618 14320 22200
rect 14844 22114 14872 22200
rect 14936 22114 14964 22222
rect 14844 22086 14964 22114
rect 14648 21344 14700 21350
rect 14648 21286 14700 21292
rect 14292 20590 14412 20618
rect 14384 20534 14412 20590
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14372 20528 14424 20534
rect 14200 20454 14320 20482
rect 14372 20470 14424 20476
rect 13740 20318 13860 20346
rect 13832 20262 13860 20318
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 12438 17504 12494 17513
rect 12438 17439 12494 17448
rect 12452 17270 12480 17439
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 13188 17202 13216 17682
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 12808 17060 12860 17066
rect 12808 17002 12860 17008
rect 12820 16794 12848 17002
rect 12808 16788 12860 16794
rect 12808 16730 12860 16736
rect 13188 16726 13216 17138
rect 13176 16720 13228 16726
rect 13176 16662 13228 16668
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12452 15706 12480 16050
rect 12532 15904 12584 15910
rect 12532 15846 12584 15852
rect 12440 15700 12492 15706
rect 12440 15642 12492 15648
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12268 14470 12388 14498
rect 12268 14346 12296 14470
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 12360 14006 12388 14350
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12452 13530 12480 15030
rect 12544 15026 12572 15846
rect 13464 15416 13492 20198
rect 13945 20156 14253 20176
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20080 14253 20100
rect 13728 19712 13780 19718
rect 13728 19654 13780 19660
rect 13820 19712 13872 19718
rect 13820 19654 13872 19660
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13542 19136 13598 19145
rect 13542 19071 13598 19080
rect 13556 18766 13584 19071
rect 13544 18760 13596 18766
rect 13544 18702 13596 18708
rect 13648 18426 13676 19314
rect 13740 18766 13768 19654
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13636 18420 13688 18426
rect 13636 18362 13688 18368
rect 13544 17808 13596 17814
rect 13544 17750 13596 17756
rect 13556 17542 13584 17750
rect 13832 17678 13860 19654
rect 13945 19068 14253 19088
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 18992 14253 19012
rect 14292 18290 14320 20454
rect 14476 19446 14504 20538
rect 14464 19440 14516 19446
rect 14464 19382 14516 19388
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14556 19168 14608 19174
rect 14556 19110 14608 19116
rect 14384 18834 14412 19110
rect 14568 18902 14596 19110
rect 14556 18896 14608 18902
rect 14462 18864 14518 18873
rect 14372 18828 14424 18834
rect 14556 18838 14608 18844
rect 14462 18799 14518 18808
rect 14372 18770 14424 18776
rect 14476 18630 14504 18799
rect 14464 18624 14516 18630
rect 14464 18566 14516 18572
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14384 18057 14412 18158
rect 14370 18048 14426 18057
rect 13945 17980 14253 18000
rect 14370 17983 14426 17992
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17904 14253 17924
rect 14280 17740 14332 17746
rect 14280 17682 14332 17688
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13636 17604 13688 17610
rect 13636 17546 13688 17552
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13556 16046 13584 16390
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13648 15638 13676 17546
rect 14292 17202 14320 17682
rect 14476 17626 14504 18566
rect 14384 17598 14504 17626
rect 14556 17672 14608 17678
rect 14556 17614 14608 17620
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13726 16824 13782 16833
rect 13726 16759 13782 16768
rect 13740 16250 13768 16759
rect 13728 16244 13780 16250
rect 13728 16186 13780 16192
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 13726 15600 13782 15609
rect 13832 15570 13860 16934
rect 13945 16892 14253 16912
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16816 14253 16836
rect 14384 16833 14412 17598
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14370 16824 14426 16833
rect 14370 16759 14426 16768
rect 14384 16454 14412 16759
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 13924 15978 13952 16390
rect 14372 16108 14424 16114
rect 14372 16050 14424 16056
rect 13912 15972 13964 15978
rect 13912 15914 13964 15920
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 13945 15804 14253 15824
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15728 14253 15748
rect 14004 15632 14056 15638
rect 14004 15574 14056 15580
rect 13726 15535 13782 15544
rect 13820 15564 13872 15570
rect 13544 15428 13596 15434
rect 13464 15388 13544 15416
rect 13544 15370 13596 15376
rect 12622 15192 12678 15201
rect 12622 15127 12678 15136
rect 12532 15020 12584 15026
rect 12532 14962 12584 14968
rect 12636 14056 12664 15127
rect 13268 14952 13320 14958
rect 13266 14920 13268 14929
rect 13320 14920 13322 14929
rect 13266 14855 13322 14864
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 12544 14028 12664 14056
rect 12992 14068 13044 14074
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 12348 13184 12400 13190
rect 12084 13144 12204 13172
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 11980 12708 12032 12714
rect 11980 12650 12032 12656
rect 12084 12442 12112 12718
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12176 12170 12204 13144
rect 12348 13126 12400 13132
rect 12360 12850 12388 13126
rect 12544 12918 12572 14028
rect 12992 14010 13044 14016
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12636 12918 12664 13874
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12728 13530 12756 13670
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12912 13394 12940 13670
rect 13004 13394 13032 14010
rect 13358 13560 13414 13569
rect 13358 13495 13414 13504
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12820 12986 12848 13126
rect 12808 12980 12860 12986
rect 12808 12922 12860 12928
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12624 12912 12676 12918
rect 12624 12854 12676 12860
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 13004 12782 13032 13330
rect 13372 13025 13400 13495
rect 13648 13433 13676 14758
rect 13740 14657 13768 15535
rect 13820 15506 13872 15512
rect 13832 15366 13860 15506
rect 13820 15360 13872 15366
rect 13820 15302 13872 15308
rect 14016 15026 14044 15574
rect 14292 15094 14320 15846
rect 14280 15088 14332 15094
rect 14280 15030 14332 15036
rect 14004 15020 14056 15026
rect 14004 14962 14056 14968
rect 14384 14906 14412 16050
rect 14476 15706 14504 17478
rect 14568 17338 14596 17614
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14568 16726 14596 17274
rect 14556 16720 14608 16726
rect 14556 16662 14608 16668
rect 14556 16448 14608 16454
rect 14556 16390 14608 16396
rect 14464 15700 14516 15706
rect 14464 15642 14516 15648
rect 14464 15564 14516 15570
rect 14464 15506 14516 15512
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 14292 14878 14412 14906
rect 13726 14648 13782 14657
rect 13726 14583 13782 14592
rect 13832 14346 13860 14826
rect 13945 14716 14253 14736
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14640 14253 14660
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 14016 14278 14044 14486
rect 14188 14476 14240 14482
rect 14292 14464 14320 14878
rect 14372 14816 14424 14822
rect 14372 14758 14424 14764
rect 14384 14482 14412 14758
rect 14240 14436 14320 14464
rect 14372 14476 14424 14482
rect 14188 14418 14240 14424
rect 14372 14418 14424 14424
rect 14096 14340 14148 14346
rect 14096 14282 14148 14288
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 14108 13870 14136 14282
rect 13728 13864 13780 13870
rect 13728 13806 13780 13812
rect 14096 13864 14148 13870
rect 14096 13806 14148 13812
rect 13634 13424 13690 13433
rect 13634 13359 13690 13368
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13358 13016 13414 13025
rect 13358 12951 13414 12960
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 12992 12776 13044 12782
rect 12992 12718 13044 12724
rect 13372 12646 13400 12786
rect 13544 12776 13596 12782
rect 13542 12744 13544 12753
rect 13596 12744 13598 12753
rect 13542 12679 13598 12688
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 12164 12164 12216 12170
rect 12164 12106 12216 12112
rect 12440 12164 12492 12170
rect 12440 12106 12492 12112
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11992 9654 12020 11698
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12256 10736 12308 10742
rect 12256 10678 12308 10684
rect 12084 10198 12112 10678
rect 12072 10192 12124 10198
rect 12072 10134 12124 10140
rect 12268 10130 12296 10678
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 12360 10305 12388 10610
rect 12346 10296 12402 10305
rect 12346 10231 12402 10240
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12164 9988 12216 9994
rect 12164 9930 12216 9936
rect 12072 9716 12124 9722
rect 12072 9658 12124 9664
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 11900 9302 12020 9330
rect 11992 8498 12020 9302
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 12084 8430 12112 9658
rect 12176 9194 12204 9930
rect 12268 9586 12296 10066
rect 12452 9654 12480 12106
rect 13542 11928 13598 11937
rect 13542 11863 13598 11872
rect 13556 11665 13584 11863
rect 13542 11656 13598 11665
rect 13542 11591 13598 11600
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13096 11218 13124 11494
rect 13648 11354 13676 13262
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13084 11212 13136 11218
rect 13084 11154 13136 11160
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12728 10266 12756 10950
rect 12820 10810 12848 10950
rect 12808 10804 12860 10810
rect 12808 10746 12860 10752
rect 12808 10532 12860 10538
rect 12808 10474 12860 10480
rect 12820 10441 12848 10474
rect 12806 10432 12862 10441
rect 12806 10367 12862 10376
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 13004 9722 13032 9862
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 13096 9586 13124 11154
rect 13740 11150 13768 13806
rect 14200 13802 14228 14418
rect 14476 14362 14504 15506
rect 14568 15366 14596 16390
rect 14556 15360 14608 15366
rect 14556 15302 14608 15308
rect 14568 15026 14596 15302
rect 14556 15020 14608 15026
rect 14556 14962 14608 14968
rect 14660 14906 14688 21286
rect 15120 20380 15148 22222
rect 15382 22200 15438 23000
rect 15934 22200 15990 23000
rect 16486 22200 16542 23000
rect 17038 22200 17094 23000
rect 17682 22200 17738 23000
rect 18234 22200 18290 23000
rect 18694 22264 18750 22273
rect 15290 20632 15346 20641
rect 15396 20602 15424 22200
rect 15842 21584 15898 21593
rect 15842 21519 15898 21528
rect 15856 21049 15884 21519
rect 15842 21040 15898 21049
rect 15842 20975 15898 20984
rect 15290 20567 15346 20576
rect 15384 20596 15436 20602
rect 15304 20534 15332 20567
rect 15384 20538 15436 20544
rect 15292 20528 15344 20534
rect 15292 20470 15344 20476
rect 15750 20496 15806 20505
rect 15750 20431 15752 20440
rect 15804 20431 15806 20440
rect 15752 20402 15804 20408
rect 15292 20392 15344 20398
rect 15120 20352 15292 20380
rect 15292 20334 15344 20340
rect 15198 20088 15254 20097
rect 15948 20058 15976 22200
rect 16500 20890 16528 22200
rect 16946 21312 17002 21321
rect 16946 21247 17002 21256
rect 16408 20862 16528 20890
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 15198 20023 15254 20032
rect 15936 20052 15988 20058
rect 15014 19952 15070 19961
rect 14832 19916 14884 19922
rect 15014 19887 15070 19896
rect 14832 19858 14884 19864
rect 14844 19378 14872 19858
rect 15028 19854 15056 19887
rect 15016 19848 15068 19854
rect 15016 19790 15068 19796
rect 15108 19848 15160 19854
rect 15108 19790 15160 19796
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14924 18624 14976 18630
rect 14924 18566 14976 18572
rect 15016 18624 15068 18630
rect 15016 18566 15068 18572
rect 14936 18426 14964 18566
rect 14924 18420 14976 18426
rect 14924 18362 14976 18368
rect 14924 18284 14976 18290
rect 14924 18226 14976 18232
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14844 16658 14872 17478
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14740 16584 14792 16590
rect 14740 16526 14792 16532
rect 14752 15570 14780 16526
rect 14936 15994 14964 18226
rect 15028 16454 15056 18566
rect 15120 18222 15148 19790
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15108 17808 15160 17814
rect 15108 17750 15160 17756
rect 15120 17270 15148 17750
rect 15108 17264 15160 17270
rect 15108 17206 15160 17212
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 14936 15966 15056 15994
rect 14924 15904 14976 15910
rect 14924 15846 14976 15852
rect 14830 15736 14886 15745
rect 14830 15671 14886 15680
rect 14740 15564 14792 15570
rect 14740 15506 14792 15512
rect 14844 15201 14872 15671
rect 14936 15570 14964 15846
rect 14924 15564 14976 15570
rect 14924 15506 14976 15512
rect 14830 15192 14886 15201
rect 14830 15127 14886 15136
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14384 14334 14504 14362
rect 14568 14878 14688 14906
rect 14278 14240 14334 14249
rect 14278 14175 14334 14184
rect 14292 14074 14320 14175
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 14188 13796 14240 13802
rect 14188 13738 14240 13744
rect 13945 13628 14253 13648
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13552 14253 13572
rect 14280 13456 14332 13462
rect 14280 13398 14332 13404
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13832 11898 13860 12582
rect 13945 12540 14253 12560
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12464 14253 12484
rect 14292 12170 14320 13398
rect 14280 12164 14332 12170
rect 14280 12106 14332 12112
rect 13912 12096 13964 12102
rect 13912 12038 13964 12044
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13924 11778 13952 12038
rect 13832 11750 13952 11778
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13832 10606 13860 11750
rect 14384 11665 14412 14334
rect 14464 14272 14516 14278
rect 14464 14214 14516 14220
rect 14476 14074 14504 14214
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14568 13546 14596 14878
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14476 13518 14596 13546
rect 14476 13190 14504 13518
rect 14660 13394 14688 14758
rect 14752 14249 14780 14962
rect 14832 14272 14884 14278
rect 14738 14240 14794 14249
rect 14832 14214 14884 14220
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14738 14175 14794 14184
rect 14740 13932 14792 13938
rect 14740 13874 14792 13880
rect 14648 13388 14700 13394
rect 14648 13330 14700 13336
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14464 13184 14516 13190
rect 14464 13126 14516 13132
rect 14568 12986 14596 13262
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14554 12744 14610 12753
rect 14554 12679 14556 12688
rect 14608 12679 14610 12688
rect 14556 12650 14608 12656
rect 14660 12434 14688 13126
rect 14752 12782 14780 13874
rect 14844 13394 14872 14214
rect 14936 14074 14964 14214
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 15028 13818 15056 15966
rect 15120 15366 15148 17206
rect 15212 16794 15240 20023
rect 15936 19994 15988 20000
rect 15658 19952 15714 19961
rect 15658 19887 15714 19896
rect 15292 19712 15344 19718
rect 15672 19689 15700 19887
rect 16224 19854 16252 20742
rect 16408 20602 16436 20862
rect 16544 20700 16852 20720
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20624 16852 20644
rect 16396 20596 16448 20602
rect 16396 20538 16448 20544
rect 16960 20466 16988 21247
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 17052 20330 17080 22200
rect 17592 21072 17644 21078
rect 17592 21014 17644 21020
rect 17132 21004 17184 21010
rect 17132 20946 17184 20952
rect 17040 20324 17092 20330
rect 17040 20266 17092 20272
rect 16120 19848 16172 19854
rect 16120 19790 16172 19796
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 15752 19712 15804 19718
rect 15292 19654 15344 19660
rect 15658 19680 15714 19689
rect 15304 18358 15332 19654
rect 15752 19654 15804 19660
rect 15658 19615 15714 19624
rect 15384 19440 15436 19446
rect 15384 19382 15436 19388
rect 15396 18766 15424 19382
rect 15384 18760 15436 18766
rect 15384 18702 15436 18708
rect 15566 18728 15622 18737
rect 15476 18692 15528 18698
rect 15764 18698 15792 19654
rect 16132 19514 16160 19790
rect 16948 19780 17000 19786
rect 16948 19722 17000 19728
rect 16544 19612 16852 19632
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19536 16852 19556
rect 16120 19508 16172 19514
rect 16120 19450 16172 19456
rect 16960 18970 16988 19722
rect 17038 19544 17094 19553
rect 17038 19479 17094 19488
rect 17052 19378 17080 19479
rect 17144 19378 17172 20946
rect 17224 20936 17276 20942
rect 17224 20878 17276 20884
rect 17236 20466 17264 20878
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 17604 20380 17632 21014
rect 17696 20534 17724 22200
rect 17866 21584 17922 21593
rect 17866 21519 17922 21528
rect 17774 21448 17830 21457
rect 17774 21383 17830 21392
rect 17684 20528 17736 20534
rect 17684 20470 17736 20476
rect 17604 20352 17724 20380
rect 17500 19916 17552 19922
rect 17500 19858 17552 19864
rect 17314 19680 17370 19689
rect 17314 19615 17370 19624
rect 17328 19514 17356 19615
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 17132 19372 17184 19378
rect 17132 19314 17184 19320
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16120 18760 16172 18766
rect 17224 18760 17276 18766
rect 16120 18702 16172 18708
rect 15566 18663 15622 18672
rect 15752 18692 15804 18698
rect 15476 18634 15528 18640
rect 15488 18426 15516 18634
rect 15476 18420 15528 18426
rect 15476 18362 15528 18368
rect 15292 18352 15344 18358
rect 15292 18294 15344 18300
rect 15474 17640 15530 17649
rect 15474 17575 15530 17584
rect 15290 17096 15346 17105
rect 15290 17031 15346 17040
rect 15200 16788 15252 16794
rect 15200 16730 15252 16736
rect 15304 16130 15332 17031
rect 15212 16102 15332 16130
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15120 13870 15148 15302
rect 14936 13790 15056 13818
rect 15108 13864 15160 13870
rect 15108 13806 15160 13812
rect 14832 13388 14884 13394
rect 14832 13330 14884 13336
rect 14936 13190 14964 13790
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 15028 13326 15056 13670
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 15212 12986 15240 16102
rect 15290 16008 15346 16017
rect 15290 15943 15346 15952
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15108 12912 15160 12918
rect 15108 12854 15160 12860
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 15016 12776 15068 12782
rect 15016 12718 15068 12724
rect 14832 12708 14884 12714
rect 14832 12650 14884 12656
rect 14476 12406 14688 12434
rect 14370 11656 14426 11665
rect 14370 11591 14426 11600
rect 13945 11452 14253 11472
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11376 14253 11396
rect 14280 11144 14332 11150
rect 14280 11086 14332 11092
rect 13268 10600 13320 10606
rect 13268 10542 13320 10548
rect 13820 10600 13872 10606
rect 13820 10542 13872 10548
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 12176 9166 12296 9194
rect 12164 9036 12216 9042
rect 12164 8978 12216 8984
rect 12176 8498 12204 8978
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 11888 8356 11940 8362
rect 11888 8298 11940 8304
rect 11900 6458 11928 8298
rect 11978 7576 12034 7585
rect 11978 7511 12034 7520
rect 11992 7313 12020 7511
rect 11978 7304 12034 7313
rect 11978 7239 12034 7248
rect 11980 6724 12032 6730
rect 11980 6666 12032 6672
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11716 5494 11836 5522
rect 11346 5468 11654 5488
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5392 11654 5412
rect 11244 5228 11296 5234
rect 11244 5170 11296 5176
rect 10876 5160 10928 5166
rect 10876 5102 10928 5108
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10704 4486 10732 4558
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10968 4480 11020 4486
rect 10968 4422 11020 4428
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 10980 4214 11008 4422
rect 10968 4208 11020 4214
rect 10968 4150 11020 4156
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10508 3936 10560 3942
rect 10508 3878 10560 3884
rect 10520 3602 10548 3878
rect 10796 3738 10824 4082
rect 10980 4078 11008 4150
rect 11072 4146 11100 4422
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10508 3596 10560 3602
rect 10508 3538 10560 3544
rect 11072 3058 11100 3946
rect 11152 3528 11204 3534
rect 11256 3516 11284 5170
rect 11346 4380 11654 4400
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4304 11654 4324
rect 11716 3618 11744 5494
rect 11794 5400 11850 5409
rect 11794 5335 11850 5344
rect 11808 5001 11836 5335
rect 11794 4992 11850 5001
rect 11794 4927 11850 4936
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11900 4078 11928 4490
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11992 3913 12020 6666
rect 12084 4146 12112 8366
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12176 5710 12204 7754
rect 12268 6730 12296 9166
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 12348 8832 12400 8838
rect 13096 8809 13124 8842
rect 12348 8774 12400 8780
rect 13082 8800 13138 8809
rect 12360 7410 12388 8774
rect 13082 8735 13138 8744
rect 12806 8664 12862 8673
rect 12806 8599 12862 8608
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12346 7304 12402 7313
rect 12346 7239 12402 7248
rect 12360 7206 12388 7239
rect 12348 7200 12400 7206
rect 12348 7142 12400 7148
rect 12440 7200 12492 7206
rect 12440 7142 12492 7148
rect 12452 7041 12480 7142
rect 12438 7032 12494 7041
rect 12348 6996 12400 7002
rect 12438 6967 12494 6976
rect 12348 6938 12400 6944
rect 12360 6905 12388 6938
rect 12346 6896 12402 6905
rect 12346 6831 12402 6840
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12348 6724 12400 6730
rect 12348 6666 12400 6672
rect 12254 6624 12310 6633
rect 12254 6559 12310 6568
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12268 5574 12296 6559
rect 12256 5568 12308 5574
rect 12256 5510 12308 5516
rect 12162 4312 12218 4321
rect 12268 4282 12296 5510
rect 12360 5302 12388 6666
rect 12544 6458 12572 7686
rect 12636 7546 12664 8434
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12624 7540 12676 7546
rect 12624 7482 12676 7488
rect 12728 7206 12756 7822
rect 12820 7818 12848 8599
rect 13096 7954 13124 8735
rect 13084 7948 13136 7954
rect 13084 7890 13136 7896
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12532 6452 12584 6458
rect 12532 6394 12584 6400
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12348 5296 12400 5302
rect 12348 5238 12400 5244
rect 12360 4690 12388 5238
rect 12348 4684 12400 4690
rect 12348 4626 12400 4632
rect 12162 4247 12218 4256
rect 12256 4276 12308 4282
rect 12072 4140 12124 4146
rect 12072 4082 12124 4088
rect 11978 3904 12034 3913
rect 11978 3839 12034 3848
rect 11992 3641 12020 3839
rect 11624 3590 11744 3618
rect 11978 3632 12034 3641
rect 11624 3534 11652 3590
rect 11978 3567 12034 3576
rect 11204 3488 11284 3516
rect 11612 3528 11664 3534
rect 11152 3470 11204 3476
rect 11612 3470 11664 3476
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 11346 3292 11654 3312
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3216 11654 3236
rect 11716 3194 11744 3402
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11256 3058 11284 3130
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 11796 2848 11848 2854
rect 11796 2790 11848 2796
rect 11808 2650 11836 2790
rect 11796 2644 11848 2650
rect 11796 2586 11848 2592
rect 11704 2576 11756 2582
rect 11702 2544 11704 2553
rect 11756 2544 11758 2553
rect 10416 2508 10468 2514
rect 11702 2479 11758 2488
rect 10416 2450 10468 2456
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10980 1970 11008 2246
rect 10968 1964 11020 1970
rect 10968 1906 11020 1912
rect 11164 1766 11192 2382
rect 11346 2204 11654 2224
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2128 11654 2148
rect 10876 1760 10928 1766
rect 10876 1702 10928 1708
rect 11152 1760 11204 1766
rect 11152 1702 11204 1708
rect 10244 870 10364 898
rect 10244 762 10272 870
rect 10336 800 10364 870
rect 10888 800 10916 1702
rect 11428 1556 11480 1562
rect 11428 1498 11480 1504
rect 11440 800 11468 1498
rect 11900 1222 11928 2994
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 12084 1601 12112 2246
rect 12176 2038 12204 4247
rect 12256 4218 12308 4224
rect 12256 4072 12308 4078
rect 12256 4014 12308 4020
rect 12346 4040 12402 4049
rect 12268 3398 12296 4014
rect 12346 3975 12402 3984
rect 12360 3641 12388 3975
rect 12346 3632 12402 3641
rect 12346 3567 12402 3576
rect 12256 3392 12308 3398
rect 12256 3334 12308 3340
rect 12532 3392 12584 3398
rect 12532 3334 12584 3340
rect 12346 3224 12402 3233
rect 12346 3159 12402 3168
rect 12360 2922 12388 3159
rect 12544 3058 12572 3334
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12348 2916 12400 2922
rect 12348 2858 12400 2864
rect 12164 2032 12216 2038
rect 12164 1974 12216 1980
rect 12256 2032 12308 2038
rect 12256 1974 12308 1980
rect 12268 1698 12296 1974
rect 12256 1692 12308 1698
rect 12256 1634 12308 1640
rect 12070 1592 12126 1601
rect 12452 1562 12480 2926
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 12070 1527 12126 1536
rect 12440 1556 12492 1562
rect 12440 1498 12492 1504
rect 12072 1488 12124 1494
rect 12072 1430 12124 1436
rect 11888 1216 11940 1222
rect 11888 1158 11940 1164
rect 12084 800 12112 1430
rect 12544 1306 12572 2518
rect 12636 1465 12664 6258
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12728 5114 12756 5714
rect 12820 5574 12848 7754
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 12912 7002 12940 7278
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 13004 5778 13032 7686
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13096 6730 13124 6802
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13096 6458 13124 6666
rect 13188 6633 13216 6666
rect 13174 6624 13230 6633
rect 13174 6559 13230 6568
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13176 5840 13228 5846
rect 13176 5782 13228 5788
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12992 5568 13044 5574
rect 12992 5510 13044 5516
rect 12728 5086 12940 5114
rect 12912 5030 12940 5086
rect 12900 5024 12952 5030
rect 12900 4966 12952 4972
rect 12912 4146 12940 4966
rect 13004 4622 13032 5510
rect 12992 4616 13044 4622
rect 12992 4558 13044 4564
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13096 4282 13124 4422
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 12992 4208 13044 4214
rect 12992 4150 13044 4156
rect 12900 4140 12952 4146
rect 12900 4082 12952 4088
rect 12714 3768 12770 3777
rect 12714 3703 12716 3712
rect 12768 3703 12770 3712
rect 12716 3674 12768 3680
rect 12728 3126 12756 3674
rect 12900 3596 12952 3602
rect 12900 3538 12952 3544
rect 12808 3392 12860 3398
rect 12808 3334 12860 3340
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 12820 2825 12848 3334
rect 12912 2922 12940 3538
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 12806 2816 12862 2825
rect 12806 2751 12862 2760
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 12728 1970 12756 2382
rect 13004 2038 13032 4150
rect 13188 3602 13216 5782
rect 13280 4554 13308 10542
rect 14292 10470 14320 11086
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 13832 10266 13860 10406
rect 13945 10364 14253 10384
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10288 14253 10308
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13542 10160 13598 10169
rect 13542 10095 13544 10104
rect 13596 10095 13598 10104
rect 13544 10066 13596 10072
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 13726 9888 13782 9897
rect 13726 9823 13782 9832
rect 13636 9512 13688 9518
rect 13636 9454 13688 9460
rect 13544 9444 13596 9450
rect 13544 9386 13596 9392
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 8838 13492 9318
rect 13556 9110 13584 9386
rect 13544 9104 13596 9110
rect 13544 9046 13596 9052
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13450 7712 13506 7721
rect 13450 7647 13506 7656
rect 13464 7449 13492 7647
rect 13450 7440 13506 7449
rect 13450 7375 13506 7384
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 13372 6798 13400 7142
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13450 6624 13506 6633
rect 13450 6559 13506 6568
rect 13360 6384 13412 6390
rect 13464 6361 13492 6559
rect 13360 6326 13412 6332
rect 13450 6352 13506 6361
rect 13372 6089 13400 6326
rect 13450 6287 13506 6296
rect 13452 6112 13504 6118
rect 13358 6080 13414 6089
rect 13452 6054 13504 6060
rect 13358 6015 13414 6024
rect 13358 5536 13414 5545
rect 13358 5471 13414 5480
rect 13268 4548 13320 4554
rect 13268 4490 13320 4496
rect 13372 4060 13400 5471
rect 13464 4214 13492 6054
rect 13556 4758 13584 8434
rect 13648 8090 13676 9454
rect 13740 9353 13768 9823
rect 14016 9518 14044 9998
rect 14292 9926 14320 10406
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14384 9738 14412 11591
rect 14476 10169 14504 12406
rect 14646 12064 14702 12073
rect 14646 11999 14702 12008
rect 14554 10296 14610 10305
rect 14554 10231 14610 10240
rect 14462 10160 14518 10169
rect 14568 10130 14596 10231
rect 14462 10095 14518 10104
rect 14556 10124 14608 10130
rect 14476 9926 14504 10095
rect 14556 10066 14608 10072
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14568 9738 14596 9862
rect 14384 9722 14596 9738
rect 14384 9716 14608 9722
rect 14384 9710 14556 9716
rect 14556 9658 14608 9664
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 13820 9376 13872 9382
rect 13726 9344 13782 9353
rect 13820 9318 13872 9324
rect 13726 9279 13782 9288
rect 13726 9208 13782 9217
rect 13726 9143 13782 9152
rect 13740 9042 13768 9143
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13728 8356 13780 8362
rect 13728 8298 13780 8304
rect 13636 8084 13688 8090
rect 13636 8026 13688 8032
rect 13648 7546 13676 8026
rect 13740 7818 13768 8298
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13726 7440 13782 7449
rect 13726 7375 13782 7384
rect 13634 6896 13690 6905
rect 13634 6831 13690 6840
rect 13648 6458 13676 6831
rect 13636 6452 13688 6458
rect 13636 6394 13688 6400
rect 13740 5953 13768 7375
rect 13726 5944 13782 5953
rect 13726 5879 13782 5888
rect 13740 5710 13768 5879
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 13648 4264 13676 5238
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13556 4236 13676 4264
rect 13452 4208 13504 4214
rect 13452 4150 13504 4156
rect 13280 4032 13400 4060
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13082 3360 13138 3369
rect 13082 3295 13138 3304
rect 13096 3126 13124 3295
rect 13084 3120 13136 3126
rect 13084 3062 13136 3068
rect 12992 2032 13044 2038
rect 12992 1974 13044 1980
rect 12716 1964 12768 1970
rect 12716 1906 12768 1912
rect 13096 1902 13124 3062
rect 13280 2938 13308 4032
rect 13358 3904 13414 3913
rect 13358 3839 13414 3848
rect 13372 3534 13400 3839
rect 13556 3534 13584 4236
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13188 2910 13308 2938
rect 13188 2310 13216 2910
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 13280 2446 13308 2790
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 13372 2106 13400 2246
rect 13360 2100 13412 2106
rect 13360 2042 13412 2048
rect 13084 1896 13136 1902
rect 13084 1838 13136 1844
rect 13176 1488 13228 1494
rect 12622 1456 12678 1465
rect 13176 1430 13228 1436
rect 12622 1391 12678 1400
rect 12544 1278 12664 1306
rect 12636 800 12664 1278
rect 13188 800 13216 1430
rect 13648 1170 13676 4082
rect 13740 3738 13768 5170
rect 13728 3732 13780 3738
rect 13728 3674 13780 3680
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13740 2446 13768 3334
rect 13832 2689 13860 9318
rect 13945 9276 14253 9296
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9200 14253 9220
rect 14292 9160 14320 9522
rect 14384 9178 14412 9590
rect 14660 9568 14688 11999
rect 14740 11824 14792 11830
rect 14740 11766 14792 11772
rect 14752 10577 14780 11766
rect 14844 11354 14872 12650
rect 14832 11348 14884 11354
rect 14832 11290 14884 11296
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 14936 10742 14964 11290
rect 15028 10810 15056 12718
rect 15120 12442 15148 12854
rect 15108 12436 15160 12442
rect 15108 12378 15160 12384
rect 15200 12232 15252 12238
rect 15200 12174 15252 12180
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 15120 11150 15148 11630
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 14924 10736 14976 10742
rect 14924 10678 14976 10684
rect 15212 10606 15240 12174
rect 15304 10810 15332 15943
rect 15488 14958 15516 17575
rect 15580 16590 15608 18663
rect 15752 18634 15804 18640
rect 16028 18284 16080 18290
rect 16028 18226 16080 18232
rect 15660 16992 15712 16998
rect 15660 16934 15712 16940
rect 15568 16584 15620 16590
rect 15568 16526 15620 16532
rect 15568 16448 15620 16454
rect 15672 16436 15700 16934
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 15844 16720 15896 16726
rect 15844 16662 15896 16668
rect 15620 16408 15700 16436
rect 15568 16390 15620 16396
rect 15580 16017 15608 16390
rect 15750 16144 15806 16153
rect 15750 16079 15806 16088
rect 15566 16008 15622 16017
rect 15566 15943 15622 15952
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15568 14884 15620 14890
rect 15568 14826 15620 14832
rect 15580 14482 15608 14826
rect 15568 14476 15620 14482
rect 15568 14418 15620 14424
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15488 14006 15516 14214
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15476 14000 15528 14006
rect 15476 13942 15528 13948
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15488 12986 15516 13806
rect 15580 13297 15608 14010
rect 15566 13288 15622 13297
rect 15672 13258 15700 15370
rect 15566 13223 15622 13232
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15476 12368 15528 12374
rect 15396 12328 15476 12356
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15200 10600 15252 10606
rect 14738 10568 14794 10577
rect 15200 10542 15252 10548
rect 14738 10503 14794 10512
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14568 9540 14688 9568
rect 14462 9208 14518 9217
rect 14108 9132 14320 9160
rect 14372 9172 14424 9178
rect 14002 8664 14058 8673
rect 14002 8599 14058 8608
rect 14016 8362 14044 8599
rect 14004 8356 14056 8362
rect 14004 8298 14056 8304
rect 14108 8276 14136 9132
rect 14462 9143 14518 9152
rect 14372 9114 14424 9120
rect 14476 9110 14504 9143
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14292 8378 14320 8910
rect 14372 8832 14424 8838
rect 14370 8800 14372 8809
rect 14464 8832 14516 8838
rect 14424 8800 14426 8809
rect 14464 8774 14516 8780
rect 14370 8735 14426 8744
rect 14370 8664 14426 8673
rect 14370 8599 14426 8608
rect 14384 8498 14412 8599
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14292 8350 14412 8378
rect 14108 8248 14320 8276
rect 14384 8265 14412 8350
rect 13945 8188 14253 8208
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8112 14253 8132
rect 14188 7812 14240 7818
rect 14188 7754 14240 7760
rect 14200 7342 14228 7754
rect 14188 7336 14240 7342
rect 14188 7278 14240 7284
rect 14292 7154 14320 8248
rect 14370 8256 14426 8265
rect 14370 8191 14426 8200
rect 14476 7954 14504 8774
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14370 7168 14426 7177
rect 14292 7126 14370 7154
rect 13945 7100 14253 7120
rect 14370 7103 14426 7112
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7024 14253 7044
rect 14372 6452 14424 6458
rect 14372 6394 14424 6400
rect 14384 6089 14412 6394
rect 14568 6361 14596 9540
rect 14752 9466 14780 9998
rect 15200 9920 15252 9926
rect 15198 9888 15200 9897
rect 15252 9888 15254 9897
rect 15198 9823 15254 9832
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 14660 9438 14780 9466
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14660 7478 14688 9438
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14752 8022 14780 9318
rect 14844 8090 14872 9454
rect 15120 9432 15148 9658
rect 15304 9518 15332 10610
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15120 9404 15220 9432
rect 15192 9364 15220 9404
rect 15028 9336 15220 9364
rect 15292 9376 15344 9382
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 14740 8016 14792 8022
rect 14740 7958 14792 7964
rect 14936 7478 14964 8366
rect 15028 7546 15056 9336
rect 15292 9318 15344 9324
rect 15304 7970 15332 9318
rect 15396 9178 15424 12328
rect 15476 12310 15528 12316
rect 15672 11558 15700 13194
rect 15764 12986 15792 16079
rect 15752 12980 15804 12986
rect 15752 12922 15804 12928
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15488 9194 15516 11086
rect 15568 10532 15620 10538
rect 15568 10474 15620 10480
rect 15580 10266 15608 10474
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15384 9172 15436 9178
rect 15488 9166 15525 9194
rect 15384 9114 15436 9120
rect 15497 9058 15525 9166
rect 15488 9030 15525 9058
rect 15488 9024 15516 9030
rect 15396 8996 15516 9024
rect 15396 8090 15424 8996
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15212 7942 15332 7970
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15120 7585 15148 7822
rect 15212 7818 15240 7942
rect 15292 7880 15344 7886
rect 15292 7822 15344 7828
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15106 7576 15162 7585
rect 15016 7540 15068 7546
rect 15106 7511 15162 7520
rect 15016 7482 15068 7488
rect 14648 7472 14700 7478
rect 14648 7414 14700 7420
rect 14924 7472 14976 7478
rect 14924 7414 14976 7420
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14646 6896 14702 6905
rect 14844 6866 14872 7278
rect 14646 6831 14648 6840
rect 14700 6831 14702 6840
rect 14832 6860 14884 6866
rect 14648 6802 14700 6808
rect 14832 6802 14884 6808
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14752 6458 14780 6598
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14844 6390 14872 6802
rect 14648 6384 14700 6390
rect 14554 6352 14610 6361
rect 14832 6384 14884 6390
rect 14648 6326 14700 6332
rect 14738 6352 14794 6361
rect 14554 6287 14610 6296
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14554 6216 14610 6225
rect 14370 6080 14426 6089
rect 13945 6012 14253 6032
rect 14370 6015 14426 6024
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5936 14253 5956
rect 14280 5908 14332 5914
rect 14280 5850 14332 5856
rect 14292 5574 14320 5850
rect 14372 5772 14424 5778
rect 14372 5714 14424 5720
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 13945 4924 14253 4944
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4848 14253 4868
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14186 4584 14242 4593
rect 14108 4321 14136 4558
rect 14186 4519 14242 4528
rect 14094 4312 14150 4321
rect 14200 4282 14228 4519
rect 14292 4486 14320 5510
rect 14384 5370 14412 5714
rect 14372 5364 14424 5370
rect 14372 5306 14424 5312
rect 14384 5030 14412 5306
rect 14476 5302 14504 6190
rect 14554 6151 14610 6160
rect 14568 5574 14596 6151
rect 14660 5914 14688 6326
rect 14832 6326 14884 6332
rect 14936 6322 14964 7414
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 15014 7168 15070 7177
rect 15014 7103 15070 7112
rect 15028 6662 15056 7103
rect 15120 7002 15148 7346
rect 15108 6996 15160 7002
rect 15108 6938 15160 6944
rect 15200 6724 15252 6730
rect 15304 6712 15332 7822
rect 15252 6684 15332 6712
rect 15200 6666 15252 6672
rect 15016 6656 15068 6662
rect 15016 6598 15068 6604
rect 15198 6488 15254 6497
rect 15198 6423 15254 6432
rect 15212 6322 15240 6423
rect 14738 6287 14794 6296
rect 14924 6316 14976 6322
rect 14648 5908 14700 5914
rect 14648 5850 14700 5856
rect 14752 5794 14780 6287
rect 14924 6258 14976 6264
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 14660 5766 14780 5794
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14464 5296 14516 5302
rect 14464 5238 14516 5244
rect 14476 5166 14504 5238
rect 14464 5160 14516 5166
rect 14464 5102 14516 5108
rect 14372 5024 14424 5030
rect 14372 4966 14424 4972
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14094 4247 14150 4256
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14280 4072 14332 4078
rect 14280 4014 14332 4020
rect 14462 4040 14518 4049
rect 13945 3836 14253 3856
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3760 14253 3780
rect 14096 3664 14148 3670
rect 14096 3606 14148 3612
rect 13910 3088 13966 3097
rect 14108 3074 14136 3606
rect 14292 3194 14320 4014
rect 14372 4004 14424 4010
rect 14462 3975 14518 3984
rect 14372 3946 14424 3952
rect 14384 3738 14412 3946
rect 14476 3942 14504 3975
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14372 3732 14424 3738
rect 14372 3674 14424 3680
rect 14660 3618 14688 5766
rect 15016 5568 15068 5574
rect 15016 5510 15068 5516
rect 15028 4554 15056 5510
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 15382 5264 15438 5273
rect 15212 4690 15240 5238
rect 15382 5199 15438 5208
rect 15396 5001 15424 5199
rect 15382 4992 15438 5001
rect 15382 4927 15438 4936
rect 15476 4752 15528 4758
rect 15476 4694 15528 4700
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 14740 4548 14792 4554
rect 14740 4490 14792 4496
rect 15016 4548 15068 4554
rect 15016 4490 15068 4496
rect 14568 3590 14688 3618
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14108 3046 14412 3074
rect 13910 3023 13912 3032
rect 13964 3023 13966 3032
rect 13912 2994 13964 3000
rect 13945 2748 14253 2768
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13818 2680 13874 2689
rect 13945 2672 14253 2692
rect 13818 2615 13874 2624
rect 13728 2440 13780 2446
rect 13728 2382 13780 2388
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 14280 2304 14332 2310
rect 14280 2246 14332 2252
rect 13740 2038 13768 2246
rect 14292 2106 14320 2246
rect 14280 2100 14332 2106
rect 14280 2042 14332 2048
rect 13728 2032 13780 2038
rect 13728 1974 13780 1980
rect 14384 1170 14412 3046
rect 14464 2984 14516 2990
rect 14568 2972 14596 3590
rect 14752 3534 14780 4490
rect 15212 4010 15240 4626
rect 15290 4448 15346 4457
rect 15290 4383 15346 4392
rect 15304 4282 15332 4383
rect 15292 4276 15344 4282
rect 15292 4218 15344 4224
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15200 4004 15252 4010
rect 15200 3946 15252 3952
rect 15108 3936 15160 3942
rect 15108 3878 15160 3884
rect 14648 3528 14700 3534
rect 14648 3470 14700 3476
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14660 3058 14688 3470
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14516 2944 14596 2972
rect 15028 2961 15056 3062
rect 15014 2952 15070 2961
rect 14464 2926 14516 2932
rect 13648 1142 13768 1170
rect 13740 800 13768 1142
rect 14292 1142 14412 1170
rect 14292 800 14320 1142
rect 10060 734 10272 762
rect 10322 0 10378 800
rect 10874 0 10930 800
rect 11426 0 11482 800
rect 12070 0 12126 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13726 0 13782 800
rect 14278 0 14334 800
rect 14476 610 14504 2926
rect 15014 2887 15070 2896
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 14752 1766 14780 2450
rect 14740 1760 14792 1766
rect 14740 1702 14792 1708
rect 14832 1556 14884 1562
rect 14832 1498 14884 1504
rect 14844 800 14872 1498
rect 14936 1494 14964 2790
rect 15016 2372 15068 2378
rect 15016 2314 15068 2320
rect 15028 1737 15056 2314
rect 15014 1728 15070 1737
rect 15014 1663 15070 1672
rect 15120 1630 15148 3878
rect 15198 3768 15254 3777
rect 15198 3703 15254 3712
rect 15212 2650 15240 3703
rect 15304 3641 15332 4014
rect 15384 3936 15436 3942
rect 15384 3878 15436 3884
rect 15290 3632 15346 3641
rect 15290 3567 15346 3576
rect 15200 2644 15252 2650
rect 15200 2586 15252 2592
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15304 1902 15332 2246
rect 15292 1896 15344 1902
rect 15292 1838 15344 1844
rect 15108 1624 15160 1630
rect 15108 1566 15160 1572
rect 14924 1488 14976 1494
rect 14924 1430 14976 1436
rect 15396 800 15424 3878
rect 15488 2961 15516 4694
rect 15580 4264 15608 10202
rect 15672 7818 15700 11494
rect 15764 9602 15792 12922
rect 15856 11830 15884 16662
rect 15948 16522 15976 16730
rect 15936 16516 15988 16522
rect 15936 16458 15988 16464
rect 16040 15706 16068 18226
rect 16132 17678 16160 18702
rect 16316 18698 16528 18714
rect 17224 18702 17276 18708
rect 16316 18692 16540 18698
rect 16316 18686 16488 18692
rect 16316 18358 16344 18686
rect 16488 18634 16540 18640
rect 16396 18624 16448 18630
rect 16396 18566 16448 18572
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 17130 18592 17186 18601
rect 16408 18358 16436 18566
rect 16544 18524 16852 18544
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18448 16852 18468
rect 16304 18352 16356 18358
rect 16304 18294 16356 18300
rect 16396 18352 16448 18358
rect 16396 18294 16448 18300
rect 16408 17678 16436 18294
rect 16764 18216 16816 18222
rect 16960 18204 16988 18566
rect 17130 18527 17186 18536
rect 16816 18176 16988 18204
rect 17040 18216 17092 18222
rect 16764 18158 16816 18164
rect 17040 18158 17092 18164
rect 17052 17785 17080 18158
rect 17038 17776 17094 17785
rect 17038 17711 17094 17720
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16132 17134 16160 17614
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 16316 17270 16344 17546
rect 16544 17436 16852 17456
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17360 16852 17380
rect 16304 17264 16356 17270
rect 16304 17206 16356 17212
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16304 17128 16356 17134
rect 16304 17070 16356 17076
rect 16212 16108 16264 16114
rect 16212 16050 16264 16056
rect 16028 15700 16080 15706
rect 16028 15642 16080 15648
rect 16224 15162 16252 16050
rect 16316 16046 16344 17070
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16684 16833 16712 16934
rect 16670 16824 16726 16833
rect 16670 16759 16726 16768
rect 16776 16658 16804 17138
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16544 16348 16852 16368
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16272 16852 16292
rect 16304 16040 16356 16046
rect 16304 15982 16356 15988
rect 16316 15638 16344 15982
rect 16960 15978 16988 16458
rect 16948 15972 17000 15978
rect 16948 15914 17000 15920
rect 16304 15632 16356 15638
rect 16304 15574 16356 15580
rect 16544 15260 16852 15280
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15184 16852 15204
rect 16212 15156 16264 15162
rect 16212 15098 16264 15104
rect 17040 15088 17092 15094
rect 17040 15030 17092 15036
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16120 13864 16172 13870
rect 16120 13806 16172 13812
rect 16026 13560 16082 13569
rect 16026 13495 16082 13504
rect 15936 13184 15988 13190
rect 15936 13126 15988 13132
rect 15844 11824 15896 11830
rect 15844 11766 15896 11772
rect 15948 11150 15976 13126
rect 16040 13025 16068 13495
rect 16026 13016 16082 13025
rect 16026 12951 16082 12960
rect 16132 12170 16160 13806
rect 16224 12782 16252 14214
rect 16544 14172 16852 14192
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14096 16852 14116
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16316 12306 16344 13262
rect 16544 13084 16852 13104
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13008 16852 13028
rect 16960 12850 16988 14962
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 17052 12730 17080 15030
rect 17144 14385 17172 18527
rect 17130 14376 17186 14385
rect 17130 14311 17186 14320
rect 17236 14278 17264 18702
rect 17316 18624 17368 18630
rect 17316 18566 17368 18572
rect 17328 17202 17356 18566
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17420 18086 17448 18362
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17512 17338 17540 19858
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17604 19417 17632 19790
rect 17590 19408 17646 19417
rect 17590 19343 17646 19352
rect 17696 18465 17724 20352
rect 17788 19378 17816 21383
rect 17880 20058 17908 21519
rect 18142 21176 18198 21185
rect 18142 21111 18198 21120
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 17868 20052 17920 20058
rect 17868 19994 17920 20000
rect 18064 19666 18092 20402
rect 18156 19854 18184 21111
rect 18248 19990 18276 22200
rect 18694 22199 18750 22208
rect 18786 22200 18842 23000
rect 19338 22200 19394 23000
rect 19890 22200 19946 23000
rect 20442 22200 20498 23000
rect 20810 22672 20866 22681
rect 20810 22607 20866 22616
rect 18326 21312 18382 21321
rect 18326 21247 18382 21256
rect 18340 20058 18368 21247
rect 18420 21208 18472 21214
rect 18420 21150 18472 21156
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 18236 19984 18288 19990
rect 18236 19926 18288 19932
rect 18144 19848 18196 19854
rect 18144 19790 18196 19796
rect 18064 19638 18184 19666
rect 18052 19508 18104 19514
rect 18052 19450 18104 19456
rect 17960 19440 18012 19446
rect 18064 19417 18092 19450
rect 17960 19382 18012 19388
rect 18050 19408 18106 19417
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 17868 19372 17920 19378
rect 17868 19314 17920 19320
rect 17682 18456 17738 18465
rect 17682 18391 17738 18400
rect 17880 18306 17908 19314
rect 17972 18873 18000 19382
rect 18050 19343 18106 19352
rect 17958 18864 18014 18873
rect 17958 18799 18014 18808
rect 18052 18760 18104 18766
rect 18052 18702 18104 18708
rect 17788 18278 17908 18306
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 17696 16969 17724 17274
rect 17682 16960 17738 16969
rect 17682 16895 17738 16904
rect 17696 16590 17724 16895
rect 17788 16697 17816 18278
rect 17960 18216 18012 18222
rect 17960 18158 18012 18164
rect 17868 18148 17920 18154
rect 17868 18090 17920 18096
rect 17880 17513 17908 18090
rect 17866 17504 17922 17513
rect 17866 17439 17922 17448
rect 17972 17270 18000 18158
rect 18064 17746 18092 18702
rect 18156 18193 18184 19638
rect 18432 18766 18460 21150
rect 18510 20768 18566 20777
rect 18510 20703 18566 20712
rect 18524 19514 18552 20703
rect 18602 20088 18658 20097
rect 18602 20023 18658 20032
rect 18616 19854 18644 20023
rect 18604 19848 18656 19854
rect 18604 19790 18656 19796
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18616 18426 18644 19654
rect 18708 18970 18736 22199
rect 18800 19718 18828 22200
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18892 20058 18920 20402
rect 19352 20346 19380 22200
rect 19904 21865 19932 22200
rect 19890 21856 19946 21865
rect 19890 21791 19946 21800
rect 20456 21729 20484 22200
rect 20442 21720 20498 21729
rect 20442 21655 20498 21664
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 19522 21040 19578 21049
rect 19522 20975 19578 20984
rect 19168 20318 19380 20346
rect 18972 20256 19024 20262
rect 19168 20244 19196 20318
rect 18972 20198 19024 20204
rect 19076 20216 19196 20244
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18878 19952 18934 19961
rect 18878 19887 18934 19896
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18788 19440 18840 19446
rect 18788 19382 18840 19388
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18696 18692 18748 18698
rect 18696 18634 18748 18640
rect 18708 18426 18736 18634
rect 18604 18420 18656 18426
rect 18604 18362 18656 18368
rect 18696 18420 18748 18426
rect 18696 18362 18748 18368
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18142 18184 18198 18193
rect 18142 18119 18198 18128
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 18052 17740 18104 17746
rect 18052 17682 18104 17688
rect 18156 17678 18184 18022
rect 18248 17746 18276 18226
rect 18326 18184 18382 18193
rect 18326 18119 18382 18128
rect 18236 17740 18288 17746
rect 18236 17682 18288 17688
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 18052 17536 18104 17542
rect 18052 17478 18104 17484
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 17960 17264 18012 17270
rect 17960 17206 18012 17212
rect 18064 16794 18092 17478
rect 18156 17338 18184 17478
rect 18248 17338 18276 17682
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 18236 17332 18288 17338
rect 18236 17274 18288 17280
rect 18144 17128 18196 17134
rect 18144 17070 18196 17076
rect 18156 16833 18184 17070
rect 18142 16824 18198 16833
rect 18052 16788 18104 16794
rect 18142 16759 18198 16768
rect 18052 16730 18104 16736
rect 17774 16688 17830 16697
rect 17774 16623 17830 16632
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17592 16448 17644 16454
rect 17592 16390 17644 16396
rect 17776 16448 17828 16454
rect 17776 16390 17828 16396
rect 17604 16153 17632 16390
rect 17684 16176 17736 16182
rect 17590 16144 17646 16153
rect 17408 16108 17460 16114
rect 17684 16118 17736 16124
rect 17590 16079 17646 16088
rect 17408 16050 17460 16056
rect 17420 15638 17448 16050
rect 17408 15632 17460 15638
rect 17408 15574 17460 15580
rect 17604 15094 17632 16079
rect 17696 15706 17724 16118
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17592 15088 17644 15094
rect 17592 15030 17644 15036
rect 17592 14952 17644 14958
rect 17592 14894 17644 14900
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17224 14272 17276 14278
rect 17224 14214 17276 14220
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 16960 12702 17080 12730
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16684 12306 16712 12582
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 16672 12300 16724 12306
rect 16672 12242 16724 12248
rect 16120 12164 16172 12170
rect 16120 12106 16172 12112
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 15936 11144 15988 11150
rect 15936 11086 15988 11092
rect 16118 11112 16174 11121
rect 16118 11047 16174 11056
rect 16026 10976 16082 10985
rect 16026 10911 16082 10920
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15948 10198 15976 10610
rect 15936 10192 15988 10198
rect 16040 10169 16068 10911
rect 16132 10266 16160 11047
rect 16224 10810 16252 12038
rect 16544 11996 16852 12016
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16394 11928 16450 11937
rect 16544 11920 16852 11940
rect 16394 11863 16450 11872
rect 16408 11665 16436 11863
rect 16672 11688 16724 11694
rect 16394 11656 16450 11665
rect 16672 11630 16724 11636
rect 16394 11591 16450 11600
rect 16304 11552 16356 11558
rect 16304 11494 16356 11500
rect 16316 11286 16344 11494
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16304 11280 16356 11286
rect 16304 11222 16356 11228
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16212 10464 16264 10470
rect 16212 10406 16264 10412
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 15936 10134 15988 10140
rect 16026 10160 16082 10169
rect 16026 10095 16082 10104
rect 15844 9920 15896 9926
rect 15844 9862 15896 9868
rect 15856 9722 15884 9862
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 16132 9654 16160 10202
rect 16224 9722 16252 10406
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16120 9648 16172 9654
rect 15764 9574 15884 9602
rect 16120 9590 16172 9596
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15672 5642 15700 7754
rect 15764 5914 15792 9454
rect 15856 9382 15884 9574
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15948 9178 15976 9522
rect 16120 9512 16172 9518
rect 16120 9454 16172 9460
rect 15936 9172 15988 9178
rect 15936 9114 15988 9120
rect 16132 9058 16160 9454
rect 15856 9030 16160 9058
rect 15856 8838 15884 9030
rect 15936 8968 15988 8974
rect 15936 8910 15988 8916
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 16224 8922 16252 9658
rect 16316 9042 16344 11222
rect 16592 11082 16620 11290
rect 16684 11150 16712 11630
rect 16856 11552 16908 11558
rect 16856 11494 16908 11500
rect 16868 11257 16896 11494
rect 16854 11248 16910 11257
rect 16854 11183 16910 11192
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16408 9586 16436 10950
rect 16544 10908 16852 10928
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10832 16852 10852
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16684 10062 16712 10406
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16544 9820 16852 9840
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9744 16852 9764
rect 16960 9674 16988 12702
rect 17236 12306 17264 13874
rect 17224 12300 17276 12306
rect 17224 12242 17276 12248
rect 17328 11830 17356 14758
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 17420 13258 17448 13670
rect 17408 13252 17460 13258
rect 17408 13194 17460 13200
rect 17420 12918 17448 13194
rect 17408 12912 17460 12918
rect 17408 12854 17460 12860
rect 17420 12238 17448 12854
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17316 11824 17368 11830
rect 17316 11766 17368 11772
rect 17132 11348 17184 11354
rect 17132 11290 17184 11296
rect 17040 11212 17092 11218
rect 17040 11154 17092 11160
rect 17052 10606 17080 11154
rect 17144 11082 17172 11290
rect 17132 11076 17184 11082
rect 17132 11018 17184 11024
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17040 10600 17092 10606
rect 17040 10542 17092 10548
rect 17236 10130 17264 10950
rect 17512 10742 17540 10950
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 17224 10124 17276 10130
rect 17276 10084 17448 10112
rect 17224 10066 17276 10072
rect 16856 9648 16908 9654
rect 16960 9646 17172 9674
rect 16856 9590 16908 9596
rect 16396 9580 16448 9586
rect 16396 9522 16448 9528
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16672 9376 16724 9382
rect 16672 9318 16724 9324
rect 16592 9178 16620 9318
rect 16580 9172 16632 9178
rect 16580 9114 16632 9120
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15856 8344 15884 8774
rect 15948 8498 15976 8910
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 16040 8634 16068 8774
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 16132 8430 16160 8910
rect 16224 8894 16344 8922
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 15936 8356 15988 8362
rect 15856 8316 15936 8344
rect 15936 8298 15988 8304
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16132 8090 16160 8230
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16316 7800 16344 8894
rect 16592 8888 16620 8978
rect 16684 8974 16712 9318
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16868 8906 16896 9590
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16960 9382 16988 9522
rect 16948 9376 17000 9382
rect 16948 9318 17000 9324
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16408 8860 16620 8888
rect 16856 8900 16908 8906
rect 16408 8809 16436 8860
rect 16856 8842 16908 8848
rect 16394 8800 16450 8809
rect 16394 8735 16450 8744
rect 16544 8732 16852 8752
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8656 16852 8676
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16684 8090 16712 8434
rect 16672 8084 16724 8090
rect 16672 8026 16724 8032
rect 16132 7772 16344 7800
rect 15752 5908 15804 5914
rect 15752 5850 15804 5856
rect 15660 5636 15712 5642
rect 15660 5578 15712 5584
rect 16132 5545 16160 7772
rect 16396 7744 16448 7750
rect 16302 7712 16358 7721
rect 16396 7686 16448 7692
rect 16302 7647 16358 7656
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16224 7410 16252 7482
rect 16212 7404 16264 7410
rect 16212 7346 16264 7352
rect 16316 7177 16344 7647
rect 16302 7168 16358 7177
rect 16302 7103 16358 7112
rect 16118 5536 16174 5545
rect 16118 5471 16174 5480
rect 16028 5092 16080 5098
rect 16028 5034 16080 5040
rect 15936 5024 15988 5030
rect 15936 4966 15988 4972
rect 15948 4690 15976 4966
rect 15936 4684 15988 4690
rect 15936 4626 15988 4632
rect 15580 4236 15700 4264
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 15580 3738 15608 4082
rect 15672 4078 15700 4236
rect 15844 4208 15896 4214
rect 15844 4150 15896 4156
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15568 3732 15620 3738
rect 15568 3674 15620 3680
rect 15856 3641 15884 4150
rect 16040 3890 16068 5034
rect 16212 4820 16264 4826
rect 16212 4762 16264 4768
rect 16120 4480 16172 4486
rect 16120 4422 16172 4428
rect 16132 4282 16160 4422
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16224 4026 16252 4762
rect 15948 3862 16068 3890
rect 16132 3998 16252 4026
rect 15842 3632 15898 3641
rect 15842 3567 15898 3576
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15568 3460 15620 3466
rect 15568 3402 15620 3408
rect 15580 3040 15608 3402
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 15672 3233 15700 3334
rect 15658 3224 15714 3233
rect 15658 3159 15714 3168
rect 15752 3188 15804 3194
rect 15752 3130 15804 3136
rect 15660 3052 15712 3058
rect 15580 3012 15660 3040
rect 15660 2994 15712 3000
rect 15474 2952 15530 2961
rect 15474 2887 15530 2896
rect 15566 2680 15622 2689
rect 15566 2615 15568 2624
rect 15620 2615 15622 2624
rect 15568 2586 15620 2592
rect 15764 1290 15792 3130
rect 15856 3097 15884 3470
rect 15842 3088 15898 3097
rect 15842 3023 15898 3032
rect 15752 1284 15804 1290
rect 15752 1226 15804 1232
rect 15948 800 15976 3862
rect 16026 3496 16082 3505
rect 16026 3431 16082 3440
rect 16040 2922 16068 3431
rect 16028 2916 16080 2922
rect 16028 2858 16080 2864
rect 16040 2582 16068 2858
rect 16028 2576 16080 2582
rect 16028 2518 16080 2524
rect 16132 1834 16160 3998
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 16120 1828 16172 1834
rect 16120 1770 16172 1776
rect 16224 1358 16252 3402
rect 16408 1442 16436 7686
rect 16544 7644 16852 7664
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7568 16852 7588
rect 16960 7410 16988 8910
rect 17052 8634 17080 9522
rect 17144 9500 17172 9646
rect 17144 9472 17264 9500
rect 17236 9178 17264 9472
rect 17420 9382 17448 10084
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17314 9208 17370 9217
rect 17224 9172 17276 9178
rect 17314 9143 17370 9152
rect 17408 9172 17460 9178
rect 17224 9114 17276 9120
rect 17132 9104 17184 9110
rect 17132 9046 17184 9052
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17144 8498 17172 9046
rect 17328 8974 17356 9143
rect 17408 9114 17460 9120
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17224 8900 17276 8906
rect 17224 8842 17276 8848
rect 17236 8634 17264 8842
rect 17224 8628 17276 8634
rect 17224 8570 17276 8576
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16946 7168 17002 7177
rect 16592 6934 16620 7142
rect 16946 7103 17002 7112
rect 16580 6928 16632 6934
rect 16580 6870 16632 6876
rect 16544 6556 16852 6576
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6480 16852 6500
rect 16960 6322 16988 7103
rect 17052 6866 17080 7686
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 17224 6724 17276 6730
rect 17224 6666 17276 6672
rect 16948 6316 17000 6322
rect 16948 6258 17000 6264
rect 17132 6316 17184 6322
rect 17132 6258 17184 6264
rect 16948 6180 17000 6186
rect 16948 6122 17000 6128
rect 16544 5468 16852 5488
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5392 16852 5412
rect 16580 5296 16632 5302
rect 16580 5238 16632 5244
rect 16592 4593 16620 5238
rect 16856 4752 16908 4758
rect 16856 4694 16908 4700
rect 16868 4593 16896 4694
rect 16960 4690 16988 6122
rect 17144 5914 17172 6258
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17144 5710 17172 5850
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17040 5228 17092 5234
rect 17144 5216 17172 5646
rect 17092 5188 17172 5216
rect 17040 5170 17092 5176
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 16578 4584 16634 4593
rect 16578 4519 16634 4528
rect 16854 4584 16910 4593
rect 16854 4519 16910 4528
rect 16544 4380 16852 4400
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4304 16852 4324
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16488 3936 16540 3942
rect 16488 3878 16540 3884
rect 16500 3466 16528 3878
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 16544 3292 16852 3312
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3216 16852 3236
rect 16544 2204 16852 2224
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2128 16852 2148
rect 16408 1414 16528 1442
rect 16212 1352 16264 1358
rect 16212 1294 16264 1300
rect 16500 800 16528 1414
rect 16960 814 16988 4082
rect 17052 2774 17080 4150
rect 17144 3534 17172 5188
rect 17132 3528 17184 3534
rect 17132 3470 17184 3476
rect 17052 2746 17172 2774
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 17052 1873 17080 2246
rect 17038 1864 17094 1873
rect 17038 1799 17094 1808
rect 17038 1728 17094 1737
rect 17038 1663 17094 1672
rect 16948 808 17000 814
rect 14464 604 14516 610
rect 14464 546 14516 552
rect 14830 0 14886 800
rect 15382 0 15438 800
rect 15934 0 15990 800
rect 16486 0 16542 800
rect 17052 800 17080 1663
rect 17144 1358 17172 2746
rect 17236 1698 17264 6666
rect 17420 3126 17448 9114
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17512 8362 17540 8978
rect 17500 8356 17552 8362
rect 17500 8298 17552 8304
rect 17604 7206 17632 14894
rect 17788 14346 17816 16390
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 17868 15020 17920 15026
rect 17868 14962 17920 14968
rect 17880 14618 17908 14962
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17776 14340 17828 14346
rect 17776 14282 17828 14288
rect 17696 14062 17908 14090
rect 17696 12442 17724 14062
rect 17880 13938 17908 14062
rect 17868 13932 17920 13938
rect 17868 13874 17920 13880
rect 17776 13728 17828 13734
rect 17776 13670 17828 13676
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17788 12374 17816 13670
rect 17960 13524 18012 13530
rect 17960 13466 18012 13472
rect 17866 13424 17922 13433
rect 17866 13359 17922 13368
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17696 11694 17724 12242
rect 17880 12186 17908 13359
rect 17972 13025 18000 13466
rect 18064 13462 18092 15438
rect 18236 15428 18288 15434
rect 18156 15388 18236 15416
rect 18052 13456 18104 13462
rect 18052 13398 18104 13404
rect 17958 13016 18014 13025
rect 17958 12951 18014 12960
rect 17788 12158 17908 12186
rect 18050 12200 18106 12209
rect 17684 11688 17736 11694
rect 17684 11630 17736 11636
rect 17684 11280 17736 11286
rect 17684 11222 17736 11228
rect 17696 11014 17724 11222
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17696 8362 17724 9998
rect 17684 8356 17736 8362
rect 17684 8298 17736 8304
rect 17788 7886 17816 12158
rect 18050 12135 18106 12144
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17880 11286 17908 12038
rect 18064 11898 18092 12135
rect 18156 12102 18184 15388
rect 18236 15370 18288 15376
rect 18340 15162 18368 18119
rect 18800 16153 18828 19382
rect 18892 19378 18920 19887
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18984 19122 19012 20198
rect 19076 20040 19104 20216
rect 19143 20156 19451 20176
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20080 19451 20100
rect 19536 20040 19564 20975
rect 19798 20496 19854 20505
rect 20364 20466 20392 21082
rect 20824 20913 20852 22607
rect 20994 22200 21050 23000
rect 21546 22200 21602 23000
rect 22098 22200 22154 23000
rect 22650 22200 22706 23000
rect 20810 20904 20866 20913
rect 20810 20839 20866 20848
rect 19798 20431 19800 20440
rect 19852 20431 19854 20440
rect 20352 20460 20404 20466
rect 19800 20402 19852 20408
rect 20352 20402 20404 20408
rect 19076 20012 19380 20040
rect 19246 19952 19302 19961
rect 19246 19887 19302 19896
rect 19260 19514 19288 19887
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19352 19310 19380 20012
rect 19444 20012 19564 20040
rect 19444 19378 19472 20012
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20168 19780 20220 19786
rect 20168 19722 20220 19728
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19524 19304 19576 19310
rect 19524 19246 19576 19252
rect 19536 19174 19564 19246
rect 19524 19168 19576 19174
rect 18984 19094 19104 19122
rect 19524 19110 19576 19116
rect 18972 18624 19024 18630
rect 18972 18566 19024 18572
rect 18984 17270 19012 18566
rect 18972 17264 19024 17270
rect 18972 17206 19024 17212
rect 18880 16584 18932 16590
rect 18880 16526 18932 16532
rect 18786 16144 18842 16153
rect 18786 16079 18842 16088
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18328 15156 18380 15162
rect 18328 15098 18380 15104
rect 18236 14340 18288 14346
rect 18236 14282 18288 14288
rect 18248 13870 18276 14282
rect 18236 13864 18288 13870
rect 18236 13806 18288 13812
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18234 13288 18290 13297
rect 18234 13223 18290 13232
rect 18248 12238 18276 13223
rect 18236 12232 18288 12238
rect 18236 12174 18288 12180
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18340 11898 18368 13806
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18236 11552 18288 11558
rect 18236 11494 18288 11500
rect 17868 11280 17920 11286
rect 17868 11222 17920 11228
rect 17960 11008 18012 11014
rect 17880 10956 17960 10962
rect 17880 10950 18012 10956
rect 17880 10934 18000 10950
rect 17880 9926 17908 10934
rect 18064 10742 18092 11494
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 17960 10736 18012 10742
rect 17958 10704 17960 10713
rect 18052 10736 18104 10742
rect 18012 10704 18014 10713
rect 18052 10678 18104 10684
rect 17958 10639 18014 10648
rect 18156 10606 18184 11086
rect 18248 11082 18276 11494
rect 18432 11082 18460 15846
rect 18616 15745 18644 15846
rect 18602 15736 18658 15745
rect 18602 15671 18658 15680
rect 18696 15632 18748 15638
rect 18694 15600 18696 15609
rect 18748 15600 18750 15609
rect 18694 15535 18750 15544
rect 18786 15192 18842 15201
rect 18512 15156 18564 15162
rect 18786 15127 18842 15136
rect 18512 15098 18564 15104
rect 18524 12714 18552 15098
rect 18696 14952 18748 14958
rect 18694 14920 18696 14929
rect 18748 14920 18750 14929
rect 18694 14855 18750 14864
rect 18800 14618 18828 15127
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18892 13870 18920 16526
rect 18972 15972 19024 15978
rect 18972 15914 19024 15920
rect 18984 15434 19012 15914
rect 19076 15609 19104 19094
rect 19143 19068 19451 19088
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 18992 19451 19012
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19536 18086 19564 18702
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19143 17980 19451 18000
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17904 19451 17924
rect 19536 17746 19564 18022
rect 19524 17740 19576 17746
rect 19524 17682 19576 17688
rect 19522 17640 19578 17649
rect 19522 17575 19524 17584
rect 19576 17575 19578 17584
rect 19524 17546 19576 17552
rect 19522 17232 19578 17241
rect 19522 17167 19578 17176
rect 19143 16892 19451 16912
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16816 19451 16836
rect 19248 16652 19300 16658
rect 19248 16594 19300 16600
rect 19260 16250 19288 16594
rect 19536 16522 19564 17167
rect 19628 16590 19656 19314
rect 19708 18692 19760 18698
rect 19708 18634 19760 18640
rect 19616 16584 19668 16590
rect 19616 16526 19668 16532
rect 19524 16516 19576 16522
rect 19524 16458 19576 16464
rect 19248 16244 19300 16250
rect 19248 16186 19300 16192
rect 19143 15804 19451 15824
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15728 19451 15748
rect 19062 15600 19118 15609
rect 19062 15535 19118 15544
rect 18972 15428 19024 15434
rect 18972 15370 19024 15376
rect 19248 15360 19300 15366
rect 19248 15302 19300 15308
rect 19260 15094 19288 15302
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19248 15088 19300 15094
rect 19248 15030 19300 15036
rect 19444 15026 19472 15098
rect 19432 15020 19484 15026
rect 19484 14980 19564 15008
rect 19432 14962 19484 14968
rect 19143 14716 19451 14736
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14640 19451 14660
rect 19430 14512 19486 14521
rect 19536 14482 19564 14980
rect 19614 14648 19670 14657
rect 19614 14583 19616 14592
rect 19668 14583 19670 14592
rect 19616 14554 19668 14560
rect 19430 14447 19486 14456
rect 19524 14476 19576 14482
rect 19444 14414 19472 14447
rect 19524 14418 19576 14424
rect 19432 14408 19484 14414
rect 19432 14350 19484 14356
rect 18880 13864 18932 13870
rect 18880 13806 18932 13812
rect 18970 13696 19026 13705
rect 19026 13654 19104 13682
rect 18970 13631 19026 13640
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18604 13320 18656 13326
rect 18604 13262 18656 13268
rect 18512 12708 18564 12714
rect 18512 12650 18564 12656
rect 18616 12442 18644 13262
rect 18708 12986 18736 13330
rect 19076 13326 19104 13654
rect 19143 13628 19451 13648
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13552 19451 13572
rect 19064 13320 19116 13326
rect 19064 13262 19116 13268
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18708 12866 18736 12922
rect 18708 12838 18828 12866
rect 18800 12782 18828 12838
rect 18788 12776 18840 12782
rect 18788 12718 18840 12724
rect 18696 12708 18748 12714
rect 18696 12650 18748 12656
rect 18604 12436 18656 12442
rect 18604 12378 18656 12384
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 18420 11076 18472 11082
rect 18420 11018 18472 11024
rect 18236 10668 18288 10674
rect 18236 10610 18288 10616
rect 18144 10600 18196 10606
rect 18144 10542 18196 10548
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 17958 10024 18014 10033
rect 17958 9959 18014 9968
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17972 9654 18000 9959
rect 17960 9648 18012 9654
rect 17960 9590 18012 9596
rect 17958 9208 18014 9217
rect 17880 9166 17958 9194
rect 17880 8974 17908 9166
rect 18064 9178 18092 10406
rect 18156 10062 18184 10542
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 18156 9518 18184 9998
rect 18144 9512 18196 9518
rect 18144 9454 18196 9460
rect 17958 9143 18014 9152
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 17958 9072 18014 9081
rect 17958 9007 18014 9016
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17972 8820 18000 9007
rect 17880 8792 18000 8820
rect 17880 8265 17908 8792
rect 17958 8664 18014 8673
rect 17958 8599 18014 8608
rect 17866 8256 17922 8265
rect 17866 8191 17922 8200
rect 17972 7954 18000 8599
rect 18156 8566 18184 9454
rect 18248 9042 18276 10610
rect 18326 10432 18382 10441
rect 18326 10367 18382 10376
rect 18236 9036 18288 9042
rect 18236 8978 18288 8984
rect 18340 8906 18368 10367
rect 18418 10296 18474 10305
rect 18418 10231 18474 10240
rect 18328 8900 18380 8906
rect 18328 8842 18380 8848
rect 18234 8800 18290 8809
rect 18234 8735 18290 8744
rect 18144 8560 18196 8566
rect 18050 8528 18106 8537
rect 18144 8502 18196 8508
rect 18050 8463 18106 8472
rect 17960 7948 18012 7954
rect 17960 7890 18012 7896
rect 17776 7880 17828 7886
rect 18064 7857 18092 8463
rect 18156 8090 18184 8502
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 17776 7822 17828 7828
rect 17866 7848 17922 7857
rect 17866 7783 17922 7792
rect 18050 7848 18106 7857
rect 18050 7783 18106 7792
rect 17880 7585 17908 7783
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17866 7576 17922 7585
rect 17866 7511 17922 7520
rect 17774 7440 17830 7449
rect 17774 7375 17830 7384
rect 17592 7200 17644 7206
rect 17592 7142 17644 7148
rect 17592 6928 17644 6934
rect 17590 6896 17592 6905
rect 17644 6896 17646 6905
rect 17590 6831 17646 6840
rect 17682 6760 17738 6769
rect 17682 6695 17738 6704
rect 17696 6662 17724 6695
rect 17500 6656 17552 6662
rect 17684 6656 17736 6662
rect 17500 6598 17552 6604
rect 17590 6624 17646 6633
rect 17512 5914 17540 6598
rect 17684 6598 17736 6604
rect 17590 6559 17646 6568
rect 17500 5908 17552 5914
rect 17500 5850 17552 5856
rect 17604 3992 17632 6559
rect 17788 6440 17816 7375
rect 17958 7032 18014 7041
rect 17958 6967 18014 6976
rect 17972 6866 18000 6967
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17958 6760 18014 6769
rect 17958 6695 18014 6704
rect 17972 6458 18000 6695
rect 17696 6412 17816 6440
rect 17960 6452 18012 6458
rect 17696 4622 17724 6412
rect 17960 6394 18012 6400
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17684 4616 17736 4622
rect 17684 4558 17736 4564
rect 17696 4282 17724 4558
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17604 3964 17724 3992
rect 17590 3904 17646 3913
rect 17590 3839 17646 3848
rect 17500 3460 17552 3466
rect 17500 3402 17552 3408
rect 17408 3120 17460 3126
rect 17408 3062 17460 3068
rect 17224 1692 17276 1698
rect 17224 1634 17276 1640
rect 17132 1352 17184 1358
rect 17130 1320 17132 1329
rect 17184 1320 17186 1329
rect 17130 1255 17186 1264
rect 17512 1086 17540 3402
rect 17604 3398 17632 3839
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17590 3224 17646 3233
rect 17590 3159 17646 3168
rect 17500 1080 17552 1086
rect 17500 1022 17552 1028
rect 16948 750 17000 756
rect 17038 0 17094 800
rect 17604 678 17632 3159
rect 17696 800 17724 3964
rect 17788 1601 17816 6258
rect 18064 5370 18092 7686
rect 18248 7177 18276 8735
rect 18432 8294 18460 10231
rect 18524 9908 18552 12038
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18616 11234 18644 11698
rect 18708 11354 18736 12650
rect 18800 12306 18828 12718
rect 18788 12300 18840 12306
rect 18788 12242 18840 12248
rect 18892 11898 18920 13126
rect 18970 12744 19026 12753
rect 18970 12679 19026 12688
rect 18880 11892 18932 11898
rect 18880 11834 18932 11840
rect 18984 11762 19012 12679
rect 18972 11756 19024 11762
rect 18972 11698 19024 11704
rect 18696 11348 18748 11354
rect 18696 11290 18748 11296
rect 18616 11206 18736 11234
rect 18602 10568 18658 10577
rect 18602 10503 18658 10512
rect 18616 10062 18644 10503
rect 18604 10056 18656 10062
rect 18708 10033 18736 11206
rect 18604 9998 18656 10004
rect 18694 10024 18750 10033
rect 18694 9959 18750 9968
rect 18524 9880 18644 9908
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18420 8288 18472 8294
rect 18420 8230 18472 8236
rect 18524 8022 18552 9114
rect 18512 8016 18564 8022
rect 18512 7958 18564 7964
rect 18420 7948 18472 7954
rect 18420 7890 18472 7896
rect 18432 7546 18460 7890
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18328 7200 18380 7206
rect 18234 7168 18290 7177
rect 18328 7142 18380 7148
rect 18234 7103 18290 7112
rect 18234 6896 18290 6905
rect 18234 6831 18290 6840
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18052 5364 18104 5370
rect 18052 5306 18104 5312
rect 17866 4856 17922 4865
rect 17866 4791 17868 4800
rect 17920 4791 17922 4800
rect 17868 4762 17920 4768
rect 17868 4548 17920 4554
rect 17868 4490 17920 4496
rect 17880 4010 17908 4490
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 17866 3904 17922 3913
rect 17866 3839 17922 3848
rect 17774 1592 17830 1601
rect 17774 1527 17830 1536
rect 17880 1018 17908 3839
rect 17972 2106 18000 4422
rect 18052 4208 18104 4214
rect 18050 4176 18052 4185
rect 18104 4176 18106 4185
rect 18050 4111 18106 4120
rect 18050 4040 18106 4049
rect 18050 3975 18106 3984
rect 18064 3534 18092 3975
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18064 2650 18092 3334
rect 18052 2644 18104 2650
rect 18052 2586 18104 2592
rect 17960 2100 18012 2106
rect 17960 2042 18012 2048
rect 18156 1170 18184 6598
rect 18248 5817 18276 6831
rect 18234 5808 18290 5817
rect 18340 5778 18368 7142
rect 18432 5778 18460 7482
rect 18616 7449 18644 9880
rect 18708 9586 18736 9959
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18970 9344 19026 9353
rect 18970 9279 19026 9288
rect 18984 8906 19012 9279
rect 18696 8900 18748 8906
rect 18696 8842 18748 8848
rect 18972 8900 19024 8906
rect 18972 8842 19024 8848
rect 18708 7478 18736 8842
rect 18788 8832 18840 8838
rect 18788 8774 18840 8780
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18800 8634 18828 8774
rect 18788 8628 18840 8634
rect 18788 8570 18840 8576
rect 18892 8498 18920 8774
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18984 8401 19012 8434
rect 18970 8392 19026 8401
rect 18970 8327 19026 8336
rect 18880 8288 18932 8294
rect 18880 8230 18932 8236
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18800 7546 18828 7686
rect 18788 7540 18840 7546
rect 18788 7482 18840 7488
rect 18696 7472 18748 7478
rect 18602 7440 18658 7449
rect 18696 7414 18748 7420
rect 18602 7375 18658 7384
rect 18512 7268 18564 7274
rect 18512 7210 18564 7216
rect 18524 6118 18552 7210
rect 18892 6866 18920 8230
rect 18984 8129 19012 8230
rect 18970 8120 19026 8129
rect 18970 8055 19026 8064
rect 18972 8016 19024 8022
rect 18972 7958 19024 7964
rect 18880 6860 18932 6866
rect 18880 6802 18932 6808
rect 18604 6792 18656 6798
rect 18984 6746 19012 7958
rect 19076 7546 19104 13262
rect 19536 12918 19564 14418
rect 19616 14068 19668 14074
rect 19616 14010 19668 14016
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19143 12540 19451 12560
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12464 19451 12484
rect 19536 12306 19564 12854
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19522 12200 19578 12209
rect 19522 12135 19578 12144
rect 19143 11452 19451 11472
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11376 19451 11396
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19260 10742 19288 11086
rect 19248 10736 19300 10742
rect 19248 10678 19300 10684
rect 19143 10364 19451 10384
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10288 19451 10308
rect 19338 10160 19394 10169
rect 19338 10095 19394 10104
rect 19352 10062 19380 10095
rect 19340 10056 19392 10062
rect 19340 9998 19392 10004
rect 19536 9738 19564 12135
rect 19628 11830 19656 14010
rect 19720 12850 19748 18634
rect 19800 18352 19852 18358
rect 19984 18352 20036 18358
rect 19800 18294 19852 18300
rect 19982 18320 19984 18329
rect 20036 18320 20038 18329
rect 19812 16658 19840 18294
rect 19982 18255 20038 18264
rect 19892 17808 19944 17814
rect 19892 17750 19944 17756
rect 19984 17808 20036 17814
rect 19984 17750 20036 17756
rect 19800 16652 19852 16658
rect 19800 16594 19852 16600
rect 19800 16448 19852 16454
rect 19800 16390 19852 16396
rect 19812 15434 19840 16390
rect 19800 15428 19852 15434
rect 19800 15370 19852 15376
rect 19812 14074 19840 15370
rect 19800 14068 19852 14074
rect 19800 14010 19852 14016
rect 19904 13954 19932 17750
rect 19996 17610 20024 17750
rect 19984 17604 20036 17610
rect 19984 17546 20036 17552
rect 19984 16992 20036 16998
rect 19984 16934 20036 16940
rect 19996 16182 20024 16934
rect 20180 16726 20208 19722
rect 20548 19378 20576 19858
rect 20824 19854 20852 20839
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 21008 19242 21036 22200
rect 21560 20602 21588 22200
rect 21548 20596 21600 20602
rect 21548 20538 21600 20544
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 21100 19553 21128 20402
rect 22112 20330 22140 22200
rect 22100 20324 22152 20330
rect 22100 20266 22152 20272
rect 21270 19816 21326 19825
rect 21270 19751 21272 19760
rect 21324 19751 21326 19760
rect 21272 19722 21324 19728
rect 21086 19544 21142 19553
rect 21086 19479 21142 19488
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 20996 19236 21048 19242
rect 20996 19178 21048 19184
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 17105 20300 18566
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 20364 17678 20392 18022
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20628 17196 20680 17202
rect 20628 17138 20680 17144
rect 20258 17096 20314 17105
rect 20258 17031 20314 17040
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20168 16720 20220 16726
rect 20168 16662 20220 16668
rect 20258 16552 20314 16561
rect 20076 16516 20128 16522
rect 20258 16487 20314 16496
rect 20076 16458 20128 16464
rect 20088 16250 20116 16458
rect 20272 16454 20300 16487
rect 20260 16448 20312 16454
rect 20260 16390 20312 16396
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 20364 16250 20392 16390
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 19984 16176 20036 16182
rect 19984 16118 20036 16124
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20076 15360 20128 15366
rect 20076 15302 20128 15308
rect 19812 13926 19932 13954
rect 19984 14000 20036 14006
rect 19984 13942 20036 13948
rect 19708 12844 19760 12850
rect 19708 12786 19760 12792
rect 19812 12730 19840 13926
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19904 13394 19932 13806
rect 19892 13388 19944 13394
rect 19892 13330 19944 13336
rect 19996 13274 20024 13942
rect 19720 12702 19840 12730
rect 19904 13246 20024 13274
rect 19720 12238 19748 12702
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19904 12102 19932 13246
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19892 12096 19944 12102
rect 19892 12038 19944 12044
rect 19616 11824 19668 11830
rect 19616 11766 19668 11772
rect 19996 11694 20024 13126
rect 19800 11688 19852 11694
rect 19800 11630 19852 11636
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19536 9710 19656 9738
rect 19522 9616 19578 9625
rect 19522 9551 19578 9560
rect 19536 9450 19564 9551
rect 19524 9444 19576 9450
rect 19524 9386 19576 9392
rect 19143 9276 19451 9296
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9200 19451 9220
rect 19536 9110 19564 9386
rect 19156 9104 19208 9110
rect 19156 9046 19208 9052
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19524 9104 19576 9110
rect 19524 9046 19576 9052
rect 19168 8362 19196 9046
rect 19444 8974 19472 9046
rect 19432 8968 19484 8974
rect 19628 8922 19656 9710
rect 19812 9450 19840 11630
rect 19996 10810 20024 11630
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19800 9444 19852 9450
rect 19800 9386 19852 9392
rect 19432 8910 19484 8916
rect 19536 8894 19656 8922
rect 19156 8356 19208 8362
rect 19156 8298 19208 8304
rect 19143 8188 19451 8208
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8112 19451 8132
rect 19536 8022 19564 8894
rect 19616 8832 19668 8838
rect 19616 8774 19668 8780
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19524 8016 19576 8022
rect 19524 7958 19576 7964
rect 19524 7880 19576 7886
rect 19524 7822 19576 7828
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 19156 7404 19208 7410
rect 19156 7346 19208 7352
rect 19168 7313 19196 7346
rect 19154 7304 19210 7313
rect 19154 7239 19210 7248
rect 19143 7100 19451 7120
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7024 19451 7044
rect 19536 6882 19564 7822
rect 19444 6854 19564 6882
rect 19444 6798 19472 6854
rect 18604 6734 18656 6740
rect 18616 6497 18644 6734
rect 18892 6718 19012 6746
rect 19432 6792 19484 6798
rect 19432 6734 19484 6740
rect 18602 6488 18658 6497
rect 18602 6423 18658 6432
rect 18786 6216 18842 6225
rect 18786 6151 18842 6160
rect 18512 6112 18564 6118
rect 18512 6054 18564 6060
rect 18234 5743 18290 5752
rect 18328 5772 18380 5778
rect 18328 5714 18380 5720
rect 18420 5772 18472 5778
rect 18420 5714 18472 5720
rect 18236 5568 18288 5574
rect 18236 5510 18288 5516
rect 18248 2514 18276 5510
rect 18524 5302 18552 6054
rect 18694 5808 18750 5817
rect 18694 5743 18750 5752
rect 18512 5296 18564 5302
rect 18512 5238 18564 5244
rect 18602 5264 18658 5273
rect 18602 5199 18604 5208
rect 18656 5199 18658 5208
rect 18604 5170 18656 5176
rect 18510 5128 18566 5137
rect 18510 5063 18566 5072
rect 18420 4616 18472 4622
rect 18420 4558 18472 4564
rect 18328 4480 18380 4486
rect 18328 4422 18380 4428
rect 18340 4282 18368 4422
rect 18328 4276 18380 4282
rect 18328 4218 18380 4224
rect 18432 3602 18460 4558
rect 18420 3596 18472 3602
rect 18420 3538 18472 3544
rect 18524 3534 18552 5063
rect 18604 5024 18656 5030
rect 18604 4966 18656 4972
rect 18616 4690 18644 4966
rect 18604 4684 18656 4690
rect 18604 4626 18656 4632
rect 18512 3528 18564 3534
rect 18512 3470 18564 3476
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18328 2984 18380 2990
rect 18326 2952 18328 2961
rect 18380 2952 18382 2961
rect 18326 2887 18382 2896
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 18326 2408 18382 2417
rect 18326 2343 18328 2352
rect 18380 2343 18382 2352
rect 18328 2314 18380 2320
rect 18432 2038 18460 3402
rect 18512 2304 18564 2310
rect 18512 2246 18564 2252
rect 18420 2032 18472 2038
rect 18420 1974 18472 1980
rect 18156 1142 18276 1170
rect 17868 1012 17920 1018
rect 17868 954 17920 960
rect 17960 944 18012 950
rect 17960 886 18012 892
rect 17592 672 17644 678
rect 17592 614 17644 620
rect 17682 0 17738 800
rect 17972 241 18000 886
rect 18248 800 18276 1142
rect 18524 921 18552 2246
rect 18616 1970 18644 4626
rect 18708 3913 18736 5743
rect 18694 3904 18750 3913
rect 18694 3839 18750 3848
rect 18694 3632 18750 3641
rect 18694 3567 18750 3576
rect 18708 3074 18736 3567
rect 18800 3233 18828 6151
rect 18892 5778 18920 6718
rect 18972 6656 19024 6662
rect 18970 6624 18972 6633
rect 19024 6624 19026 6633
rect 18970 6559 19026 6568
rect 18970 6488 19026 6497
rect 18970 6423 19026 6432
rect 18984 6089 19012 6423
rect 19444 6390 19472 6734
rect 19432 6384 19484 6390
rect 19432 6326 19484 6332
rect 19064 6316 19116 6322
rect 19064 6258 19116 6264
rect 18970 6080 19026 6089
rect 18970 6015 19026 6024
rect 19076 5914 19104 6258
rect 19524 6112 19576 6118
rect 19628 6066 19656 8774
rect 19706 7984 19762 7993
rect 19706 7919 19762 7928
rect 19720 7886 19748 7919
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19576 6060 19656 6066
rect 19524 6054 19656 6060
rect 19536 6038 19656 6054
rect 19143 6012 19451 6032
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5936 19451 5956
rect 19064 5908 19116 5914
rect 19064 5850 19116 5856
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18972 5704 19024 5710
rect 18972 5646 19024 5652
rect 19338 5672 19394 5681
rect 18984 4690 19012 5646
rect 19338 5607 19340 5616
rect 19392 5607 19394 5616
rect 19340 5578 19392 5584
rect 19628 5370 19656 6038
rect 19616 5364 19668 5370
rect 19616 5306 19668 5312
rect 19062 5264 19118 5273
rect 19062 5199 19118 5208
rect 19076 4758 19104 5199
rect 19812 5114 19840 8774
rect 19904 5284 19932 9862
rect 20088 8106 20116 15302
rect 20168 14000 20220 14006
rect 20168 13942 20220 13948
rect 20180 9994 20208 13942
rect 20272 13190 20300 15642
rect 20456 15434 20484 16934
rect 20640 16794 20668 17138
rect 20628 16788 20680 16794
rect 20628 16730 20680 16736
rect 20732 16561 20760 19110
rect 20904 18760 20956 18766
rect 20904 18702 20956 18708
rect 20810 18592 20866 18601
rect 20810 18527 20866 18536
rect 20824 18426 20852 18527
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20718 16552 20774 16561
rect 20718 16487 20774 16496
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20628 15496 20680 15502
rect 20732 15473 20760 16050
rect 20628 15438 20680 15444
rect 20718 15464 20774 15473
rect 20444 15428 20496 15434
rect 20444 15370 20496 15376
rect 20640 15162 20668 15438
rect 20718 15399 20774 15408
rect 20824 15162 20852 18226
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20812 15156 20864 15162
rect 20812 15098 20864 15104
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20444 14816 20496 14822
rect 20444 14758 20496 14764
rect 20456 14482 20484 14758
rect 20444 14476 20496 14482
rect 20444 14418 20496 14424
rect 20352 14272 20404 14278
rect 20352 14214 20404 14220
rect 20364 14074 20392 14214
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20260 12980 20312 12986
rect 20260 12922 20312 12928
rect 20272 12889 20300 12922
rect 20258 12880 20314 12889
rect 20258 12815 20314 12824
rect 20258 12336 20314 12345
rect 20258 12271 20314 12280
rect 20272 10742 20300 12271
rect 20260 10736 20312 10742
rect 20260 10678 20312 10684
rect 20364 10266 20392 13874
rect 20732 13530 20760 14962
rect 20824 14482 20852 15098
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20534 13424 20590 13433
rect 20534 13359 20590 13368
rect 20720 13388 20772 13394
rect 20548 13326 20576 13359
rect 20720 13330 20772 13336
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20444 12096 20496 12102
rect 20444 12038 20496 12044
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20168 9988 20220 9994
rect 20168 9930 20220 9936
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 20180 9489 20208 9522
rect 20364 9518 20392 10202
rect 20260 9512 20312 9518
rect 20166 9480 20222 9489
rect 20260 9454 20312 9460
rect 20352 9512 20404 9518
rect 20352 9454 20404 9460
rect 20166 9415 20222 9424
rect 20272 9178 20300 9454
rect 20352 9376 20404 9382
rect 20352 9318 20404 9324
rect 20364 9178 20392 9318
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20352 9172 20404 9178
rect 20352 9114 20404 9120
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 19996 8090 20116 8106
rect 19984 8084 20116 8090
rect 20036 8078 20116 8084
rect 19984 8026 20036 8032
rect 20180 7970 20208 8910
rect 20088 7942 20208 7970
rect 19904 5256 20024 5284
rect 19892 5160 19944 5166
rect 19890 5128 19892 5137
rect 19944 5128 19946 5137
rect 19812 5086 19890 5114
rect 19890 5063 19946 5072
rect 19143 4924 19451 4944
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4848 19451 4868
rect 19064 4752 19116 4758
rect 19064 4694 19116 4700
rect 19890 4720 19946 4729
rect 18972 4684 19024 4690
rect 19890 4655 19946 4664
rect 18972 4626 19024 4632
rect 18878 4448 18934 4457
rect 18878 4383 18934 4392
rect 18786 3224 18842 3233
rect 18786 3159 18842 3168
rect 18708 3046 18828 3074
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18708 2514 18736 2790
rect 18696 2508 18748 2514
rect 18696 2450 18748 2456
rect 18604 1964 18656 1970
rect 18604 1906 18656 1912
rect 18708 1222 18736 2450
rect 18696 1216 18748 1222
rect 18696 1158 18748 1164
rect 18510 912 18566 921
rect 18510 847 18566 856
rect 18800 800 18828 3046
rect 18892 1154 18920 4383
rect 18984 4282 19012 4626
rect 19062 4584 19118 4593
rect 19062 4519 19118 4528
rect 19800 4548 19852 4554
rect 18972 4276 19024 4282
rect 18972 4218 19024 4224
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18984 3777 19012 4082
rect 18970 3768 19026 3777
rect 18970 3703 19026 3712
rect 18970 3632 19026 3641
rect 18970 3567 19026 3576
rect 18880 1148 18932 1154
rect 18880 1090 18932 1096
rect 17958 232 18014 241
rect 17958 167 18014 176
rect 18234 0 18290 800
rect 18786 0 18842 800
rect 18984 746 19012 3567
rect 19076 3398 19104 4519
rect 19800 4490 19852 4496
rect 19616 4208 19668 4214
rect 19616 4150 19668 4156
rect 19143 3836 19451 3856
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3760 19451 3780
rect 19628 3602 19656 4150
rect 19708 4004 19760 4010
rect 19708 3946 19760 3952
rect 19156 3596 19208 3602
rect 19156 3538 19208 3544
rect 19616 3596 19668 3602
rect 19616 3538 19668 3544
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 19168 3194 19196 3538
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19338 3360 19394 3369
rect 19338 3295 19394 3304
rect 19156 3188 19208 3194
rect 19156 3130 19208 3136
rect 19352 2990 19380 3295
rect 19430 3088 19486 3097
rect 19430 3023 19432 3032
rect 19484 3023 19486 3032
rect 19432 2994 19484 3000
rect 19340 2984 19392 2990
rect 19340 2926 19392 2932
rect 19064 2916 19116 2922
rect 19064 2858 19116 2864
rect 19076 921 19104 2858
rect 19143 2748 19451 2768
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2672 19451 2692
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 19260 2009 19288 2382
rect 19246 2000 19302 2009
rect 19246 1935 19302 1944
rect 19536 1902 19564 3402
rect 19616 3392 19668 3398
rect 19616 3334 19668 3340
rect 19524 1896 19576 1902
rect 19524 1838 19576 1844
rect 19340 1420 19392 1426
rect 19340 1362 19392 1368
rect 19248 1352 19300 1358
rect 19248 1294 19300 1300
rect 19260 1193 19288 1294
rect 19246 1184 19302 1193
rect 19246 1119 19302 1128
rect 19062 912 19118 921
rect 19062 847 19118 856
rect 19352 800 19380 1362
rect 19628 882 19656 3334
rect 19720 1057 19748 3946
rect 19812 3942 19840 4490
rect 19904 4146 19932 4655
rect 19892 4140 19944 4146
rect 19892 4082 19944 4088
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19812 2514 19840 3878
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 19800 2508 19852 2514
rect 19800 2450 19852 2456
rect 19706 1048 19762 1057
rect 19706 983 19762 992
rect 19616 876 19668 882
rect 19616 818 19668 824
rect 19904 800 19932 3674
rect 19996 2774 20024 5256
rect 20088 4146 20116 7942
rect 20168 7812 20220 7818
rect 20168 7754 20220 7760
rect 20180 7546 20208 7754
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 20180 6118 20208 6666
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 20088 3670 20116 3878
rect 20076 3664 20128 3670
rect 20076 3606 20128 3612
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20088 2990 20116 3470
rect 20180 3074 20208 6054
rect 20260 4208 20312 4214
rect 20260 4150 20312 4156
rect 20272 3194 20300 4150
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20260 3188 20312 3194
rect 20260 3130 20312 3136
rect 20180 3046 20300 3074
rect 20076 2984 20128 2990
rect 20076 2926 20128 2932
rect 19996 2746 20208 2774
rect 20180 1426 20208 2746
rect 20272 1766 20300 3046
rect 20364 2774 20392 4082
rect 20456 2938 20484 12038
rect 20548 6458 20576 12718
rect 20640 12646 20668 13126
rect 20628 12640 20680 12646
rect 20628 12582 20680 12588
rect 20732 12170 20760 13330
rect 20916 12782 20944 18702
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 21008 16658 21036 17138
rect 20996 16652 21048 16658
rect 20996 16594 21048 16600
rect 20996 15088 21048 15094
rect 20996 15030 21048 15036
rect 21086 15056 21142 15065
rect 21008 13870 21036 15030
rect 21086 14991 21088 15000
rect 21140 14991 21142 15000
rect 21088 14962 21140 14968
rect 21192 14362 21220 19314
rect 21284 17105 21312 19450
rect 22664 19310 22692 22200
rect 22652 19304 22704 19310
rect 22652 19246 22704 19252
rect 21548 17604 21600 17610
rect 21548 17546 21600 17552
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21270 17096 21326 17105
rect 21270 17031 21326 17040
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21100 14334 21220 14362
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 21100 13462 21128 14334
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21088 13456 21140 13462
rect 21088 13398 21140 13404
rect 21192 13297 21220 14214
rect 21284 13841 21312 14758
rect 21376 14249 21404 15302
rect 21362 14240 21418 14249
rect 21362 14175 21418 14184
rect 21270 13832 21326 13841
rect 21270 13767 21326 13776
rect 21468 13326 21496 17478
rect 21456 13320 21508 13326
rect 21178 13288 21234 13297
rect 21456 13262 21508 13268
rect 21178 13223 21234 13232
rect 20996 13184 21048 13190
rect 20996 13126 21048 13132
rect 21008 12986 21036 13126
rect 21560 12986 21588 17546
rect 22006 13968 22062 13977
rect 22062 13926 22140 13954
rect 22006 13903 22062 13912
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 21548 12980 21600 12986
rect 21548 12922 21600 12928
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20916 12442 20944 12718
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20720 12164 20772 12170
rect 20720 12106 20772 12112
rect 20732 11914 20760 12106
rect 20994 12064 21050 12073
rect 20994 11999 21050 12008
rect 20732 11886 20944 11914
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20640 10470 20668 11562
rect 20732 11121 20760 11698
rect 20718 11112 20774 11121
rect 20718 11047 20774 11056
rect 20718 10840 20774 10849
rect 20718 10775 20774 10784
rect 20628 10464 20680 10470
rect 20628 10406 20680 10412
rect 20640 10266 20668 10406
rect 20628 10260 20680 10266
rect 20628 10202 20680 10208
rect 20640 9518 20668 10202
rect 20732 10062 20760 10775
rect 20916 10470 20944 11886
rect 21008 11286 21036 11999
rect 20996 11280 21048 11286
rect 20996 11222 21048 11228
rect 21456 11280 21508 11286
rect 21456 11222 21508 11228
rect 20904 10464 20956 10470
rect 20904 10406 20956 10412
rect 21180 10464 21232 10470
rect 21180 10406 21232 10412
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20812 9920 20864 9926
rect 20812 9862 20864 9868
rect 20628 9512 20680 9518
rect 20628 9454 20680 9460
rect 20718 9480 20774 9489
rect 20718 9415 20774 9424
rect 20628 9376 20680 9382
rect 20628 9318 20680 9324
rect 20640 8090 20668 9318
rect 20732 8809 20760 9415
rect 20718 8800 20774 8809
rect 20718 8735 20774 8744
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20732 7750 20760 8502
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20536 6452 20588 6458
rect 20536 6394 20588 6400
rect 20640 6361 20668 6598
rect 20626 6352 20682 6361
rect 20548 6310 20626 6338
rect 20548 3602 20576 6310
rect 20626 6287 20682 6296
rect 20628 6248 20680 6254
rect 20628 6190 20680 6196
rect 20640 5370 20668 6190
rect 20628 5364 20680 5370
rect 20628 5306 20680 5312
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 20536 3596 20588 3602
rect 20536 3538 20588 3544
rect 20640 3505 20668 5170
rect 20732 3602 20760 7686
rect 20824 3738 20852 9862
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20916 6458 20944 9658
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21100 8945 21128 9522
rect 21086 8936 21142 8945
rect 21086 8871 21142 8880
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 21100 8537 21128 8570
rect 21086 8528 21142 8537
rect 21086 8463 21142 8472
rect 20994 7576 21050 7585
rect 20994 7511 21050 7520
rect 21008 7478 21036 7511
rect 20996 7472 21048 7478
rect 20996 7414 21048 7420
rect 20994 6488 21050 6497
rect 20904 6452 20956 6458
rect 20994 6423 21050 6432
rect 20904 6394 20956 6400
rect 21008 5710 21036 6423
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20916 4185 20944 4558
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 20902 4176 20958 4185
rect 20902 4111 20958 4120
rect 20904 4072 20956 4078
rect 20904 4014 20956 4020
rect 20916 3738 20944 4014
rect 20812 3732 20864 3738
rect 20812 3674 20864 3680
rect 20904 3732 20956 3738
rect 20904 3674 20956 3680
rect 20720 3596 20772 3602
rect 20720 3538 20772 3544
rect 20626 3496 20682 3505
rect 20626 3431 20682 3440
rect 20732 3369 20760 3538
rect 20718 3360 20774 3369
rect 20718 3295 20774 3304
rect 20628 2984 20680 2990
rect 20626 2952 20628 2961
rect 20680 2952 20682 2961
rect 20456 2910 20576 2938
rect 20364 2746 20484 2774
rect 20260 1760 20312 1766
rect 20260 1702 20312 1708
rect 20168 1420 20220 1426
rect 20168 1362 20220 1368
rect 20456 800 20484 2746
rect 20548 2582 20576 2910
rect 20626 2887 20682 2896
rect 20720 2848 20772 2854
rect 20640 2796 20720 2802
rect 20640 2790 20772 2796
rect 20640 2774 20760 2790
rect 20536 2576 20588 2582
rect 20640 2553 20668 2774
rect 20536 2518 20588 2524
rect 20626 2544 20682 2553
rect 20626 2479 20682 2488
rect 21008 800 21036 4422
rect 21100 4078 21128 8463
rect 21192 6254 21220 10406
rect 21272 9376 21324 9382
rect 21272 9318 21324 9324
rect 21180 6248 21232 6254
rect 21180 6190 21232 6196
rect 21284 4146 21312 9318
rect 21364 8900 21416 8906
rect 21364 8842 21416 8848
rect 21272 4140 21324 4146
rect 21272 4082 21324 4088
rect 21088 4072 21140 4078
rect 21088 4014 21140 4020
rect 21376 3534 21404 8842
rect 21468 5166 21496 11222
rect 21560 7274 21588 12922
rect 21638 11656 21694 11665
rect 21638 11591 21694 11600
rect 21652 11082 21680 11591
rect 21640 11076 21692 11082
rect 21640 11018 21692 11024
rect 21548 7268 21600 7274
rect 21548 7210 21600 7216
rect 21456 5160 21508 5166
rect 21456 5102 21508 5108
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 21364 3528 21416 3534
rect 21364 3470 21416 3476
rect 21088 2440 21140 2446
rect 21088 2382 21140 2388
rect 21364 2440 21416 2446
rect 21364 2382 21416 2388
rect 18972 740 19024 746
rect 18972 682 19024 688
rect 19338 0 19394 800
rect 19890 0 19946 800
rect 20442 0 20498 800
rect 20994 0 21050 800
rect 21100 610 21128 2382
rect 21376 1601 21404 2382
rect 21362 1592 21418 1601
rect 21362 1527 21418 1536
rect 21560 800 21588 3946
rect 21652 3505 21680 11018
rect 22008 7472 22060 7478
rect 22008 7414 22060 7420
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 21638 3496 21694 3505
rect 21638 3431 21694 3440
rect 21088 604 21140 610
rect 21088 546 21140 552
rect 21546 0 21602 800
rect 21836 649 21864 5646
rect 22020 2553 22048 7414
rect 22112 3466 22140 13926
rect 22284 7268 22336 7274
rect 22284 7210 22336 7216
rect 22100 3460 22152 3466
rect 22100 3402 22152 3408
rect 22100 2848 22152 2854
rect 22100 2790 22152 2796
rect 22006 2544 22062 2553
rect 22006 2479 22062 2488
rect 22112 800 22140 2790
rect 22296 2378 22324 7210
rect 22652 2916 22704 2922
rect 22652 2858 22704 2864
rect 22284 2372 22336 2378
rect 22284 2314 22336 2320
rect 22664 800 22692 2858
rect 21822 640 21878 649
rect 21822 575 21878 584
rect 22098 0 22154 800
rect 22650 0 22706 800
<< via2 >>
rect 1582 19760 1638 19816
rect 1490 17176 1546 17232
rect 1398 5752 1454 5808
rect 2134 18420 2190 18456
rect 2134 18400 2136 18420
rect 2136 18400 2188 18420
rect 2188 18400 2190 18420
rect 2410 19216 2466 19272
rect 2410 18572 2412 18592
rect 2412 18572 2464 18592
rect 2464 18572 2466 18592
rect 2410 18536 2466 18572
rect 2870 19760 2926 19816
rect 2594 18400 2650 18456
rect 2962 17720 3018 17776
rect 4342 21392 4398 21448
rect 3882 20440 3938 20496
rect 3238 19352 3294 19408
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3514 17620 3516 17640
rect 3516 17620 3568 17640
rect 3568 17620 3570 17640
rect 3514 17584 3570 17620
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3330 15000 3386 15056
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 4066 19080 4122 19136
rect 4066 18828 4122 18864
rect 4066 18808 4068 18828
rect 4068 18808 4120 18828
rect 4120 18808 4122 18828
rect 3238 13776 3294 13832
rect 2042 5616 2098 5672
rect 1858 2352 1914 2408
rect 1582 856 1638 912
rect 2318 4120 2374 4176
rect 2226 1944 2282 2000
rect 2594 4140 2650 4176
rect 2594 4120 2596 4140
rect 2596 4120 2648 4140
rect 2648 4120 2650 4140
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3238 5616 3294 5672
rect 2686 1808 2742 1864
rect 3054 3984 3110 4040
rect 2778 1536 2834 1592
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 4526 20032 4582 20088
rect 4158 14320 4214 14376
rect 3974 11736 4030 11792
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 4802 19896 4858 19952
rect 4802 19624 4858 19680
rect 5170 20984 5226 21040
rect 5078 20304 5134 20360
rect 5722 21120 5778 21176
rect 4894 19216 4950 19272
rect 4802 17176 4858 17232
rect 5078 18964 5134 19000
rect 5078 18944 5080 18964
rect 5080 18944 5132 18964
rect 5132 18944 5134 18964
rect 4986 17584 5042 17640
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 2042 584 2098 640
rect 3882 3576 3938 3632
rect 4066 3848 4122 3904
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 3974 1400 4030 1456
rect 4434 5652 4436 5672
rect 4436 5652 4488 5672
rect 4488 5652 4490 5672
rect 4434 5616 4490 5652
rect 4986 16788 5042 16824
rect 4986 16768 4988 16788
rect 4988 16768 5040 16788
rect 5040 16768 5042 16788
rect 5170 17876 5226 17912
rect 5170 17856 5172 17876
rect 5172 17856 5224 17876
rect 5224 17856 5226 17876
rect 5354 18964 5410 19000
rect 5354 18944 5356 18964
rect 5356 18944 5408 18964
rect 5408 18944 5410 18964
rect 5354 18708 5356 18728
rect 5356 18708 5408 18728
rect 5408 18708 5410 18728
rect 5354 18672 5410 18708
rect 5354 17992 5410 18048
rect 5078 16632 5134 16688
rect 4986 16496 5042 16552
rect 5354 17076 5356 17096
rect 5356 17076 5408 17096
rect 5408 17076 5410 17096
rect 5354 17040 5410 17076
rect 6734 21256 6790 21312
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6090 19796 6092 19816
rect 6092 19796 6144 19816
rect 6144 19796 6146 19816
rect 5630 15988 5632 16008
rect 5632 15988 5684 16008
rect 5684 15988 5686 16008
rect 5630 15952 5686 15988
rect 5630 15816 5686 15872
rect 4802 6860 4858 6896
rect 4802 6840 4804 6860
rect 4804 6840 4856 6860
rect 4856 6840 4858 6860
rect 4802 4156 4804 4176
rect 4804 4156 4856 4176
rect 4856 4156 4858 4176
rect 4802 4120 4858 4156
rect 4710 3712 4766 3768
rect 4894 3576 4950 3632
rect 4894 3476 4896 3496
rect 4896 3476 4948 3496
rect 4948 3476 4950 3496
rect 4894 3440 4950 3476
rect 4986 3304 5042 3360
rect 4802 2760 4858 2816
rect 4894 2488 4950 2544
rect 5262 6976 5318 7032
rect 5262 3440 5318 3496
rect 5262 2896 5318 2952
rect 6090 19760 6146 19796
rect 6550 19760 6606 19816
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 5906 18264 5962 18320
rect 5446 5244 5448 5264
rect 5448 5244 5500 5264
rect 5500 5244 5502 5264
rect 5446 5208 5502 5244
rect 5446 4820 5502 4856
rect 5446 4800 5448 4820
rect 5448 4800 5500 4820
rect 5500 4800 5502 4820
rect 5538 4120 5594 4176
rect 5446 4004 5502 4040
rect 5446 3984 5448 4004
rect 5448 3984 5500 4004
rect 5500 3984 5502 4004
rect 6458 19080 6514 19136
rect 6090 18944 6146 19000
rect 6826 20576 6882 20632
rect 6918 20440 6974 20496
rect 6550 18536 6606 18592
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6550 17332 6606 17368
rect 6550 17312 6552 17332
rect 6552 17312 6604 17332
rect 6604 17312 6606 17332
rect 6550 16496 6606 16552
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 7010 19896 7066 19952
rect 6918 19372 6974 19408
rect 6918 19352 6920 19372
rect 6920 19352 6972 19372
rect 6972 19352 6974 19372
rect 6826 19080 6882 19136
rect 6826 18672 6882 18728
rect 6918 18400 6974 18456
rect 6826 18148 6882 18184
rect 6826 18128 6828 18148
rect 6828 18128 6880 18148
rect 6880 18128 6882 18148
rect 7286 18672 7342 18728
rect 8482 21664 8538 21720
rect 7746 20204 7748 20224
rect 7748 20204 7800 20224
rect 7800 20204 7802 20224
rect 7746 20168 7802 20204
rect 6734 16360 6790 16416
rect 6642 16224 6698 16280
rect 6458 16088 6514 16144
rect 6550 15952 6606 16008
rect 6182 15428 6238 15464
rect 6182 15408 6184 15428
rect 6184 15408 6236 15428
rect 6236 15408 6238 15428
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6458 14592 6514 14648
rect 6642 15816 6698 15872
rect 5906 9868 5908 9888
rect 5908 9868 5960 9888
rect 5960 9868 5962 9888
rect 5906 9832 5962 9868
rect 5814 5888 5870 5944
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 6642 14456 6698 14512
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6918 15272 6974 15328
rect 6826 11600 6882 11656
rect 7470 17992 7526 18048
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6550 8900 6606 8936
rect 6550 8880 6552 8900
rect 6552 8880 6604 8900
rect 6604 8880 6606 8900
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6550 7828 6552 7848
rect 6552 7828 6604 7848
rect 6604 7828 6606 7848
rect 6550 7792 6606 7828
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 5998 5752 6054 5808
rect 5722 5480 5778 5536
rect 6550 6196 6552 6216
rect 6552 6196 6604 6216
rect 6604 6196 6606 6216
rect 6550 6160 6606 6196
rect 6734 9832 6790 9888
rect 6826 9424 6882 9480
rect 7194 13368 7250 13424
rect 7194 13132 7196 13152
rect 7196 13132 7248 13152
rect 7248 13132 7250 13152
rect 7194 13096 7250 13132
rect 7562 17448 7618 17504
rect 7562 17176 7618 17232
rect 7286 12824 7342 12880
rect 6734 6704 6790 6760
rect 6734 6452 6790 6488
rect 6734 6432 6736 6452
rect 6736 6432 6788 6452
rect 6788 6432 6790 6452
rect 6550 5616 6606 5672
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 5906 5344 5962 5400
rect 5722 3984 5778 4040
rect 5722 3712 5778 3768
rect 5446 3032 5502 3088
rect 7102 9580 7158 9616
rect 7102 9560 7104 9580
rect 7104 9560 7156 9580
rect 7156 9560 7158 9580
rect 6918 7928 6974 7984
rect 6458 4528 6514 4584
rect 6550 4428 6552 4448
rect 6552 4428 6604 4448
rect 6604 4428 6606 4448
rect 6550 4392 6606 4428
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6274 3712 6330 3768
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 5906 2644 5962 2680
rect 5906 2624 5908 2644
rect 5908 2624 5960 2644
rect 5960 2624 5962 2644
rect 6274 2624 6330 2680
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 6550 1672 6606 1728
rect 6734 4936 6790 4992
rect 6826 4156 6828 4176
rect 6828 4156 6880 4176
rect 6880 4156 6882 4176
rect 6826 4120 6882 4156
rect 7102 7384 7158 7440
rect 7286 9152 7342 9208
rect 8206 19352 8262 19408
rect 8574 20032 8630 20088
rect 8022 19080 8078 19136
rect 8206 17992 8262 18048
rect 8022 17176 8078 17232
rect 7746 12688 7802 12744
rect 7654 12316 7656 12336
rect 7656 12316 7708 12336
rect 7708 12316 7710 12336
rect 7654 12280 7710 12316
rect 7654 12144 7710 12200
rect 7654 10784 7710 10840
rect 7746 10532 7802 10568
rect 7746 10512 7748 10532
rect 7748 10512 7800 10532
rect 7800 10512 7802 10532
rect 7562 8780 7564 8800
rect 7564 8780 7616 8800
rect 7616 8780 7618 8800
rect 7562 8744 7618 8780
rect 7286 8336 7342 8392
rect 7378 7520 7434 7576
rect 7470 7248 7526 7304
rect 7746 8472 7802 8528
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 9586 21800 9642 21856
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8574 17992 8630 18048
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8022 14864 8078 14920
rect 8114 12980 8170 13016
rect 8114 12960 8116 12980
rect 8116 12960 8168 12980
rect 8168 12960 8170 12980
rect 8114 11736 8170 11792
rect 7930 9988 7986 10024
rect 7930 9968 7932 9988
rect 7932 9968 7984 9988
rect 7984 9968 7986 9988
rect 8114 11192 8170 11248
rect 8482 15000 8538 15056
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 9402 18808 9458 18864
rect 9402 18536 9458 18592
rect 9770 20984 9826 21040
rect 9954 20984 10010 21040
rect 10230 20576 10286 20632
rect 9586 19080 9642 19136
rect 9494 18400 9550 18456
rect 9862 18400 9918 18456
rect 9402 17992 9458 18048
rect 9402 17856 9458 17912
rect 9402 17448 9458 17504
rect 9770 17448 9826 17504
rect 9770 17332 9826 17368
rect 9770 17312 9772 17332
rect 9772 17312 9824 17332
rect 9824 17312 9826 17332
rect 9218 15544 9274 15600
rect 9770 16360 9826 16416
rect 9770 16088 9826 16144
rect 9402 15136 9458 15192
rect 8574 13268 8576 13288
rect 8576 13268 8628 13288
rect 8628 13268 8630 13288
rect 8574 13232 8630 13268
rect 8574 12280 8630 12336
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 9402 14864 9458 14920
rect 10414 21936 10470 21992
rect 10414 21120 10470 21176
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11794 20576 11850 20632
rect 10782 20032 10838 20088
rect 10046 16768 10102 16824
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 9126 11872 9182 11928
rect 9126 11464 9182 11520
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8298 10648 8354 10704
rect 8114 10104 8170 10160
rect 8390 9580 8446 9616
rect 8390 9560 8392 9580
rect 8392 9560 8444 9580
rect 8444 9560 8446 9580
rect 8574 11056 8630 11112
rect 9126 10376 9182 10432
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 9126 10240 9182 10296
rect 9126 9832 9182 9888
rect 8666 9696 8722 9752
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8666 9016 8722 9072
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 7194 6024 7250 6080
rect 7286 5752 7342 5808
rect 7470 6296 7526 6352
rect 6826 3984 6882 4040
rect 6734 3340 6736 3360
rect 6736 3340 6788 3360
rect 6788 3340 6790 3360
rect 6734 3304 6790 3340
rect 6734 3168 6790 3224
rect 6826 2624 6882 2680
rect 7654 5208 7710 5264
rect 7654 4684 7710 4720
rect 7654 4664 7656 4684
rect 7656 4664 7708 4684
rect 7708 4664 7710 4684
rect 7286 2644 7342 2680
rect 7286 2624 7288 2644
rect 7288 2624 7340 2644
rect 7340 2624 7342 2644
rect 7010 1264 7066 1320
rect 8390 6704 8446 6760
rect 8206 5616 8262 5672
rect 7838 720 7894 776
rect 8022 5344 8078 5400
rect 8114 5072 8170 5128
rect 8022 2760 8078 2816
rect 9126 7520 9182 7576
rect 9126 7112 9182 7168
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 9402 12552 9458 12608
rect 9678 13368 9734 13424
rect 9586 12960 9642 13016
rect 9586 12552 9642 12608
rect 9310 6296 9366 6352
rect 8574 5888 8630 5944
rect 9218 6024 9274 6080
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 9218 5888 9274 5944
rect 8482 4528 8538 4584
rect 8298 3168 8354 3224
rect 9126 5636 9182 5672
rect 9126 5616 9128 5636
rect 9128 5616 9180 5636
rect 9180 5616 9182 5636
rect 9126 4936 9182 4992
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 9310 5616 9366 5672
rect 10322 17484 10324 17504
rect 10324 17484 10376 17504
rect 10376 17484 10378 17504
rect 10322 17448 10378 17484
rect 10322 17176 10378 17232
rect 10322 16360 10378 16416
rect 10322 16224 10378 16280
rect 10322 15952 10378 16008
rect 10046 15272 10102 15328
rect 10782 19488 10838 19544
rect 10874 19080 10930 19136
rect 10966 18400 11022 18456
rect 11794 20304 11850 20360
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11334 17992 11390 18048
rect 11242 17756 11244 17776
rect 11244 17756 11296 17776
rect 11296 17756 11298 17776
rect 11242 17720 11298 17756
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 10782 16632 10838 16688
rect 11702 16632 11758 16688
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 10782 14728 10838 14784
rect 10782 14320 10838 14376
rect 10966 14340 11022 14376
rect 10966 14320 10968 14340
rect 10968 14320 11020 14340
rect 11020 14320 11022 14340
rect 11886 15544 11942 15600
rect 12162 19216 12218 19272
rect 13082 20032 13138 20088
rect 13082 19760 13138 19816
rect 12070 17312 12126 17368
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 10414 13776 10470 13832
rect 10046 12824 10102 12880
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11794 13096 11850 13152
rect 11794 12552 11850 12608
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11150 10784 11206 10840
rect 10322 9696 10378 9752
rect 9494 6296 9550 6352
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 10782 9288 10838 9344
rect 9862 6976 9918 7032
rect 9310 4800 9366 4856
rect 8758 4528 8814 4584
rect 8666 3984 8722 4040
rect 9402 4548 9458 4584
rect 9402 4528 9404 4548
rect 9404 4528 9456 4548
rect 9456 4528 9458 4548
rect 9310 4256 9366 4312
rect 9218 3848 9274 3904
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 8298 1264 8354 1320
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 8942 1536 8998 1592
rect 9586 3168 9642 3224
rect 9586 2896 9642 2952
rect 9954 3984 10010 4040
rect 9770 3476 9772 3496
rect 9772 3476 9824 3496
rect 9824 3476 9826 3496
rect 9770 3440 9826 3476
rect 9954 3304 10010 3360
rect 9402 2644 9458 2680
rect 9402 2624 9404 2644
rect 9404 2624 9456 2644
rect 9456 2624 9458 2644
rect 9218 2488 9274 2544
rect 9586 2624 9642 2680
rect 9494 2080 9550 2136
rect 10598 7384 10654 7440
rect 10598 6432 10654 6488
rect 10966 8472 11022 8528
rect 11058 7656 11114 7712
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11242 8472 11298 8528
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11058 6332 11060 6352
rect 11060 6332 11112 6352
rect 11112 6332 11114 6352
rect 10414 6024 10470 6080
rect 11058 6296 11114 6332
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 14186 20984 14242 21040
rect 12438 17448 12494 17504
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 13542 19080 13598 19136
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 14462 18808 14518 18864
rect 14370 17992 14426 18048
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13726 16768 13782 16824
rect 13726 15544 13782 15600
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 14370 16768 14426 16824
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 12622 15136 12678 15192
rect 13266 14900 13268 14920
rect 13268 14900 13320 14920
rect 13320 14900 13322 14920
rect 13266 14864 13322 14900
rect 13358 13504 13414 13560
rect 13726 14592 13782 14648
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13634 13368 13690 13424
rect 13358 12960 13414 13016
rect 13542 12724 13544 12744
rect 13544 12724 13596 12744
rect 13596 12724 13598 12744
rect 13542 12688 13598 12724
rect 12346 10240 12402 10296
rect 13542 11872 13598 11928
rect 13542 11600 13598 11656
rect 12806 10376 12862 10432
rect 18694 22208 18750 22264
rect 15290 20576 15346 20632
rect 15842 21528 15898 21584
rect 15842 20984 15898 21040
rect 15750 20460 15806 20496
rect 15750 20440 15752 20460
rect 15752 20440 15804 20460
rect 15804 20440 15806 20460
rect 15198 20032 15254 20088
rect 16946 21256 17002 21312
rect 15014 19896 15070 19952
rect 14830 15680 14886 15736
rect 14830 15136 14886 15192
rect 14278 14184 14334 14240
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 14738 14184 14794 14240
rect 14554 12708 14610 12744
rect 14554 12688 14556 12708
rect 14556 12688 14608 12708
rect 14608 12688 14610 12708
rect 15658 19896 15714 19952
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 15658 19624 15714 19680
rect 15566 18672 15622 18728
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 17038 19488 17094 19544
rect 17866 21528 17922 21584
rect 17774 21392 17830 21448
rect 17314 19624 17370 19680
rect 15474 17584 15530 17640
rect 15290 17040 15346 17096
rect 15290 15952 15346 16008
rect 14370 11600 14426 11656
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 11978 7520 12034 7576
rect 11978 7248 12034 7304
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11794 5344 11850 5400
rect 11794 4936 11850 4992
rect 13082 8744 13138 8800
rect 12806 8608 12862 8664
rect 12346 7248 12402 7304
rect 12438 6976 12494 7032
rect 12346 6840 12402 6896
rect 12254 6568 12310 6624
rect 12162 4256 12218 4312
rect 11978 3848 12034 3904
rect 11978 3576 12034 3632
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11702 2524 11704 2544
rect 11704 2524 11756 2544
rect 11756 2524 11758 2544
rect 11702 2488 11758 2524
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12346 3984 12402 4040
rect 12346 3576 12402 3632
rect 12346 3168 12402 3224
rect 12070 1536 12126 1592
rect 13174 6568 13230 6624
rect 12714 3732 12770 3768
rect 12714 3712 12716 3732
rect 12716 3712 12768 3732
rect 12768 3712 12770 3732
rect 12806 2760 12862 2816
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13542 10124 13598 10160
rect 13542 10104 13544 10124
rect 13544 10104 13596 10124
rect 13596 10104 13598 10124
rect 13726 9832 13782 9888
rect 13450 7656 13506 7712
rect 13450 7384 13506 7440
rect 13450 6568 13506 6624
rect 13450 6296 13506 6352
rect 13358 6024 13414 6080
rect 13358 5480 13414 5536
rect 14646 12008 14702 12064
rect 14554 10240 14610 10296
rect 14462 10104 14518 10160
rect 13726 9288 13782 9344
rect 13726 9152 13782 9208
rect 13726 7384 13782 7440
rect 13634 6840 13690 6896
rect 13726 5888 13782 5944
rect 13082 3304 13138 3360
rect 13358 3848 13414 3904
rect 12622 1400 12678 1456
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 15750 16088 15806 16144
rect 15566 15952 15622 16008
rect 15566 13232 15622 13288
rect 14738 10512 14794 10568
rect 14002 8608 14058 8664
rect 14462 9152 14518 9208
rect 14370 8780 14372 8800
rect 14372 8780 14424 8800
rect 14424 8780 14426 8800
rect 14370 8744 14426 8780
rect 14370 8608 14426 8664
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 14370 8200 14426 8256
rect 14370 7112 14426 7168
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 15198 9868 15200 9888
rect 15200 9868 15252 9888
rect 15252 9868 15254 9888
rect 15198 9832 15254 9868
rect 15106 7520 15162 7576
rect 14646 6860 14702 6896
rect 14646 6840 14648 6860
rect 14648 6840 14700 6860
rect 14700 6840 14702 6860
rect 14554 6296 14610 6352
rect 14370 6024 14426 6080
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 14186 4528 14242 4584
rect 14094 4256 14150 4312
rect 14554 6160 14610 6216
rect 14738 6296 14794 6352
rect 15014 7112 15070 7168
rect 15198 6432 15254 6488
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 13910 3052 13966 3088
rect 13910 3032 13912 3052
rect 13912 3032 13964 3052
rect 13964 3032 13966 3052
rect 14462 3984 14518 4040
rect 15382 5208 15438 5264
rect 15382 4936 15438 4992
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 13818 2624 13874 2680
rect 15290 4392 15346 4448
rect 15014 2896 15070 2952
rect 15014 1672 15070 1728
rect 15198 3712 15254 3768
rect 15290 3576 15346 3632
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 17130 18536 17186 18592
rect 17038 17720 17094 17776
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16670 16768 16726 16824
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16026 13504 16082 13560
rect 16026 12960 16082 13016
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 17130 14320 17186 14376
rect 17590 19352 17646 19408
rect 18142 21120 18198 21176
rect 20810 22616 20866 22672
rect 18326 21256 18382 21312
rect 17682 18400 17738 18456
rect 18050 19352 18106 19408
rect 17958 18808 18014 18864
rect 17682 16904 17738 16960
rect 17866 17448 17922 17504
rect 18510 20712 18566 20768
rect 18602 20032 18658 20088
rect 19890 21800 19946 21856
rect 20442 21664 20498 21720
rect 19522 20984 19578 21040
rect 18878 19896 18934 19952
rect 18142 18128 18198 18184
rect 18326 18128 18382 18184
rect 18142 16768 18198 16824
rect 17774 16632 17830 16688
rect 17590 16088 17646 16144
rect 16118 11056 16174 11112
rect 16026 10920 16082 10976
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16394 11872 16450 11928
rect 16394 11600 16450 11656
rect 16026 10104 16082 10160
rect 16854 11192 16910 11248
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16394 8744 16450 8800
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16302 7656 16358 7712
rect 16302 7112 16358 7168
rect 16118 5480 16174 5536
rect 15842 3576 15898 3632
rect 15658 3168 15714 3224
rect 15474 2896 15530 2952
rect 15566 2644 15622 2680
rect 15566 2624 15568 2644
rect 15568 2624 15620 2644
rect 15620 2624 15622 2644
rect 15842 3032 15898 3088
rect 16026 3440 16082 3496
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 17314 9152 17370 9208
rect 16946 7112 17002 7168
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16578 4528 16634 4584
rect 16854 4528 16910 4584
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 17038 1808 17094 1864
rect 17038 1672 17094 1728
rect 17866 13368 17922 13424
rect 17958 12960 18014 13016
rect 18050 12144 18106 12200
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19798 20460 19854 20496
rect 20810 20848 20866 20904
rect 19798 20440 19800 20460
rect 19800 20440 19852 20460
rect 19852 20440 19854 20460
rect 19246 19896 19302 19952
rect 18786 16088 18842 16144
rect 18234 13232 18290 13288
rect 17958 10684 17960 10704
rect 17960 10684 18012 10704
rect 18012 10684 18014 10704
rect 17958 10648 18014 10684
rect 18602 15680 18658 15736
rect 18694 15580 18696 15600
rect 18696 15580 18748 15600
rect 18748 15580 18750 15600
rect 18694 15544 18750 15580
rect 18786 15136 18842 15192
rect 18694 14900 18696 14920
rect 18696 14900 18748 14920
rect 18748 14900 18750 14920
rect 18694 14864 18750 14900
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19522 17604 19578 17640
rect 19522 17584 19524 17604
rect 19524 17584 19576 17604
rect 19576 17584 19578 17604
rect 19522 17176 19578 17232
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19062 15544 19118 15600
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19430 14456 19486 14512
rect 19614 14612 19670 14648
rect 19614 14592 19616 14612
rect 19616 14592 19668 14612
rect 19668 14592 19670 14612
rect 18970 13640 19026 13696
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 17958 9968 18014 10024
rect 17958 9152 18014 9208
rect 17958 9016 18014 9072
rect 17958 8608 18014 8664
rect 17866 8200 17922 8256
rect 18326 10376 18382 10432
rect 18418 10240 18474 10296
rect 18234 8744 18290 8800
rect 18050 8472 18106 8528
rect 17866 7792 17922 7848
rect 18050 7792 18106 7848
rect 17866 7520 17922 7576
rect 17774 7384 17830 7440
rect 17590 6876 17592 6896
rect 17592 6876 17644 6896
rect 17644 6876 17646 6896
rect 17590 6840 17646 6876
rect 17682 6704 17738 6760
rect 17590 6568 17646 6624
rect 17958 6976 18014 7032
rect 17958 6704 18014 6760
rect 17590 3848 17646 3904
rect 17130 1300 17132 1320
rect 17132 1300 17184 1320
rect 17184 1300 17186 1320
rect 17130 1264 17186 1300
rect 17590 3168 17646 3224
rect 18970 12688 19026 12744
rect 18602 10512 18658 10568
rect 18694 9968 18750 10024
rect 18234 7112 18290 7168
rect 18234 6840 18290 6896
rect 17866 4820 17922 4856
rect 17866 4800 17868 4820
rect 17868 4800 17920 4820
rect 17920 4800 17922 4820
rect 17866 3848 17922 3904
rect 17774 1536 17830 1592
rect 18050 4156 18052 4176
rect 18052 4156 18104 4176
rect 18104 4156 18106 4176
rect 18050 4120 18106 4156
rect 18050 3984 18106 4040
rect 18234 5752 18290 5808
rect 18970 9288 19026 9344
rect 18970 8336 19026 8392
rect 18602 7384 18658 7440
rect 18970 8064 19026 8120
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19522 12144 19578 12200
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19338 10104 19394 10160
rect 19982 18300 19984 18320
rect 19984 18300 20036 18320
rect 20036 18300 20038 18320
rect 19982 18264 20038 18300
rect 21270 19780 21326 19816
rect 21270 19760 21272 19780
rect 21272 19760 21324 19780
rect 21324 19760 21326 19780
rect 21086 19488 21142 19544
rect 20258 17040 20314 17096
rect 20258 16496 20314 16552
rect 19522 9560 19578 9616
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19154 7248 19210 7304
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 18602 6432 18658 6488
rect 18786 6160 18842 6216
rect 18694 5752 18750 5808
rect 18602 5228 18658 5264
rect 18602 5208 18604 5228
rect 18604 5208 18656 5228
rect 18656 5208 18658 5228
rect 18510 5072 18566 5128
rect 18326 2932 18328 2952
rect 18328 2932 18380 2952
rect 18380 2932 18382 2952
rect 18326 2896 18382 2932
rect 18326 2372 18382 2408
rect 18326 2352 18328 2372
rect 18328 2352 18380 2372
rect 18380 2352 18382 2372
rect 18694 3848 18750 3904
rect 18694 3576 18750 3632
rect 18970 6604 18972 6624
rect 18972 6604 19024 6624
rect 19024 6604 19026 6624
rect 18970 6568 19026 6604
rect 18970 6432 19026 6488
rect 18970 6024 19026 6080
rect 19706 7928 19762 7984
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19338 5636 19394 5672
rect 19338 5616 19340 5636
rect 19340 5616 19392 5636
rect 19392 5616 19394 5636
rect 19062 5208 19118 5264
rect 20810 18536 20866 18592
rect 20718 16496 20774 16552
rect 20718 15408 20774 15464
rect 20258 12824 20314 12880
rect 20258 12280 20314 12336
rect 20534 13368 20590 13424
rect 20166 9424 20222 9480
rect 19890 5108 19892 5128
rect 19892 5108 19944 5128
rect 19944 5108 19946 5128
rect 19890 5072 19946 5108
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19890 4664 19946 4720
rect 18878 4392 18934 4448
rect 18786 3168 18842 3224
rect 18510 856 18566 912
rect 19062 4528 19118 4584
rect 18970 3712 19026 3768
rect 18970 3576 19026 3632
rect 17958 176 18014 232
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19338 3304 19394 3360
rect 19430 3052 19486 3088
rect 19430 3032 19432 3052
rect 19432 3032 19484 3052
rect 19484 3032 19486 3052
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 19246 1944 19302 2000
rect 19246 1128 19302 1184
rect 19062 856 19118 912
rect 19706 992 19762 1048
rect 21086 15020 21142 15056
rect 21086 15000 21088 15020
rect 21088 15000 21140 15020
rect 21140 15000 21142 15020
rect 21270 17040 21326 17096
rect 21362 14184 21418 14240
rect 21270 13776 21326 13832
rect 21178 13232 21234 13288
rect 22006 13912 22062 13968
rect 20994 12008 21050 12064
rect 20718 11056 20774 11112
rect 20718 10784 20774 10840
rect 20718 9424 20774 9480
rect 20718 8744 20774 8800
rect 20626 6296 20682 6352
rect 21086 8880 21142 8936
rect 21086 8472 21142 8528
rect 20994 7520 21050 7576
rect 20994 6432 21050 6488
rect 20902 4120 20958 4176
rect 20626 3440 20682 3496
rect 20718 3304 20774 3360
rect 20626 2932 20628 2952
rect 20628 2932 20680 2952
rect 20680 2932 20682 2952
rect 20626 2896 20682 2932
rect 20626 2488 20682 2544
rect 21638 11600 21694 11656
rect 21362 1536 21418 1592
rect 21638 3440 21694 3496
rect 22006 2488 22062 2544
rect 21822 584 21878 640
<< metal3 >>
rect 20805 22674 20871 22677
rect 22200 22674 23000 22704
rect 20805 22672 23000 22674
rect 20805 22616 20810 22672
rect 20866 22616 23000 22672
rect 20805 22614 23000 22616
rect 20805 22611 20871 22614
rect 22200 22584 23000 22614
rect 18689 22266 18755 22269
rect 22200 22266 23000 22296
rect 18689 22264 23000 22266
rect 18689 22208 18694 22264
rect 18750 22208 23000 22264
rect 18689 22206 23000 22208
rect 18689 22203 18755 22206
rect 22200 22176 23000 22206
rect 5022 21932 5028 21996
rect 5092 21994 5098 21996
rect 10409 21994 10475 21997
rect 5092 21992 10475 21994
rect 5092 21936 10414 21992
rect 10470 21936 10475 21992
rect 5092 21934 10475 21936
rect 5092 21932 5098 21934
rect 10409 21931 10475 21934
rect 9581 21858 9647 21861
rect 19885 21858 19951 21861
rect 9581 21856 19951 21858
rect 9581 21800 9586 21856
rect 9642 21800 19890 21856
rect 19946 21800 19951 21856
rect 9581 21798 19951 21800
rect 9581 21795 9647 21798
rect 19885 21795 19951 21798
rect 8477 21722 8543 21725
rect 20437 21722 20503 21725
rect 22200 21722 23000 21752
rect 8477 21720 20503 21722
rect 8477 21664 8482 21720
rect 8538 21664 20442 21720
rect 20498 21664 20503 21720
rect 8477 21662 20503 21664
rect 8477 21659 8543 21662
rect 20437 21659 20503 21662
rect 20670 21662 23000 21722
rect 5390 21524 5396 21588
rect 5460 21586 5466 21588
rect 15837 21586 15903 21589
rect 5460 21584 15903 21586
rect 5460 21528 15842 21584
rect 15898 21528 15903 21584
rect 5460 21526 15903 21528
rect 5460 21524 5466 21526
rect 15837 21523 15903 21526
rect 17861 21586 17927 21589
rect 20670 21586 20730 21662
rect 22200 21632 23000 21662
rect 17861 21584 20730 21586
rect 17861 21528 17866 21584
rect 17922 21528 20730 21584
rect 17861 21526 20730 21528
rect 17861 21523 17927 21526
rect 4337 21450 4403 21453
rect 17769 21450 17835 21453
rect 4337 21448 17835 21450
rect 4337 21392 4342 21448
rect 4398 21392 17774 21448
rect 17830 21392 17835 21448
rect 4337 21390 17835 21392
rect 4337 21387 4403 21390
rect 17769 21387 17835 21390
rect 6729 21314 6795 21317
rect 16941 21314 17007 21317
rect 6729 21312 17007 21314
rect 6729 21256 6734 21312
rect 6790 21256 16946 21312
rect 17002 21256 17007 21312
rect 6729 21254 17007 21256
rect 6729 21251 6795 21254
rect 16941 21251 17007 21254
rect 18321 21314 18387 21317
rect 22200 21314 23000 21344
rect 18321 21312 23000 21314
rect 18321 21256 18326 21312
rect 18382 21256 23000 21312
rect 18321 21254 23000 21256
rect 18321 21251 18387 21254
rect 22200 21224 23000 21254
rect 5717 21178 5783 21181
rect 10409 21178 10475 21181
rect 18137 21178 18203 21181
rect 5717 21176 10242 21178
rect 5717 21120 5722 21176
rect 5778 21120 10242 21176
rect 5717 21118 10242 21120
rect 5717 21115 5783 21118
rect 5165 21042 5231 21045
rect 9765 21042 9831 21045
rect 9949 21042 10015 21045
rect 5165 21040 10015 21042
rect 5165 20984 5170 21040
rect 5226 20984 9770 21040
rect 9826 20984 9954 21040
rect 10010 20984 10015 21040
rect 5165 20982 10015 20984
rect 10182 21042 10242 21118
rect 10409 21176 18203 21178
rect 10409 21120 10414 21176
rect 10470 21120 18142 21176
rect 18198 21120 18203 21176
rect 10409 21118 18203 21120
rect 10409 21115 10475 21118
rect 18137 21115 18203 21118
rect 14181 21042 14247 21045
rect 10182 21040 14247 21042
rect 10182 20984 14186 21040
rect 14242 20984 14247 21040
rect 10182 20982 14247 20984
rect 5165 20979 5231 20982
rect 9765 20979 9831 20982
rect 9949 20979 10015 20982
rect 14181 20979 14247 20982
rect 15837 21042 15903 21045
rect 19517 21042 19583 21045
rect 15837 21040 19583 21042
rect 15837 20984 15842 21040
rect 15898 20984 19522 21040
rect 19578 20984 19583 21040
rect 15837 20982 19583 20984
rect 15837 20979 15903 20982
rect 19517 20979 19583 20982
rect 2262 20844 2268 20908
rect 2332 20906 2338 20908
rect 20805 20906 20871 20909
rect 2332 20904 20871 20906
rect 2332 20848 20810 20904
rect 20866 20848 20871 20904
rect 2332 20846 20871 20848
rect 2332 20844 2338 20846
rect 20805 20843 20871 20846
rect 18505 20770 18571 20773
rect 22200 20770 23000 20800
rect 18505 20768 23000 20770
rect 18505 20712 18510 20768
rect 18566 20712 23000 20768
rect 18505 20710 23000 20712
rect 18505 20707 18571 20710
rect 6142 20704 6462 20705
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 20639 6462 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 16538 20704 16858 20705
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 22200 20680 23000 20710
rect 16538 20639 16858 20640
rect 6821 20634 6887 20637
rect 10225 20634 10291 20637
rect 6686 20632 10291 20634
rect 6686 20576 6826 20632
rect 6882 20576 10230 20632
rect 10286 20576 10291 20632
rect 6686 20574 10291 20576
rect 3877 20498 3943 20501
rect 6686 20498 6746 20574
rect 6821 20571 6887 20574
rect 10225 20571 10291 20574
rect 11789 20634 11855 20637
rect 15285 20634 15351 20637
rect 11789 20632 15351 20634
rect 11789 20576 11794 20632
rect 11850 20576 15290 20632
rect 15346 20576 15351 20632
rect 11789 20574 15351 20576
rect 11789 20571 11855 20574
rect 15285 20571 15351 20574
rect 3877 20496 6746 20498
rect 3877 20440 3882 20496
rect 3938 20440 6746 20496
rect 3877 20438 6746 20440
rect 6913 20498 6979 20501
rect 15745 20498 15811 20501
rect 19793 20498 19859 20501
rect 6913 20496 15811 20498
rect 6913 20440 6918 20496
rect 6974 20440 15750 20496
rect 15806 20440 15811 20496
rect 6913 20438 15811 20440
rect 3877 20435 3943 20438
rect 6913 20435 6979 20438
rect 15745 20435 15811 20438
rect 15886 20496 19859 20498
rect 15886 20440 19798 20496
rect 19854 20440 19859 20496
rect 15886 20438 19859 20440
rect 5073 20362 5139 20365
rect 11789 20362 11855 20365
rect 5073 20360 11855 20362
rect 5073 20304 5078 20360
rect 5134 20304 11794 20360
rect 11850 20304 11855 20360
rect 5073 20302 11855 20304
rect 5073 20299 5139 20302
rect 11789 20299 11855 20302
rect 13670 20300 13676 20364
rect 13740 20362 13746 20364
rect 15886 20362 15946 20438
rect 19793 20435 19859 20438
rect 22200 20362 23000 20392
rect 13740 20302 15946 20362
rect 19014 20302 23000 20362
rect 13740 20300 13746 20302
rect 7230 20164 7236 20228
rect 7300 20226 7306 20228
rect 7741 20226 7807 20229
rect 7300 20224 7807 20226
rect 7300 20168 7746 20224
rect 7802 20168 7807 20224
rect 7300 20166 7807 20168
rect 7300 20164 7306 20166
rect 7741 20163 7807 20166
rect 3543 20160 3863 20161
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 20095 3863 20096
rect 8741 20160 9061 20161
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 20095 9061 20096
rect 13939 20160 14259 20161
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 20095 14259 20096
rect 4521 20090 4587 20093
rect 8569 20090 8635 20093
rect 4521 20088 8635 20090
rect 4521 20032 4526 20088
rect 4582 20032 8574 20088
rect 8630 20032 8635 20088
rect 4521 20030 8635 20032
rect 4521 20027 4587 20030
rect 8569 20027 8635 20030
rect 10777 20090 10843 20093
rect 13077 20090 13143 20093
rect 10777 20088 13143 20090
rect 10777 20032 10782 20088
rect 10838 20032 13082 20088
rect 13138 20032 13143 20088
rect 10777 20030 13143 20032
rect 10777 20027 10843 20030
rect 13077 20027 13143 20030
rect 15193 20090 15259 20093
rect 18597 20090 18663 20093
rect 15193 20088 18663 20090
rect 15193 20032 15198 20088
rect 15254 20032 18602 20088
rect 18658 20032 18663 20088
rect 15193 20030 18663 20032
rect 15193 20027 15259 20030
rect 18597 20027 18663 20030
rect 4797 19954 4863 19957
rect 2730 19952 4863 19954
rect 2730 19896 4802 19952
rect 4858 19896 4863 19952
rect 2730 19894 4863 19896
rect 1577 19818 1643 19821
rect 2730 19818 2790 19894
rect 4797 19891 4863 19894
rect 7005 19954 7071 19957
rect 15009 19954 15075 19957
rect 7005 19952 15075 19954
rect 7005 19896 7010 19952
rect 7066 19896 15014 19952
rect 15070 19896 15075 19952
rect 7005 19894 15075 19896
rect 7005 19891 7071 19894
rect 15009 19891 15075 19894
rect 15653 19954 15719 19957
rect 18873 19954 18939 19957
rect 15653 19952 18939 19954
rect 15653 19896 15658 19952
rect 15714 19896 18878 19952
rect 18934 19896 18939 19952
rect 15653 19894 18939 19896
rect 19014 19954 19074 20302
rect 22200 20272 23000 20302
rect 19137 20160 19457 20161
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 20095 19457 20096
rect 19241 19954 19307 19957
rect 19014 19952 19307 19954
rect 19014 19896 19246 19952
rect 19302 19896 19307 19952
rect 19014 19894 19307 19896
rect 15653 19891 15719 19894
rect 18873 19891 18939 19894
rect 19241 19891 19307 19894
rect 1577 19816 2790 19818
rect 1577 19760 1582 19816
rect 1638 19760 2790 19816
rect 1577 19758 2790 19760
rect 2865 19818 2931 19821
rect 6085 19818 6151 19821
rect 2865 19816 6151 19818
rect 2865 19760 2870 19816
rect 2926 19760 6090 19816
rect 6146 19760 6151 19816
rect 2865 19758 6151 19760
rect 1577 19755 1643 19758
rect 2865 19755 2931 19758
rect 6085 19755 6151 19758
rect 6545 19818 6611 19821
rect 13077 19818 13143 19821
rect 21265 19818 21331 19821
rect 22200 19818 23000 19848
rect 6545 19816 12450 19818
rect 6545 19760 6550 19816
rect 6606 19760 12450 19816
rect 6545 19758 12450 19760
rect 6545 19755 6611 19758
rect 4797 19684 4863 19685
rect 4797 19682 4844 19684
rect 2454 19622 2790 19682
rect 4752 19680 4844 19682
rect 4752 19624 4802 19680
rect 4752 19622 4844 19624
rect 2454 19277 2514 19622
rect 2730 19546 2790 19622
rect 4797 19620 4844 19622
rect 4908 19620 4914 19684
rect 12390 19682 12450 19758
rect 13077 19816 21331 19818
rect 13077 19760 13082 19816
rect 13138 19760 21270 19816
rect 21326 19760 21331 19816
rect 13077 19758 21331 19760
rect 13077 19755 13143 19758
rect 21265 19755 21331 19758
rect 21406 19758 23000 19818
rect 15653 19682 15719 19685
rect 12390 19680 15719 19682
rect 12390 19624 15658 19680
rect 15714 19624 15719 19680
rect 12390 19622 15719 19624
rect 4797 19619 4863 19620
rect 15653 19619 15719 19622
rect 17309 19682 17375 19685
rect 21406 19682 21466 19758
rect 22200 19728 23000 19758
rect 17309 19680 21466 19682
rect 17309 19624 17314 19680
rect 17370 19624 21466 19680
rect 17309 19622 21466 19624
rect 17309 19619 17375 19622
rect 6142 19616 6462 19617
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 19551 6462 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 16538 19616 16858 19617
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 19551 16858 19552
rect 5942 19546 5948 19548
rect 2730 19486 5948 19546
rect 5942 19484 5948 19486
rect 6012 19484 6018 19548
rect 7230 19484 7236 19548
rect 7300 19546 7306 19548
rect 10777 19546 10843 19549
rect 7300 19544 10843 19546
rect 7300 19488 10782 19544
rect 10838 19488 10843 19544
rect 7300 19486 10843 19488
rect 7300 19484 7306 19486
rect 10777 19483 10843 19486
rect 17033 19546 17099 19549
rect 17166 19546 17172 19548
rect 17033 19544 17172 19546
rect 17033 19488 17038 19544
rect 17094 19488 17172 19544
rect 17033 19486 17172 19488
rect 17033 19483 17099 19486
rect 17166 19484 17172 19486
rect 17236 19484 17242 19548
rect 20662 19484 20668 19548
rect 20732 19546 20738 19548
rect 21081 19546 21147 19549
rect 20732 19544 21147 19546
rect 20732 19488 21086 19544
rect 21142 19488 21147 19544
rect 20732 19486 21147 19488
rect 20732 19484 20738 19486
rect 21081 19483 21147 19486
rect 3233 19410 3299 19413
rect 6913 19410 6979 19413
rect 7782 19410 7788 19412
rect 3233 19408 7788 19410
rect 3233 19352 3238 19408
rect 3294 19352 6918 19408
rect 6974 19352 7788 19408
rect 3233 19350 7788 19352
rect 3233 19347 3299 19350
rect 6913 19347 6979 19350
rect 7782 19348 7788 19350
rect 7852 19348 7858 19412
rect 8201 19410 8267 19413
rect 17585 19410 17651 19413
rect 8201 19408 17651 19410
rect 8201 19352 8206 19408
rect 8262 19352 17590 19408
rect 17646 19352 17651 19408
rect 8201 19350 17651 19352
rect 8201 19347 8267 19350
rect 17585 19347 17651 19350
rect 18045 19410 18111 19413
rect 22200 19410 23000 19440
rect 18045 19408 23000 19410
rect 18045 19352 18050 19408
rect 18106 19352 23000 19408
rect 18045 19350 23000 19352
rect 18045 19347 18111 19350
rect 22200 19320 23000 19350
rect 2405 19272 2514 19277
rect 2405 19216 2410 19272
rect 2466 19216 2514 19272
rect 2405 19214 2514 19216
rect 4889 19274 4955 19277
rect 12157 19274 12223 19277
rect 4889 19272 12450 19274
rect 4889 19216 4894 19272
rect 4950 19216 12162 19272
rect 12218 19216 12450 19272
rect 4889 19214 12450 19216
rect 2405 19211 2471 19214
rect 4889 19211 4955 19214
rect 12157 19211 12223 19214
rect 4061 19138 4127 19141
rect 6453 19138 6519 19141
rect 4061 19136 6519 19138
rect 4061 19080 4066 19136
rect 4122 19080 6458 19136
rect 6514 19080 6519 19136
rect 4061 19078 6519 19080
rect 4061 19075 4127 19078
rect 6453 19075 6519 19078
rect 6821 19138 6887 19141
rect 8017 19138 8083 19141
rect 6821 19136 8083 19138
rect 6821 19080 6826 19136
rect 6882 19080 8022 19136
rect 8078 19080 8083 19136
rect 6821 19078 8083 19080
rect 6821 19075 6887 19078
rect 8017 19075 8083 19078
rect 9254 19076 9260 19140
rect 9324 19138 9330 19140
rect 9581 19138 9647 19141
rect 10869 19140 10935 19141
rect 10869 19138 10916 19140
rect 9324 19136 9647 19138
rect 9324 19080 9586 19136
rect 9642 19080 9647 19136
rect 9324 19078 9647 19080
rect 10824 19136 10916 19138
rect 10824 19080 10874 19136
rect 10824 19078 10916 19080
rect 9324 19076 9330 19078
rect 9581 19075 9647 19078
rect 10869 19076 10916 19078
rect 10980 19076 10986 19140
rect 12198 19076 12204 19140
rect 12268 19138 12274 19140
rect 12390 19138 12450 19214
rect 13537 19138 13603 19141
rect 12268 19136 13603 19138
rect 12268 19080 13542 19136
rect 13598 19080 13603 19136
rect 12268 19078 13603 19080
rect 12268 19076 12274 19078
rect 10869 19075 10935 19076
rect 13537 19075 13603 19078
rect 3543 19072 3863 19073
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 19007 3863 19008
rect 8741 19072 9061 19073
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 19007 9061 19008
rect 13939 19072 14259 19073
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 19007 14259 19008
rect 19137 19072 19457 19073
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 19007 19457 19008
rect 5073 19004 5139 19005
rect 5022 18940 5028 19004
rect 5092 19002 5139 19004
rect 5349 19004 5415 19005
rect 5349 19002 5396 19004
rect 5092 19000 5184 19002
rect 5134 18944 5184 19000
rect 5092 18942 5184 18944
rect 5304 19000 5396 19002
rect 5304 18944 5354 19000
rect 5304 18942 5396 18944
rect 5092 18940 5139 18942
rect 5073 18939 5139 18940
rect 5349 18940 5396 18942
rect 5460 18940 5466 19004
rect 5942 18940 5948 19004
rect 6012 19002 6018 19004
rect 6085 19002 6151 19005
rect 6012 19000 6151 19002
rect 6012 18944 6090 19000
rect 6146 18944 6151 19000
rect 6012 18942 6151 18944
rect 6012 18940 6018 18942
rect 5349 18939 5415 18940
rect 6085 18939 6151 18942
rect 9262 18942 13876 19002
rect 4061 18866 4127 18869
rect 9262 18866 9322 18942
rect 4061 18864 9322 18866
rect 4061 18808 4066 18864
rect 4122 18808 9322 18864
rect 4061 18806 9322 18808
rect 9397 18866 9463 18869
rect 13670 18866 13676 18868
rect 9397 18864 13676 18866
rect 9397 18808 9402 18864
rect 9458 18808 13676 18864
rect 9397 18806 13676 18808
rect 4061 18803 4127 18806
rect 9397 18803 9463 18806
rect 13670 18804 13676 18806
rect 13740 18804 13746 18868
rect 13816 18866 13876 18942
rect 14457 18866 14523 18869
rect 13816 18864 14523 18866
rect 13816 18808 14462 18864
rect 14518 18808 14523 18864
rect 13816 18806 14523 18808
rect 14457 18803 14523 18806
rect 17953 18866 18019 18869
rect 22200 18866 23000 18896
rect 17953 18864 23000 18866
rect 17953 18808 17958 18864
rect 18014 18808 23000 18864
rect 17953 18806 23000 18808
rect 17953 18803 18019 18806
rect 22200 18776 23000 18806
rect 5349 18730 5415 18733
rect 5758 18730 5764 18732
rect 2730 18728 5764 18730
rect 2730 18672 5354 18728
rect 5410 18672 5764 18728
rect 2730 18670 5764 18672
rect 2405 18594 2471 18597
rect 2730 18594 2790 18670
rect 5349 18667 5415 18670
rect 5758 18668 5764 18670
rect 5828 18668 5834 18732
rect 6821 18730 6887 18733
rect 5904 18728 6887 18730
rect 5904 18672 6826 18728
rect 6882 18672 6887 18728
rect 5904 18670 6887 18672
rect 2405 18592 2790 18594
rect 2405 18536 2410 18592
rect 2466 18536 2790 18592
rect 2405 18534 2790 18536
rect 2405 18531 2471 18534
rect 2129 18458 2195 18461
rect 2262 18458 2268 18460
rect 2129 18456 2268 18458
rect 2129 18400 2134 18456
rect 2190 18400 2268 18456
rect 2129 18398 2268 18400
rect 2129 18395 2195 18398
rect 2262 18396 2268 18398
rect 2332 18396 2338 18460
rect 2589 18458 2655 18461
rect 5904 18458 5964 18670
rect 6821 18667 6887 18670
rect 7281 18730 7347 18733
rect 15561 18730 15627 18733
rect 7281 18728 15627 18730
rect 7281 18672 7286 18728
rect 7342 18672 15566 18728
rect 15622 18672 15627 18728
rect 7281 18670 15627 18672
rect 7281 18667 7347 18670
rect 15561 18667 15627 18670
rect 6545 18594 6611 18597
rect 9397 18594 9463 18597
rect 6545 18592 9463 18594
rect 6545 18536 6550 18592
rect 6606 18536 9402 18592
rect 9458 18536 9463 18592
rect 6545 18534 9463 18536
rect 6545 18531 6611 18534
rect 9397 18531 9463 18534
rect 17125 18594 17191 18597
rect 20805 18594 20871 18597
rect 17125 18592 20871 18594
rect 17125 18536 17130 18592
rect 17186 18536 20810 18592
rect 20866 18536 20871 18592
rect 17125 18534 20871 18536
rect 17125 18531 17191 18534
rect 20805 18531 20871 18534
rect 6142 18528 6462 18529
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 18463 6462 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 16538 18528 16858 18529
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 18463 16858 18464
rect 2589 18456 5964 18458
rect 2589 18400 2594 18456
rect 2650 18400 5964 18456
rect 2589 18398 5964 18400
rect 6913 18458 6979 18461
rect 9489 18458 9555 18461
rect 9857 18458 9923 18461
rect 10961 18458 11027 18461
rect 6913 18456 11027 18458
rect 6913 18400 6918 18456
rect 6974 18400 9494 18456
rect 9550 18400 9862 18456
rect 9918 18400 10966 18456
rect 11022 18400 11027 18456
rect 6913 18398 11027 18400
rect 2589 18395 2655 18398
rect 6913 18395 6979 18398
rect 9489 18395 9555 18398
rect 9857 18395 9923 18398
rect 10961 18395 11027 18398
rect 17677 18458 17743 18461
rect 22200 18458 23000 18488
rect 17677 18456 23000 18458
rect 17677 18400 17682 18456
rect 17738 18400 23000 18456
rect 17677 18398 23000 18400
rect 17677 18395 17743 18398
rect 22200 18368 23000 18398
rect 5901 18322 5967 18325
rect 19977 18322 20043 18325
rect 5901 18320 20043 18322
rect 5901 18264 5906 18320
rect 5962 18264 19982 18320
rect 20038 18264 20043 18320
rect 5901 18262 20043 18264
rect 5901 18259 5967 18262
rect 19977 18259 20043 18262
rect 6821 18186 6887 18189
rect 18137 18186 18203 18189
rect 6821 18184 18203 18186
rect 6821 18128 6826 18184
rect 6882 18128 18142 18184
rect 18198 18128 18203 18184
rect 6821 18126 18203 18128
rect 6821 18123 6887 18126
rect 18137 18123 18203 18126
rect 18321 18186 18387 18189
rect 18321 18184 19626 18186
rect 18321 18128 18326 18184
rect 18382 18128 19626 18184
rect 18321 18126 19626 18128
rect 18321 18123 18387 18126
rect 5349 18050 5415 18053
rect 7465 18050 7531 18053
rect 8201 18050 8267 18053
rect 8569 18050 8635 18053
rect 5349 18048 8267 18050
rect 5349 17992 5354 18048
rect 5410 17992 7470 18048
rect 7526 17992 8206 18048
rect 8262 17992 8267 18048
rect 5349 17990 8267 17992
rect 5349 17987 5415 17990
rect 7465 17987 7531 17990
rect 8201 17987 8267 17990
rect 8526 18048 8635 18050
rect 8526 17992 8574 18048
rect 8630 17992 8635 18048
rect 8526 17987 8635 17992
rect 9397 18050 9463 18053
rect 11329 18050 11395 18053
rect 9397 18048 11395 18050
rect 9397 17992 9402 18048
rect 9458 17992 11334 18048
rect 11390 17992 11395 18048
rect 9397 17990 11395 17992
rect 9397 17987 9463 17990
rect 11329 17987 11395 17990
rect 14365 18050 14431 18053
rect 17534 18050 17540 18052
rect 14365 18048 17540 18050
rect 14365 17992 14370 18048
rect 14426 17992 17540 18048
rect 14365 17990 17540 17992
rect 14365 17987 14431 17990
rect 17534 17988 17540 17990
rect 17604 17988 17610 18052
rect 19566 18050 19626 18126
rect 22200 18050 23000 18080
rect 19566 17990 23000 18050
rect 3543 17984 3863 17985
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 17919 3863 17920
rect 5165 17914 5231 17917
rect 8526 17914 8586 17987
rect 8741 17984 9061 17985
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 17919 9061 17920
rect 13939 17984 14259 17985
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 17919 14259 17920
rect 19137 17984 19457 17985
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 22200 17960 23000 17990
rect 19137 17919 19457 17920
rect 5165 17912 8586 17914
rect 5165 17856 5170 17912
rect 5226 17856 8586 17912
rect 5165 17854 8586 17856
rect 9397 17914 9463 17917
rect 9397 17912 12450 17914
rect 9397 17856 9402 17912
rect 9458 17856 12450 17912
rect 9397 17854 12450 17856
rect 5165 17851 5231 17854
rect 9397 17851 9463 17854
rect 2957 17778 3023 17781
rect 11237 17778 11303 17781
rect 2957 17776 11303 17778
rect 2957 17720 2962 17776
rect 3018 17720 11242 17776
rect 11298 17720 11303 17776
rect 2957 17718 11303 17720
rect 12390 17778 12450 17854
rect 17033 17778 17099 17781
rect 12390 17776 17099 17778
rect 12390 17720 17038 17776
rect 17094 17720 17099 17776
rect 12390 17718 17099 17720
rect 2957 17715 3023 17718
rect 11237 17715 11303 17718
rect 17033 17715 17099 17718
rect 3509 17642 3575 17645
rect 4981 17642 5047 17645
rect 15469 17642 15535 17645
rect 19517 17642 19583 17645
rect 3509 17640 15535 17642
rect 3509 17584 3514 17640
rect 3570 17584 4986 17640
rect 5042 17584 15474 17640
rect 15530 17584 15535 17640
rect 3509 17582 15535 17584
rect 3509 17579 3575 17582
rect 4981 17579 5047 17582
rect 15469 17579 15535 17582
rect 15656 17640 19583 17642
rect 15656 17584 19522 17640
rect 19578 17584 19583 17640
rect 15656 17582 19583 17584
rect 7557 17506 7623 17509
rect 9397 17506 9463 17509
rect 7557 17504 9463 17506
rect 7557 17448 7562 17504
rect 7618 17448 9402 17504
rect 9458 17448 9463 17504
rect 7557 17446 9463 17448
rect 7557 17443 7623 17446
rect 9397 17443 9463 17446
rect 9765 17506 9831 17509
rect 10317 17506 10383 17509
rect 9765 17504 10383 17506
rect 9765 17448 9770 17504
rect 9826 17448 10322 17504
rect 10378 17448 10383 17504
rect 9765 17446 10383 17448
rect 9765 17443 9831 17446
rect 10317 17443 10383 17446
rect 12433 17506 12499 17509
rect 15656 17506 15716 17582
rect 19517 17579 19583 17582
rect 12433 17504 15716 17506
rect 12433 17448 12438 17504
rect 12494 17448 15716 17504
rect 12433 17446 15716 17448
rect 17861 17506 17927 17509
rect 22200 17506 23000 17536
rect 17861 17504 23000 17506
rect 17861 17448 17866 17504
rect 17922 17448 23000 17504
rect 17861 17446 23000 17448
rect 12433 17443 12499 17446
rect 17861 17443 17927 17446
rect 6142 17440 6462 17441
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 17375 6462 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 16538 17440 16858 17441
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 22200 17416 23000 17446
rect 16538 17375 16858 17376
rect 6545 17370 6611 17373
rect 9765 17370 9831 17373
rect 6545 17368 9831 17370
rect 6545 17312 6550 17368
rect 6606 17312 9770 17368
rect 9826 17312 9831 17368
rect 6545 17310 9831 17312
rect 6545 17307 6611 17310
rect 9765 17307 9831 17310
rect 12065 17370 12131 17373
rect 12065 17368 16314 17370
rect 12065 17312 12070 17368
rect 12126 17312 16314 17368
rect 12065 17310 16314 17312
rect 12065 17307 12131 17310
rect 0 17234 800 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 800 17174
rect 1485 17171 1551 17174
rect 4797 17234 4863 17237
rect 7557 17234 7623 17237
rect 4797 17232 7623 17234
rect 4797 17176 4802 17232
rect 4858 17176 7562 17232
rect 7618 17176 7623 17232
rect 4797 17174 7623 17176
rect 4797 17171 4863 17174
rect 7557 17171 7623 17174
rect 8017 17234 8083 17237
rect 9254 17234 9260 17236
rect 8017 17232 9260 17234
rect 8017 17176 8022 17232
rect 8078 17176 9260 17232
rect 8017 17174 9260 17176
rect 8017 17171 8083 17174
rect 9254 17172 9260 17174
rect 9324 17172 9330 17236
rect 10317 17234 10383 17237
rect 16254 17234 16314 17310
rect 19517 17234 19583 17237
rect 10317 17232 16130 17234
rect 10317 17176 10322 17232
rect 10378 17176 16130 17232
rect 10317 17174 16130 17176
rect 16254 17232 19583 17234
rect 16254 17176 19522 17232
rect 19578 17176 19583 17232
rect 16254 17174 19583 17176
rect 10317 17171 10383 17174
rect 5349 17098 5415 17101
rect 15285 17098 15351 17101
rect 16070 17098 16130 17174
rect 19517 17171 19583 17174
rect 20253 17098 20319 17101
rect 5349 17096 15946 17098
rect 5349 17040 5354 17096
rect 5410 17040 15290 17096
rect 15346 17040 15946 17096
rect 5349 17038 15946 17040
rect 16070 17096 20319 17098
rect 16070 17040 20258 17096
rect 20314 17040 20319 17096
rect 16070 17038 20319 17040
rect 5349 17035 5415 17038
rect 15285 17035 15351 17038
rect 15886 16962 15946 17038
rect 20253 17035 20319 17038
rect 21265 17098 21331 17101
rect 22200 17098 23000 17128
rect 21265 17096 23000 17098
rect 21265 17040 21270 17096
rect 21326 17040 23000 17096
rect 21265 17038 23000 17040
rect 21265 17035 21331 17038
rect 22200 17008 23000 17038
rect 17677 16962 17743 16965
rect 15886 16960 17743 16962
rect 15886 16904 17682 16960
rect 17738 16904 17743 16960
rect 15886 16902 17743 16904
rect 17677 16899 17743 16902
rect 3543 16896 3863 16897
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 16831 3863 16832
rect 8741 16896 9061 16897
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 16831 9061 16832
rect 13939 16896 14259 16897
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 16831 14259 16832
rect 19137 16896 19457 16897
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 16831 19457 16832
rect 4981 16828 5047 16829
rect 4981 16826 5028 16828
rect 4936 16824 5028 16826
rect 4936 16768 4986 16824
rect 4936 16766 5028 16768
rect 4981 16764 5028 16766
rect 5092 16764 5098 16828
rect 10041 16826 10107 16829
rect 13721 16826 13787 16829
rect 10041 16824 13787 16826
rect 10041 16768 10046 16824
rect 10102 16768 13726 16824
rect 13782 16768 13787 16824
rect 10041 16766 13787 16768
rect 4981 16763 5047 16764
rect 10041 16763 10107 16766
rect 13721 16763 13787 16766
rect 14365 16826 14431 16829
rect 16665 16826 16731 16829
rect 18137 16826 18203 16829
rect 14365 16824 18203 16826
rect 14365 16768 14370 16824
rect 14426 16768 16670 16824
rect 16726 16768 18142 16824
rect 18198 16768 18203 16824
rect 14365 16766 18203 16768
rect 14365 16763 14431 16766
rect 16665 16763 16731 16766
rect 18137 16763 18203 16766
rect 5073 16690 5139 16693
rect 8518 16690 8524 16692
rect 5073 16688 8524 16690
rect 5073 16632 5078 16688
rect 5134 16632 8524 16688
rect 5073 16630 8524 16632
rect 5073 16627 5139 16630
rect 8518 16628 8524 16630
rect 8588 16690 8594 16692
rect 10777 16690 10843 16693
rect 8588 16688 10843 16690
rect 8588 16632 10782 16688
rect 10838 16632 10843 16688
rect 8588 16630 10843 16632
rect 8588 16628 8594 16630
rect 10777 16627 10843 16630
rect 11697 16690 11763 16693
rect 17769 16690 17835 16693
rect 11697 16688 17835 16690
rect 11697 16632 11702 16688
rect 11758 16632 17774 16688
rect 17830 16632 17835 16688
rect 11697 16630 17835 16632
rect 11697 16627 11763 16630
rect 17769 16627 17835 16630
rect 4838 16492 4844 16556
rect 4908 16554 4914 16556
rect 4981 16554 5047 16557
rect 4908 16552 5047 16554
rect 4908 16496 4986 16552
rect 5042 16496 5047 16552
rect 4908 16494 5047 16496
rect 4908 16492 4914 16494
rect 4981 16491 5047 16494
rect 6545 16554 6611 16557
rect 6862 16554 6868 16556
rect 6545 16552 6868 16554
rect 6545 16496 6550 16552
rect 6606 16496 6868 16552
rect 6545 16494 6868 16496
rect 6545 16491 6611 16494
rect 6862 16492 6868 16494
rect 6932 16492 6938 16556
rect 20253 16554 20319 16557
rect 9446 16552 20319 16554
rect 9446 16496 20258 16552
rect 20314 16496 20319 16552
rect 9446 16494 20319 16496
rect 6729 16418 6795 16421
rect 9446 16418 9506 16494
rect 20253 16491 20319 16494
rect 20713 16554 20779 16557
rect 22200 16554 23000 16584
rect 20713 16552 23000 16554
rect 20713 16496 20718 16552
rect 20774 16496 23000 16552
rect 20713 16494 23000 16496
rect 20713 16491 20779 16494
rect 22200 16464 23000 16494
rect 6729 16416 9506 16418
rect 6729 16360 6734 16416
rect 6790 16360 9506 16416
rect 6729 16358 9506 16360
rect 9765 16418 9831 16421
rect 10317 16418 10383 16421
rect 9765 16416 10383 16418
rect 9765 16360 9770 16416
rect 9826 16360 10322 16416
rect 10378 16360 10383 16416
rect 9765 16358 10383 16360
rect 6729 16355 6795 16358
rect 9765 16355 9831 16358
rect 10317 16355 10383 16358
rect 6142 16352 6462 16353
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 16287 6462 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 16538 16352 16858 16353
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 16287 16858 16288
rect 6637 16282 6703 16285
rect 10317 16282 10383 16285
rect 6637 16280 10383 16282
rect 6637 16224 6642 16280
rect 6698 16224 10322 16280
rect 10378 16224 10383 16280
rect 6637 16222 10383 16224
rect 6637 16219 6703 16222
rect 10317 16219 10383 16222
rect 6453 16146 6519 16149
rect 9765 16146 9831 16149
rect 15745 16146 15811 16149
rect 17585 16146 17651 16149
rect 6453 16144 9831 16146
rect 6453 16088 6458 16144
rect 6514 16088 9770 16144
rect 9826 16088 9831 16144
rect 6453 16086 9831 16088
rect 6453 16083 6519 16086
rect 9765 16083 9831 16086
rect 10182 16144 17651 16146
rect 10182 16088 15750 16144
rect 15806 16088 17590 16144
rect 17646 16088 17651 16144
rect 10182 16086 17651 16088
rect 5625 16010 5691 16013
rect 6545 16010 6611 16013
rect 10182 16010 10242 16086
rect 15745 16083 15811 16086
rect 17585 16083 17651 16086
rect 18781 16146 18847 16149
rect 22200 16146 23000 16176
rect 18781 16144 23000 16146
rect 18781 16088 18786 16144
rect 18842 16088 23000 16144
rect 18781 16086 23000 16088
rect 18781 16083 18847 16086
rect 22200 16056 23000 16086
rect 5625 16008 10242 16010
rect 5625 15952 5630 16008
rect 5686 15952 6550 16008
rect 6606 15952 10242 16008
rect 5625 15950 10242 15952
rect 10317 16010 10383 16013
rect 15285 16010 15351 16013
rect 15561 16010 15627 16013
rect 10317 16008 15627 16010
rect 10317 15952 10322 16008
rect 10378 15952 15290 16008
rect 15346 15952 15566 16008
rect 15622 15952 15627 16008
rect 10317 15950 15627 15952
rect 5625 15947 5691 15950
rect 6545 15947 6611 15950
rect 10317 15947 10383 15950
rect 15285 15947 15351 15950
rect 15561 15947 15627 15950
rect 5625 15874 5691 15877
rect 6637 15874 6703 15877
rect 5625 15872 6703 15874
rect 5625 15816 5630 15872
rect 5686 15816 6642 15872
rect 6698 15816 6703 15872
rect 5625 15814 6703 15816
rect 5625 15811 5691 15814
rect 6637 15811 6703 15814
rect 3543 15808 3863 15809
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 15743 3863 15744
rect 8741 15808 9061 15809
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 15743 9061 15744
rect 13939 15808 14259 15809
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 15743 14259 15744
rect 19137 15808 19457 15809
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 15743 19457 15744
rect 14825 15738 14891 15741
rect 18597 15738 18663 15741
rect 14825 15736 18663 15738
rect 14825 15680 14830 15736
rect 14886 15680 18602 15736
rect 18658 15680 18663 15736
rect 14825 15678 18663 15680
rect 14825 15675 14891 15678
rect 18597 15675 18663 15678
rect 9213 15602 9279 15605
rect 11881 15602 11947 15605
rect 9213 15600 11947 15602
rect 9213 15544 9218 15600
rect 9274 15544 11886 15600
rect 11942 15544 11947 15600
rect 9213 15542 11947 15544
rect 9213 15539 9279 15542
rect 11881 15539 11947 15542
rect 13721 15602 13787 15605
rect 18689 15602 18755 15605
rect 13721 15600 18755 15602
rect 13721 15544 13726 15600
rect 13782 15544 18694 15600
rect 18750 15544 18755 15600
rect 13721 15542 18755 15544
rect 13721 15539 13787 15542
rect 18689 15539 18755 15542
rect 19057 15602 19123 15605
rect 22200 15602 23000 15632
rect 19057 15600 23000 15602
rect 19057 15544 19062 15600
rect 19118 15544 23000 15600
rect 19057 15542 23000 15544
rect 19057 15539 19123 15542
rect 22200 15512 23000 15542
rect 6177 15466 6243 15469
rect 20713 15466 20779 15469
rect 6177 15464 20779 15466
rect 6177 15408 6182 15464
rect 6238 15408 20718 15464
rect 20774 15408 20779 15464
rect 6177 15406 20779 15408
rect 6177 15403 6243 15406
rect 20713 15403 20779 15406
rect 6913 15330 6979 15333
rect 10041 15330 10107 15333
rect 6913 15328 10107 15330
rect 6913 15272 6918 15328
rect 6974 15272 10046 15328
rect 10102 15272 10107 15328
rect 6913 15270 10107 15272
rect 6913 15267 6979 15270
rect 10041 15267 10107 15270
rect 6142 15264 6462 15265
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 15199 6462 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 16538 15264 16858 15265
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 15199 16858 15200
rect 9397 15194 9463 15197
rect 8342 15192 9463 15194
rect 8342 15136 9402 15192
rect 9458 15136 9463 15192
rect 8342 15134 9463 15136
rect 3325 15058 3391 15061
rect 8342 15058 8402 15134
rect 9397 15131 9463 15134
rect 12617 15194 12683 15197
rect 14825 15194 14891 15197
rect 12617 15192 14891 15194
rect 12617 15136 12622 15192
rect 12678 15136 14830 15192
rect 14886 15136 14891 15192
rect 12617 15134 14891 15136
rect 12617 15131 12683 15134
rect 14825 15131 14891 15134
rect 18781 15194 18847 15197
rect 22200 15194 23000 15224
rect 18781 15192 23000 15194
rect 18781 15136 18786 15192
rect 18842 15136 23000 15192
rect 18781 15134 23000 15136
rect 18781 15131 18847 15134
rect 22200 15104 23000 15134
rect 3325 15056 8402 15058
rect 3325 15000 3330 15056
rect 3386 15000 8402 15056
rect 3325 14998 8402 15000
rect 8477 15058 8543 15061
rect 21081 15058 21147 15061
rect 8477 15056 21147 15058
rect 8477 15000 8482 15056
rect 8538 15000 21086 15056
rect 21142 15000 21147 15056
rect 8477 14998 21147 15000
rect 3325 14995 3391 14998
rect 8477 14995 8543 14998
rect 21081 14995 21147 14998
rect 8017 14922 8083 14925
rect 9397 14922 9463 14925
rect 13261 14922 13327 14925
rect 18689 14922 18755 14925
rect 8017 14920 9322 14922
rect 8017 14864 8022 14920
rect 8078 14864 9322 14920
rect 8017 14862 9322 14864
rect 8017 14859 8083 14862
rect 3543 14720 3863 14721
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 14655 3863 14656
rect 8741 14720 9061 14721
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 14655 9061 14656
rect 6453 14650 6519 14653
rect 9262 14650 9322 14862
rect 9397 14920 13327 14922
rect 9397 14864 9402 14920
rect 9458 14864 13266 14920
rect 13322 14864 13327 14920
rect 9397 14862 13327 14864
rect 9397 14859 9463 14862
rect 13261 14859 13327 14862
rect 13494 14920 18755 14922
rect 13494 14864 18694 14920
rect 18750 14864 18755 14920
rect 13494 14862 18755 14864
rect 10777 14786 10843 14789
rect 10910 14786 10916 14788
rect 10777 14784 10916 14786
rect 10777 14728 10782 14784
rect 10838 14728 10916 14784
rect 10777 14726 10916 14728
rect 10777 14723 10843 14726
rect 10910 14724 10916 14726
rect 10980 14786 10986 14788
rect 13494 14786 13554 14862
rect 18689 14859 18755 14862
rect 10980 14726 13554 14786
rect 10980 14724 10986 14726
rect 13939 14720 14259 14721
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 14655 14259 14656
rect 19137 14720 19457 14721
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 14655 19457 14656
rect 13721 14650 13787 14653
rect 6453 14648 6562 14650
rect 6453 14592 6458 14648
rect 6514 14592 6562 14648
rect 6453 14587 6562 14592
rect 9262 14648 13787 14650
rect 9262 14592 13726 14648
rect 13782 14592 13787 14648
rect 9262 14590 13787 14592
rect 13721 14587 13787 14590
rect 19609 14650 19675 14653
rect 22200 14650 23000 14680
rect 19609 14648 23000 14650
rect 19609 14592 19614 14648
rect 19670 14592 23000 14648
rect 19609 14590 23000 14592
rect 19609 14587 19675 14590
rect 4153 14378 4219 14381
rect 6502 14378 6562 14587
rect 22200 14560 23000 14590
rect 6637 14514 6703 14517
rect 19425 14514 19491 14517
rect 6637 14512 19491 14514
rect 6637 14456 6642 14512
rect 6698 14456 19430 14512
rect 19486 14456 19491 14512
rect 6637 14454 19491 14456
rect 6637 14451 6703 14454
rect 19425 14451 19491 14454
rect 10777 14378 10843 14381
rect 4153 14376 10843 14378
rect 4153 14320 4158 14376
rect 4214 14320 10782 14376
rect 10838 14320 10843 14376
rect 4153 14318 10843 14320
rect 4153 14315 4219 14318
rect 10777 14315 10843 14318
rect 10961 14378 11027 14381
rect 17125 14378 17191 14381
rect 10961 14376 17191 14378
rect 10961 14320 10966 14376
rect 11022 14320 17130 14376
rect 17186 14320 17191 14376
rect 10961 14318 17191 14320
rect 10961 14315 11027 14318
rect 17125 14315 17191 14318
rect 5942 14180 5948 14244
rect 6012 14180 6018 14244
rect 14273 14242 14339 14245
rect 14733 14244 14799 14245
rect 14733 14242 14780 14244
rect 14273 14240 14780 14242
rect 14844 14242 14850 14244
rect 21357 14242 21423 14245
rect 22200 14242 23000 14272
rect 14273 14184 14278 14240
rect 14334 14184 14738 14240
rect 14273 14182 14780 14184
rect 5950 13970 6010 14180
rect 14273 14179 14339 14182
rect 14733 14180 14780 14182
rect 14844 14182 14926 14242
rect 21357 14240 23000 14242
rect 21357 14184 21362 14240
rect 21418 14184 23000 14240
rect 21357 14182 23000 14184
rect 14844 14180 14850 14182
rect 14733 14179 14799 14180
rect 21357 14179 21423 14182
rect 6142 14176 6462 14177
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 14111 6462 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 16538 14176 16858 14177
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 22200 14152 23000 14182
rect 16538 14111 16858 14112
rect 15694 14106 15700 14108
rect 11838 14046 15700 14106
rect 11838 13970 11898 14046
rect 15694 14044 15700 14046
rect 15764 14044 15770 14108
rect 22001 13970 22067 13973
rect 5950 13910 11898 13970
rect 13126 13968 22067 13970
rect 13126 13912 22006 13968
rect 22062 13912 22067 13968
rect 13126 13910 22067 13912
rect 3233 13834 3299 13837
rect 10409 13834 10475 13837
rect 13126 13834 13186 13910
rect 22001 13907 22067 13910
rect 21265 13834 21331 13837
rect 22200 13834 23000 13864
rect 3233 13832 13186 13834
rect 3233 13776 3238 13832
rect 3294 13776 10414 13832
rect 10470 13776 13186 13832
rect 3233 13774 13186 13776
rect 13678 13774 14474 13834
rect 3233 13771 3299 13774
rect 10409 13771 10475 13774
rect 13678 13698 13738 13774
rect 13494 13638 13738 13698
rect 14414 13698 14474 13774
rect 21265 13832 23000 13834
rect 21265 13776 21270 13832
rect 21326 13776 23000 13832
rect 21265 13774 23000 13776
rect 21265 13771 21331 13774
rect 22200 13744 23000 13774
rect 18965 13698 19031 13701
rect 14414 13696 19031 13698
rect 14414 13640 18970 13696
rect 19026 13640 19031 13696
rect 14414 13638 19031 13640
rect 3543 13632 3863 13633
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 13567 3863 13568
rect 8741 13632 9061 13633
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 13567 9061 13568
rect 12198 13562 12204 13564
rect 9124 13502 12204 13562
rect 7189 13426 7255 13429
rect 9124 13426 9184 13502
rect 12198 13500 12204 13502
rect 12268 13562 12274 13564
rect 13353 13562 13419 13565
rect 12268 13560 13419 13562
rect 12268 13504 13358 13560
rect 13414 13504 13419 13560
rect 12268 13502 13419 13504
rect 12268 13500 12274 13502
rect 13353 13499 13419 13502
rect 7189 13424 9184 13426
rect 7189 13368 7194 13424
rect 7250 13368 9184 13424
rect 7189 13366 9184 13368
rect 9673 13426 9739 13429
rect 13494 13426 13554 13638
rect 18965 13635 19031 13638
rect 13939 13632 14259 13633
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 13567 14259 13568
rect 19137 13632 19457 13633
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 13567 19457 13568
rect 16021 13562 16087 13565
rect 16021 13560 19074 13562
rect 16021 13504 16026 13560
rect 16082 13504 19074 13560
rect 16021 13502 19074 13504
rect 16021 13499 16087 13502
rect 9673 13424 13554 13426
rect 9673 13368 9678 13424
rect 9734 13368 13554 13424
rect 9673 13366 13554 13368
rect 13629 13426 13695 13429
rect 17861 13426 17927 13429
rect 13629 13424 17927 13426
rect 13629 13368 13634 13424
rect 13690 13368 17866 13424
rect 17922 13368 17927 13424
rect 13629 13366 17927 13368
rect 19014 13426 19074 13502
rect 20529 13426 20595 13429
rect 19014 13424 20595 13426
rect 19014 13368 20534 13424
rect 20590 13368 20595 13424
rect 19014 13366 20595 13368
rect 7189 13363 7255 13366
rect 9673 13363 9739 13366
rect 13629 13363 13695 13366
rect 17861 13363 17927 13366
rect 20529 13363 20595 13366
rect 8569 13290 8635 13293
rect 15561 13290 15627 13293
rect 18229 13290 18295 13293
rect 8569 13288 15627 13290
rect 8569 13232 8574 13288
rect 8630 13232 15566 13288
rect 15622 13232 15627 13288
rect 8569 13230 15627 13232
rect 8569 13227 8635 13230
rect 15561 13227 15627 13230
rect 15702 13288 18295 13290
rect 15702 13232 18234 13288
rect 18290 13232 18295 13288
rect 15702 13230 18295 13232
rect 6862 13092 6868 13156
rect 6932 13154 6938 13156
rect 7189 13154 7255 13157
rect 6932 13152 7255 13154
rect 6932 13096 7194 13152
rect 7250 13096 7255 13152
rect 6932 13094 7255 13096
rect 6932 13092 6938 13094
rect 7189 13091 7255 13094
rect 11789 13154 11855 13157
rect 15702 13154 15762 13230
rect 18229 13227 18295 13230
rect 21173 13290 21239 13293
rect 22200 13290 23000 13320
rect 21173 13288 23000 13290
rect 21173 13232 21178 13288
rect 21234 13232 23000 13288
rect 21173 13230 23000 13232
rect 21173 13227 21239 13230
rect 22200 13200 23000 13230
rect 11789 13152 15762 13154
rect 11789 13096 11794 13152
rect 11850 13096 15762 13152
rect 11789 13094 15762 13096
rect 11789 13091 11855 13094
rect 6142 13088 6462 13089
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 13023 6462 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 16538 13088 16858 13089
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 13023 16858 13024
rect 8109 13018 8175 13021
rect 9581 13018 9647 13021
rect 8109 13016 9647 13018
rect 8109 12960 8114 13016
rect 8170 12960 9586 13016
rect 9642 12960 9647 13016
rect 8109 12958 9647 12960
rect 8109 12955 8175 12958
rect 9581 12955 9647 12958
rect 13353 13018 13419 13021
rect 16021 13018 16087 13021
rect 13353 13016 16087 13018
rect 13353 12960 13358 13016
rect 13414 12960 16026 13016
rect 16082 12960 16087 13016
rect 13353 12958 16087 12960
rect 13353 12955 13419 12958
rect 16021 12955 16087 12958
rect 17953 13018 18019 13021
rect 17953 13016 20546 13018
rect 17953 12960 17958 13016
rect 18014 12960 20546 13016
rect 17953 12958 20546 12960
rect 17953 12955 18019 12958
rect 7281 12882 7347 12885
rect 8518 12882 8524 12884
rect 7281 12880 8524 12882
rect 7281 12824 7286 12880
rect 7342 12824 8524 12880
rect 7281 12822 8524 12824
rect 7281 12819 7347 12822
rect 8518 12820 8524 12822
rect 8588 12820 8594 12884
rect 10041 12882 10107 12885
rect 20253 12882 20319 12885
rect 10041 12880 20319 12882
rect 10041 12824 10046 12880
rect 10102 12824 20258 12880
rect 20314 12824 20319 12880
rect 10041 12822 20319 12824
rect 20486 12882 20546 12958
rect 22200 12882 23000 12912
rect 20486 12822 23000 12882
rect 10041 12819 10107 12822
rect 20253 12819 20319 12822
rect 22200 12792 23000 12822
rect 7741 12746 7807 12749
rect 13537 12746 13603 12749
rect 7741 12744 13603 12746
rect 7741 12688 7746 12744
rect 7802 12688 13542 12744
rect 13598 12688 13603 12744
rect 7741 12686 13603 12688
rect 7741 12683 7807 12686
rect 13537 12683 13603 12686
rect 14549 12746 14615 12749
rect 18965 12746 19031 12749
rect 14549 12744 19031 12746
rect 14549 12688 14554 12744
rect 14610 12688 18970 12744
rect 19026 12688 19031 12744
rect 14549 12686 19031 12688
rect 14549 12683 14615 12686
rect 18965 12683 19031 12686
rect 9397 12610 9463 12613
rect 9581 12610 9647 12613
rect 11789 12610 11855 12613
rect 9397 12608 11855 12610
rect 9397 12552 9402 12608
rect 9458 12552 9586 12608
rect 9642 12552 11794 12608
rect 11850 12552 11855 12608
rect 9397 12550 11855 12552
rect 9397 12547 9463 12550
rect 9581 12547 9647 12550
rect 11789 12547 11855 12550
rect 3543 12544 3863 12545
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 12479 3863 12480
rect 8741 12544 9061 12545
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 12479 9061 12480
rect 13939 12544 14259 12545
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 12479 14259 12480
rect 19137 12544 19457 12545
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 12479 19457 12480
rect 7649 12338 7715 12341
rect 8334 12338 8340 12340
rect 7649 12336 8340 12338
rect 7649 12280 7654 12336
rect 7710 12280 8340 12336
rect 7649 12278 8340 12280
rect 7649 12275 7715 12278
rect 8334 12276 8340 12278
rect 8404 12276 8410 12340
rect 8569 12338 8635 12341
rect 20253 12338 20319 12341
rect 22200 12338 23000 12368
rect 8569 12336 20319 12338
rect 8569 12280 8574 12336
rect 8630 12280 20258 12336
rect 20314 12280 20319 12336
rect 8569 12278 20319 12280
rect 8569 12275 8635 12278
rect 20253 12275 20319 12278
rect 20486 12278 23000 12338
rect 7649 12202 7715 12205
rect 18045 12202 18111 12205
rect 19517 12202 19583 12205
rect 20486 12202 20546 12278
rect 22200 12248 23000 12278
rect 7649 12200 17970 12202
rect 7649 12144 7654 12200
rect 7710 12144 17970 12200
rect 7649 12142 17970 12144
rect 7649 12139 7715 12142
rect 14641 12066 14707 12069
rect 14774 12066 14780 12068
rect 14641 12064 14780 12066
rect 14641 12008 14646 12064
rect 14702 12008 14780 12064
rect 14641 12006 14780 12008
rect 14641 12003 14707 12006
rect 14774 12004 14780 12006
rect 14844 12004 14850 12068
rect 17910 12066 17970 12142
rect 18045 12200 20546 12202
rect 18045 12144 18050 12200
rect 18106 12144 19522 12200
rect 19578 12144 20546 12200
rect 18045 12142 20546 12144
rect 18045 12139 18111 12142
rect 19517 12139 19583 12142
rect 20989 12066 21055 12069
rect 17910 12064 21055 12066
rect 17910 12008 20994 12064
rect 21050 12008 21055 12064
rect 17910 12006 21055 12008
rect 20989 12003 21055 12006
rect 6142 12000 6462 12001
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 11935 6462 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 16538 12000 16858 12001
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 11935 16858 11936
rect 9121 11930 9187 11933
rect 7974 11928 9187 11930
rect 7974 11872 9126 11928
rect 9182 11872 9187 11928
rect 7974 11870 9187 11872
rect 3969 11794 4035 11797
rect 7974 11794 8034 11870
rect 9121 11867 9187 11870
rect 13537 11930 13603 11933
rect 16389 11930 16455 11933
rect 22200 11930 23000 11960
rect 13537 11928 16455 11930
rect 13537 11872 13542 11928
rect 13598 11872 16394 11928
rect 16450 11872 16455 11928
rect 13537 11870 16455 11872
rect 13537 11867 13603 11870
rect 16389 11867 16455 11870
rect 16990 11870 23000 11930
rect 3969 11792 8034 11794
rect 3969 11736 3974 11792
rect 4030 11736 8034 11792
rect 3969 11734 8034 11736
rect 8109 11794 8175 11797
rect 16990 11794 17050 11870
rect 22200 11840 23000 11870
rect 8109 11792 17050 11794
rect 8109 11736 8114 11792
rect 8170 11736 17050 11792
rect 8109 11734 17050 11736
rect 3969 11731 4035 11734
rect 8109 11731 8175 11734
rect 6821 11658 6887 11661
rect 13537 11658 13603 11661
rect 14365 11658 14431 11661
rect 6821 11656 13603 11658
rect 6821 11600 6826 11656
rect 6882 11600 13542 11656
rect 13598 11600 13603 11656
rect 6821 11598 13603 11600
rect 6821 11595 6887 11598
rect 13537 11595 13603 11598
rect 13816 11656 14431 11658
rect 13816 11600 14370 11656
rect 14426 11600 14431 11656
rect 13816 11598 14431 11600
rect 9121 11522 9187 11525
rect 13816 11522 13876 11598
rect 14365 11595 14431 11598
rect 16389 11658 16455 11661
rect 21633 11658 21699 11661
rect 16389 11656 21699 11658
rect 16389 11600 16394 11656
rect 16450 11600 21638 11656
rect 21694 11600 21699 11656
rect 16389 11598 21699 11600
rect 16389 11595 16455 11598
rect 21633 11595 21699 11598
rect 9121 11520 13876 11522
rect 9121 11464 9126 11520
rect 9182 11464 13876 11520
rect 9121 11462 13876 11464
rect 9121 11459 9187 11462
rect 3543 11456 3863 11457
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 11391 3863 11392
rect 8741 11456 9061 11457
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 11391 9061 11392
rect 13939 11456 14259 11457
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 11391 14259 11392
rect 19137 11456 19457 11457
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 11391 19457 11392
rect 22200 11386 23000 11416
rect 19566 11326 23000 11386
rect 8109 11250 8175 11253
rect 16849 11250 16915 11253
rect 19566 11250 19626 11326
rect 22200 11296 23000 11326
rect 8109 11248 16682 11250
rect 8109 11192 8114 11248
rect 8170 11192 16682 11248
rect 8109 11190 16682 11192
rect 8109 11187 8175 11190
rect 8569 11114 8635 11117
rect 16113 11114 16179 11117
rect 8569 11112 16179 11114
rect 8569 11056 8574 11112
rect 8630 11056 16118 11112
rect 16174 11056 16179 11112
rect 8569 11054 16179 11056
rect 16622 11114 16682 11190
rect 16849 11248 19626 11250
rect 16849 11192 16854 11248
rect 16910 11192 19626 11248
rect 16849 11190 19626 11192
rect 16849 11187 16915 11190
rect 20713 11114 20779 11117
rect 16622 11112 20779 11114
rect 16622 11056 20718 11112
rect 20774 11056 20779 11112
rect 16622 11054 20779 11056
rect 8569 11051 8635 11054
rect 16113 11051 16179 11054
rect 20713 11051 20779 11054
rect 16021 10978 16087 10981
rect 22200 10978 23000 11008
rect 12390 10976 16087 10978
rect 12390 10920 16026 10976
rect 16082 10920 16087 10976
rect 12390 10918 16087 10920
rect 6142 10912 6462 10913
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 10847 6462 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 7649 10842 7715 10845
rect 11145 10842 11211 10845
rect 12390 10842 12450 10918
rect 16021 10915 16087 10918
rect 16990 10918 23000 10978
rect 16538 10912 16858 10913
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 10847 16858 10848
rect 7649 10840 11211 10842
rect 7649 10784 7654 10840
rect 7710 10784 11150 10840
rect 11206 10784 11211 10840
rect 7649 10782 11211 10784
rect 7649 10779 7715 10782
rect 11145 10779 11211 10782
rect 11792 10782 12450 10842
rect 8293 10706 8359 10709
rect 11792 10706 11852 10782
rect 8293 10704 11852 10706
rect 8293 10648 8298 10704
rect 8354 10648 11852 10704
rect 8293 10646 11852 10648
rect 8293 10643 8359 10646
rect 12014 10644 12020 10708
rect 12084 10706 12090 10708
rect 16990 10706 17050 10918
rect 22200 10888 23000 10918
rect 20713 10842 20779 10845
rect 12084 10646 17050 10706
rect 17542 10840 20779 10842
rect 17542 10784 20718 10840
rect 20774 10784 20779 10840
rect 17542 10782 20779 10784
rect 12084 10644 12090 10646
rect 7741 10570 7807 10573
rect 14733 10570 14799 10573
rect 17542 10570 17602 10782
rect 20713 10779 20779 10782
rect 17953 10706 18019 10709
rect 17953 10704 19626 10706
rect 17953 10648 17958 10704
rect 18014 10648 19626 10704
rect 17953 10646 19626 10648
rect 17953 10643 18019 10646
rect 7741 10568 14658 10570
rect 7741 10512 7746 10568
rect 7802 10512 14658 10568
rect 7741 10510 14658 10512
rect 7741 10507 7807 10510
rect 9121 10434 9187 10437
rect 12801 10434 12867 10437
rect 9121 10432 12867 10434
rect 9121 10376 9126 10432
rect 9182 10376 12806 10432
rect 12862 10376 12867 10432
rect 9121 10374 12867 10376
rect 14598 10434 14658 10510
rect 14733 10568 17602 10570
rect 14733 10512 14738 10568
rect 14794 10512 17602 10568
rect 14733 10510 17602 10512
rect 14733 10507 14799 10510
rect 17902 10508 17908 10572
rect 17972 10570 17978 10572
rect 18597 10570 18663 10573
rect 17972 10568 18663 10570
rect 17972 10512 18602 10568
rect 18658 10512 18663 10568
rect 17972 10510 18663 10512
rect 17972 10508 17978 10510
rect 18597 10507 18663 10510
rect 18321 10434 18387 10437
rect 14598 10432 18387 10434
rect 14598 10376 18326 10432
rect 18382 10376 18387 10432
rect 14598 10374 18387 10376
rect 19566 10434 19626 10646
rect 22200 10434 23000 10464
rect 19566 10374 23000 10434
rect 9121 10371 9187 10374
rect 12801 10371 12867 10374
rect 18321 10371 18387 10374
rect 3543 10368 3863 10369
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 10303 3863 10304
rect 8741 10368 9061 10369
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 10303 9061 10304
rect 13939 10368 14259 10369
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 10303 14259 10304
rect 19137 10368 19457 10369
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 22200 10344 23000 10374
rect 19137 10303 19457 10304
rect 9121 10298 9187 10301
rect 12341 10298 12407 10301
rect 14549 10298 14615 10301
rect 18413 10298 18479 10301
rect 9121 10296 12266 10298
rect 9121 10240 9126 10296
rect 9182 10240 12266 10296
rect 9121 10238 12266 10240
rect 9121 10235 9187 10238
rect 8109 10162 8175 10165
rect 9622 10162 9628 10164
rect 8109 10160 9628 10162
rect 8109 10104 8114 10160
rect 8170 10104 9628 10160
rect 8109 10102 9628 10104
rect 8109 10099 8175 10102
rect 9622 10100 9628 10102
rect 9692 10100 9698 10164
rect 9806 10100 9812 10164
rect 9876 10162 9882 10164
rect 12014 10162 12020 10164
rect 9876 10102 12020 10162
rect 9876 10100 9882 10102
rect 12014 10100 12020 10102
rect 12084 10100 12090 10164
rect 12206 10162 12266 10238
rect 12341 10296 13876 10298
rect 12341 10240 12346 10296
rect 12402 10240 13876 10296
rect 12341 10238 13876 10240
rect 12341 10235 12407 10238
rect 13537 10162 13603 10165
rect 12206 10160 13603 10162
rect 12206 10104 13542 10160
rect 13598 10104 13603 10160
rect 12206 10102 13603 10104
rect 13816 10162 13876 10238
rect 14549 10296 18479 10298
rect 14549 10240 14554 10296
rect 14610 10240 18418 10296
rect 18474 10240 18479 10296
rect 14549 10238 18479 10240
rect 14549 10235 14615 10238
rect 18413 10235 18479 10238
rect 14457 10162 14523 10165
rect 13816 10160 14523 10162
rect 13816 10104 14462 10160
rect 14518 10104 14523 10160
rect 13816 10102 14523 10104
rect 13537 10099 13603 10102
rect 14457 10099 14523 10102
rect 16021 10162 16087 10165
rect 19333 10162 19399 10165
rect 16021 10160 19399 10162
rect 16021 10104 16026 10160
rect 16082 10104 19338 10160
rect 19394 10104 19399 10160
rect 16021 10102 19399 10104
rect 16021 10099 16087 10102
rect 19333 10099 19399 10102
rect 7925 10026 7991 10029
rect 9622 10026 9628 10028
rect 7925 10024 9628 10026
rect 7925 9968 7930 10024
rect 7986 9968 9628 10024
rect 7925 9966 9628 9968
rect 7925 9963 7991 9966
rect 9622 9964 9628 9966
rect 9692 9964 9698 10028
rect 17953 10026 18019 10029
rect 9768 10024 18019 10026
rect 9768 9968 17958 10024
rect 18014 9968 18019 10024
rect 9768 9966 18019 9968
rect 4102 9828 4108 9892
rect 4172 9890 4178 9892
rect 5901 9890 5967 9893
rect 4172 9888 5967 9890
rect 4172 9832 5906 9888
rect 5962 9832 5967 9888
rect 4172 9830 5967 9832
rect 4172 9828 4178 9830
rect 5901 9827 5967 9830
rect 6729 9890 6795 9893
rect 9121 9890 9187 9893
rect 6729 9888 9187 9890
rect 6729 9832 6734 9888
rect 6790 9832 9126 9888
rect 9182 9832 9187 9888
rect 6729 9830 9187 9832
rect 6729 9827 6795 9830
rect 9121 9827 9187 9830
rect 9622 9828 9628 9892
rect 9692 9890 9698 9892
rect 9768 9890 9828 9966
rect 17953 9963 18019 9966
rect 18689 10026 18755 10029
rect 22200 10026 23000 10056
rect 18689 10024 23000 10026
rect 18689 9968 18694 10024
rect 18750 9968 23000 10024
rect 18689 9966 23000 9968
rect 18689 9963 18755 9966
rect 22200 9936 23000 9966
rect 9692 9830 9828 9890
rect 13721 9890 13787 9893
rect 15193 9890 15259 9893
rect 13721 9888 15259 9890
rect 13721 9832 13726 9888
rect 13782 9832 15198 9888
rect 15254 9832 15259 9888
rect 13721 9830 15259 9832
rect 9692 9828 9698 9830
rect 13721 9827 13787 9830
rect 15193 9827 15259 9830
rect 6142 9824 6462 9825
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 9759 6462 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 16538 9824 16858 9825
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 9759 16858 9760
rect 8661 9754 8727 9757
rect 10317 9754 10383 9757
rect 8661 9752 10383 9754
rect 8661 9696 8666 9752
rect 8722 9696 10322 9752
rect 10378 9696 10383 9752
rect 8661 9694 10383 9696
rect 8661 9691 8727 9694
rect 10317 9691 10383 9694
rect 5206 9556 5212 9620
rect 5276 9618 5282 9620
rect 7097 9618 7163 9621
rect 7230 9618 7236 9620
rect 5276 9616 7236 9618
rect 5276 9560 7102 9616
rect 7158 9560 7236 9616
rect 5276 9558 7236 9560
rect 5276 9556 5282 9558
rect 7097 9555 7163 9558
rect 7230 9556 7236 9558
rect 7300 9556 7306 9620
rect 8385 9618 8451 9621
rect 19517 9618 19583 9621
rect 8385 9616 19583 9618
rect 8385 9560 8390 9616
rect 8446 9560 19522 9616
rect 19578 9560 19583 9616
rect 8385 9558 19583 9560
rect 8385 9555 8451 9558
rect 19517 9555 19583 9558
rect 6821 9482 6887 9485
rect 20161 9482 20227 9485
rect 6821 9480 20227 9482
rect 6821 9424 6826 9480
rect 6882 9424 20166 9480
rect 20222 9424 20227 9480
rect 6821 9422 20227 9424
rect 6821 9419 6887 9422
rect 20161 9419 20227 9422
rect 20713 9482 20779 9485
rect 22200 9482 23000 9512
rect 20713 9480 23000 9482
rect 20713 9424 20718 9480
rect 20774 9424 23000 9480
rect 20713 9422 23000 9424
rect 20713 9419 20779 9422
rect 22200 9392 23000 9422
rect 10777 9346 10843 9349
rect 13721 9346 13787 9349
rect 10777 9344 13787 9346
rect 10777 9288 10782 9344
rect 10838 9288 13726 9344
rect 13782 9288 13787 9344
rect 10777 9286 13787 9288
rect 10777 9283 10843 9286
rect 13721 9283 13787 9286
rect 14590 9284 14596 9348
rect 14660 9346 14666 9348
rect 18965 9346 19031 9349
rect 14660 9344 19031 9346
rect 14660 9288 18970 9344
rect 19026 9288 19031 9344
rect 14660 9286 19031 9288
rect 14660 9284 14666 9286
rect 18965 9283 19031 9286
rect 3543 9280 3863 9281
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 9215 3863 9216
rect 8741 9280 9061 9281
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 9215 9061 9216
rect 13939 9280 14259 9281
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 9215 14259 9216
rect 19137 9280 19457 9281
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 9215 19457 9216
rect 7281 9210 7347 9213
rect 8150 9210 8156 9212
rect 7281 9208 8156 9210
rect 7281 9152 7286 9208
rect 7342 9152 8156 9208
rect 7281 9150 8156 9152
rect 7281 9147 7347 9150
rect 8150 9148 8156 9150
rect 8220 9148 8226 9212
rect 13721 9210 13787 9213
rect 9630 9208 13787 9210
rect 9630 9152 13726 9208
rect 13782 9152 13787 9208
rect 9630 9150 13787 9152
rect 8661 9074 8727 9077
rect 9630 9074 9690 9150
rect 13721 9147 13787 9150
rect 14457 9210 14523 9213
rect 14457 9208 17096 9210
rect 14457 9152 14462 9208
rect 14518 9152 17096 9208
rect 14457 9150 17096 9152
rect 14457 9147 14523 9150
rect 8661 9072 9690 9074
rect 8661 9016 8666 9072
rect 8722 9016 9690 9072
rect 8661 9014 9690 9016
rect 17036 9074 17096 9150
rect 17166 9148 17172 9212
rect 17236 9210 17242 9212
rect 17309 9210 17375 9213
rect 17953 9210 18019 9213
rect 17236 9208 17375 9210
rect 17236 9152 17314 9208
rect 17370 9152 17375 9208
rect 17236 9150 17375 9152
rect 17236 9148 17242 9150
rect 17309 9147 17375 9150
rect 17772 9208 18019 9210
rect 17772 9152 17958 9208
rect 18014 9152 18019 9208
rect 17772 9150 18019 9152
rect 17772 9074 17832 9150
rect 17953 9147 18019 9150
rect 17036 9014 17832 9074
rect 17953 9074 18019 9077
rect 22200 9074 23000 9104
rect 17953 9072 23000 9074
rect 17953 9016 17958 9072
rect 18014 9016 23000 9072
rect 17953 9014 23000 9016
rect 8661 9011 8727 9014
rect 17953 9011 18019 9014
rect 22200 8984 23000 9014
rect 5574 8876 5580 8940
rect 5644 8938 5650 8940
rect 6545 8938 6611 8941
rect 21081 8938 21147 8941
rect 5644 8936 21147 8938
rect 5644 8880 6550 8936
rect 6606 8880 21086 8936
rect 21142 8880 21147 8936
rect 5644 8878 21147 8880
rect 5644 8876 5650 8878
rect 6545 8875 6611 8878
rect 21081 8875 21147 8878
rect 7230 8740 7236 8804
rect 7300 8802 7306 8804
rect 7557 8802 7623 8805
rect 7300 8800 7623 8802
rect 7300 8744 7562 8800
rect 7618 8744 7623 8800
rect 7300 8742 7623 8744
rect 7300 8740 7306 8742
rect 7557 8739 7623 8742
rect 13077 8802 13143 8805
rect 14365 8802 14431 8805
rect 16389 8802 16455 8805
rect 13077 8800 16455 8802
rect 13077 8744 13082 8800
rect 13138 8744 14370 8800
rect 14426 8744 16394 8800
rect 16450 8744 16455 8800
rect 13077 8742 16455 8744
rect 13077 8739 13143 8742
rect 14365 8739 14431 8742
rect 16389 8739 16455 8742
rect 18229 8802 18295 8805
rect 20713 8802 20779 8805
rect 18229 8800 20779 8802
rect 18229 8744 18234 8800
rect 18290 8744 20718 8800
rect 20774 8744 20779 8800
rect 18229 8742 20779 8744
rect 18229 8739 18295 8742
rect 20713 8739 20779 8742
rect 6142 8736 6462 8737
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 8671 6462 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 16538 8736 16858 8737
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 8671 16858 8672
rect 12801 8666 12867 8669
rect 13997 8666 14063 8669
rect 12801 8664 14063 8666
rect 12801 8608 12806 8664
rect 12862 8608 14002 8664
rect 14058 8608 14063 8664
rect 12801 8606 14063 8608
rect 12801 8603 12867 8606
rect 13997 8603 14063 8606
rect 14365 8666 14431 8669
rect 17953 8666 18019 8669
rect 22200 8666 23000 8696
rect 14365 8664 16130 8666
rect 14365 8608 14370 8664
rect 14426 8608 16130 8664
rect 14365 8606 16130 8608
rect 14365 8603 14431 8606
rect 7741 8532 7807 8533
rect 7741 8530 7788 8532
rect 7660 8528 7788 8530
rect 7852 8530 7858 8532
rect 10961 8530 11027 8533
rect 7852 8528 11027 8530
rect 7660 8472 7746 8528
rect 7852 8472 10966 8528
rect 11022 8472 11027 8528
rect 7660 8470 7788 8472
rect 7741 8468 7788 8470
rect 7852 8470 11027 8472
rect 7852 8468 7858 8470
rect 7741 8467 7807 8468
rect 10961 8467 11027 8470
rect 11237 8530 11303 8533
rect 14590 8530 14596 8532
rect 11237 8528 14596 8530
rect 11237 8472 11242 8528
rect 11298 8472 14596 8528
rect 11237 8470 14596 8472
rect 11237 8467 11303 8470
rect 14590 8468 14596 8470
rect 14660 8468 14666 8532
rect 16070 8530 16130 8606
rect 17953 8664 23000 8666
rect 17953 8608 17958 8664
rect 18014 8608 23000 8664
rect 17953 8606 23000 8608
rect 17953 8603 18019 8606
rect 22200 8576 23000 8606
rect 18045 8530 18111 8533
rect 16070 8528 18111 8530
rect 16070 8472 18050 8528
rect 18106 8472 18111 8528
rect 16070 8470 18111 8472
rect 18045 8467 18111 8470
rect 18822 8468 18828 8532
rect 18892 8530 18898 8532
rect 21081 8530 21147 8533
rect 18892 8528 21147 8530
rect 18892 8472 21086 8528
rect 21142 8472 21147 8528
rect 18892 8470 21147 8472
rect 18892 8468 18898 8470
rect 21081 8467 21147 8470
rect 7281 8394 7347 8397
rect 18965 8394 19031 8397
rect 7281 8392 19031 8394
rect 7281 8336 7286 8392
rect 7342 8336 18970 8392
rect 19026 8336 19031 8392
rect 7281 8334 19031 8336
rect 7281 8331 7347 8334
rect 18965 8331 19031 8334
rect 14365 8258 14431 8261
rect 17861 8258 17927 8261
rect 14365 8256 17927 8258
rect 14365 8200 14370 8256
rect 14426 8200 17866 8256
rect 17922 8200 17927 8256
rect 14365 8198 17927 8200
rect 14365 8195 14431 8198
rect 17861 8195 17927 8198
rect 3543 8192 3863 8193
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 8127 3863 8128
rect 8741 8192 9061 8193
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 8127 9061 8128
rect 13939 8192 14259 8193
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 8127 14259 8128
rect 19137 8192 19457 8193
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 8127 19457 8128
rect 18270 8060 18276 8124
rect 18340 8122 18346 8124
rect 18965 8122 19031 8125
rect 22200 8122 23000 8152
rect 18340 8120 19031 8122
rect 18340 8064 18970 8120
rect 19026 8064 19031 8120
rect 18340 8062 19031 8064
rect 18340 8060 18346 8062
rect 18965 8059 19031 8062
rect 19934 8062 23000 8122
rect 6913 7986 6979 7989
rect 19701 7986 19767 7989
rect 6913 7984 19767 7986
rect 6913 7928 6918 7984
rect 6974 7928 19706 7984
rect 19762 7928 19767 7984
rect 6913 7926 19767 7928
rect 6913 7923 6979 7926
rect 19701 7923 19767 7926
rect 6545 7850 6611 7853
rect 17861 7850 17927 7853
rect 6545 7848 17927 7850
rect 6545 7792 6550 7848
rect 6606 7792 17866 7848
rect 17922 7792 17927 7848
rect 6545 7790 17927 7792
rect 6545 7787 6611 7790
rect 17861 7787 17927 7790
rect 18045 7850 18111 7853
rect 19934 7850 19994 8062
rect 22200 8032 23000 8062
rect 18045 7848 19994 7850
rect 18045 7792 18050 7848
rect 18106 7792 19994 7848
rect 18045 7790 19994 7792
rect 18045 7787 18111 7790
rect 7598 7652 7604 7716
rect 7668 7714 7674 7716
rect 11053 7714 11119 7717
rect 7668 7712 11119 7714
rect 7668 7656 11058 7712
rect 11114 7656 11119 7712
rect 7668 7654 11119 7656
rect 7668 7652 7674 7654
rect 11053 7651 11119 7654
rect 13445 7714 13511 7717
rect 16297 7714 16363 7717
rect 22200 7714 23000 7744
rect 13445 7712 16363 7714
rect 13445 7656 13450 7712
rect 13506 7656 16302 7712
rect 16358 7656 16363 7712
rect 13445 7654 16363 7656
rect 13445 7651 13511 7654
rect 16297 7651 16363 7654
rect 16990 7654 23000 7714
rect 6142 7648 6462 7649
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 7583 6462 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 16538 7648 16858 7649
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 7583 16858 7584
rect 7373 7578 7439 7581
rect 9121 7578 9187 7581
rect 7373 7576 9187 7578
rect 7373 7520 7378 7576
rect 7434 7520 9126 7576
rect 9182 7520 9187 7576
rect 7373 7518 9187 7520
rect 7373 7515 7439 7518
rect 9121 7515 9187 7518
rect 11973 7578 12039 7581
rect 15101 7578 15167 7581
rect 11973 7576 15167 7578
rect 11973 7520 11978 7576
rect 12034 7520 15106 7576
rect 15162 7520 15167 7576
rect 11973 7518 15167 7520
rect 11973 7515 12039 7518
rect 15101 7515 15167 7518
rect 4470 7380 4476 7444
rect 4540 7442 4546 7444
rect 7097 7442 7163 7445
rect 7598 7442 7604 7444
rect 4540 7440 7604 7442
rect 4540 7384 7102 7440
rect 7158 7384 7604 7440
rect 4540 7382 7604 7384
rect 4540 7380 4546 7382
rect 7097 7379 7163 7382
rect 7598 7380 7604 7382
rect 7668 7380 7674 7444
rect 10593 7442 10659 7445
rect 13445 7442 13511 7445
rect 10593 7440 13511 7442
rect 10593 7384 10598 7440
rect 10654 7384 13450 7440
rect 13506 7384 13511 7440
rect 10593 7382 13511 7384
rect 10593 7379 10659 7382
rect 13445 7379 13511 7382
rect 13721 7442 13787 7445
rect 16990 7442 17050 7654
rect 22200 7624 23000 7654
rect 17861 7578 17927 7581
rect 20989 7578 21055 7581
rect 17861 7576 21055 7578
rect 17861 7520 17866 7576
rect 17922 7520 20994 7576
rect 21050 7520 21055 7576
rect 17861 7518 21055 7520
rect 17861 7515 17927 7518
rect 20989 7515 21055 7518
rect 13721 7440 17050 7442
rect 13721 7384 13726 7440
rect 13782 7384 17050 7440
rect 13721 7382 17050 7384
rect 17769 7442 17835 7445
rect 18597 7442 18663 7445
rect 17769 7440 18663 7442
rect 17769 7384 17774 7440
rect 17830 7384 18602 7440
rect 18658 7384 18663 7440
rect 17769 7382 18663 7384
rect 13721 7379 13787 7382
rect 17769 7379 17835 7382
rect 18597 7379 18663 7382
rect 7465 7306 7531 7309
rect 11973 7306 12039 7309
rect 7465 7304 12039 7306
rect 7465 7248 7470 7304
rect 7526 7248 11978 7304
rect 12034 7248 12039 7304
rect 7465 7246 12039 7248
rect 7465 7243 7531 7246
rect 11973 7243 12039 7246
rect 12341 7306 12407 7309
rect 19149 7306 19215 7309
rect 12341 7304 19215 7306
rect 12341 7248 12346 7304
rect 12402 7248 19154 7304
rect 19210 7248 19215 7304
rect 12341 7246 19215 7248
rect 12341 7243 12407 7246
rect 19149 7243 19215 7246
rect 9121 7170 9187 7173
rect 14365 7170 14431 7173
rect 15009 7170 15075 7173
rect 9121 7168 13876 7170
rect 9121 7112 9126 7168
rect 9182 7112 13876 7168
rect 9121 7110 13876 7112
rect 9121 7107 9187 7110
rect 3543 7104 3863 7105
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 7039 3863 7040
rect 8741 7104 9061 7105
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 7039 9061 7040
rect 5257 7034 5323 7037
rect 8150 7034 8156 7036
rect 5257 7032 8156 7034
rect 5257 6976 5262 7032
rect 5318 6976 8156 7032
rect 5257 6974 8156 6976
rect 5257 6971 5323 6974
rect 8150 6972 8156 6974
rect 8220 6972 8226 7036
rect 9857 7034 9923 7037
rect 12433 7034 12499 7037
rect 9857 7032 12499 7034
rect 9857 6976 9862 7032
rect 9918 6976 12438 7032
rect 12494 6976 12499 7032
rect 9857 6974 12499 6976
rect 9857 6971 9923 6974
rect 12433 6971 12499 6974
rect 4797 6900 4863 6901
rect 4797 6898 4844 6900
rect 4752 6896 4844 6898
rect 4752 6840 4802 6896
rect 4752 6838 4844 6840
rect 4797 6836 4844 6838
rect 4908 6836 4914 6900
rect 12341 6898 12407 6901
rect 13629 6898 13695 6901
rect 6870 6838 12082 6898
rect 4797 6835 4863 6836
rect 6729 6762 6795 6765
rect 6870 6762 6930 6838
rect 6729 6760 6930 6762
rect 6729 6704 6734 6760
rect 6790 6704 6930 6760
rect 6729 6702 6930 6704
rect 8385 6762 8451 6765
rect 12022 6762 12082 6838
rect 12341 6896 13695 6898
rect 12341 6840 12346 6896
rect 12402 6840 13634 6896
rect 13690 6840 13695 6896
rect 12341 6838 13695 6840
rect 13816 6898 13876 7110
rect 14365 7168 15075 7170
rect 14365 7112 14370 7168
rect 14426 7112 15014 7168
rect 15070 7112 15075 7168
rect 14365 7110 15075 7112
rect 14365 7107 14431 7110
rect 15009 7107 15075 7110
rect 16297 7170 16363 7173
rect 16941 7170 17007 7173
rect 18229 7170 18295 7173
rect 22200 7170 23000 7200
rect 16297 7168 18295 7170
rect 16297 7112 16302 7168
rect 16358 7112 16946 7168
rect 17002 7112 18234 7168
rect 18290 7112 18295 7168
rect 16297 7110 18295 7112
rect 16297 7107 16363 7110
rect 16941 7107 17007 7110
rect 18229 7107 18295 7110
rect 19566 7110 23000 7170
rect 13939 7104 14259 7105
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 7039 14259 7040
rect 19137 7104 19457 7105
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 7039 19457 7040
rect 17953 7034 18019 7037
rect 14414 7032 18019 7034
rect 14414 6976 17958 7032
rect 18014 6976 18019 7032
rect 14414 6974 18019 6976
rect 14414 6898 14474 6974
rect 17953 6971 18019 6974
rect 13816 6838 14474 6898
rect 14641 6898 14707 6901
rect 17585 6898 17651 6901
rect 14641 6896 17651 6898
rect 14641 6840 14646 6896
rect 14702 6840 17590 6896
rect 17646 6840 17651 6896
rect 14641 6838 17651 6840
rect 12341 6835 12407 6838
rect 13629 6835 13695 6838
rect 14641 6835 14707 6838
rect 17585 6835 17651 6838
rect 18229 6898 18295 6901
rect 19566 6898 19626 7110
rect 22200 7080 23000 7110
rect 18229 6896 19626 6898
rect 18229 6840 18234 6896
rect 18290 6840 19626 6896
rect 18229 6838 19626 6840
rect 18229 6835 18295 6838
rect 17677 6762 17743 6765
rect 8385 6760 11852 6762
rect 8385 6704 8390 6760
rect 8446 6704 11852 6760
rect 8385 6702 11852 6704
rect 12022 6760 17743 6762
rect 12022 6704 17682 6760
rect 17738 6704 17743 6760
rect 12022 6702 17743 6704
rect 6729 6699 6795 6702
rect 8385 6699 8451 6702
rect 6142 6560 6462 6561
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 6495 6462 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 6729 6490 6795 6493
rect 10593 6490 10659 6493
rect 6729 6488 10659 6490
rect 6729 6432 6734 6488
rect 6790 6432 10598 6488
rect 10654 6432 10659 6488
rect 6729 6430 10659 6432
rect 11792 6490 11852 6702
rect 17677 6699 17743 6702
rect 17953 6762 18019 6765
rect 22200 6762 23000 6792
rect 17953 6760 23000 6762
rect 17953 6704 17958 6760
rect 18014 6704 23000 6760
rect 17953 6702 23000 6704
rect 17953 6699 18019 6702
rect 22200 6672 23000 6702
rect 12249 6626 12315 6629
rect 13169 6626 13235 6629
rect 12249 6624 13235 6626
rect 12249 6568 12254 6624
rect 12310 6568 13174 6624
rect 13230 6568 13235 6624
rect 12249 6566 13235 6568
rect 12249 6563 12315 6566
rect 13169 6563 13235 6566
rect 13445 6626 13511 6629
rect 17585 6626 17651 6629
rect 18965 6626 19031 6629
rect 13445 6624 16452 6626
rect 13445 6568 13450 6624
rect 13506 6568 16452 6624
rect 13445 6566 16452 6568
rect 13445 6563 13511 6566
rect 15193 6490 15259 6493
rect 11792 6488 15259 6490
rect 11792 6432 15198 6488
rect 15254 6432 15259 6488
rect 11792 6430 15259 6432
rect 6729 6427 6795 6430
rect 10593 6427 10659 6430
rect 15193 6427 15259 6430
rect 7465 6354 7531 6357
rect 9305 6354 9371 6357
rect 9489 6354 9555 6357
rect 7465 6352 9555 6354
rect 7465 6296 7470 6352
rect 7526 6296 9310 6352
rect 9366 6296 9494 6352
rect 9550 6296 9555 6352
rect 7465 6294 9555 6296
rect 7465 6291 7531 6294
rect 9305 6291 9371 6294
rect 9489 6291 9555 6294
rect 11053 6354 11119 6357
rect 13445 6354 13511 6357
rect 11053 6352 13511 6354
rect 11053 6296 11058 6352
rect 11114 6296 13450 6352
rect 13506 6296 13511 6352
rect 11053 6294 13511 6296
rect 11053 6291 11119 6294
rect 13445 6291 13511 6294
rect 14549 6354 14615 6357
rect 14733 6354 14799 6357
rect 14549 6352 14799 6354
rect 14549 6296 14554 6352
rect 14610 6296 14738 6352
rect 14794 6296 14799 6352
rect 14549 6294 14799 6296
rect 16392 6354 16452 6566
rect 17585 6624 19031 6626
rect 17585 6568 17590 6624
rect 17646 6568 18970 6624
rect 19026 6568 19031 6624
rect 17585 6566 19031 6568
rect 17585 6563 17651 6566
rect 18965 6563 19031 6566
rect 16538 6560 16858 6561
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 6495 16858 6496
rect 17902 6428 17908 6492
rect 17972 6490 17978 6492
rect 18597 6490 18663 6493
rect 17972 6488 18663 6490
rect 17972 6432 18602 6488
rect 18658 6432 18663 6488
rect 17972 6430 18663 6432
rect 17972 6428 17978 6430
rect 18597 6427 18663 6430
rect 18965 6490 19031 6493
rect 20989 6490 21055 6493
rect 18965 6488 21055 6490
rect 18965 6432 18970 6488
rect 19026 6432 20994 6488
rect 21050 6432 21055 6488
rect 18965 6430 21055 6432
rect 18965 6427 19031 6430
rect 20989 6427 21055 6430
rect 20621 6354 20687 6357
rect 16392 6352 20687 6354
rect 16392 6296 20626 6352
rect 20682 6296 20687 6352
rect 16392 6294 20687 6296
rect 14549 6291 14615 6294
rect 14733 6291 14799 6294
rect 20621 6291 20687 6294
rect 6545 6218 6611 6221
rect 14549 6218 14615 6221
rect 6545 6216 14615 6218
rect 6545 6160 6550 6216
rect 6606 6160 14554 6216
rect 14610 6160 14615 6216
rect 6545 6158 14615 6160
rect 6545 6155 6611 6158
rect 14549 6155 14615 6158
rect 18781 6218 18847 6221
rect 22200 6218 23000 6248
rect 18781 6216 23000 6218
rect 18781 6160 18786 6216
rect 18842 6160 23000 6216
rect 18781 6158 23000 6160
rect 18781 6155 18847 6158
rect 22200 6128 23000 6158
rect 7189 6082 7255 6085
rect 9213 6084 9279 6085
rect 7966 6082 7972 6084
rect 7189 6080 7972 6082
rect 7189 6024 7194 6080
rect 7250 6024 7972 6080
rect 7189 6022 7972 6024
rect 7189 6019 7255 6022
rect 7966 6020 7972 6022
rect 8036 6020 8042 6084
rect 9213 6080 9260 6084
rect 9324 6082 9330 6084
rect 10409 6082 10475 6085
rect 13353 6082 13419 6085
rect 9213 6024 9218 6080
rect 9213 6020 9260 6024
rect 9324 6022 9370 6082
rect 10409 6080 13419 6082
rect 10409 6024 10414 6080
rect 10470 6024 13358 6080
rect 13414 6024 13419 6080
rect 10409 6022 13419 6024
rect 9324 6020 9330 6022
rect 9213 6019 9279 6020
rect 10409 6019 10475 6022
rect 13353 6019 13419 6022
rect 14365 6082 14431 6085
rect 18965 6082 19031 6085
rect 14365 6080 19031 6082
rect 14365 6024 14370 6080
rect 14426 6024 18970 6080
rect 19026 6024 19031 6080
rect 14365 6022 19031 6024
rect 14365 6019 14431 6022
rect 18965 6019 19031 6022
rect 3543 6016 3863 6017
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 5951 3863 5952
rect 8741 6016 9061 6017
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 5951 9061 5952
rect 13939 6016 14259 6017
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 5951 14259 5952
rect 19137 6016 19457 6017
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 5951 19457 5952
rect 5809 5946 5875 5949
rect 8569 5946 8635 5949
rect 5809 5944 8635 5946
rect 5809 5888 5814 5944
rect 5870 5888 8574 5944
rect 8630 5888 8635 5944
rect 5809 5886 8635 5888
rect 5809 5883 5875 5886
rect 8569 5883 8635 5886
rect 9213 5946 9279 5949
rect 13721 5946 13787 5949
rect 9213 5944 13787 5946
rect 9213 5888 9218 5944
rect 9274 5888 13726 5944
rect 13782 5888 13787 5944
rect 9213 5886 13787 5888
rect 9213 5883 9279 5886
rect 13721 5883 13787 5886
rect 0 5810 800 5840
rect 1393 5810 1459 5813
rect 0 5808 1459 5810
rect 0 5752 1398 5808
rect 1454 5752 1459 5808
rect 0 5750 1459 5752
rect 0 5720 800 5750
rect 1393 5747 1459 5750
rect 5993 5810 6059 5813
rect 7281 5810 7347 5813
rect 18229 5810 18295 5813
rect 5993 5808 7160 5810
rect 5993 5752 5998 5808
rect 6054 5752 7160 5808
rect 5993 5750 7160 5752
rect 5993 5747 6059 5750
rect 2037 5674 2103 5677
rect 3233 5674 3299 5677
rect 4429 5674 4495 5677
rect 6545 5674 6611 5677
rect 2037 5672 6611 5674
rect 2037 5616 2042 5672
rect 2098 5616 3238 5672
rect 3294 5616 4434 5672
rect 4490 5616 6550 5672
rect 6606 5616 6611 5672
rect 2037 5614 6611 5616
rect 7100 5674 7160 5750
rect 7281 5808 18295 5810
rect 7281 5752 7286 5808
rect 7342 5752 18234 5808
rect 18290 5752 18295 5808
rect 7281 5750 18295 5752
rect 7281 5747 7347 5750
rect 18229 5747 18295 5750
rect 18689 5810 18755 5813
rect 22200 5810 23000 5840
rect 18689 5808 23000 5810
rect 18689 5752 18694 5808
rect 18750 5752 23000 5808
rect 18689 5750 23000 5752
rect 18689 5747 18755 5750
rect 22200 5720 23000 5750
rect 8201 5674 8267 5677
rect 9121 5674 9187 5677
rect 7100 5672 9187 5674
rect 7100 5616 8206 5672
rect 8262 5616 9126 5672
rect 9182 5616 9187 5672
rect 7100 5614 9187 5616
rect 2037 5611 2103 5614
rect 3233 5611 3299 5614
rect 4429 5611 4495 5614
rect 6545 5611 6611 5614
rect 8201 5611 8267 5614
rect 9121 5611 9187 5614
rect 9305 5674 9371 5677
rect 19333 5674 19399 5677
rect 9305 5672 19399 5674
rect 9305 5616 9310 5672
rect 9366 5616 19338 5672
rect 19394 5616 19399 5672
rect 9305 5614 19399 5616
rect 9305 5611 9371 5614
rect 19333 5611 19399 5614
rect 5717 5538 5783 5541
rect 5942 5538 5948 5540
rect 5717 5536 5948 5538
rect 5717 5480 5722 5536
rect 5778 5480 5948 5536
rect 5717 5478 5948 5480
rect 5717 5475 5783 5478
rect 5942 5476 5948 5478
rect 6012 5476 6018 5540
rect 13353 5538 13419 5541
rect 16113 5538 16179 5541
rect 13353 5536 16179 5538
rect 13353 5480 13358 5536
rect 13414 5480 16118 5536
rect 16174 5480 16179 5536
rect 13353 5478 16179 5480
rect 13353 5475 13419 5478
rect 16113 5475 16179 5478
rect 6142 5472 6462 5473
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 5407 6462 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 16538 5472 16858 5473
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 5407 16858 5408
rect 5390 5340 5396 5404
rect 5460 5402 5466 5404
rect 5901 5402 5967 5405
rect 8017 5402 8083 5405
rect 5460 5400 5967 5402
rect 5460 5344 5906 5400
rect 5962 5344 5967 5400
rect 5460 5342 5967 5344
rect 5460 5340 5466 5342
rect 5901 5339 5967 5342
rect 7422 5400 8083 5402
rect 7422 5344 8022 5400
rect 8078 5344 8083 5400
rect 7422 5342 8083 5344
rect 5441 5266 5507 5269
rect 7422 5266 7482 5342
rect 8017 5339 8083 5342
rect 11789 5402 11855 5405
rect 11789 5400 15578 5402
rect 11789 5344 11794 5400
rect 11850 5344 15578 5400
rect 11789 5342 15578 5344
rect 11789 5339 11855 5342
rect 5441 5264 7482 5266
rect 5441 5208 5446 5264
rect 5502 5208 7482 5264
rect 5441 5206 7482 5208
rect 7649 5266 7715 5269
rect 15377 5266 15443 5269
rect 7649 5264 15443 5266
rect 7649 5208 7654 5264
rect 7710 5208 15382 5264
rect 15438 5208 15443 5264
rect 7649 5206 15443 5208
rect 15518 5266 15578 5342
rect 18597 5266 18663 5269
rect 15518 5264 18663 5266
rect 15518 5208 18602 5264
rect 18658 5208 18663 5264
rect 15518 5206 18663 5208
rect 5441 5203 5507 5206
rect 7649 5203 7715 5206
rect 15377 5203 15443 5206
rect 18597 5203 18663 5206
rect 19057 5266 19123 5269
rect 22200 5266 23000 5296
rect 19057 5264 23000 5266
rect 19057 5208 19062 5264
rect 19118 5208 23000 5264
rect 19057 5206 23000 5208
rect 19057 5203 19123 5206
rect 22200 5176 23000 5206
rect 8109 5130 8175 5133
rect 18505 5130 18571 5133
rect 19885 5130 19951 5133
rect 8109 5128 18571 5130
rect 8109 5072 8114 5128
rect 8170 5072 18510 5128
rect 18566 5072 18571 5128
rect 8109 5070 18571 5072
rect 8109 5067 8175 5070
rect 18505 5067 18571 5070
rect 19014 5128 19951 5130
rect 19014 5072 19890 5128
rect 19946 5072 19951 5128
rect 19014 5070 19951 5072
rect 5758 4932 5764 4996
rect 5828 4994 5834 4996
rect 6729 4994 6795 4997
rect 5828 4992 6795 4994
rect 5828 4936 6734 4992
rect 6790 4936 6795 4992
rect 5828 4934 6795 4936
rect 5828 4932 5834 4934
rect 6729 4931 6795 4934
rect 9121 4994 9187 4997
rect 11789 4994 11855 4997
rect 9121 4992 11855 4994
rect 9121 4936 9126 4992
rect 9182 4936 11794 4992
rect 11850 4936 11855 4992
rect 9121 4934 11855 4936
rect 9121 4931 9187 4934
rect 11789 4931 11855 4934
rect 15377 4994 15443 4997
rect 19014 4994 19074 5070
rect 19885 5067 19951 5070
rect 15377 4992 19074 4994
rect 15377 4936 15382 4992
rect 15438 4936 19074 4992
rect 15377 4934 19074 4936
rect 15377 4931 15443 4934
rect 3543 4928 3863 4929
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 4863 3863 4864
rect 8741 4928 9061 4929
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 4863 9061 4864
rect 13939 4928 14259 4929
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 4863 14259 4864
rect 19137 4928 19457 4929
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 4863 19457 4864
rect 5441 4858 5507 4861
rect 7782 4858 7788 4860
rect 5441 4856 7788 4858
rect 5441 4800 5446 4856
rect 5502 4800 7788 4856
rect 5441 4798 7788 4800
rect 5441 4795 5507 4798
rect 7782 4796 7788 4798
rect 7852 4796 7858 4860
rect 9305 4858 9371 4861
rect 9305 4856 12450 4858
rect 9305 4800 9310 4856
rect 9366 4800 12450 4856
rect 9305 4798 12450 4800
rect 9305 4795 9371 4798
rect 7649 4722 7715 4725
rect 12390 4722 12450 4798
rect 17534 4796 17540 4860
rect 17604 4858 17610 4860
rect 17861 4858 17927 4861
rect 22200 4858 23000 4888
rect 17604 4856 17927 4858
rect 17604 4800 17866 4856
rect 17922 4800 17927 4856
rect 17604 4798 17927 4800
rect 17604 4796 17610 4798
rect 17861 4795 17927 4798
rect 20486 4798 23000 4858
rect 19885 4722 19951 4725
rect 7649 4720 12082 4722
rect 7649 4664 7654 4720
rect 7710 4664 12082 4720
rect 7649 4662 12082 4664
rect 12390 4720 19951 4722
rect 12390 4664 19890 4720
rect 19946 4664 19951 4720
rect 12390 4662 19951 4664
rect 7649 4659 7715 4662
rect 6453 4586 6519 4589
rect 7414 4586 7420 4588
rect 6453 4584 7420 4586
rect 6453 4528 6458 4584
rect 6514 4528 7420 4584
rect 6453 4526 7420 4528
rect 6453 4523 6519 4526
rect 7414 4524 7420 4526
rect 7484 4524 7490 4588
rect 8477 4586 8543 4589
rect 8753 4586 8819 4589
rect 8477 4584 8819 4586
rect 8477 4528 8482 4584
rect 8538 4528 8758 4584
rect 8814 4528 8819 4584
rect 8477 4526 8819 4528
rect 8477 4523 8543 4526
rect 8753 4523 8819 4526
rect 9397 4586 9463 4589
rect 12022 4586 12082 4662
rect 19885 4659 19951 4662
rect 14181 4586 14247 4589
rect 16573 4586 16639 4589
rect 9397 4584 11852 4586
rect 9397 4528 9402 4584
rect 9458 4528 11852 4584
rect 9397 4526 11852 4528
rect 12022 4584 14247 4586
rect 12022 4528 14186 4584
rect 14242 4528 14247 4584
rect 12022 4526 14247 4528
rect 9397 4523 9463 4526
rect 6545 4450 6611 4453
rect 8518 4450 8524 4452
rect 6545 4448 8524 4450
rect 6545 4392 6550 4448
rect 6606 4392 8524 4448
rect 6545 4390 8524 4392
rect 6545 4387 6611 4390
rect 8518 4388 8524 4390
rect 8588 4388 8594 4452
rect 11792 4450 11852 4526
rect 14181 4523 14247 4526
rect 14782 4584 16639 4586
rect 14782 4528 16578 4584
rect 16634 4528 16639 4584
rect 14782 4526 16639 4528
rect 14782 4450 14842 4526
rect 16573 4523 16639 4526
rect 16849 4586 16915 4589
rect 17166 4586 17172 4588
rect 16849 4584 17172 4586
rect 16849 4528 16854 4584
rect 16910 4528 17172 4584
rect 16849 4526 17172 4528
rect 16849 4523 16915 4526
rect 17166 4524 17172 4526
rect 17236 4524 17242 4588
rect 19057 4586 19123 4589
rect 20486 4586 20546 4798
rect 22200 4768 23000 4798
rect 19057 4584 20546 4586
rect 19057 4528 19062 4584
rect 19118 4528 20546 4584
rect 19057 4526 20546 4528
rect 19057 4523 19123 4526
rect 11792 4390 14842 4450
rect 15142 4388 15148 4452
rect 15212 4450 15218 4452
rect 15285 4450 15351 4453
rect 15212 4448 15351 4450
rect 15212 4392 15290 4448
rect 15346 4392 15351 4448
rect 15212 4390 15351 4392
rect 15212 4388 15218 4390
rect 15285 4387 15351 4390
rect 18873 4450 18939 4453
rect 22200 4450 23000 4480
rect 18873 4448 23000 4450
rect 18873 4392 18878 4448
rect 18934 4392 23000 4448
rect 18873 4390 23000 4392
rect 18873 4387 18939 4390
rect 6142 4384 6462 4385
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 4319 6462 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 16538 4384 16858 4385
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 22200 4360 23000 4390
rect 16538 4319 16858 4320
rect 9305 4314 9371 4317
rect 6686 4312 9371 4314
rect 6686 4256 9310 4312
rect 9366 4256 9371 4312
rect 6686 4254 9371 4256
rect 2313 4178 2379 4181
rect 2589 4178 2655 4181
rect 4797 4178 4863 4181
rect 2313 4176 2514 4178
rect 2313 4120 2318 4176
rect 2374 4120 2514 4176
rect 2313 4118 2514 4120
rect 2313 4115 2379 4118
rect 2454 4042 2514 4118
rect 2589 4176 4863 4178
rect 2589 4120 2594 4176
rect 2650 4120 4802 4176
rect 4858 4120 4863 4176
rect 2589 4118 4863 4120
rect 2589 4115 2655 4118
rect 4797 4115 4863 4118
rect 5533 4178 5599 4181
rect 6686 4178 6746 4254
rect 9305 4251 9371 4254
rect 12157 4314 12223 4317
rect 14089 4314 14155 4317
rect 12157 4312 14155 4314
rect 12157 4256 12162 4312
rect 12218 4256 14094 4312
rect 14150 4256 14155 4312
rect 12157 4254 14155 4256
rect 12157 4251 12223 4254
rect 14089 4251 14155 4254
rect 5533 4176 6746 4178
rect 5533 4120 5538 4176
rect 5594 4120 6746 4176
rect 5533 4118 6746 4120
rect 6821 4178 6887 4181
rect 6821 4176 17418 4178
rect 6821 4120 6826 4176
rect 6882 4120 17418 4176
rect 6821 4118 17418 4120
rect 5533 4115 5599 4118
rect 6821 4115 6887 4118
rect 3049 4042 3115 4045
rect 5441 4042 5507 4045
rect 2454 3982 2790 4042
rect 2730 3498 2790 3982
rect 3049 4040 5507 4042
rect 3049 3984 3054 4040
rect 3110 3984 5446 4040
rect 5502 3984 5507 4040
rect 3049 3982 5507 3984
rect 3049 3979 3115 3982
rect 5441 3979 5507 3982
rect 5574 3980 5580 4044
rect 5644 4042 5650 4044
rect 5717 4042 5783 4045
rect 6821 4044 6887 4045
rect 6821 4042 6868 4044
rect 5644 4040 5783 4042
rect 5644 3984 5722 4040
rect 5778 3984 5783 4040
rect 5644 3982 5783 3984
rect 6776 4040 6868 4042
rect 6776 3984 6826 4040
rect 6776 3982 6868 3984
rect 5644 3980 5650 3982
rect 5717 3979 5783 3982
rect 6821 3980 6868 3982
rect 6932 3980 6938 4044
rect 8661 4042 8727 4045
rect 8526 4040 8727 4042
rect 8526 3984 8666 4040
rect 8722 3984 8727 4040
rect 8526 3982 8727 3984
rect 6821 3979 6887 3980
rect 4061 3906 4127 3909
rect 8526 3906 8586 3982
rect 8661 3979 8727 3982
rect 9949 4042 10015 4045
rect 12341 4042 12407 4045
rect 14457 4044 14523 4045
rect 9949 4040 12407 4042
rect 9949 3984 9954 4040
rect 10010 3984 12346 4040
rect 12402 3984 12407 4040
rect 9949 3982 12407 3984
rect 9949 3979 10015 3982
rect 12341 3979 12407 3982
rect 14406 3980 14412 4044
rect 14476 4042 14523 4044
rect 17358 4042 17418 4118
rect 17534 4116 17540 4180
rect 17604 4178 17610 4180
rect 18045 4178 18111 4181
rect 17604 4176 18111 4178
rect 17604 4120 18050 4176
rect 18106 4120 18111 4176
rect 17604 4118 18111 4120
rect 17604 4116 17610 4118
rect 18045 4115 18111 4118
rect 20662 4116 20668 4180
rect 20732 4178 20738 4180
rect 20897 4178 20963 4181
rect 20732 4176 20963 4178
rect 20732 4120 20902 4176
rect 20958 4120 20963 4176
rect 20732 4118 20963 4120
rect 20732 4116 20738 4118
rect 20897 4115 20963 4118
rect 18045 4042 18111 4045
rect 14476 4040 14568 4042
rect 14518 3984 14568 4040
rect 14476 3982 14568 3984
rect 17358 4040 18111 4042
rect 17358 3984 18050 4040
rect 18106 3984 18111 4040
rect 17358 3982 18111 3984
rect 14476 3980 14523 3982
rect 14457 3979 14523 3980
rect 18045 3979 18111 3982
rect 4061 3904 8586 3906
rect 4061 3848 4066 3904
rect 4122 3848 8586 3904
rect 4061 3846 8586 3848
rect 9213 3906 9279 3909
rect 9438 3906 9444 3908
rect 9213 3904 9444 3906
rect 9213 3848 9218 3904
rect 9274 3848 9444 3904
rect 9213 3846 9444 3848
rect 4061 3843 4127 3846
rect 9213 3843 9279 3846
rect 9438 3844 9444 3846
rect 9508 3844 9514 3908
rect 11973 3906 12039 3909
rect 13353 3906 13419 3909
rect 11973 3904 13419 3906
rect 11973 3848 11978 3904
rect 12034 3848 13358 3904
rect 13414 3848 13419 3904
rect 11973 3846 13419 3848
rect 11973 3843 12039 3846
rect 13353 3843 13419 3846
rect 16246 3844 16252 3908
rect 16316 3906 16322 3908
rect 17585 3906 17651 3909
rect 16316 3904 17651 3906
rect 16316 3848 17590 3904
rect 17646 3848 17651 3904
rect 16316 3846 17651 3848
rect 16316 3844 16322 3846
rect 17585 3843 17651 3846
rect 17861 3906 17927 3909
rect 18689 3906 18755 3909
rect 22200 3906 23000 3936
rect 17861 3904 18755 3906
rect 17861 3848 17866 3904
rect 17922 3848 18694 3904
rect 18750 3848 18755 3904
rect 17861 3846 18755 3848
rect 17861 3843 17927 3846
rect 18689 3843 18755 3846
rect 20624 3846 23000 3906
rect 3543 3840 3863 3841
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 3775 3863 3776
rect 8741 3840 9061 3841
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 3775 9061 3776
rect 13939 3840 14259 3841
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 3775 14259 3776
rect 19137 3840 19457 3841
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 3775 19457 3776
rect 4705 3770 4771 3773
rect 5717 3770 5783 3773
rect 4705 3768 5783 3770
rect 4705 3712 4710 3768
rect 4766 3712 5722 3768
rect 5778 3712 5783 3768
rect 4705 3710 5783 3712
rect 4705 3707 4771 3710
rect 5717 3707 5783 3710
rect 6269 3770 6335 3773
rect 6862 3770 6868 3772
rect 6269 3768 6868 3770
rect 6269 3712 6274 3768
rect 6330 3712 6868 3768
rect 6269 3710 6868 3712
rect 6269 3707 6335 3710
rect 6862 3708 6868 3710
rect 6932 3708 6938 3772
rect 12709 3770 12775 3773
rect 9216 3768 12775 3770
rect 9216 3712 12714 3768
rect 12770 3712 12775 3768
rect 9216 3710 12775 3712
rect 3877 3634 3943 3637
rect 4102 3634 4108 3636
rect 3877 3632 4108 3634
rect 3877 3576 3882 3632
rect 3938 3576 4108 3632
rect 3877 3574 4108 3576
rect 3877 3571 3943 3574
rect 4102 3572 4108 3574
rect 4172 3572 4178 3636
rect 4889 3634 4955 3637
rect 9216 3634 9276 3710
rect 12709 3707 12775 3710
rect 15193 3770 15259 3773
rect 18965 3770 19031 3773
rect 15193 3768 19031 3770
rect 15193 3712 15198 3768
rect 15254 3712 18970 3768
rect 19026 3712 19031 3768
rect 15193 3710 19031 3712
rect 15193 3707 15259 3710
rect 18965 3707 19031 3710
rect 11973 3634 12039 3637
rect 4889 3632 9276 3634
rect 4889 3576 4894 3632
rect 4950 3576 9276 3632
rect 4889 3574 9276 3576
rect 9400 3632 12039 3634
rect 9400 3576 11978 3632
rect 12034 3576 12039 3632
rect 9400 3574 12039 3576
rect 4889 3571 4955 3574
rect 4470 3498 4476 3500
rect 2730 3438 4476 3498
rect 4470 3436 4476 3438
rect 4540 3498 4546 3500
rect 4889 3498 4955 3501
rect 5257 3500 5323 3501
rect 4540 3496 4955 3498
rect 4540 3440 4894 3496
rect 4950 3440 4955 3496
rect 4540 3438 4955 3440
rect 4540 3436 4546 3438
rect 4889 3435 4955 3438
rect 5206 3436 5212 3500
rect 5276 3498 5323 3500
rect 9400 3498 9460 3574
rect 11973 3571 12039 3574
rect 12341 3634 12407 3637
rect 15285 3634 15351 3637
rect 12341 3632 15351 3634
rect 12341 3576 12346 3632
rect 12402 3576 15290 3632
rect 15346 3576 15351 3632
rect 12341 3574 15351 3576
rect 12341 3571 12407 3574
rect 15285 3571 15351 3574
rect 15837 3634 15903 3637
rect 18689 3634 18755 3637
rect 15837 3632 18755 3634
rect 15837 3576 15842 3632
rect 15898 3576 18694 3632
rect 18750 3576 18755 3632
rect 15837 3574 18755 3576
rect 15837 3571 15903 3574
rect 18689 3571 18755 3574
rect 18965 3634 19031 3637
rect 20624 3634 20684 3846
rect 22200 3816 23000 3846
rect 18965 3632 20684 3634
rect 18965 3576 18970 3632
rect 19026 3576 20684 3632
rect 18965 3574 20684 3576
rect 18965 3571 19031 3574
rect 5276 3496 5368 3498
rect 5318 3440 5368 3496
rect 5276 3438 5368 3440
rect 5582 3438 9460 3498
rect 9765 3498 9831 3501
rect 16021 3498 16087 3501
rect 20621 3498 20687 3501
rect 9765 3496 16087 3498
rect 9765 3440 9770 3496
rect 9826 3440 16026 3496
rect 16082 3440 16087 3496
rect 9765 3438 16087 3440
rect 5276 3436 5323 3438
rect 5257 3435 5323 3436
rect 4981 3362 5047 3365
rect 5582 3362 5642 3438
rect 9765 3435 9831 3438
rect 16021 3435 16087 3438
rect 16254 3496 20687 3498
rect 16254 3440 20626 3496
rect 20682 3440 20687 3496
rect 16254 3438 20687 3440
rect 4981 3360 5642 3362
rect 4981 3304 4986 3360
rect 5042 3304 5642 3360
rect 4981 3302 5642 3304
rect 6729 3362 6795 3365
rect 9949 3362 10015 3365
rect 6729 3360 10015 3362
rect 6729 3304 6734 3360
rect 6790 3304 9954 3360
rect 10010 3304 10015 3360
rect 6729 3302 10015 3304
rect 4981 3299 5047 3302
rect 6729 3299 6795 3302
rect 9949 3299 10015 3302
rect 13077 3362 13143 3365
rect 16254 3362 16314 3438
rect 20621 3435 20687 3438
rect 21633 3498 21699 3501
rect 22200 3498 23000 3528
rect 21633 3496 23000 3498
rect 21633 3440 21638 3496
rect 21694 3440 23000 3496
rect 21633 3438 23000 3440
rect 21633 3435 21699 3438
rect 22200 3408 23000 3438
rect 13077 3360 16314 3362
rect 13077 3304 13082 3360
rect 13138 3304 16314 3360
rect 13077 3302 16314 3304
rect 19333 3362 19399 3365
rect 20713 3362 20779 3365
rect 19333 3360 20779 3362
rect 19333 3304 19338 3360
rect 19394 3304 20718 3360
rect 20774 3304 20779 3360
rect 19333 3302 20779 3304
rect 13077 3299 13143 3302
rect 19333 3299 19399 3302
rect 20713 3299 20779 3302
rect 6142 3296 6462 3297
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 3231 6462 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 16538 3296 16858 3297
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 3231 16858 3232
rect 6729 3226 6795 3229
rect 7230 3226 7236 3228
rect 6729 3224 7236 3226
rect 6729 3168 6734 3224
rect 6790 3168 7236 3224
rect 6729 3166 7236 3168
rect 6729 3163 6795 3166
rect 7230 3164 7236 3166
rect 7300 3164 7306 3228
rect 8293 3226 8359 3229
rect 9581 3226 9647 3229
rect 8293 3224 9647 3226
rect 8293 3168 8298 3224
rect 8354 3168 9586 3224
rect 9642 3168 9647 3224
rect 8293 3166 9647 3168
rect 8293 3163 8359 3166
rect 9581 3163 9647 3166
rect 12341 3226 12407 3229
rect 15653 3226 15719 3229
rect 12341 3224 15719 3226
rect 12341 3168 12346 3224
rect 12402 3168 15658 3224
rect 15714 3168 15719 3224
rect 12341 3166 15719 3168
rect 12341 3163 12407 3166
rect 15653 3163 15719 3166
rect 17585 3226 17651 3229
rect 18781 3226 18847 3229
rect 17585 3224 18847 3226
rect 17585 3168 17590 3224
rect 17646 3168 18786 3224
rect 18842 3168 18847 3224
rect 17585 3166 18847 3168
rect 17585 3163 17651 3166
rect 18781 3163 18847 3166
rect 5441 3090 5507 3093
rect 13905 3090 13971 3093
rect 5441 3088 13971 3090
rect 5441 3032 5446 3088
rect 5502 3032 13910 3088
rect 13966 3032 13971 3088
rect 5441 3030 13971 3032
rect 5441 3027 5507 3030
rect 13905 3027 13971 3030
rect 15837 3090 15903 3093
rect 19425 3090 19491 3093
rect 15837 3088 19491 3090
rect 15837 3032 15842 3088
rect 15898 3032 19430 3088
rect 19486 3032 19491 3088
rect 15837 3030 19491 3032
rect 15837 3027 15903 3030
rect 19425 3027 19491 3030
rect 5257 2954 5323 2957
rect 9581 2954 9647 2957
rect 15009 2954 15075 2957
rect 5257 2952 9276 2954
rect 5257 2896 5262 2952
rect 5318 2896 9276 2952
rect 5257 2894 9276 2896
rect 5257 2891 5323 2894
rect 4797 2818 4863 2821
rect 8017 2818 8083 2821
rect 4797 2816 8083 2818
rect 4797 2760 4802 2816
rect 4858 2760 8022 2816
rect 8078 2760 8083 2816
rect 4797 2758 8083 2760
rect 9216 2818 9276 2894
rect 9581 2952 15075 2954
rect 9581 2896 9586 2952
rect 9642 2896 15014 2952
rect 15070 2896 15075 2952
rect 9581 2894 15075 2896
rect 9581 2891 9647 2894
rect 15009 2891 15075 2894
rect 15469 2954 15535 2957
rect 18321 2954 18387 2957
rect 15469 2952 18387 2954
rect 15469 2896 15474 2952
rect 15530 2896 18326 2952
rect 18382 2896 18387 2952
rect 15469 2894 18387 2896
rect 15469 2891 15535 2894
rect 18321 2891 18387 2894
rect 20621 2954 20687 2957
rect 22200 2954 23000 2984
rect 20621 2952 23000 2954
rect 20621 2896 20626 2952
rect 20682 2896 23000 2952
rect 20621 2894 23000 2896
rect 20621 2891 20687 2894
rect 22200 2864 23000 2894
rect 12801 2818 12867 2821
rect 9216 2816 12867 2818
rect 9216 2760 12806 2816
rect 12862 2760 12867 2816
rect 9216 2758 12867 2760
rect 4797 2755 4863 2758
rect 8017 2755 8083 2758
rect 12801 2755 12867 2758
rect 3543 2752 3863 2753
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2687 3863 2688
rect 8741 2752 9061 2753
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2687 9061 2688
rect 13939 2752 14259 2753
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2687 14259 2688
rect 19137 2752 19457 2753
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2687 19457 2688
rect 5901 2684 5967 2685
rect 5901 2682 5948 2684
rect 5856 2680 5948 2682
rect 5856 2624 5906 2680
rect 5856 2622 5948 2624
rect 5901 2620 5948 2622
rect 6012 2620 6018 2684
rect 6269 2682 6335 2685
rect 6821 2682 6887 2685
rect 6269 2680 6887 2682
rect 6269 2624 6274 2680
rect 6330 2624 6826 2680
rect 6882 2624 6887 2680
rect 6269 2622 6887 2624
rect 5901 2619 5967 2620
rect 6269 2619 6335 2622
rect 6821 2619 6887 2622
rect 7281 2682 7347 2685
rect 7966 2682 7972 2684
rect 7281 2680 7972 2682
rect 7281 2624 7286 2680
rect 7342 2624 7972 2680
rect 7281 2622 7972 2624
rect 7281 2619 7347 2622
rect 7966 2620 7972 2622
rect 8036 2620 8042 2684
rect 9254 2620 9260 2684
rect 9324 2682 9330 2684
rect 9397 2682 9463 2685
rect 9324 2680 9463 2682
rect 9324 2624 9402 2680
rect 9458 2624 9463 2680
rect 9324 2622 9463 2624
rect 9324 2620 9330 2622
rect 9397 2619 9463 2622
rect 9581 2682 9647 2685
rect 13813 2682 13879 2685
rect 9581 2680 13879 2682
rect 9581 2624 9586 2680
rect 9642 2624 13818 2680
rect 13874 2624 13879 2680
rect 9581 2622 13879 2624
rect 9581 2619 9647 2622
rect 13813 2619 13879 2622
rect 15561 2682 15627 2685
rect 15694 2682 15700 2684
rect 15561 2680 15700 2682
rect 15561 2624 15566 2680
rect 15622 2624 15700 2680
rect 15561 2622 15700 2624
rect 15561 2619 15627 2622
rect 15694 2620 15700 2622
rect 15764 2620 15770 2684
rect 4889 2546 4955 2549
rect 9213 2546 9279 2549
rect 4889 2544 9279 2546
rect 4889 2488 4894 2544
rect 4950 2488 9218 2544
rect 9274 2488 9279 2544
rect 4889 2486 9279 2488
rect 4889 2483 4955 2486
rect 9213 2483 9279 2486
rect 11697 2546 11763 2549
rect 20621 2546 20687 2549
rect 11697 2544 20687 2546
rect 11697 2488 11702 2544
rect 11758 2488 20626 2544
rect 20682 2488 20687 2544
rect 11697 2486 20687 2488
rect 11697 2483 11763 2486
rect 20621 2483 20687 2486
rect 22001 2546 22067 2549
rect 22200 2546 23000 2576
rect 22001 2544 23000 2546
rect 22001 2488 22006 2544
rect 22062 2488 23000 2544
rect 22001 2486 23000 2488
rect 22001 2483 22067 2486
rect 22200 2456 23000 2486
rect 1853 2410 1919 2413
rect 18321 2410 18387 2413
rect 1853 2408 18387 2410
rect 1853 2352 1858 2408
rect 1914 2352 18326 2408
rect 18382 2352 18387 2408
rect 1853 2350 18387 2352
rect 1853 2347 1919 2350
rect 18321 2347 18387 2350
rect 6142 2208 6462 2209
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2143 6462 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 16538 2208 16858 2209
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2143 16858 2144
rect 9489 2140 9555 2141
rect 9438 2076 9444 2140
rect 9508 2138 9555 2140
rect 9508 2136 9600 2138
rect 9550 2080 9600 2136
rect 9508 2078 9600 2080
rect 9508 2076 9555 2078
rect 9489 2075 9555 2076
rect 2221 2002 2287 2005
rect 19241 2002 19307 2005
rect 22200 2002 23000 2032
rect 2221 2000 23000 2002
rect 2221 1944 2226 2000
rect 2282 1944 19246 2000
rect 19302 1944 23000 2000
rect 2221 1942 23000 1944
rect 2221 1939 2287 1942
rect 19241 1939 19307 1942
rect 22200 1912 23000 1942
rect 2681 1866 2747 1869
rect 17033 1866 17099 1869
rect 2681 1864 17099 1866
rect 2681 1808 2686 1864
rect 2742 1808 17038 1864
rect 17094 1808 17099 1864
rect 2681 1806 17099 1808
rect 2681 1803 2747 1806
rect 17033 1803 17099 1806
rect 6545 1730 6611 1733
rect 15009 1730 15075 1733
rect 6545 1728 15075 1730
rect 6545 1672 6550 1728
rect 6606 1672 15014 1728
rect 15070 1672 15075 1728
rect 6545 1670 15075 1672
rect 6545 1667 6611 1670
rect 15009 1667 15075 1670
rect 17033 1730 17099 1733
rect 18270 1730 18276 1732
rect 17033 1728 18276 1730
rect 17033 1672 17038 1728
rect 17094 1672 18276 1728
rect 17033 1670 18276 1672
rect 17033 1667 17099 1670
rect 18270 1668 18276 1670
rect 18340 1668 18346 1732
rect 2773 1594 2839 1597
rect 8937 1594 9003 1597
rect 2773 1592 9003 1594
rect 2773 1536 2778 1592
rect 2834 1536 8942 1592
rect 8998 1536 9003 1592
rect 2773 1534 9003 1536
rect 2773 1531 2839 1534
rect 8937 1531 9003 1534
rect 12065 1594 12131 1597
rect 17769 1594 17835 1597
rect 21357 1594 21423 1597
rect 22200 1594 23000 1624
rect 12065 1592 17835 1594
rect 12065 1536 12070 1592
rect 12126 1536 17774 1592
rect 17830 1536 17835 1592
rect 12065 1534 17835 1536
rect 12065 1531 12131 1534
rect 17769 1531 17835 1534
rect 18646 1592 23000 1594
rect 18646 1536 21362 1592
rect 21418 1536 23000 1592
rect 18646 1534 23000 1536
rect 3969 1458 4035 1461
rect 12617 1458 12683 1461
rect 3969 1456 12683 1458
rect 3969 1400 3974 1456
rect 4030 1400 12622 1456
rect 12678 1400 12683 1456
rect 3969 1398 12683 1400
rect 3969 1395 4035 1398
rect 12617 1395 12683 1398
rect 5390 1260 5396 1324
rect 5460 1322 5466 1324
rect 7005 1322 7071 1325
rect 5460 1320 7071 1322
rect 5460 1264 7010 1320
rect 7066 1264 7071 1320
rect 5460 1262 7071 1264
rect 5460 1260 5466 1262
rect 7005 1259 7071 1262
rect 8293 1322 8359 1325
rect 17125 1322 17191 1325
rect 8293 1320 17191 1322
rect 8293 1264 8298 1320
rect 8354 1264 17130 1320
rect 17186 1264 17191 1320
rect 8293 1262 17191 1264
rect 8293 1259 8359 1262
rect 17125 1259 17191 1262
rect 8150 1124 8156 1188
rect 8220 1186 8226 1188
rect 18646 1186 18706 1534
rect 21357 1531 21423 1534
rect 22200 1504 23000 1534
rect 8220 1126 18706 1186
rect 19241 1186 19307 1189
rect 19241 1184 19994 1186
rect 19241 1128 19246 1184
rect 19302 1128 19994 1184
rect 19241 1126 19994 1128
rect 8220 1124 8226 1126
rect 19241 1123 19307 1126
rect 7414 988 7420 1052
rect 7484 1050 7490 1052
rect 19701 1050 19767 1053
rect 7484 1048 19767 1050
rect 7484 992 19706 1048
rect 19762 992 19767 1048
rect 7484 990 19767 992
rect 19934 1050 19994 1126
rect 22200 1050 23000 1080
rect 19934 990 23000 1050
rect 7484 988 7490 990
rect 19701 987 19767 990
rect 22200 960 23000 990
rect 1577 914 1643 917
rect 18505 914 18571 917
rect 19057 914 19123 917
rect 1577 912 18571 914
rect 1577 856 1582 912
rect 1638 856 18510 912
rect 18566 856 18571 912
rect 1577 854 18571 856
rect 1577 851 1643 854
rect 18505 851 18571 854
rect 18646 912 19123 914
rect 18646 856 19062 912
rect 19118 856 19123 912
rect 18646 854 19123 856
rect 7833 778 7899 781
rect 18646 778 18706 854
rect 19057 851 19123 854
rect 7833 776 18706 778
rect 7833 720 7838 776
rect 7894 720 18706 776
rect 7833 718 18706 720
rect 7833 715 7899 718
rect 2037 642 2103 645
rect 17534 642 17540 644
rect 2037 640 17540 642
rect 2037 584 2042 640
rect 2098 584 17540 640
rect 2037 582 17540 584
rect 2037 579 2103 582
rect 17534 580 17540 582
rect 17604 580 17610 644
rect 21817 642 21883 645
rect 22200 642 23000 672
rect 21817 640 23000 642
rect 21817 584 21822 640
rect 21878 584 23000 640
rect 21817 582 23000 584
rect 21817 579 21883 582
rect 22200 552 23000 582
rect 17953 234 18019 237
rect 22200 234 23000 264
rect 17953 232 23000 234
rect 17953 176 17958 232
rect 18014 176 23000 232
rect 17953 174 23000 176
rect 17953 171 18019 174
rect 22200 144 23000 174
<< via3 >>
rect 5028 21932 5092 21996
rect 5396 21524 5460 21588
rect 2268 20844 2332 20908
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 13676 20300 13740 20364
rect 7236 20164 7300 20228
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 4844 19680 4908 19684
rect 4844 19624 4858 19680
rect 4858 19624 4908 19680
rect 4844 19620 4908 19624
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 5948 19484 6012 19548
rect 7236 19484 7300 19548
rect 17172 19484 17236 19548
rect 20668 19484 20732 19548
rect 7788 19348 7852 19412
rect 9260 19076 9324 19140
rect 10916 19136 10980 19140
rect 10916 19080 10930 19136
rect 10930 19080 10980 19136
rect 10916 19076 10980 19080
rect 12204 19076 12268 19140
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 5028 19000 5092 19004
rect 5028 18944 5078 19000
rect 5078 18944 5092 19000
rect 5028 18940 5092 18944
rect 5396 19000 5460 19004
rect 5396 18944 5410 19000
rect 5410 18944 5460 19000
rect 5396 18940 5460 18944
rect 5948 18940 6012 19004
rect 13676 18804 13740 18868
rect 5764 18668 5828 18732
rect 2268 18396 2332 18460
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 17540 17988 17604 18052
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 9260 17172 9324 17236
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 5028 16824 5092 16828
rect 5028 16768 5042 16824
rect 5042 16768 5092 16824
rect 5028 16764 5092 16768
rect 8524 16628 8588 16692
rect 4844 16492 4908 16556
rect 6868 16492 6932 16556
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 10916 14724 10980 14788
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 5948 14180 6012 14244
rect 14780 14240 14844 14244
rect 14780 14184 14794 14240
rect 14794 14184 14844 14240
rect 14780 14180 14844 14184
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 15700 14044 15764 14108
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 12204 13500 12268 13564
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 6868 13092 6932 13156
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 8524 12820 8588 12884
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 8340 12276 8404 12340
rect 14780 12004 14844 12068
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 12020 10644 12084 10708
rect 17908 10508 17972 10572
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 9628 10100 9692 10164
rect 9812 10100 9876 10164
rect 12020 10100 12084 10164
rect 9628 9964 9692 10028
rect 4108 9828 4172 9892
rect 9628 9828 9692 9892
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 5212 9556 5276 9620
rect 7236 9556 7300 9620
rect 14596 9284 14660 9348
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 8156 9148 8220 9212
rect 17172 9148 17236 9212
rect 5580 8876 5644 8940
rect 7236 8740 7300 8804
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 7788 8528 7852 8532
rect 7788 8472 7802 8528
rect 7802 8472 7852 8528
rect 7788 8468 7852 8472
rect 14596 8468 14660 8532
rect 18828 8468 18892 8532
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 18276 8060 18340 8124
rect 7604 7652 7668 7716
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 4476 7380 4540 7444
rect 7604 7380 7668 7444
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 8156 6972 8220 7036
rect 4844 6896 4908 6900
rect 4844 6840 4858 6896
rect 4858 6840 4908 6896
rect 4844 6836 4908 6840
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 17908 6428 17972 6492
rect 7972 6020 8036 6084
rect 9260 6080 9324 6084
rect 9260 6024 9274 6080
rect 9274 6024 9324 6080
rect 9260 6020 9324 6024
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 5948 5476 6012 5540
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 5396 5340 5460 5404
rect 5764 4932 5828 4996
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 7788 4796 7852 4860
rect 17540 4796 17604 4860
rect 7420 4524 7484 4588
rect 8524 4388 8588 4452
rect 17172 4524 17236 4588
rect 15148 4388 15212 4452
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 5580 3980 5644 4044
rect 6868 4040 6932 4044
rect 6868 3984 6882 4040
rect 6882 3984 6932 4040
rect 6868 3980 6932 3984
rect 14412 4040 14476 4044
rect 17540 4116 17604 4180
rect 20668 4116 20732 4180
rect 14412 3984 14462 4040
rect 14462 3984 14476 4040
rect 14412 3980 14476 3984
rect 9444 3844 9508 3908
rect 16252 3844 16316 3908
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 6868 3708 6932 3772
rect 4108 3572 4172 3636
rect 4476 3436 4540 3500
rect 5212 3496 5276 3500
rect 5212 3440 5262 3496
rect 5262 3440 5276 3496
rect 5212 3436 5276 3440
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 7236 3164 7300 3228
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 5948 2680 6012 2684
rect 5948 2624 5962 2680
rect 5962 2624 6012 2680
rect 5948 2620 6012 2624
rect 7972 2620 8036 2684
rect 9260 2620 9324 2684
rect 15700 2620 15764 2684
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 9444 2136 9508 2140
rect 9444 2080 9494 2136
rect 9494 2080 9508 2136
rect 9444 2076 9508 2080
rect 18276 1668 18340 1732
rect 5396 1260 5460 1324
rect 8156 1124 8220 1188
rect 7420 988 7484 1052
rect 17540 580 17604 644
<< metal4 >>
rect 5027 21996 5093 21997
rect 5027 21932 5028 21996
rect 5092 21932 5093 21996
rect 5027 21931 5093 21932
rect 2267 20908 2333 20909
rect 2267 20844 2268 20908
rect 2332 20844 2333 20908
rect 2267 20843 2333 20844
rect 2270 18461 2330 20843
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 4843 19684 4909 19685
rect 4843 19620 4844 19684
rect 4908 19620 4909 19684
rect 4843 19619 4909 19620
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 2267 18460 2333 18461
rect 2267 18396 2268 18460
rect 2332 18396 2333 18460
rect 2267 18395 2333 18396
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 4846 16557 4906 19619
rect 5030 19005 5090 21931
rect 5395 21588 5461 21589
rect 5395 21524 5396 21588
rect 5460 21524 5461 21588
rect 5395 21523 5461 21524
rect 5398 19005 5458 21523
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 7235 20228 7301 20229
rect 7235 20164 7236 20228
rect 7300 20164 7301 20228
rect 7235 20163 7301 20164
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 5947 19548 6013 19549
rect 5947 19484 5948 19548
rect 6012 19484 6013 19548
rect 5947 19483 6013 19484
rect 5950 19005 6010 19483
rect 5027 19004 5093 19005
rect 5027 18940 5028 19004
rect 5092 18940 5093 19004
rect 5027 18939 5093 18940
rect 5395 19004 5461 19005
rect 5395 18940 5396 19004
rect 5460 18940 5461 19004
rect 5395 18939 5461 18940
rect 5947 19004 6013 19005
rect 5947 18940 5948 19004
rect 6012 18940 6013 19004
rect 5947 18939 6013 18940
rect 5763 18732 5829 18733
rect 5763 18668 5764 18732
rect 5828 18668 5829 18732
rect 5763 18667 5829 18668
rect 5027 16828 5093 16829
rect 5027 16764 5028 16828
rect 5092 16764 5093 16828
rect 5027 16763 5093 16764
rect 4843 16556 4909 16557
rect 4843 16492 4844 16556
rect 4908 16492 4909 16556
rect 4843 16491 4909 16492
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 5030 12698 5090 16763
rect 5766 14058 5826 18667
rect 5950 14245 6010 18939
rect 6142 18528 6462 19552
rect 7238 19549 7298 20163
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 7235 19548 7301 19549
rect 7235 19484 7236 19548
rect 7300 19484 7301 19548
rect 7235 19483 7301 19484
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6867 16492 6868 16542
rect 6932 16492 6933 16542
rect 6867 16491 6933 16492
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 5947 14244 6013 14245
rect 5947 14180 5948 14244
rect 6012 14180 6013 14244
rect 5947 14179 6013 14180
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6867 13156 6933 13157
rect 6867 13092 6868 13156
rect 6932 13092 6933 13156
rect 6867 13091 6933 13092
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 4107 9892 4173 9893
rect 4107 9828 4108 9892
rect 4172 9828 4173 9892
rect 4107 9827 4173 9828
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 4110 3637 4170 9827
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 5211 9620 5277 9621
rect 5211 9556 5212 9620
rect 5276 9556 5277 9620
rect 5211 9555 5277 9556
rect 4475 7444 4541 7445
rect 4475 7380 4476 7444
rect 4540 7380 4541 7444
rect 4475 7379 4541 7380
rect 4107 3636 4173 3637
rect 4107 3572 4108 3636
rect 4172 3572 4173 3636
rect 4107 3571 4173 3572
rect 4478 3501 4538 7379
rect 4846 6901 4906 7022
rect 4843 6900 4909 6901
rect 4843 6836 4844 6900
rect 4908 6836 4909 6900
rect 4843 6835 4909 6836
rect 5214 3501 5274 9555
rect 5579 8940 5645 8941
rect 5579 8876 5580 8940
rect 5644 8876 5645 8940
rect 5579 8875 5645 8876
rect 5582 7170 5642 8875
rect 5398 7110 5642 7170
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 5398 5810 5458 7110
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 5398 5750 5642 5810
rect 5395 5404 5461 5405
rect 5395 5340 5396 5404
rect 5460 5340 5461 5404
rect 5395 5339 5461 5340
rect 4475 3500 4541 3501
rect 4475 3436 4476 3500
rect 4540 3436 4541 3500
rect 4475 3435 4541 3436
rect 5211 3500 5277 3501
rect 5211 3436 5212 3500
rect 5276 3436 5277 3500
rect 5211 3435 5277 3436
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 5398 1325 5458 5339
rect 5582 4045 5642 5750
rect 5766 4997 5826 6342
rect 5947 5540 6013 5541
rect 5947 5476 5948 5540
rect 6012 5476 6013 5540
rect 5947 5475 6013 5476
rect 5763 4996 5829 4997
rect 5763 4932 5764 4996
rect 5828 4932 5829 4996
rect 5763 4931 5829 4932
rect 5579 4044 5645 4045
rect 5579 3980 5580 4044
rect 5644 3980 5645 4044
rect 5579 3979 5645 3980
rect 5950 2685 6010 5475
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6870 4045 6930 13091
rect 7238 12450 7298 19483
rect 7787 19412 7853 19413
rect 7787 19348 7788 19412
rect 7852 19348 7853 19412
rect 7787 19347 7853 19348
rect 7238 12390 7666 12450
rect 7238 9621 7298 10422
rect 7235 9620 7301 9621
rect 7235 9556 7236 9620
rect 7300 9556 7301 9620
rect 7235 9555 7301 9556
rect 7235 8804 7301 8805
rect 7235 8740 7236 8804
rect 7300 8740 7301 8804
rect 7235 8739 7301 8740
rect 6867 4044 6933 4045
rect 6867 3980 6868 4044
rect 6932 3980 6933 4044
rect 6867 3979 6933 3980
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 5947 2684 6013 2685
rect 5947 2620 5948 2684
rect 6012 2620 6013 2684
rect 5947 2619 6013 2620
rect 6142 2208 6462 3232
rect 7238 3229 7298 8739
rect 7606 7717 7666 12390
rect 7790 8533 7850 19347
rect 8741 19072 9061 20096
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 13675 20364 13741 20365
rect 13675 20300 13676 20364
rect 13740 20300 13741 20364
rect 13675 20299 13741 20300
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 9259 19140 9325 19141
rect 9259 19076 9260 19140
rect 9324 19076 9325 19140
rect 9259 19075 9325 19076
rect 10915 19140 10981 19141
rect 10915 19076 10916 19140
rect 10980 19076 10981 19140
rect 10915 19075 10981 19076
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8342 12341 8402 17902
rect 8741 16896 9061 17920
rect 9262 17237 9322 19075
rect 9259 17236 9325 17237
rect 9259 17172 9260 17236
rect 9324 17172 9325 17236
rect 9259 17171 9325 17172
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8523 16692 8589 16693
rect 8523 16628 8524 16692
rect 8588 16628 8589 16692
rect 8523 16627 8589 16628
rect 8526 12885 8586 16627
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 10918 14789 10978 19075
rect 11340 18528 11660 19552
rect 12203 19140 12269 19141
rect 12203 19076 12204 19140
rect 12268 19076 12269 19140
rect 12203 19075 12269 19076
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 10915 14788 10981 14789
rect 10915 14724 10916 14788
rect 10980 14724 10981 14788
rect 10915 14723 10981 14724
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8523 12884 8589 12885
rect 8523 12820 8524 12884
rect 8588 12820 8589 12884
rect 8523 12819 8589 12820
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8339 12340 8405 12341
rect 8339 12276 8340 12340
rect 8404 12276 8405 12340
rect 8339 12275 8405 12276
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 12206 13565 12266 19075
rect 13678 18869 13738 20299
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13675 18868 13741 18869
rect 13675 18804 13676 18868
rect 13740 18804 13741 18868
rect 13675 18803 13741 18804
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 17171 19548 17237 19549
rect 17171 19484 17172 19548
rect 17236 19484 17237 19548
rect 17171 19483 17237 19484
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 17174 18138 17234 19483
rect 19137 19072 19457 20096
rect 20667 19548 20733 19549
rect 20667 19484 20668 19548
rect 20732 19484 20733 19548
rect 20667 19483 20733 19484
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 17539 18052 17605 18053
rect 17539 17988 17540 18052
rect 17604 17988 17605 18052
rect 17539 17987 17605 17988
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 14779 14244 14845 14245
rect 14779 14180 14780 14244
rect 14844 14180 14845 14244
rect 14779 14179 14845 14180
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 12203 13564 12269 13565
rect 12203 13500 12204 13564
rect 12268 13500 12269 13564
rect 12203 13499 12269 13500
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 9627 10164 9693 10165
rect 9627 10100 9628 10164
rect 9692 10162 9693 10164
rect 9811 10164 9877 10165
rect 9811 10162 9812 10164
rect 9692 10102 9812 10162
rect 9692 10100 9693 10102
rect 9627 10099 9693 10100
rect 9811 10100 9812 10102
rect 9876 10100 9877 10164
rect 9811 10099 9877 10100
rect 9627 10028 9693 10029
rect 9627 9964 9628 10028
rect 9692 9964 9693 10028
rect 9627 9963 9693 9964
rect 9630 9893 9690 9963
rect 9627 9892 9693 9893
rect 9627 9828 9628 9892
rect 9692 9828 9693 9892
rect 9627 9827 9693 9828
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 7787 8532 7853 8533
rect 7787 8468 7788 8532
rect 7852 8468 7853 8532
rect 7787 8467 7853 8468
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 7603 7716 7669 7717
rect 7603 7652 7604 7716
rect 7668 7652 7669 7716
rect 7603 7651 7669 7652
rect 7606 7445 7666 7651
rect 7603 7444 7669 7445
rect 7603 7380 7604 7444
rect 7668 7380 7669 7444
rect 7603 7379 7669 7380
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8155 7036 8221 7037
rect 8155 6972 8156 7036
rect 8220 6972 8221 7036
rect 8155 6971 8221 6972
rect 7971 6084 8037 6085
rect 7971 6020 7972 6084
rect 8036 6020 8037 6084
rect 7971 6019 8037 6020
rect 7787 4860 7853 4861
rect 7787 4796 7788 4860
rect 7852 4796 7853 4860
rect 7787 4795 7853 4796
rect 7419 4588 7485 4589
rect 7419 4524 7420 4588
rect 7484 4524 7485 4588
rect 7419 4523 7485 4524
rect 7235 3228 7301 3229
rect 7235 3164 7236 3228
rect 7300 3164 7301 3228
rect 7235 3163 7301 3164
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 5395 1324 5461 1325
rect 5395 1260 5396 1324
rect 5460 1260 5461 1324
rect 5395 1259 5461 1260
rect 7422 1053 7482 4523
rect 7790 2498 7850 4795
rect 7974 2685 8034 6019
rect 7971 2684 8037 2685
rect 7971 2620 7972 2684
rect 8036 2620 8037 2684
rect 7971 2619 8037 2620
rect 8158 1189 8218 6971
rect 8741 6016 9061 7040
rect 11340 9824 11660 10848
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 12019 10708 12085 10709
rect 12019 10644 12020 10708
rect 12084 10644 12085 10708
rect 12019 10643 12085 10644
rect 12022 10165 12082 10643
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 12019 10164 12085 10165
rect 12019 10100 12020 10164
rect 12084 10100 12085 10164
rect 12019 10099 12085 10100
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 9259 6084 9325 6085
rect 9259 6020 9260 6084
rect 9324 6020 9325 6084
rect 9259 6019 9325 6020
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 9262 2685 9322 6019
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 9443 3908 9509 3909
rect 9443 3844 9444 3908
rect 9508 3844 9509 3908
rect 9443 3843 9509 3844
rect 9259 2684 9325 2685
rect 9259 2620 9260 2684
rect 9324 2620 9325 2684
rect 9259 2619 9325 2620
rect 9446 2141 9506 3843
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 9443 2140 9509 2141
rect 9443 2076 9444 2140
rect 9508 2076 9509 2140
rect 11340 2128 11660 2144
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 14414 4045 14474 12462
rect 14782 12069 14842 14179
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 15699 14108 15765 14109
rect 15699 14044 15700 14108
rect 15764 14044 15765 14108
rect 15699 14043 15765 14044
rect 14779 12068 14845 12069
rect 14779 12004 14780 12068
rect 14844 12004 14845 12068
rect 14779 12003 14845 12004
rect 14595 9348 14661 9349
rect 14595 9284 14596 9348
rect 14660 9284 14661 9348
rect 14595 9283 14661 9284
rect 14598 8533 14658 9283
rect 14595 8532 14661 8533
rect 14595 8468 14596 8532
rect 14660 8468 14661 8532
rect 14595 8467 14661 8468
rect 14411 4044 14477 4045
rect 14411 3980 14412 4044
rect 14476 3980 14477 4044
rect 14411 3979 14477 3980
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 15702 2685 15762 14043
rect 16254 3909 16314 13822
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 17542 4861 17602 17987
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 20670 16778 20730 19483
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 18827 8532 18893 8533
rect 18827 8468 18828 8532
rect 18892 8468 18893 8532
rect 18827 8467 18893 8468
rect 18275 8124 18341 8125
rect 18275 8060 18276 8124
rect 18340 8060 18341 8124
rect 18275 8059 18341 8060
rect 17539 4860 17605 4861
rect 17539 4796 17540 4860
rect 17604 4796 17605 4860
rect 17539 4795 17605 4796
rect 17171 4588 17237 4589
rect 17171 4524 17172 4588
rect 17236 4524 17237 4588
rect 17171 4523 17237 4524
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16251 3908 16317 3909
rect 16251 3844 16252 3908
rect 16316 3844 16317 3908
rect 16251 3843 16317 3844
rect 16538 3296 16858 4320
rect 17174 3858 17234 4523
rect 17539 4180 17605 4181
rect 17539 4116 17540 4180
rect 17604 4116 17605 4180
rect 17539 4115 17605 4116
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 15699 2684 15765 2685
rect 15699 2620 15700 2684
rect 15764 2620 15765 2684
rect 15699 2619 15765 2620
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 9443 2075 9509 2076
rect 8155 1188 8221 1189
rect 8155 1124 8156 1188
rect 8220 1124 8221 1188
rect 8155 1123 8221 1124
rect 7419 1052 7485 1053
rect 7419 988 7420 1052
rect 7484 988 7485 1052
rect 7419 987 7485 988
rect 17542 645 17602 4115
rect 18278 1733 18338 8059
rect 18830 7258 18890 8467
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 20667 4180 20733 4181
rect 20667 4116 20668 4180
rect 20732 4116 20733 4180
rect 20667 4115 20733 4116
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 20670 2498 20730 4115
rect 18275 1732 18341 1733
rect 18275 1668 18276 1732
rect 18340 1668 18341 1732
rect 18275 1667 18341 1668
rect 17539 644 17605 645
rect 17539 580 17540 644
rect 17604 580 17605 644
rect 17539 579 17605 580
<< via4 >>
rect 6782 16556 7018 16778
rect 6782 16542 6868 16556
rect 6868 16542 6932 16556
rect 6932 16542 7018 16556
rect 5678 13822 5914 14058
rect 4942 12462 5178 12698
rect 4758 7022 4994 7258
rect 5678 6342 5914 6578
rect 7150 10422 7386 10658
rect 6782 3772 7018 3858
rect 6782 3708 6868 3772
rect 6868 3708 6932 3772
rect 6932 3708 7018 3772
rect 6782 3622 7018 3708
rect 8254 17902 8490 18138
rect 8070 9212 8306 9298
rect 8070 9148 8156 9212
rect 8156 9148 8220 9212
rect 8220 9148 8306 9212
rect 8070 9062 8306 9148
rect 17086 17902 17322 18138
rect 7702 2262 7938 2498
rect 14326 12462 14562 12698
rect 8438 4452 8674 4538
rect 8438 4388 8524 4452
rect 8524 4388 8588 4452
rect 8588 4388 8674 4452
rect 8438 4302 8674 4388
rect 15062 4452 15298 4538
rect 15062 4388 15148 4452
rect 15148 4388 15212 4452
rect 15212 4388 15298 4452
rect 15062 4302 15298 4388
rect 16166 13822 16402 14058
rect 17086 9212 17322 9298
rect 17086 9148 17172 9212
rect 17172 9148 17236 9212
rect 17236 9148 17322 9212
rect 17086 9062 17322 9148
rect 20582 16542 20818 16778
rect 17822 10572 18058 10658
rect 17822 10508 17908 10572
rect 17908 10508 17972 10572
rect 17972 10508 18058 10572
rect 17822 10422 18058 10508
rect 17822 6492 18058 6578
rect 17822 6428 17908 6492
rect 17908 6428 17972 6492
rect 17972 6428 18058 6492
rect 17822 6342 18058 6428
rect 17086 3622 17322 3858
rect 18742 7022 18978 7258
rect 20582 2262 20818 2498
<< metal5 >>
rect 8212 18138 17364 18180
rect 8212 17902 8254 18138
rect 8490 17902 17086 18138
rect 17322 17902 17364 18138
rect 8212 17860 17364 17902
rect 6740 16778 20860 16820
rect 6740 16542 6782 16778
rect 7018 16542 20582 16778
rect 20818 16542 20860 16778
rect 6740 16500 20860 16542
rect 5636 14058 16444 14100
rect 5636 13822 5678 14058
rect 5914 13822 16166 14058
rect 16402 13822 16444 14058
rect 5636 13780 16444 13822
rect 4900 12698 14604 12740
rect 4900 12462 4942 12698
rect 5178 12462 14326 12698
rect 14562 12462 14604 12698
rect 4900 12420 14604 12462
rect 7108 10658 18100 10700
rect 7108 10422 7150 10658
rect 7386 10422 17822 10658
rect 18058 10422 18100 10658
rect 7108 10380 18100 10422
rect 8028 9298 17364 9340
rect 8028 9062 8070 9298
rect 8306 9062 17086 9298
rect 17322 9062 17364 9298
rect 8028 9020 17364 9062
rect 4716 7258 19020 7300
rect 4716 7022 4758 7258
rect 4994 7022 18742 7258
rect 18978 7022 19020 7258
rect 4716 6980 19020 7022
rect 5636 6578 18100 6620
rect 5636 6342 5678 6578
rect 5914 6342 17822 6578
rect 18058 6342 18100 6578
rect 5636 6300 18100 6342
rect 8396 4538 15340 4580
rect 8396 4302 8438 4538
rect 8674 4302 15062 4538
rect 15298 4302 15340 4538
rect 8396 4260 15340 4302
rect 6740 3858 17364 3900
rect 6740 3622 6782 3858
rect 7018 3622 17086 3858
rect 17322 3622 17364 3858
rect 6740 3580 17364 3622
rect 7660 2498 20860 2540
rect 7660 2262 7702 2498
rect 7938 2262 20582 2498
rect 20818 2262 20860 2498
rect 7660 2220 20860 2262
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3128 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1649977179
transform -1 0 4508 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform 1 0 3772 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1649977179
transform 1 0 3312 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1649977179
transform -1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform -1 0 3404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1649977179
transform -1 0 1656 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1649977179
transform 1 0 4416 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1649977179
transform -1 0 2392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1649977179
transform -1 0 1932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1649977179
transform -1 0 2300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1649977179
transform 1 0 3036 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1649977179
transform 1 0 4048 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1649977179
transform -1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1649977179
transform 1 0 4232 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1649977179
transform -1 0 3312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1649977179
transform -1 0 2944 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1649977179
transform -1 0 3128 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1649977179
transform -1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform -1 0 4048 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1649977179
transform -1 0 1564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1649977179
transform -1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1649977179
transform 1 0 5796 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1649977179
transform -1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1649977179
transform 1 0 4048 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1649977179
transform -1 0 1656 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1649977179
transform -1 0 5336 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1649977179
transform -1 0 4968 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold45_A
timestamp 1649977179
transform -1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 1564 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 2024 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 2760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 10764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 17940 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 6992 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 7176 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 7544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 7544 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 19412 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 6624 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 3772 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 5336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 4140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 3404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 4968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 5704 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 5980 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 3128 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 2668 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 4876 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 3128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 2024 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 2392 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 2024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 2392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 3588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 4232 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 2760 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 5704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 2392 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 2024 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 3496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 1932 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 3680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 2668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 3036 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 1840 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 3404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 4968 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 2300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 2024 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 2024 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 2576 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 2760 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 3128 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 1840 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 4416 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 3864 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 2576 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 5244 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 4232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 5336 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 2300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 6624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 6256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 6900 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform -1 0 1564 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6808 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6532 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7176 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 16836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6900 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 4968 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 1564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 4692 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8004 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7636 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8004 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9384 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16192 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 16836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5612 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10580 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 12512 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5520 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 5244 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5152 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 7728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4692 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 5612 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 5152 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 4508 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 4140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5520 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 4600 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4416 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4324 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 4140 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5612 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 4784 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6440 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7360 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6716 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 3036 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.sky130_fd_sc_hd__buf_4_0__A
timestamp 1649977179
transform -1 0 5060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1649977179
transform -1 0 2392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 1932 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.sky130_fd_sc_hd__buf_4_0__A
timestamp 1649977179
transform -1 0 2760 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.sky130_fd_sc_hd__buf_4_0__A
timestamp 1649977179
transform -1 0 5244 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5520 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5152 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6164 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7728 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 7544 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 14720 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 15272 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6808 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 6624 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 6900 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 4600 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 7268 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1649977179
transform -1 0 2116 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1649977179
transform -1 0 2760 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1649977179
transform -1 0 5612 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output97_A
timestamp 1649977179
transform 1 0 6992 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output98_A
timestamp 1649977179
transform -1 0 6532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output99_A
timestamp 1649977179
transform 1 0 6440 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output112_A
timestamp 1649977179
transform 1 0 6624 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 2208 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1649977179
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32
timestamp 1649977179
transform 1 0 4048 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42
timestamp 1649977179
transform 1 0 4968 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48
timestamp 1649977179
transform 1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1649977179
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64
timestamp 1649977179
transform 1 0 6992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70
timestamp 1649977179
transform 1 0 7544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76
timestamp 1649977179
transform 1 0 8096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_87
timestamp 1649977179
transform 1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_93
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_105
timestamp 1649977179
transform 1 0 10764 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_127
timestamp 1649977179
transform 1 0 12788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1649977179
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_144
timestamp 1649977179
transform 1 0 14352 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_155
timestamp 1649977179
transform 1 0 15364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1649977179
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_178
timestamp 1649977179
transform 1 0 17480 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_183
timestamp 1649977179
transform 1 0 17940 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1649977179
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_6
timestamp 1649977179
transform 1 0 1656 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_11
timestamp 1649977179
transform 1 0 2116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_16
timestamp 1649977179
transform 1 0 2576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_21
timestamp 1649977179
transform 1 0 3036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_26
timestamp 1649977179
transform 1 0 3496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_32 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4048 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_44
timestamp 1649977179
transform 1 0 5152 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_49
timestamp 1649977179
transform 1 0 5612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1649977179
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_63
timestamp 1649977179
transform 1 0 6900 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_68
timestamp 1649977179
transform 1 0 7360 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_74
timestamp 1649977179
transform 1 0 7912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_80
timestamp 1649977179
transform 1 0 8464 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_90
timestamp 1649977179
transform 1 0 9384 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_100
timestamp 1649977179
transform 1 0 10304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_113 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_122
timestamp 1649977179
transform 1 0 12328 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_133
timestamp 1649977179
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_144
timestamp 1649977179
transform 1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_171
timestamp 1649977179
transform 1 0 16836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_189
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1649977179
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1649977179
transform 1 0 20332 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1649977179
transform 1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_5
timestamp 1649977179
transform 1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_9
timestamp 1649977179
transform 1 0 1932 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_13
timestamp 1649977179
transform 1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_17
timestamp 1649977179
transform 1 0 2668 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_21
timestamp 1649977179
transform 1 0 3036 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_34
timestamp 1649977179
transform 1 0 4232 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_39
timestamp 1649977179
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_44
timestamp 1649977179
transform 1 0 5152 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_49
timestamp 1649977179
transform 1 0 5612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_54
timestamp 1649977179
transform 1 0 6072 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_59
timestamp 1649977179
transform 1 0 6532 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_64
timestamp 1649977179
transform 1 0 6992 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_69
timestamp 1649977179
transform 1 0 7452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_75
timestamp 1649977179
transform 1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1649977179
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_95
timestamp 1649977179
transform 1 0 9844 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_106
timestamp 1649977179
transform 1 0 10856 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_124
timestamp 1649977179
transform 1 0 12512 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_128
timestamp 1649977179
transform 1 0 12880 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_157
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1649977179
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_208
timestamp 1649977179
transform 1 0 20240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_219
timestamp 1649977179
transform 1 0 21252 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_5
timestamp 1649977179
transform 1 0 1564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_9
timestamp 1649977179
transform 1 0 1932 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_13
timestamp 1649977179
transform 1 0 2300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1649977179
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_21
timestamp 1649977179
transform 1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_25
timestamp 1649977179
transform 1 0 3404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_29
timestamp 1649977179
transform 1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_34
timestamp 1649977179
transform 1 0 4232 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1649977179
transform 1 0 5152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_49
timestamp 1649977179
transform 1 0 5612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1649977179
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_63
timestamp 1649977179
transform 1 0 6900 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_68
timestamp 1649977179
transform 1 0 7360 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_73
timestamp 1649977179
transform 1 0 7820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_78
timestamp 1649977179
transform 1 0 8280 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_83
timestamp 1649977179
transform 1 0 8740 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 1649977179
transform 1 0 9292 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_99
timestamp 1649977179
transform 1 0 10212 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1649977179
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1649977179
transform 1 0 12420 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_134
timestamp 1649977179
transform 1 0 13432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_147
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_158
timestamp 1649977179
transform 1 0 15640 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_173
timestamp 1649977179
transform 1 0 17020 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 1649977179
transform 1 0 18032 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_202
timestamp 1649977179
transform 1 0 19688 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_208
timestamp 1649977179
transform 1 0 20240 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1649977179
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_6
timestamp 1649977179
transform 1 0 1656 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_10
timestamp 1649977179
transform 1 0 2024 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_14
timestamp 1649977179
transform 1 0 2392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_18
timestamp 1649977179
transform 1 0 2760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_22
timestamp 1649977179
transform 1 0 3128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1649977179
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_34
timestamp 1649977179
transform 1 0 4232 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_38
timestamp 1649977179
transform 1 0 4600 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_42
timestamp 1649977179
transform 1 0 4968 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_47
timestamp 1649977179
transform 1 0 5428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_52
timestamp 1649977179
transform 1 0 5888 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_57
timestamp 1649977179
transform 1 0 6348 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_62
timestamp 1649977179
transform 1 0 6808 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_67
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_72
timestamp 1649977179
transform 1 0 7728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_87
timestamp 1649977179
transform 1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_105
timestamp 1649977179
transform 1 0 10764 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_123
timestamp 1649977179
transform 1 0 12420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_134
timestamp 1649977179
transform 1 0 13432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_145
timestamp 1649977179
transform 1 0 14444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 1649977179
transform 1 0 15640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_169
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_180
timestamp 1649977179
transform 1 0 17664 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_191
timestamp 1649977179
transform 1 0 18676 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_213
timestamp 1649977179
transform 1 0 20700 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1649977179
transform 1 0 21252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_5
timestamp 1649977179
transform 1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_9
timestamp 1649977179
transform 1 0 1932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_13
timestamp 1649977179
transform 1 0 2300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_17
timestamp 1649977179
transform 1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_21
timestamp 1649977179
transform 1 0 3036 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_25
timestamp 1649977179
transform 1 0 3404 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_29
timestamp 1649977179
transform 1 0 3772 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_33
timestamp 1649977179
transform 1 0 4140 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_37
timestamp 1649977179
transform 1 0 4508 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_41
timestamp 1649977179
transform 1 0 4876 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_45
timestamp 1649977179
transform 1 0 5244 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_49
timestamp 1649977179
transform 1 0 5612 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1649977179
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_62
timestamp 1649977179
transform 1 0 6808 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_67
timestamp 1649977179
transform 1 0 7268 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_72
timestamp 1649977179
transform 1 0 7728 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_77
timestamp 1649977179
transform 1 0 8188 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_87
timestamp 1649977179
transform 1 0 9108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_97
timestamp 1649977179
transform 1 0 10028 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_129
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_147
timestamp 1649977179
transform 1 0 14628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1649977179
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1649977179
transform 1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_194
timestamp 1649977179
transform 1 0 18952 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_198
timestamp 1649977179
transform 1 0 19320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_208
timestamp 1649977179
transform 1 0 20240 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1649977179
transform 1 0 21436 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_6
timestamp 1649977179
transform 1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_10
timestamp 1649977179
transform 1 0 2024 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_14
timestamp 1649977179
transform 1 0 2392 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_18
timestamp 1649977179
transform 1 0 2760 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_22
timestamp 1649977179
transform 1 0 3128 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1649977179
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_34
timestamp 1649977179
transform 1 0 4232 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_38
timestamp 1649977179
transform 1 0 4600 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_42
timestamp 1649977179
transform 1 0 4968 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_46
timestamp 1649977179
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_50
timestamp 1649977179
transform 1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_54
timestamp 1649977179
transform 1 0 6072 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 1649977179
transform 1 0 6532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_95
timestamp 1649977179
transform 1 0 9844 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_99
timestamp 1649977179
transform 1 0 10212 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1649977179
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_152
timestamp 1649977179
transform 1 0 15088 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_156
timestamp 1649977179
transform 1 0 15456 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_178
timestamp 1649977179
transform 1 0 17480 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_191
timestamp 1649977179
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_213
timestamp 1649977179
transform 1 0 20700 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 1649977179
transform 1 0 21252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1649977179
transform 1 0 1656 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_10
timestamp 1649977179
transform 1 0 2024 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_7_14 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2392 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_20
timestamp 1649977179
transform 1 0 2944 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_23
timestamp 1649977179
transform 1 0 3220 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_31
timestamp 1649977179
transform 1 0 3956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_35
timestamp 1649977179
transform 1 0 4324 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_38
timestamp 1649977179
transform 1 0 4600 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_42
timestamp 1649977179
transform 1 0 4968 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_46
timestamp 1649977179
transform 1 0 5336 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_50
timestamp 1649977179
transform 1 0 5704 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_60
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_65
timestamp 1649977179
transform 1 0 7084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_70
timestamp 1649977179
transform 1 0 7544 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_88
timestamp 1649977179
transform 1 0 9200 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_98
timestamp 1649977179
transform 1 0 10120 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1649977179
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_122
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_128
timestamp 1649977179
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_146
timestamp 1649977179
transform 1 0 14536 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_172
timestamp 1649977179
transform 1 0 16928 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_190
timestamp 1649977179
transform 1 0 18584 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_208
timestamp 1649977179
transform 1 0 20240 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_220
timestamp 1649977179
transform 1 0 21344 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1564 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_17 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1649977179
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_34
timestamp 1649977179
transform 1 0 4232 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_38
timestamp 1649977179
transform 1 0 4600 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_45
timestamp 1649977179
transform 1 0 5244 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_49
timestamp 1649977179
transform 1 0 5612 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_57
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_61
timestamp 1649977179
transform 1 0 6716 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_71
timestamp 1649977179
transform 1 0 7636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_87
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_98
timestamp 1649977179
transform 1 0 10120 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_127
timestamp 1649977179
transform 1 0 12788 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1649977179
transform 1 0 14352 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_155
timestamp 1649977179
transform 1 0 15364 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_166
timestamp 1649977179
transform 1 0 16376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_188
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_215
timestamp 1649977179
transform 1 0 20884 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_43
timestamp 1649977179
transform 1 0 5060 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_46
timestamp 1649977179
transform 1 0 5336 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_50
timestamp 1649977179
transform 1 0 5704 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_61
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_65
timestamp 1649977179
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_83
timestamp 1649977179
transform 1 0 8740 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1649977179
transform 1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1649977179
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_121
timestamp 1649977179
transform 1 0 12236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_132
timestamp 1649977179
transform 1 0 13248 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_144
timestamp 1649977179
transform 1 0 14352 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_148
timestamp 1649977179
transform 1 0 14720 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1649977179
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_172
timestamp 1649977179
transform 1 0 16928 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_190
timestamp 1649977179
transform 1 0 18584 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_201
timestamp 1649977179
transform 1 0 19596 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_212
timestamp 1649977179
transform 1 0 20608 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_216
timestamp 1649977179
transform 1 0 20976 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1649977179
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_56
timestamp 1649977179
transform 1 0 6256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_60
timestamp 1649977179
transform 1 0 6624 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_64
timestamp 1649977179
transform 1 0 6992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_68
timestamp 1649977179
transform 1 0 7360 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_78
timestamp 1649977179
transform 1 0 8280 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_89
timestamp 1649977179
transform 1 0 9292 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_99
timestamp 1649977179
transform 1 0 10212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_132
timestamp 1649977179
transform 1 0 13248 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1649977179
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_150
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_156
timestamp 1649977179
transform 1 0 15456 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_178
timestamp 1649977179
transform 1 0 17480 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1649977179
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_199
timestamp 1649977179
transform 1 0 19412 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_217
timestamp 1649977179
transform 1 0 21068 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_62
timestamp 1649977179
transform 1 0 6808 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 1649977179
transform 1 0 7176 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_70
timestamp 1649977179
transform 1 0 7544 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_74
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_79
timestamp 1649977179
transform 1 0 8372 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_89
timestamp 1649977179
transform 1 0 9292 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_107
timestamp 1649977179
transform 1 0 10948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_122
timestamp 1649977179
transform 1 0 12328 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_140
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_145
timestamp 1649977179
transform 1 0 14444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_171
timestamp 1649977179
transform 1 0 16836 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_182
timestamp 1649977179
transform 1 0 17848 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_199
timestamp 1649977179
transform 1 0 19412 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1649977179
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_57
timestamp 1649977179
transform 1 0 6348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_60
timestamp 1649977179
transform 1 0 6624 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_64
timestamp 1649977179
transform 1 0 6992 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_68
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_72
timestamp 1649977179
transform 1 0 7728 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_88
timestamp 1649977179
transform 1 0 9200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_99
timestamp 1649977179
transform 1 0 10212 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_110
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_114
timestamp 1649977179
transform 1 0 11592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_118
timestamp 1649977179
transform 1 0 11960 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_160
timestamp 1649977179
transform 1 0 15824 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_171
timestamp 1649977179
transform 1 0 16836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_182
timestamp 1649977179
transform 1 0 17848 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_193
timestamp 1649977179
transform 1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_206
timestamp 1649977179
transform 1 0 20056 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_217
timestamp 1649977179
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_62
timestamp 1649977179
transform 1 0 6808 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_66
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_70
timestamp 1649977179
transform 1 0 7544 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_80
timestamp 1649977179
transform 1 0 8464 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_90
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_121
timestamp 1649977179
transform 1 0 12236 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_131
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_142
timestamp 1649977179
transform 1 0 14168 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_153
timestamp 1649977179
transform 1 0 15180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_179
timestamp 1649977179
transform 1 0 17572 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_183
timestamp 1649977179
transform 1 0 17940 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_201
timestamp 1649977179
transform 1 0 19596 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_212
timestamp 1649977179
transform 1 0 20608 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_216
timestamp 1649977179
transform 1 0 20976 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_59
timestamp 1649977179
transform 1 0 6532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_63
timestamp 1649977179
transform 1 0 6900 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_67
timestamp 1649977179
transform 1 0 7268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_72
timestamp 1649977179
transform 1 0 7728 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1649977179
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_99
timestamp 1649977179
transform 1 0 10212 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_119
timestamp 1649977179
transform 1 0 12052 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_123
timestamp 1649977179
transform 1 0 12420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_134
timestamp 1649977179
transform 1 0 13432 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1649977179
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_150
timestamp 1649977179
transform 1 0 14904 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_161
timestamp 1649977179
transform 1 0 15916 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_169
timestamp 1649977179
transform 1 0 16652 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_187
timestamp 1649977179
transform 1 0 18308 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_213
timestamp 1649977179
transform 1 0 20700 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_219
timestamp 1649977179
transform 1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_60
timestamp 1649977179
transform 1 0 6624 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_64
timestamp 1649977179
transform 1 0 6992 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_68
timestamp 1649977179
transform 1 0 7360 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_73
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 1649977179
transform 1 0 8280 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_88
timestamp 1649977179
transform 1 0 9200 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_99
timestamp 1649977179
transform 1 0 10212 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_131
timestamp 1649977179
transform 1 0 13156 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 1649977179
transform 1 0 13616 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_147
timestamp 1649977179
transform 1 0 14628 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1649977179
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_164
timestamp 1649977179
transform 1 0 16192 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_185
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_203
timestamp 1649977179
transform 1 0 19780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_63
timestamp 1649977179
transform 1 0 6900 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_67
timestamp 1649977179
transform 1 0 7268 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_72
timestamp 1649977179
transform 1 0 7728 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_87
timestamp 1649977179
transform 1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_92
timestamp 1649977179
transform 1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_110
timestamp 1649977179
transform 1 0 11224 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_132
timestamp 1649977179
transform 1 0 13248 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1649977179
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_147
timestamp 1649977179
transform 1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_176
timestamp 1649977179
transform 1 0 17296 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_187
timestamp 1649977179
transform 1 0 18308 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_214
timestamp 1649977179
transform 1 0 20792 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_65
timestamp 1649977179
transform 1 0 7084 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_74
timestamp 1649977179
transform 1 0 7912 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_84
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_102
timestamp 1649977179
transform 1 0 10488 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_106
timestamp 1649977179
transform 1 0 10856 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_131
timestamp 1649977179
transform 1 0 13156 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_135
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_185
timestamp 1649977179
transform 1 0 18124 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_196
timestamp 1649977179
transform 1 0 19136 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_207
timestamp 1649977179
transform 1 0 20148 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_218
timestamp 1649977179
transform 1 0 21160 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_222
timestamp 1649977179
transform 1 0 21528 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_72
timestamp 1649977179
transform 1 0 7728 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_101
timestamp 1649977179
transform 1 0 10396 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_106
timestamp 1649977179
transform 1 0 10856 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_110
timestamp 1649977179
transform 1 0 11224 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_120
timestamp 1649977179
transform 1 0 12144 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_168
timestamp 1649977179
transform 1 0 16560 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_181
timestamp 1649977179
transform 1 0 17756 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_200
timestamp 1649977179
transform 1 0 19504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_219
timestamp 1649977179
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_77
timestamp 1649977179
transform 1 0 8188 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_82
timestamp 1649977179
transform 1 0 8648 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_101
timestamp 1649977179
transform 1 0 10396 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_117
timestamp 1649977179
transform 1 0 11868 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_121
timestamp 1649977179
transform 1 0 12236 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_131
timestamp 1649977179
transform 1 0 13156 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_141
timestamp 1649977179
transform 1 0 14076 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_145
timestamp 1649977179
transform 1 0 14444 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_155
timestamp 1649977179
transform 1 0 15364 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1649977179
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_185
timestamp 1649977179
transform 1 0 18124 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_206
timestamp 1649977179
transform 1 0 20056 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1649977179
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_69
timestamp 1649977179
transform 1 0 7452 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_73
timestamp 1649977179
transform 1 0 7820 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1649977179
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_95
timestamp 1649977179
transform 1 0 9844 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_99
timestamp 1649977179
transform 1 0 10212 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_132
timestamp 1649977179
transform 1 0 13248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_137
timestamp 1649977179
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_144
timestamp 1649977179
transform 1 0 14352 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_155
timestamp 1649977179
transform 1 0 15364 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_178
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_188
timestamp 1649977179
transform 1 0 18400 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1649977179
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1649977179
transform 1 0 20056 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_217
timestamp 1649977179
transform 1 0 21068 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_65
timestamp 1649977179
transform 1 0 7084 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_70
timestamp 1649977179
transform 1 0 7544 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_74
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_79
timestamp 1649977179
transform 1 0 8372 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_89
timestamp 1649977179
transform 1 0 9292 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1649977179
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_129
timestamp 1649977179
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_133
timestamp 1649977179
transform 1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_138
timestamp 1649977179
transform 1 0 13800 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_160
timestamp 1649977179
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_165
timestamp 1649977179
transform 1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_185
timestamp 1649977179
transform 1 0 18124 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1649977179
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_207
timestamp 1649977179
transform 1 0 20148 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_218
timestamp 1649977179
transform 1 0 21160 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_222
timestamp 1649977179
transform 1 0 21528 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_63
timestamp 1649977179
transform 1 0 6900 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_67
timestamp 1649977179
transform 1 0 7268 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_72
timestamp 1649977179
transform 1 0 7728 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1649977179
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_115
timestamp 1649977179
transform 1 0 11684 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_120
timestamp 1649977179
transform 1 0 12144 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_150
timestamp 1649977179
transform 1 0 14904 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_161
timestamp 1649977179
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_166
timestamp 1649977179
transform 1 0 16376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_186
timestamp 1649977179
transform 1 0 18216 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1649977179
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_203
timestamp 1649977179
transform 1 0 19780 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_214
timestamp 1649977179
transform 1 0 20792 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_220
timestamp 1649977179
transform 1 0 21344 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_60
timestamp 1649977179
transform 1 0 6624 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_65
timestamp 1649977179
transform 1 0 7084 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_70
timestamp 1649977179
transform 1 0 7544 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_88
timestamp 1649977179
transform 1 0 9200 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_92
timestamp 1649977179
transform 1 0 9568 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1649977179
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_122
timestamp 1649977179
transform 1 0 12328 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_127
timestamp 1649977179
transform 1 0 12788 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_138
timestamp 1649977179
transform 1 0 13800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_156
timestamp 1649977179
transform 1 0 15456 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1649977179
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_177
timestamp 1649977179
transform 1 0 17388 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_186
timestamp 1649977179
transform 1 0 18216 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_197
timestamp 1649977179
transform 1 0 19228 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_215
timestamp 1649977179
transform 1 0 20884 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1649977179
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_51
timestamp 1649977179
transform 1 0 5796 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_56
timestamp 1649977179
transform 1 0 6256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_61
timestamp 1649977179
transform 1 0 6716 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_71
timestamp 1649977179
transform 1 0 7636 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1649977179
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_94
timestamp 1649977179
transform 1 0 9752 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_99
timestamp 1649977179
transform 1 0 10212 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_132
timestamp 1649977179
transform 1 0 13248 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1649977179
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_151
timestamp 1649977179
transform 1 0 14996 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_156
timestamp 1649977179
transform 1 0 15456 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_178
timestamp 1649977179
transform 1 0 17480 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1649977179
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_213
timestamp 1649977179
transform 1 0 20700 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_42
timestamp 1649977179
transform 1 0 4968 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_46
timestamp 1649977179
transform 1 0 5336 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_50
timestamp 1649977179
transform 1 0 5704 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1649977179
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_67
timestamp 1649977179
transform 1 0 7268 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_85
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_89
timestamp 1649977179
transform 1 0 9292 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_99
timestamp 1649977179
transform 1 0 10212 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1649977179
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_116
timestamp 1649977179
transform 1 0 11776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_127
timestamp 1649977179
transform 1 0 12788 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_138
timestamp 1649977179
transform 1 0 13800 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_148
timestamp 1649977179
transform 1 0 14720 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_178
timestamp 1649977179
transform 1 0 17480 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_196
timestamp 1649977179
transform 1 0 19136 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_207
timestamp 1649977179
transform 1 0 20148 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_218
timestamp 1649977179
transform 1 0 21160 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_222
timestamp 1649977179
transform 1 0 21528 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_10
timestamp 1649977179
transform 1 0 2024 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_16
timestamp 1649977179
transform 1 0 2576 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_33
timestamp 1649977179
transform 1 0 4140 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_36
timestamp 1649977179
transform 1 0 4416 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_40
timestamp 1649977179
transform 1 0 4784 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_43
timestamp 1649977179
transform 1 0 5060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_47
timestamp 1649977179
transform 1 0 5428 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_51
timestamp 1649977179
transform 1 0 5796 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_56
timestamp 1649977179
transform 1 0 6256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_61
timestamp 1649977179
transform 1 0 6716 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_79
timestamp 1649977179
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_115
timestamp 1649977179
transform 1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1649977179
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_150
timestamp 1649977179
transform 1 0 14904 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_162
timestamp 1649977179
transform 1 0 16008 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_173
timestamp 1649977179
transform 1 0 17020 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_184
timestamp 1649977179
transform 1 0 18032 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1649977179
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1649977179
transform 1 0 20056 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_217
timestamp 1649977179
transform 1 0 21068 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_5
timestamp 1649977179
transform 1 0 1564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_10
timestamp 1649977179
transform 1 0 2024 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_14
timestamp 1649977179
transform 1 0 2392 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_18
timestamp 1649977179
transform 1 0 2760 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_22
timestamp 1649977179
transform 1 0 3128 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_26
timestamp 1649977179
transform 1 0 3496 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_30
timestamp 1649977179
transform 1 0 3864 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_34
timestamp 1649977179
transform 1 0 4232 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_42
timestamp 1649977179
transform 1 0 4968 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_46
timestamp 1649977179
transform 1 0 5336 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_50
timestamp 1649977179
transform 1 0 5704 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_61
timestamp 1649977179
transform 1 0 6716 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_71
timestamp 1649977179
transform 1 0 7636 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_89
timestamp 1649977179
transform 1 0 9292 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_101
timestamp 1649977179
transform 1 0 10396 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1649977179
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_122
timestamp 1649977179
transform 1 0 12328 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_126
timestamp 1649977179
transform 1 0 12696 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_144
timestamp 1649977179
transform 1 0 14352 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_162
timestamp 1649977179
transform 1 0 16008 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1649977179
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_171
timestamp 1649977179
transform 1 0 16836 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_189
timestamp 1649977179
transform 1 0 18492 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_207
timestamp 1649977179
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1649977179
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_11
timestamp 1649977179
transform 1 0 2116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_18
timestamp 1649977179
transform 1 0 2760 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_22
timestamp 1649977179
transform 1 0 3128 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1649977179
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_33
timestamp 1649977179
transform 1 0 4140 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_37
timestamp 1649977179
transform 1 0 4508 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_45
timestamp 1649977179
transform 1 0 5244 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_49
timestamp 1649977179
transform 1 0 5612 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 1649977179
transform 1 0 6900 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 1649977179
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_101
timestamp 1649977179
transform 1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_112
timestamp 1649977179
transform 1 0 11408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_122
timestamp 1649977179
transform 1 0 12328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_127
timestamp 1649977179
transform 1 0 12788 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1649977179
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_150
timestamp 1649977179
transform 1 0 14904 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_160
timestamp 1649977179
transform 1 0 15824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_179
timestamp 1649977179
transform 1 0 17572 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_190
timestamp 1649977179
transform 1 0 18584 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1649977179
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_206
timestamp 1649977179
transform 1 0 20056 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_217
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_8
timestamp 1649977179
transform 1 0 1840 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_12
timestamp 1649977179
transform 1 0 2208 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_16
timestamp 1649977179
transform 1 0 2576 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_20
timestamp 1649977179
transform 1 0 2944 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_24
timestamp 1649977179
transform 1 0 3312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_28
timestamp 1649977179
transform 1 0 3680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_32
timestamp 1649977179
transform 1 0 4048 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_36
timestamp 1649977179
transform 1 0 4416 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_40
timestamp 1649977179
transform 1 0 4784 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_44
timestamp 1649977179
transform 1 0 5152 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_49
timestamp 1649977179
transform 1 0 5612 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_63
timestamp 1649977179
transform 1 0 6900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_68
timestamp 1649977179
transform 1 0 7360 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_79
timestamp 1649977179
transform 1 0 8372 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_83
timestamp 1649977179
transform 1 0 8740 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_88
timestamp 1649977179
transform 1 0 9200 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_99
timestamp 1649977179
transform 1 0 10212 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1649977179
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_122
timestamp 1649977179
transform 1 0 12328 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_130
timestamp 1649977179
transform 1 0 13064 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_140
timestamp 1649977179
transform 1 0 13984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_146
timestamp 1649977179
transform 1 0 14536 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_157
timestamp 1649977179
transform 1 0 15548 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_179
timestamp 1649977179
transform 1 0 17572 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_199
timestamp 1649977179
transform 1 0 19412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_210
timestamp 1649977179
transform 1 0 20424 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_6
timestamp 1649977179
transform 1 0 1656 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_10
timestamp 1649977179
transform 1 0 2024 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_14
timestamp 1649977179
transform 1 0 2392 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_18
timestamp 1649977179
transform 1 0 2760 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_22
timestamp 1649977179
transform 1 0 3128 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1649977179
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_33
timestamp 1649977179
transform 1 0 4140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_37
timestamp 1649977179
transform 1 0 4508 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_42
timestamp 1649977179
transform 1 0 4968 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_47
timestamp 1649977179
transform 1 0 5428 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_52
timestamp 1649977179
transform 1 0 5888 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_57
timestamp 1649977179
transform 1 0 6348 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_62
timestamp 1649977179
transform 1 0 6808 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_67
timestamp 1649977179
transform 1 0 7268 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_72
timestamp 1649977179
transform 1 0 7728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1649977179
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_104
timestamp 1649977179
transform 1 0 10672 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_115
timestamp 1649977179
transform 1 0 11684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_151
timestamp 1649977179
transform 1 0 14996 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_171
timestamp 1649977179
transform 1 0 16836 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 1649977179
transform 1 0 17296 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_186
timestamp 1649977179
transform 1 0 18216 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1649977179
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_206
timestamp 1649977179
transform 1 0 20056 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_211
timestamp 1649977179
transform 1 0 20516 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_5
timestamp 1649977179
transform 1 0 1564 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_9
timestamp 1649977179
transform 1 0 1932 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_13
timestamp 1649977179
transform 1 0 2300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_17
timestamp 1649977179
transform 1 0 2668 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_21
timestamp 1649977179
transform 1 0 3036 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_25
timestamp 1649977179
transform 1 0 3404 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_29
timestamp 1649977179
transform 1 0 3772 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_34
timestamp 1649977179
transform 1 0 4232 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_44
timestamp 1649977179
transform 1 0 5152 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_49
timestamp 1649977179
transform 1 0 5612 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_54
timestamp 1649977179
transform 1 0 6072 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_61
timestamp 1649977179
transform 1 0 6716 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_66
timestamp 1649977179
transform 1 0 7176 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_71
timestamp 1649977179
transform 1 0 7636 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_76
timestamp 1649977179
transform 1 0 8096 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_86
timestamp 1649977179
transform 1 0 9016 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_92
timestamp 1649977179
transform 1 0 9568 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1649977179
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_122
timestamp 1649977179
transform 1 0 12328 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_128
timestamp 1649977179
transform 1 0 12880 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_146
timestamp 1649977179
transform 1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1649977179
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_173
timestamp 1649977179
transform 1 0 17020 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1649977179
transform 1 0 17572 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_185
timestamp 1649977179
transform 1 0 18124 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_191
timestamp 1649977179
transform 1 0 18676 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1649977179
transform 1 0 19228 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1649977179
transform 1 0 19780 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_215
timestamp 1649977179
transform 1 0 20884 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_9
timestamp 1649977179
transform 1 0 1932 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_20
timestamp 1649977179
transform 1 0 2944 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1649977179
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_31
timestamp 1649977179
transform 1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_36
timestamp 1649977179
transform 1 0 4416 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_46
timestamp 1649977179
transform 1 0 5336 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_51
timestamp 1649977179
transform 1 0 5796 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_56
timestamp 1649977179
transform 1 0 6256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_61
timestamp 1649977179
transform 1 0 6716 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_66
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_71
timestamp 1649977179
transform 1 0 7636 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_76
timestamp 1649977179
transform 1 0 8096 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1649977179
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_88
timestamp 1649977179
transform 1 0 9200 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_94
timestamp 1649977179
transform 1 0 9752 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_105
timestamp 1649977179
transform 1 0 10764 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_123
timestamp 1649977179
transform 1 0 12420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1649977179
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_145
timestamp 1649977179
transform 1 0 14444 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_156
timestamp 1649977179
transform 1 0 15456 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_161
timestamp 1649977179
transform 1 0 15916 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_171
timestamp 1649977179
transform 1 0 16836 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_183
timestamp 1649977179
transform 1 0 17940 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1649977179
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_201
timestamp 1649977179
transform 1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_217
timestamp 1649977179
transform 1 0 21068 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_8
timestamp 1649977179
transform 1 0 1840 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_14
timestamp 1649977179
transform 1 0 2392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_19
timestamp 1649977179
transform 1 0 2852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_26
timestamp 1649977179
transform 1 0 3496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_32
timestamp 1649977179
transform 1 0 4048 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_38
timestamp 1649977179
transform 1 0 4600 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_42
timestamp 1649977179
transform 1 0 4968 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_48
timestamp 1649977179
transform 1 0 5520 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1649977179
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_63
timestamp 1649977179
transform 1 0 6900 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_75
timestamp 1649977179
transform 1 0 8004 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_91
timestamp 1649977179
transform 1 0 9476 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_99
timestamp 1649977179
transform 1 0 10212 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1649977179
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_123
timestamp 1649977179
transform 1 0 12420 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_133
timestamp 1649977179
transform 1 0 13340 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_138
timestamp 1649977179
transform 1 0 13800 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_145
timestamp 1649977179
transform 1 0 14444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_151
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_157
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1649977179
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_173
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1649977179
transform 1 0 17572 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_185
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1649977179
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_195
timestamp 1649977179
transform 1 0 19044 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_201
timestamp 1649977179
transform 1 0 19596 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_207
timestamp 1649977179
transform 1 0 20148 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_213
timestamp 1649977179
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _066_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7728 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1649977179
transform -1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1649977179
transform -1 0 18952 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1649977179
transform -1 0 6716 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform -1 0 7084 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform -1 0 13800 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform -1 0 11224 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform -1 0 15456 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform -1 0 16376 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform 1 0 11868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform -1 0 8556 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform -1 0 7268 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform -1 0 7728 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform -1 0 5428 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform -1 0 11776 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform -1 0 4968 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform -1 0 8188 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform -1 0 4692 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform -1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform -1 0 6072 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform -1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform -1 0 8188 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform -1 0 6992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform -1 0 4232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform -1 0 5612 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform -1 0 7268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform -1 0 7820 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform -1 0 6072 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform -1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform -1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform -1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform -1 0 5152 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 3496 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform -1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform -1 0 5428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform -1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform -1 0 5888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform -1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform -1 0 7176 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform -1 0 7452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform -1 0 8096 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1649977179
transform -1 0 9016 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 6256 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1649977179
transform -1 0 7176 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1649977179
transform -1 0 6716 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1649977179
transform -1 0 6808 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1649977179
transform -1 0 5152 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1649977179
transform -1 0 6900 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1649977179
transform -1 0 18952 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1649977179
transform -1 0 13800 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1649977179
transform -1 0 5796 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1649977179
transform -1 0 12788 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1649977179
transform -1 0 7636 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1649977179
transform -1 0 5336 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1649977179
transform -1 0 4416 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1649977179
transform -1 0 4876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1649977179
transform -1 0 6072 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1649977179
transform -1 0 6348 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15916 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 12236 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 12236 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 15640 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 12236 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 12236 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 15640 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 15640 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9844 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold2 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15824 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold3
timestamp 1649977179
transform 1 0 8464 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1649977179
transform -1 0 21068 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1649977179
transform -1 0 9384 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1649977179
transform -1 0 18952 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1649977179
transform -1 0 8464 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1649977179
transform -1 0 18216 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1649977179
transform -1 0 8648 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1649977179
transform -1 0 21436 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1649977179
transform -1 0 13156 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1649977179
transform 1 0 13340 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1649977179
transform -1 0 10304 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1649977179
transform 1 0 13248 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1649977179
transform -1 0 8648 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1649977179
transform -1 0 17480 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1649977179
transform 1 0 16100 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1649977179
transform 1 0 6900 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1649977179
transform -1 0 8832 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1649977179
transform -1 0 9384 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold22
timestamp 1649977179
transform -1 0 21436 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1649977179
transform -1 0 12236 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1649977179
transform -1 0 9292 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1649977179
transform -1 0 11224 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1649977179
transform -1 0 10212 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1649977179
transform 1 0 11592 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1649977179
transform 1 0 11592 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1649977179
transform -1 0 12328 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1649977179
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1649977179
transform 1 0 7544 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1649977179
transform -1 0 10120 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1649977179
transform -1 0 20056 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1649977179
transform -1 0 9108 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1649977179
transform -1 0 12788 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1649977179
transform -1 0 6900 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1649977179
transform -1 0 10212 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1649977179
transform -1 0 14720 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1649977179
transform -1 0 10028 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1649977179
transform -1 0 8648 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1649977179
transform 1 0 7912 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1649977179
transform -1 0 7636 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1649977179
transform -1 0 8648 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1649977179
transform -1 0 7636 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 4876 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 11960 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 16928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 14628 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 16192 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 8372 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 7728 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 8188 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 16376 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 7820 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 6348 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 6808 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 7268 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 7728 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform -1 0 11224 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 7544 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input24 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 6532 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform 1 0 7636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform -1 0 6992 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1649977179
transform -1 0 7912 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1649977179
transform 1 0 9844 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1649977179
transform -1 0 9292 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform -1 0 7544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1649977179
transform 1 0 3128 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform 1 0 3680 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1649977179
transform 1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 3496 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1649977179
transform -1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1649977179
transform 1 0 5704 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 2944 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1649977179
transform 1 0 6532 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform -1 0 4048 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1649977179
transform 1 0 7636 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1649977179
transform 1 0 8188 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1649977179
transform 1 0 9108 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform -1 0 8096 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform 1 0 9844 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1649977179
transform 1 0 10396 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform -1 0 7636 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform -1 0 2484 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1649977179
transform 1 0 2024 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform -1 0 2852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1649977179
transform 1 0 3128 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1649977179
transform 1 0 3128 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1649977179
transform 1 0 4232 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform -1 0 4232 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input61
timestamp 1649977179
transform 1 0 5152 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input62
timestamp 1649977179
transform 1 0 5704 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1649977179
transform -1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1649977179
transform -1 0 21252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1649977179
transform -1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1649977179
transform -1 0 21436 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1649977179
transform -1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1649977179
transform 1 0 1564 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17112 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18584 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16376 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14904 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15824 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12144 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12512 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14536 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12788 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9292 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12420 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 13156 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14904 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18768 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 19412 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19596 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19780 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20056 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18216 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12328 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13984 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16376 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10212 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11868 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12880 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16008 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8372 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 9200 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8556 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7820 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9200 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9752 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10948 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11868 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13064 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14720 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15364 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16100 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17020 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17940 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18676 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17664 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20700 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19412 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10212 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10948 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10396 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9016 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11040 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14628 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15916 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18216 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16928 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6716 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7728 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8740 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10948 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11040 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10580 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11684 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11684 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12328 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16284 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18308 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18124 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 19780 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19320 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 19780 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18768 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 19412 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 19780 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17848 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l2_in_1__155 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17940 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16560 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17020 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16008 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_3.mux_l2_in_1__158
timestamp 1649977179
transform -1 0 9292 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14352 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17572 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13524 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15364 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12972 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15548 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l2_in_1__160
timestamp 1649977179
transform -1 0 14352 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12420 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13340 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11592 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12604 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_1__161
timestamp 1649977179
transform -1 0 9292 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10856 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10396 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7084 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15640 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform -1 0 15640 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16652 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15088 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_17.mux_l2_in_1__156
timestamp 1649977179
transform -1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16836 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13800 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13340 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15364 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l2_in_1__157
timestamp 1649977179
transform -1 0 8648 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform -1 0 13800 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1649977179
transform -1 0 21252 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_33.mux_l1_in_1__159
timestamp 1649977179
transform -1 0 13616 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1649977179
transform -1 0 20332 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20424 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 19320 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 17940 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18308 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 17756 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_0.mux_l2_in_1__162
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 18308 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8372 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13800 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 14812 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1649977179
transform 1 0 15548 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1649977179
transform 1 0 15088 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_2.mux_l1_in_3__135
timestamp 1649977179
transform -1 0 13800 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14996 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15364 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18676 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10028 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10396 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 17664 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_4.mux_l1_in_3__145
timestamp 1649977179
transform 1 0 13432 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1649977179
transform 1 0 12420 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10212 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12788 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12972 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12788 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13800 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14168 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_2_
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_6.mux_l1_in_3__146
timestamp 1649977179
transform -1 0 7360 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_3_
timestamp 1649977179
transform -1 0 16008 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16192 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20240 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7268 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_8.mux_l2_in_1__147
timestamp 1649977179
transform -1 0 6716 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9200 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8096 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8372 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_10.mux_l2_in_1__163
timestamp 1649977179
transform -1 0 9200 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9568 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10212 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9936 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10764 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_12.mux_l2_in_1__164
timestamp 1649977179
transform 1 0 15640 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10856 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9200 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13616 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14996 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15456 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_14.mux_l2_in_1__165
timestamp 1649977179
transform -1 0 6072 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14720 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7728 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 17572 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_16.mux_l1_in_1__133
timestamp 1649977179
transform -1 0 7544 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18584 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_1_
timestamp 1649977179
transform -1 0 20424 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_18.mux_l1_in_1__134
timestamp 1649977179
transform -1 0 5612 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20240 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13800 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1649977179
transform -1 0 20148 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20332 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_20.mux_l1_in_1__136
timestamp 1649977179
transform -1 0 6256 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20240 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6716 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1649977179
transform -1 0 19228 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_1_
timestamp 1649977179
transform 1 0 20332 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_22.mux_l1_in_1__137
timestamp 1649977179
transform -1 0 16652 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19964 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 17020 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12144 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12420 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_24.mux_l2_in_1__138
timestamp 1649977179
transform -1 0 11040 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10948 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11408 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9844 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_26.mux_l2_in_0__139
timestamp 1649977179
transform -1 0 8648 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10580 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10212 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_28.mux_l2_in_0__140
timestamp 1649977179
transform 1 0 10948 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10212 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 11592 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14352 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_30.mux_l2_in_0__141
timestamp 1649977179
transform -1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13800 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 5336 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17480 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_32.mux_l2_in_0__142
timestamp 1649977179
transform -1 0 6900 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17572 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_34.mux_l2_in_0__143
timestamp 1649977179
transform -1 0 6072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6440 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18032 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_36.mux_l2_in_0__144
timestamp 1649977179
transform -1 0 14352 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8372 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10212 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10304 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9016 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10120 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8648 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_0.mux_l2_in_1__148
timestamp 1649977179
transform -1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12420 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_2.mux_l2_in_1__150
timestamp 1649977179
transform -1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10212 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10396 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15088 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12604 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_4.mux_l2_in_1__153
timestamp 1649977179
transform 1 0 13432 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 11224 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13248 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 13432 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16468 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17480 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15732 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14628 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_8.mux_l2_in_1__154
timestamp 1649977179
transform -1 0 16284 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15732 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14536 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18860 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18032 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_16.mux_l2_in_1__149
timestamp 1649977179
transform -1 0 8648 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17020 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16744 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20240 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19780 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20332 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_24.mux_l2_in_1__151
timestamp 1649977179
transform -1 0 8280 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19320 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9292 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20608 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20516 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1649977179
transform -1 0 21068 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_32.mux_l2_in_1__152
timestamp 1649977179
transform -1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1649977179
transform 1 0 20240 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7452 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output72 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform 1 0 20976 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 17848 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 9568 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 12512 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform 1 0 17204 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 19412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 18308 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 18124 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform 1 0 17572 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 18584 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform 1 0 21068 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 19412 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 18584 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 16008 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 21068 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform 1 0 18584 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform 1 0 12512 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform 1 0 18584 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform 1 0 20884 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 20884 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform 1 0 8280 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform 1 0 18676 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform 1 0 18584 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform 1 0 8280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform 1 0 8096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform 1 0 19872 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform 1 0 18584 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform 1 0 15088 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform 1 0 14168 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1649977179
transform 1 0 12696 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform 1 0 9384 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform 1 0 8280 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform 1 0 19780 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform 1 0 14628 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform 1 0 17204 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform 1 0 15732 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform 1 0 17020 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform 1 0 18308 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21068 0 1 19584
box -38 -48 1142 592
<< labels >>
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 0 nsew ground input
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 0 nsew ground input
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 0 nsew ground input
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 1 nsew power input
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 1 nsew power input
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 1 nsew power input
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 1 nsew power input
rlabel metal2 s 294 0 350 800 6 bottom_left_grid_pin_1_
port 2 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 ccff_tail
port 4 nsew signal tristate
rlabel metal3 s 22200 3816 23000 3936 6 chanx_right_in[0]
port 5 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[10]
port 6 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[11]
port 7 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[12]
port 8 nsew signal input
rlabel metal3 s 22200 9936 23000 10056 6 chanx_right_in[13]
port 9 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[14]
port 10 nsew signal input
rlabel metal3 s 22200 10888 23000 11008 6 chanx_right_in[15]
port 11 nsew signal input
rlabel metal3 s 22200 11296 23000 11416 6 chanx_right_in[16]
port 12 nsew signal input
rlabel metal3 s 22200 11840 23000 11960 6 chanx_right_in[17]
port 13 nsew signal input
rlabel metal3 s 22200 12248 23000 12368 6 chanx_right_in[18]
port 14 nsew signal input
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_in[19]
port 15 nsew signal input
rlabel metal3 s 22200 4360 23000 4480 6 chanx_right_in[1]
port 16 nsew signal input
rlabel metal3 s 22200 4768 23000 4888 6 chanx_right_in[2]
port 17 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[3]
port 18 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 chanx_right_in[4]
port 19 nsew signal input
rlabel metal3 s 22200 6128 23000 6248 6 chanx_right_in[5]
port 20 nsew signal input
rlabel metal3 s 22200 6672 23000 6792 6 chanx_right_in[6]
port 21 nsew signal input
rlabel metal3 s 22200 7080 23000 7200 6 chanx_right_in[7]
port 22 nsew signal input
rlabel metal3 s 22200 7624 23000 7744 6 chanx_right_in[8]
port 23 nsew signal input
rlabel metal3 s 22200 8032 23000 8152 6 chanx_right_in[9]
port 24 nsew signal input
rlabel metal3 s 22200 13200 23000 13320 6 chanx_right_out[0]
port 25 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[10]
port 26 nsew signal tristate
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[11]
port 27 nsew signal tristate
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[12]
port 28 nsew signal tristate
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[13]
port 29 nsew signal tristate
rlabel metal3 s 22200 19728 23000 19848 6 chanx_right_out[14]
port 30 nsew signal tristate
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[15]
port 31 nsew signal tristate
rlabel metal3 s 22200 20680 23000 20800 6 chanx_right_out[16]
port 32 nsew signal tristate
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[17]
port 33 nsew signal tristate
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[18]
port 34 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 chanx_right_out[19]
port 35 nsew signal tristate
rlabel metal3 s 22200 13744 23000 13864 6 chanx_right_out[1]
port 36 nsew signal tristate
rlabel metal3 s 22200 14152 23000 14272 6 chanx_right_out[2]
port 37 nsew signal tristate
rlabel metal3 s 22200 14560 23000 14680 6 chanx_right_out[3]
port 38 nsew signal tristate
rlabel metal3 s 22200 15104 23000 15224 6 chanx_right_out[4]
port 39 nsew signal tristate
rlabel metal3 s 22200 15512 23000 15632 6 chanx_right_out[5]
port 40 nsew signal tristate
rlabel metal3 s 22200 16056 23000 16176 6 chanx_right_out[6]
port 41 nsew signal tristate
rlabel metal3 s 22200 16464 23000 16584 6 chanx_right_out[7]
port 42 nsew signal tristate
rlabel metal3 s 22200 17008 23000 17128 6 chanx_right_out[8]
port 43 nsew signal tristate
rlabel metal3 s 22200 17416 23000 17536 6 chanx_right_out[9]
port 44 nsew signal tristate
rlabel metal2 s 846 0 902 800 6 chany_bottom_in[0]
port 45 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[10]
port 46 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 chany_bottom_in[11]
port 47 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 chany_bottom_in[12]
port 48 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[13]
port 49 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_in[14]
port 50 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[15]
port 51 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[16]
port 52 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[17]
port 53 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_in[18]
port 54 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[19]
port 55 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_in[1]
port 56 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 chany_bottom_in[2]
port 57 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 chany_bottom_in[3]
port 58 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 chany_bottom_in[4]
port 59 nsew signal input
rlabel metal2 s 3606 0 3662 800 6 chany_bottom_in[5]
port 60 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_in[6]
port 61 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 chany_bottom_in[7]
port 62 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 chany_bottom_in[8]
port 63 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 chany_bottom_in[9]
port 64 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 chany_bottom_out[0]
port 65 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[10]
port 66 nsew signal tristate
rlabel metal2 s 18234 0 18290 800 6 chany_bottom_out[11]
port 67 nsew signal tristate
rlabel metal2 s 18786 0 18842 800 6 chany_bottom_out[12]
port 68 nsew signal tristate
rlabel metal2 s 19338 0 19394 800 6 chany_bottom_out[13]
port 69 nsew signal tristate
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_out[14]
port 70 nsew signal tristate
rlabel metal2 s 20442 0 20498 800 6 chany_bottom_out[15]
port 71 nsew signal tristate
rlabel metal2 s 20994 0 21050 800 6 chany_bottom_out[16]
port 72 nsew signal tristate
rlabel metal2 s 21546 0 21602 800 6 chany_bottom_out[17]
port 73 nsew signal tristate
rlabel metal2 s 22098 0 22154 800 6 chany_bottom_out[18]
port 74 nsew signal tristate
rlabel metal2 s 22650 0 22706 800 6 chany_bottom_out[19]
port 75 nsew signal tristate
rlabel metal2 s 12622 0 12678 800 6 chany_bottom_out[1]
port 76 nsew signal tristate
rlabel metal2 s 13174 0 13230 800 6 chany_bottom_out[2]
port 77 nsew signal tristate
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_out[3]
port 78 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 chany_bottom_out[4]
port 79 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 chany_bottom_out[5]
port 80 nsew signal tristate
rlabel metal2 s 15382 0 15438 800 6 chany_bottom_out[6]
port 81 nsew signal tristate
rlabel metal2 s 15934 0 15990 800 6 chany_bottom_out[7]
port 82 nsew signal tristate
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_out[8]
port 83 nsew signal tristate
rlabel metal2 s 17038 0 17094 800 6 chany_bottom_out[9]
port 84 nsew signal tristate
rlabel metal2 s 846 22200 902 23000 6 chany_top_in[0]
port 85 nsew signal input
rlabel metal2 s 6458 22200 6514 23000 6 chany_top_in[10]
port 86 nsew signal input
rlabel metal2 s 7010 22200 7066 23000 6 chany_top_in[11]
port 87 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[12]
port 88 nsew signal input
rlabel metal2 s 8114 22200 8170 23000 6 chany_top_in[13]
port 89 nsew signal input
rlabel metal2 s 8666 22200 8722 23000 6 chany_top_in[14]
port 90 nsew signal input
rlabel metal2 s 9218 22200 9274 23000 6 chany_top_in[15]
port 91 nsew signal input
rlabel metal2 s 9770 22200 9826 23000 6 chany_top_in[16]
port 92 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[17]
port 93 nsew signal input
rlabel metal2 s 10874 22200 10930 23000 6 chany_top_in[18]
port 94 nsew signal input
rlabel metal2 s 11426 22200 11482 23000 6 chany_top_in[19]
port 95 nsew signal input
rlabel metal2 s 1398 22200 1454 23000 6 chany_top_in[1]
port 96 nsew signal input
rlabel metal2 s 1950 22200 2006 23000 6 chany_top_in[2]
port 97 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 chany_top_in[3]
port 98 nsew signal input
rlabel metal2 s 3054 22200 3110 23000 6 chany_top_in[4]
port 99 nsew signal input
rlabel metal2 s 3606 22200 3662 23000 6 chany_top_in[5]
port 100 nsew signal input
rlabel metal2 s 4158 22200 4214 23000 6 chany_top_in[6]
port 101 nsew signal input
rlabel metal2 s 4710 22200 4766 23000 6 chany_top_in[7]
port 102 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[8]
port 103 nsew signal input
rlabel metal2 s 5814 22200 5870 23000 6 chany_top_in[9]
port 104 nsew signal input
rlabel metal2 s 12070 22200 12126 23000 6 chany_top_out[0]
port 105 nsew signal tristate
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 106 nsew signal tristate
rlabel metal2 s 18234 22200 18290 23000 6 chany_top_out[11]
port 107 nsew signal tristate
rlabel metal2 s 18786 22200 18842 23000 6 chany_top_out[12]
port 108 nsew signal tristate
rlabel metal2 s 19338 22200 19394 23000 6 chany_top_out[13]
port 109 nsew signal tristate
rlabel metal2 s 19890 22200 19946 23000 6 chany_top_out[14]
port 110 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[15]
port 111 nsew signal tristate
rlabel metal2 s 20994 22200 21050 23000 6 chany_top_out[16]
port 112 nsew signal tristate
rlabel metal2 s 21546 22200 21602 23000 6 chany_top_out[17]
port 113 nsew signal tristate
rlabel metal2 s 22098 22200 22154 23000 6 chany_top_out[18]
port 114 nsew signal tristate
rlabel metal2 s 22650 22200 22706 23000 6 chany_top_out[19]
port 115 nsew signal tristate
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_out[1]
port 116 nsew signal tristate
rlabel metal2 s 13174 22200 13230 23000 6 chany_top_out[2]
port 117 nsew signal tristate
rlabel metal2 s 13726 22200 13782 23000 6 chany_top_out[3]
port 118 nsew signal tristate
rlabel metal2 s 14278 22200 14334 23000 6 chany_top_out[4]
port 119 nsew signal tristate
rlabel metal2 s 14830 22200 14886 23000 6 chany_top_out[5]
port 120 nsew signal tristate
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[6]
port 121 nsew signal tristate
rlabel metal2 s 15934 22200 15990 23000 6 chany_top_out[7]
port 122 nsew signal tristate
rlabel metal2 s 16486 22200 16542 23000 6 chany_top_out[8]
port 123 nsew signal tristate
rlabel metal2 s 17038 22200 17094 23000 6 chany_top_out[9]
port 124 nsew signal tristate
rlabel metal3 s 22200 22584 23000 22704 6 prog_clk_0_E_in
port 125 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_34_
port 126 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_35_
port 127 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_36_
port 128 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_37_
port 129 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_38_
port 130 nsew signal input
rlabel metal3 s 22200 2456 23000 2576 6 right_bottom_grid_pin_39_
port 131 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_40_
port 132 nsew signal input
rlabel metal3 s 22200 3408 23000 3528 6 right_bottom_grid_pin_41_
port 133 nsew signal input
rlabel metal2 s 294 22200 350 23000 6 top_left_grid_pin_1_
port 134 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
