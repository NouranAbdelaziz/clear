VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sb_2__2_
  CLASS BLOCK ;
  FOREIGN sb_2__2_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 115.000 BY 115.000 ;
  PIN SC_IN_BOT
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END SC_IN_BOT
  PIN SC_OUT_BOT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END SC_OUT_BOT
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 30.710 10.640 32.310 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.700 10.640 58.300 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.690 10.640 84.290 103.600 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 17.715 10.640 19.315 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.705 10.640 45.305 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.695 10.640 71.295 103.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 95.685 10.640 97.285 103.600 ;
    END
  END VPWR
  PIN bottom_left_grid_pin_42_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 4.000 ;
    END
  END bottom_left_grid_pin_42_
  PIN bottom_left_grid_pin_43_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END bottom_left_grid_pin_43_
  PIN bottom_left_grid_pin_44_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END bottom_left_grid_pin_44_
  PIN bottom_left_grid_pin_45_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END bottom_left_grid_pin_45_
  PIN bottom_left_grid_pin_46_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END bottom_left_grid_pin_46_
  PIN bottom_left_grid_pin_47_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 0.000 12.330 4.000 ;
    END
  END bottom_left_grid_pin_47_
  PIN bottom_left_grid_pin_48_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END bottom_left_grid_pin_48_
  PIN bottom_left_grid_pin_49_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END bottom_left_grid_pin_49_
  PIN bottom_right_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END bottom_right_grid_pin_1_
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 28.600 115.000 29.200 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 111.000 85.720 115.000 86.320 ;
    END
  END ccff_tail
  PIN chanx_left_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END chanx_left_in[0]
  PIN chanx_left_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END chanx_left_in[10]
  PIN chanx_left_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END chanx_left_in[11]
  PIN chanx_left_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.960 4.000 47.560 ;
    END
  END chanx_left_in[12]
  PIN chanx_left_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END chanx_left_in[13]
  PIN chanx_left_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END chanx_left_in[14]
  PIN chanx_left_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END chanx_left_in[15]
  PIN chanx_left_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 56.480 4.000 57.080 ;
    END
  END chanx_left_in[16]
  PIN chanx_left_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END chanx_left_in[17]
  PIN chanx_left_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END chanx_left_in[18]
  PIN chanx_left_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END chanx_left_in[19]
  PIN chanx_left_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END chanx_left_in[1]
  PIN chanx_left_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END chanx_left_in[2]
  PIN chanx_left_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END chanx_left_in[3]
  PIN chanx_left_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END chanx_left_in[4]
  PIN chanx_left_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END chanx_left_in[5]
  PIN chanx_left_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END chanx_left_in[6]
  PIN chanx_left_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END chanx_left_in[7]
  PIN chanx_left_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END chanx_left_in[8]
  PIN chanx_left_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END chanx_left_in[9]
  PIN chanx_left_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END chanx_left_out[0]
  PIN chanx_left_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END chanx_left_out[10]
  PIN chanx_left_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END chanx_left_out[11]
  PIN chanx_left_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END chanx_left_out[12]
  PIN chanx_left_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END chanx_left_out[13]
  PIN chanx_left_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END chanx_left_out[14]
  PIN chanx_left_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.360 4.000 101.960 ;
    END
  END chanx_left_out[15]
  PIN chanx_left_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 103.400 4.000 104.000 ;
    END
  END chanx_left_out[16]
  PIN chanx_left_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.120 4.000 106.720 ;
    END
  END chanx_left_out[17]
  PIN chanx_left_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.160 4.000 108.760 ;
    END
  END chanx_left_out[18]
  PIN chanx_left_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.880 4.000 111.480 ;
    END
  END chanx_left_out[19]
  PIN chanx_left_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END chanx_left_out[1]
  PIN chanx_left_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END chanx_left_out[2]
  PIN chanx_left_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.800 4.000 73.400 ;
    END
  END chanx_left_out[3]
  PIN chanx_left_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END chanx_left_out[4]
  PIN chanx_left_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END chanx_left_out[5]
  PIN chanx_left_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END chanx_left_out[6]
  PIN chanx_left_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 82.320 4.000 82.920 ;
    END
  END chanx_left_out[7]
  PIN chanx_left_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END chanx_left_out[8]
  PIN chanx_left_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END chanx_left_out[9]
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 4.000 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 0.000 60.630 4.000 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 0.000 27.510 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.330 0.000 89.610 4.000 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.370 0.000 100.650 4.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.510 0.000 104.790 4.000 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.390 0.000 71.670 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END chany_bottom_out[9]
  PIN left_bottom_grid_pin_34_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 0.720 4.000 1.320 ;
    END
  END left_bottom_grid_pin_34_
  PIN left_bottom_grid_pin_35_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END left_bottom_grid_pin_35_
  PIN left_bottom_grid_pin_36_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END left_bottom_grid_pin_36_
  PIN left_bottom_grid_pin_37_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END left_bottom_grid_pin_37_
  PIN left_bottom_grid_pin_38_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END left_bottom_grid_pin_38_
  PIN left_bottom_grid_pin_39_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END left_bottom_grid_pin_39_
  PIN left_bottom_grid_pin_40_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END left_bottom_grid_pin_40_
  PIN left_bottom_grid_pin_41_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END left_bottom_grid_pin_41_
  PIN left_top_grid_pin_1_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END left_top_grid_pin_1_
  PIN prog_clk_0_S_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 0.000 113.990 4.000 ;
    END
  END prog_clk_0_S_in
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 109.480 103.445 ;
      LAYER met1 ;
        RECT 0.990 6.500 114.010 104.000 ;
      LAYER met2 ;
        RECT 1.020 4.280 113.980 113.405 ;
        RECT 1.570 0.835 2.570 4.280 ;
        RECT 3.410 0.835 4.870 4.280 ;
        RECT 5.710 0.835 7.170 4.280 ;
        RECT 8.010 0.835 9.470 4.280 ;
        RECT 10.310 0.835 11.770 4.280 ;
        RECT 12.610 0.835 13.610 4.280 ;
        RECT 14.450 0.835 15.910 4.280 ;
        RECT 16.750 0.835 18.210 4.280 ;
        RECT 19.050 0.835 20.510 4.280 ;
        RECT 21.350 0.835 22.810 4.280 ;
        RECT 23.650 0.835 24.650 4.280 ;
        RECT 25.490 0.835 26.950 4.280 ;
        RECT 27.790 0.835 29.250 4.280 ;
        RECT 30.090 0.835 31.550 4.280 ;
        RECT 32.390 0.835 33.850 4.280 ;
        RECT 34.690 0.835 35.690 4.280 ;
        RECT 36.530 0.835 37.990 4.280 ;
        RECT 38.830 0.835 40.290 4.280 ;
        RECT 41.130 0.835 42.590 4.280 ;
        RECT 43.430 0.835 44.890 4.280 ;
        RECT 45.730 0.835 46.730 4.280 ;
        RECT 47.570 0.835 49.030 4.280 ;
        RECT 49.870 0.835 51.330 4.280 ;
        RECT 52.170 0.835 53.630 4.280 ;
        RECT 54.470 0.835 55.930 4.280 ;
        RECT 56.770 0.835 58.230 4.280 ;
        RECT 59.070 0.835 60.070 4.280 ;
        RECT 60.910 0.835 62.370 4.280 ;
        RECT 63.210 0.835 64.670 4.280 ;
        RECT 65.510 0.835 66.970 4.280 ;
        RECT 67.810 0.835 69.270 4.280 ;
        RECT 70.110 0.835 71.110 4.280 ;
        RECT 71.950 0.835 73.410 4.280 ;
        RECT 74.250 0.835 75.710 4.280 ;
        RECT 76.550 0.835 78.010 4.280 ;
        RECT 78.850 0.835 80.310 4.280 ;
        RECT 81.150 0.835 82.150 4.280 ;
        RECT 82.990 0.835 84.450 4.280 ;
        RECT 85.290 0.835 86.750 4.280 ;
        RECT 87.590 0.835 89.050 4.280 ;
        RECT 89.890 0.835 91.350 4.280 ;
        RECT 92.190 0.835 93.190 4.280 ;
        RECT 94.030 0.835 95.490 4.280 ;
        RECT 96.330 0.835 97.790 4.280 ;
        RECT 98.630 0.835 100.090 4.280 ;
        RECT 100.930 0.835 102.390 4.280 ;
        RECT 103.230 0.835 104.230 4.280 ;
        RECT 105.070 0.835 106.530 4.280 ;
        RECT 107.370 0.835 108.830 4.280 ;
        RECT 109.670 0.835 111.130 4.280 ;
        RECT 111.970 0.835 113.430 4.280 ;
      LAYER met3 ;
        RECT 4.400 112.520 111.000 113.385 ;
        RECT 3.990 111.880 111.000 112.520 ;
        RECT 4.400 110.480 111.000 111.880 ;
        RECT 3.990 109.160 111.000 110.480 ;
        RECT 4.400 107.760 111.000 109.160 ;
        RECT 3.990 107.120 111.000 107.760 ;
        RECT 4.400 105.720 111.000 107.120 ;
        RECT 3.990 104.400 111.000 105.720 ;
        RECT 4.400 103.000 111.000 104.400 ;
        RECT 3.990 102.360 111.000 103.000 ;
        RECT 4.400 100.960 111.000 102.360 ;
        RECT 3.990 99.640 111.000 100.960 ;
        RECT 4.400 98.240 111.000 99.640 ;
        RECT 3.990 97.600 111.000 98.240 ;
        RECT 4.400 96.200 111.000 97.600 ;
        RECT 3.990 94.880 111.000 96.200 ;
        RECT 4.400 93.480 111.000 94.880 ;
        RECT 3.990 92.840 111.000 93.480 ;
        RECT 4.400 91.440 111.000 92.840 ;
        RECT 3.990 90.800 111.000 91.440 ;
        RECT 4.400 89.400 111.000 90.800 ;
        RECT 3.990 88.080 111.000 89.400 ;
        RECT 4.400 86.720 111.000 88.080 ;
        RECT 4.400 86.680 110.600 86.720 ;
        RECT 3.990 86.040 110.600 86.680 ;
        RECT 4.400 85.320 110.600 86.040 ;
        RECT 4.400 84.640 111.000 85.320 ;
        RECT 3.990 83.320 111.000 84.640 ;
        RECT 4.400 81.920 111.000 83.320 ;
        RECT 3.990 81.280 111.000 81.920 ;
        RECT 4.400 79.880 111.000 81.280 ;
        RECT 3.990 78.560 111.000 79.880 ;
        RECT 4.400 77.160 111.000 78.560 ;
        RECT 3.990 76.520 111.000 77.160 ;
        RECT 4.400 75.120 111.000 76.520 ;
        RECT 3.990 73.800 111.000 75.120 ;
        RECT 4.400 72.400 111.000 73.800 ;
        RECT 3.990 71.760 111.000 72.400 ;
        RECT 4.400 70.360 111.000 71.760 ;
        RECT 3.990 69.720 111.000 70.360 ;
        RECT 4.400 68.320 111.000 69.720 ;
        RECT 3.990 67.000 111.000 68.320 ;
        RECT 4.400 65.600 111.000 67.000 ;
        RECT 3.990 64.960 111.000 65.600 ;
        RECT 4.400 63.560 111.000 64.960 ;
        RECT 3.990 62.240 111.000 63.560 ;
        RECT 4.400 60.840 111.000 62.240 ;
        RECT 3.990 60.200 111.000 60.840 ;
        RECT 4.400 58.800 111.000 60.200 ;
        RECT 3.990 57.480 111.000 58.800 ;
        RECT 4.400 56.080 111.000 57.480 ;
        RECT 3.990 55.440 111.000 56.080 ;
        RECT 4.400 54.040 111.000 55.440 ;
        RECT 3.990 52.720 111.000 54.040 ;
        RECT 4.400 51.320 111.000 52.720 ;
        RECT 3.990 50.680 111.000 51.320 ;
        RECT 4.400 49.280 111.000 50.680 ;
        RECT 3.990 47.960 111.000 49.280 ;
        RECT 4.400 46.560 111.000 47.960 ;
        RECT 3.990 45.920 111.000 46.560 ;
        RECT 4.400 44.520 111.000 45.920 ;
        RECT 3.990 43.880 111.000 44.520 ;
        RECT 4.400 42.480 111.000 43.880 ;
        RECT 3.990 41.160 111.000 42.480 ;
        RECT 4.400 39.760 111.000 41.160 ;
        RECT 3.990 39.120 111.000 39.760 ;
        RECT 4.400 37.720 111.000 39.120 ;
        RECT 3.990 36.400 111.000 37.720 ;
        RECT 4.400 35.000 111.000 36.400 ;
        RECT 3.990 34.360 111.000 35.000 ;
        RECT 4.400 32.960 111.000 34.360 ;
        RECT 3.990 31.640 111.000 32.960 ;
        RECT 4.400 30.240 111.000 31.640 ;
        RECT 3.990 29.600 111.000 30.240 ;
        RECT 4.400 28.200 110.600 29.600 ;
        RECT 3.990 26.880 111.000 28.200 ;
        RECT 4.400 25.480 111.000 26.880 ;
        RECT 3.990 24.840 111.000 25.480 ;
        RECT 4.400 23.440 111.000 24.840 ;
        RECT 3.990 22.800 111.000 23.440 ;
        RECT 4.400 21.400 111.000 22.800 ;
        RECT 3.990 20.080 111.000 21.400 ;
        RECT 4.400 18.680 111.000 20.080 ;
        RECT 3.990 18.040 111.000 18.680 ;
        RECT 4.400 16.640 111.000 18.040 ;
        RECT 3.990 15.320 111.000 16.640 ;
        RECT 4.400 13.920 111.000 15.320 ;
        RECT 3.990 13.280 111.000 13.920 ;
        RECT 4.400 11.880 111.000 13.280 ;
        RECT 3.990 10.560 111.000 11.880 ;
        RECT 4.400 9.160 111.000 10.560 ;
        RECT 3.990 8.520 111.000 9.160 ;
        RECT 4.400 7.120 111.000 8.520 ;
        RECT 3.990 5.800 111.000 7.120 ;
        RECT 4.400 4.400 111.000 5.800 ;
        RECT 3.990 3.760 111.000 4.400 ;
        RECT 4.400 2.360 111.000 3.760 ;
        RECT 3.990 1.720 111.000 2.360 ;
        RECT 4.400 0.855 111.000 1.720 ;
      LAYER met4 ;
        RECT 8.575 10.240 17.315 88.225 ;
        RECT 19.715 10.240 30.310 88.225 ;
        RECT 32.710 10.240 43.305 88.225 ;
        RECT 45.705 10.240 56.300 88.225 ;
        RECT 58.700 10.240 69.295 88.225 ;
        RECT 71.695 10.240 82.290 88.225 ;
        RECT 84.690 10.240 95.285 88.225 ;
        RECT 97.685 10.240 101.825 88.225 ;
        RECT 8.575 4.935 101.825 10.240 ;
      LAYER met5 ;
        RECT 19.900 17.900 73.020 19.500 ;
  END
END sb_2__2_
END LIBRARY

