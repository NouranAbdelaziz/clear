magic
tech sky130A
magscale 1 2
timestamp 1650891705
<< viali >>
rect 2145 17221 2179 17255
rect 2421 17153 2455 17187
rect 5365 16201 5399 16235
rect 4905 16133 4939 16167
rect 5181 16065 5215 16099
rect 3709 15861 3743 15895
rect 3433 15657 3467 15691
rect 4445 15657 4479 15691
rect 4997 15657 5031 15691
rect 7021 15657 7055 15691
rect 7665 15657 7699 15691
rect 5181 15589 5215 15623
rect 3985 15521 4019 15555
rect 7389 15521 7423 15555
rect 3617 15453 3651 15487
rect 4261 15453 4295 15487
rect 4629 15453 4663 15487
rect 4813 15453 4847 15487
rect 6469 15453 6503 15487
rect 7297 15385 7331 15419
rect 5549 15317 5583 15351
rect 6285 15317 6319 15351
rect 7757 15317 7791 15351
rect 8033 15317 8067 15351
rect 3065 15113 3099 15147
rect 3249 15113 3283 15147
rect 3617 15113 3651 15147
rect 4077 15113 4111 15147
rect 4445 15113 4479 15147
rect 5089 15113 5123 15147
rect 6009 15113 6043 15147
rect 6377 15113 6411 15147
rect 7849 15113 7883 15147
rect 6929 15045 6963 15079
rect 3433 14977 3467 15011
rect 3801 14977 3835 15011
rect 4261 14977 4295 15011
rect 4629 14977 4663 15011
rect 5181 14977 5215 15011
rect 5457 14977 5491 15011
rect 6193 14977 6227 15011
rect 7665 14977 7699 15011
rect 8033 14977 8067 15011
rect 2881 14909 2915 14943
rect 4813 14909 4847 14943
rect 5825 14909 5859 14943
rect 7021 14909 7055 14943
rect 7113 14909 7147 14943
rect 5641 14841 5675 14875
rect 7481 14841 7515 14875
rect 2605 14773 2639 14807
rect 6561 14773 6595 14807
rect 8217 14773 8251 14807
rect 8493 14773 8527 14807
rect 8677 14773 8711 14807
rect 8861 14773 8895 14807
rect 5273 14569 5307 14603
rect 7205 14569 7239 14603
rect 8125 14569 8159 14603
rect 8493 14569 8527 14603
rect 9781 14569 9815 14603
rect 2605 14501 2639 14535
rect 3341 14501 3375 14535
rect 3617 14501 3651 14535
rect 4905 14501 4939 14535
rect 6377 14501 6411 14535
rect 9045 14501 9079 14535
rect 9413 14501 9447 14535
rect 1961 14433 1995 14467
rect 2237 14433 2271 14467
rect 2881 14433 2915 14467
rect 3065 14433 3099 14467
rect 6101 14433 6135 14467
rect 6929 14433 6963 14467
rect 7757 14433 7791 14467
rect 9137 14433 9171 14467
rect 2513 14365 2547 14399
rect 3801 14365 3835 14399
rect 4537 14365 4571 14399
rect 5089 14365 5123 14399
rect 5457 14365 5491 14399
rect 5917 14365 5951 14399
rect 6837 14365 6871 14399
rect 7665 14365 7699 14399
rect 8309 14365 8343 14399
rect 8677 14365 8711 14399
rect 9597 14365 9631 14399
rect 3157 14297 3191 14331
rect 3985 14297 4019 14331
rect 6745 14297 6779 14331
rect 7573 14297 7607 14331
rect 1685 14229 1719 14263
rect 4353 14229 4387 14263
rect 4721 14229 4755 14263
rect 5549 14229 5583 14263
rect 6009 14229 6043 14263
rect 1501 14025 1535 14059
rect 3801 14025 3835 14059
rect 5917 14025 5951 14059
rect 8861 14025 8895 14059
rect 9229 14025 9263 14059
rect 10057 14025 10091 14059
rect 1685 13957 1719 13991
rect 2789 13957 2823 13991
rect 3617 13957 3651 13991
rect 4169 13957 4203 13991
rect 4261 13957 4295 13991
rect 6653 13957 6687 13991
rect 8493 13957 8527 13991
rect 9873 13957 9907 13991
rect 1869 13889 1903 13923
rect 2421 13889 2455 13923
rect 3065 13889 3099 13923
rect 3249 13889 3283 13923
rect 4997 13889 5031 13923
rect 5089 13889 5123 13923
rect 5825 13889 5859 13923
rect 9045 13889 9079 13923
rect 9413 13889 9447 13923
rect 9597 13889 9631 13923
rect 2145 13821 2179 13855
rect 3433 13821 3467 13855
rect 4353 13821 4387 13855
rect 5273 13821 5307 13855
rect 6101 13821 6135 13855
rect 8217 13821 8251 13855
rect 9689 13821 9723 13855
rect 4629 13685 4663 13719
rect 5457 13685 5491 13719
rect 6469 13685 6503 13719
rect 2697 13481 2731 13515
rect 3801 13481 3835 13515
rect 4813 13481 4847 13515
rect 6469 13481 6503 13515
rect 8585 13481 8619 13515
rect 9045 13481 9079 13515
rect 9505 13481 9539 13515
rect 10517 13481 10551 13515
rect 10701 13481 10735 13515
rect 10241 13413 10275 13447
rect 1685 13345 1719 13379
rect 3525 13345 3559 13379
rect 4445 13345 4479 13379
rect 5457 13345 5491 13379
rect 5917 13345 5951 13379
rect 6745 13345 6779 13379
rect 7573 13345 7607 13379
rect 1961 13277 1995 13311
rect 2513 13277 2547 13311
rect 3341 13277 3375 13311
rect 6101 13277 6135 13311
rect 6929 13277 6963 13311
rect 7757 13277 7791 13311
rect 8769 13277 8803 13311
rect 9229 13277 9263 13311
rect 9689 13277 9723 13311
rect 10057 13277 10091 13311
rect 10885 13277 10919 13311
rect 2237 13209 2271 13243
rect 4261 13209 4295 13243
rect 5365 13209 5399 13243
rect 6837 13209 6871 13243
rect 8217 13209 8251 13243
rect 10425 13209 10459 13243
rect 2881 13141 2915 13175
rect 3249 13141 3283 13175
rect 4169 13141 4203 13175
rect 4905 13141 4939 13175
rect 5273 13141 5307 13175
rect 6009 13141 6043 13175
rect 7297 13141 7331 13175
rect 7665 13141 7699 13175
rect 8125 13141 8159 13175
rect 9781 13141 9815 13175
rect 1685 12937 1719 12971
rect 2145 12937 2179 12971
rect 2329 12937 2363 12971
rect 3065 12937 3099 12971
rect 4629 12937 4663 12971
rect 5733 12937 5767 12971
rect 6561 12937 6595 12971
rect 8493 12937 8527 12971
rect 9321 12937 9355 12971
rect 9689 12937 9723 12971
rect 7297 12869 7331 12903
rect 9781 12869 9815 12903
rect 10609 12869 10643 12903
rect 10885 12869 10919 12903
rect 1777 12801 1811 12835
rect 4353 12801 4387 12835
rect 4997 12801 5031 12835
rect 5089 12801 5123 12835
rect 5825 12801 5859 12835
rect 6745 12801 6779 12835
rect 7205 12801 7239 12835
rect 8033 12801 8067 12835
rect 8861 12801 8895 12835
rect 10793 12801 10827 12835
rect 1593 12733 1627 12767
rect 5273 12733 5307 12767
rect 5641 12733 5675 12767
rect 7481 12733 7515 12767
rect 7757 12733 7791 12767
rect 7941 12733 7975 12767
rect 8953 12733 8987 12767
rect 9045 12733 9079 12767
rect 9873 12733 9907 12767
rect 11069 12733 11103 12767
rect 6193 12665 6227 12699
rect 8401 12665 8435 12699
rect 10149 12665 10183 12699
rect 11345 12665 11379 12699
rect 11621 12665 11655 12699
rect 11805 12665 11839 12699
rect 11989 12665 12023 12699
rect 2513 12597 2547 12631
rect 4537 12597 4571 12631
rect 6837 12597 6871 12631
rect 10333 12597 10367 12631
rect 2881 12393 2915 12427
rect 5273 12393 5307 12427
rect 8585 12393 8619 12427
rect 9781 12393 9815 12427
rect 11437 12393 11471 12427
rect 11989 12393 12023 12427
rect 12909 12393 12943 12427
rect 14289 12393 14323 12427
rect 5549 12325 5583 12359
rect 10793 12325 10827 12359
rect 11713 12325 11747 12359
rect 12265 12325 12299 12359
rect 1685 12257 1719 12291
rect 2237 12257 2271 12291
rect 2329 12257 2363 12291
rect 3341 12257 3375 12291
rect 3433 12257 3467 12291
rect 9505 12257 9539 12291
rect 10333 12257 10367 12291
rect 11253 12257 11287 12291
rect 12541 12257 12575 12291
rect 14473 12257 14507 12291
rect 1961 12189 1995 12223
rect 2421 12189 2455 12223
rect 3801 12189 3835 12223
rect 4629 12189 4663 12223
rect 5457 12189 5491 12223
rect 6662 12189 6696 12223
rect 6929 12189 6963 12223
rect 7021 12189 7055 12223
rect 7277 12189 7311 12223
rect 8769 12189 8803 12223
rect 9321 12189 9355 12223
rect 9413 12189 9447 12223
rect 10241 12189 10275 12223
rect 10609 12189 10643 12223
rect 10149 12121 10183 12155
rect 11621 12121 11655 12155
rect 14933 12121 14967 12155
rect 2789 12053 2823 12087
rect 3249 12053 3283 12087
rect 5089 12053 5123 12087
rect 8401 12053 8435 12087
rect 8953 12053 8987 12087
rect 10977 12053 11011 12087
rect 12081 12053 12115 12087
rect 12633 12053 12667 12087
rect 13461 12053 13495 12087
rect 14105 12053 14139 12087
rect 15301 12053 15335 12087
rect 1777 11849 1811 11883
rect 2237 11849 2271 11883
rect 2697 11849 2731 11883
rect 3065 11849 3099 11883
rect 3893 11849 3927 11883
rect 4721 11849 4755 11883
rect 9045 11849 9079 11883
rect 11529 11849 11563 11883
rect 12541 11849 12575 11883
rect 14565 11849 14599 11883
rect 14841 11849 14875 11883
rect 3433 11781 3467 11815
rect 3525 11781 3559 11815
rect 8309 11781 8343 11815
rect 10701 11781 10735 11815
rect 10793 11781 10827 11815
rect 11897 11781 11931 11815
rect 13185 11781 13219 11815
rect 15393 11781 15427 11815
rect 1869 11713 1903 11747
rect 4261 11713 4295 11747
rect 4353 11713 4387 11747
rect 5069 11713 5103 11747
rect 6633 11713 6667 11747
rect 8217 11713 8251 11747
rect 8953 11713 8987 11747
rect 9873 11713 9907 11747
rect 11161 11713 11195 11747
rect 12081 11713 12115 11747
rect 14749 11713 14783 11747
rect 1593 11645 1627 11679
rect 2513 11645 2547 11679
rect 2605 11645 2639 11679
rect 3341 11645 3375 11679
rect 4169 11645 4203 11679
rect 4813 11645 4847 11679
rect 6377 11645 6411 11679
rect 8401 11645 8435 11679
rect 8769 11645 8803 11679
rect 9965 11645 9999 11679
rect 10149 11645 10183 11679
rect 10885 11645 10919 11679
rect 11805 11645 11839 11679
rect 12265 11645 12299 11679
rect 12633 11645 12667 11679
rect 13829 11645 13863 11679
rect 15025 11645 15059 11679
rect 6193 11577 6227 11611
rect 7849 11577 7883 11611
rect 9505 11577 9539 11611
rect 14013 11577 14047 11611
rect 14381 11577 14415 11611
rect 7757 11509 7791 11543
rect 9413 11509 9447 11543
rect 10333 11509 10367 11543
rect 12817 11509 12851 11543
rect 13093 11509 13127 11543
rect 13369 11509 13403 11543
rect 13645 11509 13679 11543
rect 14197 11509 14231 11543
rect 15301 11509 15335 11543
rect 15577 11509 15611 11543
rect 4629 11305 4663 11339
rect 7665 11305 7699 11339
rect 8953 11305 8987 11339
rect 10609 11305 10643 11339
rect 12449 11305 12483 11339
rect 12725 11305 12759 11339
rect 12909 11305 12943 11339
rect 13185 11305 13219 11339
rect 14289 11305 14323 11339
rect 14565 11305 14599 11339
rect 15485 11305 15519 11339
rect 2789 11237 2823 11271
rect 6193 11237 6227 11271
rect 9781 11237 9815 11271
rect 14933 11237 14967 11271
rect 1685 11169 1719 11203
rect 2237 11169 2271 11203
rect 3341 11169 3375 11203
rect 3525 11169 3559 11203
rect 4077 11169 4111 11203
rect 4169 11169 4203 11203
rect 8217 11169 8251 11203
rect 8677 11169 8711 11203
rect 9413 11169 9447 11203
rect 9505 11169 9539 11203
rect 10333 11169 10367 11203
rect 11161 11169 11195 11203
rect 11989 11169 12023 11203
rect 13737 11169 13771 11203
rect 1961 11101 1995 11135
rect 2421 11101 2455 11135
rect 6101 11101 6135 11135
rect 7573 11101 7607 11135
rect 9321 11101 9355 11135
rect 10149 11101 10183 11135
rect 10241 11101 10275 11135
rect 11897 11101 11931 11135
rect 13369 11101 13403 11135
rect 14197 11101 14231 11135
rect 2329 11033 2363 11067
rect 3249 11033 3283 11067
rect 5834 11033 5868 11067
rect 7328 11033 7362 11067
rect 10977 11033 11011 11067
rect 11069 11033 11103 11067
rect 12265 11033 12299 11067
rect 15025 11033 15059 11067
rect 15577 11033 15611 11067
rect 2881 10965 2915 10999
rect 4261 10965 4295 10999
rect 4721 10965 4755 10999
rect 8033 10965 8067 10999
rect 8125 10965 8159 10999
rect 11437 10965 11471 10999
rect 11805 10965 11839 10999
rect 13001 10965 13035 10999
rect 13553 10965 13587 10999
rect 14749 10965 14783 10999
rect 15209 10965 15243 10999
rect 1593 10761 1627 10795
rect 1961 10761 1995 10795
rect 2421 10761 2455 10795
rect 9689 10761 9723 10795
rect 10885 10761 10919 10795
rect 10977 10761 11011 10795
rect 11529 10761 11563 10795
rect 11989 10761 12023 10795
rect 12725 10761 12759 10795
rect 14013 10761 14047 10795
rect 14105 10761 14139 10795
rect 14289 10761 14323 10795
rect 15301 10761 15335 10795
rect 15485 10761 15519 10795
rect 2789 10693 2823 10727
rect 5948 10693 5982 10727
rect 7849 10693 7883 10727
rect 13737 10693 13771 10727
rect 14841 10693 14875 10727
rect 2053 10625 2087 10659
rect 2881 10625 2915 10659
rect 3341 10625 3375 10659
rect 3608 10625 3642 10659
rect 6644 10625 6678 10659
rect 10057 10625 10091 10659
rect 11897 10625 11931 10659
rect 13174 10625 13208 10659
rect 14473 10625 14507 10659
rect 1869 10557 1903 10591
rect 2697 10557 2731 10591
rect 6193 10557 6227 10591
rect 6377 10557 6411 10591
rect 9505 10557 9539 10591
rect 10149 10557 10183 10591
rect 10241 10557 10275 10591
rect 11069 10557 11103 10591
rect 12081 10557 12115 10591
rect 12817 10557 12851 10591
rect 13001 10557 13035 10591
rect 13369 10557 13403 10591
rect 15025 10557 15059 10591
rect 3249 10489 3283 10523
rect 15577 10489 15611 10523
rect 4721 10421 4755 10455
rect 4813 10421 4847 10455
rect 7757 10421 7791 10455
rect 10517 10421 10551 10455
rect 12357 10421 12391 10455
rect 14749 10421 14783 10455
rect 10333 10217 10367 10251
rect 11253 10217 11287 10251
rect 14289 10217 14323 10251
rect 15669 10217 15703 10251
rect 2145 10149 2179 10183
rect 3617 10149 3651 10183
rect 7389 10149 7423 10183
rect 10425 10149 10459 10183
rect 14473 10149 14507 10183
rect 15209 10149 15243 10183
rect 1593 10081 1627 10115
rect 1685 10081 1719 10115
rect 5181 10081 5215 10115
rect 7297 10081 7331 10115
rect 8769 10081 8803 10115
rect 10885 10081 10919 10115
rect 10977 10081 11011 10115
rect 11897 10081 11931 10115
rect 12633 10081 12667 10115
rect 13461 10081 13495 10115
rect 15025 10081 15059 10115
rect 2237 10013 2271 10047
rect 8953 10013 8987 10047
rect 12449 10013 12483 10047
rect 13277 10013 13311 10047
rect 13737 10013 13771 10047
rect 14657 10013 14691 10047
rect 2504 9945 2538 9979
rect 4914 9945 4948 9979
rect 5273 9945 5307 9979
rect 8502 9945 8536 9979
rect 9198 9945 9232 9979
rect 11621 9945 11655 9979
rect 13369 9945 13403 9979
rect 15393 9945 15427 9979
rect 1777 9877 1811 9911
rect 3801 9877 3835 9911
rect 6561 9877 6595 9911
rect 10793 9877 10827 9911
rect 11713 9877 11747 9911
rect 12081 9877 12115 9911
rect 12541 9877 12575 9911
rect 12909 9877 12943 9911
rect 14105 9877 14139 9911
rect 14841 9877 14875 9911
rect 4721 9673 4755 9707
rect 6193 9673 6227 9707
rect 7849 9673 7883 9707
rect 12725 9673 12759 9707
rect 14381 9673 14415 9707
rect 14841 9673 14875 9707
rect 15301 9673 15335 9707
rect 1777 9605 1811 9639
rect 9588 9605 9622 9639
rect 11069 9605 11103 9639
rect 11897 9605 11931 9639
rect 13553 9605 13587 9639
rect 1501 9537 1535 9571
rect 2982 9537 3016 9571
rect 3249 9537 3283 9571
rect 3341 9537 3375 9571
rect 3597 9537 3631 9571
rect 4813 9537 4847 9571
rect 5069 9537 5103 9571
rect 6377 9537 6411 9571
rect 6644 9537 6678 9571
rect 8962 9537 8996 9571
rect 9229 9537 9263 9571
rect 9321 9537 9355 9571
rect 10793 9537 10827 9571
rect 12817 9537 12851 9571
rect 14473 9537 14507 9571
rect 15209 9537 15243 9571
rect 11989 9469 12023 9503
rect 12081 9469 12115 9503
rect 12909 9469 12943 9503
rect 13645 9469 13679 9503
rect 13829 9469 13863 9503
rect 14565 9469 14599 9503
rect 15393 9469 15427 9503
rect 1869 9401 1903 9435
rect 7757 9401 7791 9435
rect 12357 9401 12391 9435
rect 10701 9333 10735 9367
rect 11529 9333 11563 9367
rect 13185 9333 13219 9367
rect 14013 9333 14047 9367
rect 8953 9129 8987 9163
rect 10425 9129 10459 9163
rect 11253 9129 11287 9163
rect 12081 9129 12115 9163
rect 14933 9129 14967 9163
rect 2145 9061 2179 9095
rect 3617 9061 3651 9095
rect 5917 9061 5951 9095
rect 12909 9061 12943 9095
rect 14105 9061 14139 9095
rect 1593 8993 1627 9027
rect 1685 8993 1719 9027
rect 2237 8993 2271 9027
rect 3985 8993 4019 9027
rect 10977 8993 11011 9027
rect 11897 8993 11931 9027
rect 12725 8993 12759 9027
rect 13369 8993 13403 9027
rect 13553 8993 13587 9027
rect 14565 8993 14599 9027
rect 14657 8993 14691 9027
rect 15393 8993 15427 9027
rect 15485 8993 15519 9027
rect 2493 8925 2527 8959
rect 3801 8925 3835 8959
rect 5558 8925 5592 8959
rect 5825 8925 5859 8959
rect 7297 8925 7331 8959
rect 7389 8925 7423 8959
rect 10333 8925 10367 8959
rect 10885 8925 10919 8959
rect 11621 8925 11655 8959
rect 12449 8925 12483 8959
rect 7030 8857 7064 8891
rect 7634 8857 7668 8891
rect 10088 8857 10122 8891
rect 11713 8857 11747 8891
rect 12541 8857 12575 8891
rect 13277 8857 13311 8891
rect 14473 8857 14507 8891
rect 1777 8789 1811 8823
rect 4445 8789 4479 8823
rect 8769 8789 8803 8823
rect 10793 8789 10827 8823
rect 13737 8789 13771 8823
rect 15301 8789 15335 8823
rect 1869 8585 1903 8619
rect 4813 8585 4847 8619
rect 7757 8585 7791 8619
rect 9137 8585 9171 8619
rect 11529 8585 11563 8619
rect 11989 8585 12023 8619
rect 12357 8585 12391 8619
rect 13185 8585 13219 8619
rect 13553 8585 13587 8619
rect 15209 8585 15243 8619
rect 15301 8585 15335 8619
rect 3004 8517 3038 8551
rect 6622 8517 6656 8551
rect 11161 8517 11195 8551
rect 13645 8517 13679 8551
rect 1777 8449 1811 8483
rect 3249 8449 3283 8483
rect 4454 8449 4488 8483
rect 4721 8449 4755 8483
rect 5926 8449 5960 8483
rect 7849 8449 7883 8483
rect 9689 8449 9723 8483
rect 9945 8449 9979 8483
rect 11897 8449 11931 8483
rect 12725 8449 12759 8483
rect 12817 8449 12851 8483
rect 14381 8449 14415 8483
rect 6193 8381 6227 8415
rect 6377 8381 6411 8415
rect 12173 8381 12207 8415
rect 12909 8381 12943 8415
rect 13829 8381 13863 8415
rect 14473 8381 14507 8415
rect 14657 8381 14691 8415
rect 15485 8381 15519 8415
rect 1593 8313 1627 8347
rect 3341 8313 3375 8347
rect 11069 8245 11103 8279
rect 14013 8245 14047 8279
rect 14841 8245 14875 8279
rect 1869 8041 1903 8075
rect 4813 8041 4847 8075
rect 8953 8041 8987 8075
rect 4445 7973 4479 8007
rect 14105 7973 14139 8007
rect 8493 7905 8527 7939
rect 12357 7905 12391 7939
rect 12449 7905 12483 7939
rect 12909 7905 12943 7939
rect 13829 7905 13863 7939
rect 14749 7905 14783 7939
rect 15485 7905 15519 7939
rect 3617 7837 3651 7871
rect 3985 7837 4019 7871
rect 4261 7837 4295 7871
rect 6377 7837 6411 7871
rect 7941 7837 7975 7871
rect 8769 7837 8803 7871
rect 10333 7837 10367 7871
rect 10425 7837 10459 7871
rect 3157 7769 3191 7803
rect 6285 7769 6319 7803
rect 10066 7769 10100 7803
rect 10692 7769 10726 7803
rect 12265 7769 12299 7803
rect 14565 7769 14599 7803
rect 15393 7769 15427 7803
rect 3433 7701 3467 7735
rect 11805 7701 11839 7735
rect 11897 7701 11931 7735
rect 13001 7701 13035 7735
rect 13093 7701 13127 7735
rect 13461 7701 13495 7735
rect 13553 7701 13587 7735
rect 14473 7701 14507 7735
rect 14933 7701 14967 7735
rect 15301 7701 15335 7735
rect 3341 7497 3375 7531
rect 4813 7497 4847 7531
rect 11161 7497 11195 7531
rect 12357 7497 12391 7531
rect 13553 7497 13587 7531
rect 14381 7497 14415 7531
rect 5948 7429 5982 7463
rect 11897 7429 11931 7463
rect 12817 7429 12851 7463
rect 15209 7429 15243 7463
rect 1501 7361 1535 7395
rect 1869 7361 1903 7395
rect 2136 7361 2170 7395
rect 4465 7361 4499 7395
rect 4721 7361 4755 7395
rect 7490 7361 7524 7395
rect 7849 7361 7883 7395
rect 9597 7361 9631 7395
rect 9689 7361 9723 7395
rect 9956 7361 9990 7395
rect 11989 7361 12023 7395
rect 12725 7361 12759 7395
rect 13461 7361 13495 7395
rect 14473 7361 14507 7395
rect 6193 7293 6227 7327
rect 7757 7293 7791 7327
rect 12173 7293 12207 7327
rect 12909 7293 12943 7327
rect 13277 7293 13311 7327
rect 14657 7293 14691 7327
rect 15301 7293 15335 7327
rect 15393 7293 15427 7327
rect 3249 7225 3283 7259
rect 11529 7225 11563 7259
rect 14013 7225 14047 7259
rect 1685 7157 1719 7191
rect 6377 7157 6411 7191
rect 11069 7157 11103 7191
rect 13921 7157 13955 7191
rect 14841 7157 14875 7191
rect 12081 6953 12115 6987
rect 5917 6885 5951 6919
rect 11253 6885 11287 6919
rect 1593 6817 1627 6851
rect 3985 6817 4019 6851
rect 5825 6817 5859 6851
rect 8769 6817 8803 6851
rect 10609 6817 10643 6851
rect 11897 6817 11931 6851
rect 12633 6817 12667 6851
rect 13369 6817 13403 6851
rect 13461 6817 13495 6851
rect 13921 6817 13955 6851
rect 14657 6817 14691 6851
rect 15393 6817 15427 6851
rect 15577 6817 15611 6851
rect 1777 6749 1811 6783
rect 3617 6749 3651 6783
rect 4261 6749 4295 6783
rect 7297 6749 7331 6783
rect 10333 6749 10367 6783
rect 11621 6749 11655 6783
rect 12449 6749 12483 6783
rect 13277 6749 13311 6783
rect 3372 6681 3406 6715
rect 5558 6681 5592 6715
rect 7030 6681 7064 6715
rect 8524 6681 8558 6715
rect 10088 6681 10122 6715
rect 10793 6681 10827 6715
rect 12541 6681 12575 6715
rect 1685 6613 1719 6647
rect 2145 6613 2179 6647
rect 2237 6613 2271 6647
rect 4445 6613 4479 6647
rect 7389 6613 7423 6647
rect 8953 6613 8987 6647
rect 10701 6613 10735 6647
rect 11161 6613 11195 6647
rect 11713 6613 11747 6647
rect 12909 6613 12943 6647
rect 14105 6613 14139 6647
rect 14473 6613 14507 6647
rect 14565 6613 14599 6647
rect 14933 6613 14967 6647
rect 15301 6613 15335 6647
rect 1593 6409 1627 6443
rect 4721 6409 4755 6443
rect 7757 6409 7791 6443
rect 12633 6409 12667 6443
rect 12725 6409 12759 6443
rect 13093 6409 13127 6443
rect 13553 6409 13587 6443
rect 14013 6409 14047 6443
rect 9566 6341 9600 6375
rect 13645 6341 13679 6375
rect 1777 6273 1811 6307
rect 1869 6273 1903 6307
rect 2136 6273 2170 6307
rect 3341 6273 3375 6307
rect 3608 6273 3642 6307
rect 4813 6273 4847 6307
rect 5080 6273 5114 6307
rect 6377 6273 6411 6307
rect 6644 6273 6678 6307
rect 7849 6273 7883 6307
rect 8116 6273 8150 6307
rect 11253 6273 11287 6307
rect 11897 6273 11931 6307
rect 11989 6273 12023 6307
rect 14381 6273 14415 6307
rect 9321 6205 9355 6239
rect 10977 6205 11011 6239
rect 12081 6205 12115 6239
rect 12541 6205 12575 6239
rect 13829 6205 13863 6239
rect 14473 6205 14507 6239
rect 14565 6205 14599 6239
rect 14841 6205 14875 6239
rect 9229 6137 9263 6171
rect 11529 6137 11563 6171
rect 15301 6137 15335 6171
rect 15577 6137 15611 6171
rect 3249 6069 3283 6103
rect 6193 6069 6227 6103
rect 10701 6069 10735 6103
rect 13185 6069 13219 6103
rect 15209 6069 15243 6103
rect 3433 5865 3467 5899
rect 5181 5865 5215 5899
rect 10517 5865 10551 5899
rect 14749 5865 14783 5899
rect 15485 5865 15519 5899
rect 8493 5797 8527 5831
rect 14841 5797 14875 5831
rect 15301 5797 15335 5831
rect 9045 5729 9079 5763
rect 9229 5729 9263 5763
rect 9873 5729 9907 5763
rect 10701 5729 10735 5763
rect 10885 5729 10919 5763
rect 11529 5729 11563 5763
rect 12909 5729 12943 5763
rect 13645 5729 13679 5763
rect 14381 5729 14415 5763
rect 3617 5661 3651 5695
rect 3801 5661 3835 5695
rect 5273 5661 5307 5695
rect 7113 5661 7147 5695
rect 8769 5661 8803 5695
rect 10149 5661 10183 5695
rect 11805 5661 11839 5695
rect 12633 5661 12667 5695
rect 13553 5661 13587 5695
rect 14565 5661 14599 5695
rect 3157 5593 3191 5627
rect 4068 5593 4102 5627
rect 7380 5593 7414 5627
rect 15025 5593 15059 5627
rect 15669 5593 15703 5627
rect 1869 5525 1903 5559
rect 6561 5525 6595 5559
rect 9321 5525 9355 5559
rect 9689 5525 9723 5559
rect 10057 5525 10091 5559
rect 10977 5525 11011 5559
rect 11345 5525 11379 5559
rect 11713 5525 11747 5559
rect 12173 5525 12207 5559
rect 12265 5525 12299 5559
rect 12725 5525 12759 5559
rect 13093 5525 13127 5559
rect 13461 5525 13495 5559
rect 1777 5321 1811 5355
rect 2145 5321 2179 5355
rect 4353 5321 4387 5355
rect 4813 5321 4847 5355
rect 10517 5321 10551 5355
rect 10609 5321 10643 5355
rect 11069 5321 11103 5355
rect 11529 5321 11563 5355
rect 11989 5321 12023 5355
rect 13461 5321 13495 5355
rect 13553 5321 13587 5355
rect 13921 5321 13955 5355
rect 15393 5321 15427 5355
rect 3893 5253 3927 5287
rect 5926 5253 5960 5287
rect 7512 5253 7546 5287
rect 9689 5253 9723 5287
rect 12633 5253 12667 5287
rect 14013 5253 14047 5287
rect 14473 5253 14507 5287
rect 15209 5253 15243 5287
rect 2237 5185 2271 5219
rect 2493 5185 2527 5219
rect 4261 5185 4295 5219
rect 7757 5185 7791 5219
rect 7849 5185 7883 5219
rect 8116 5185 8150 5219
rect 11253 5185 11287 5219
rect 11897 5185 11931 5219
rect 12725 5185 12759 5219
rect 14289 5185 14323 5219
rect 1593 5117 1627 5151
rect 1685 5117 1719 5151
rect 4169 5117 4203 5151
rect 6193 5117 6227 5151
rect 9781 5117 9815 5151
rect 9873 5117 9907 5151
rect 10701 5117 10735 5151
rect 12173 5117 12207 5151
rect 12449 5117 12483 5151
rect 13369 5117 13403 5151
rect 14565 5117 14599 5151
rect 15025 5117 15059 5151
rect 6377 5049 6411 5083
rect 9321 5049 9355 5083
rect 14749 5049 14783 5083
rect 3617 4981 3651 5015
rect 4721 4981 4755 5015
rect 9229 4981 9263 5015
rect 10149 4981 10183 5015
rect 13093 4981 13127 5015
rect 15577 4981 15611 5015
rect 5181 4777 5215 4811
rect 8769 4777 8803 4811
rect 13001 4777 13035 4811
rect 14841 4777 14875 4811
rect 14933 4777 14967 4811
rect 15577 4777 15611 4811
rect 7113 4709 7147 4743
rect 13553 4709 13587 4743
rect 14197 4709 14231 4743
rect 1593 4641 1627 4675
rect 1869 4641 1903 4675
rect 9045 4641 9079 4675
rect 9873 4641 9907 4675
rect 10057 4641 10091 4675
rect 10793 4641 10827 4675
rect 10885 4641 10919 4675
rect 11529 4641 11563 4675
rect 11713 4641 11747 4675
rect 12357 4641 12391 4675
rect 15209 4641 15243 4675
rect 2136 4573 2170 4607
rect 3617 4573 3651 4607
rect 3801 4573 3835 4607
rect 7021 4573 7055 4607
rect 8493 4573 8527 4607
rect 9321 4573 9355 4607
rect 10149 4573 10183 4607
rect 10977 4573 11011 4607
rect 12633 4573 12667 4607
rect 13369 4573 13403 4607
rect 13737 4573 13771 4607
rect 14381 4573 14415 4607
rect 4068 4505 4102 4539
rect 5273 4505 5307 4539
rect 8226 4505 8260 4539
rect 14473 4505 14507 4539
rect 15301 4505 15335 4539
rect 1777 4437 1811 4471
rect 3249 4437 3283 4471
rect 3433 4437 3467 4471
rect 9229 4437 9263 4471
rect 9689 4437 9723 4471
rect 10517 4437 10551 4471
rect 11345 4437 11379 4471
rect 11805 4437 11839 4471
rect 12173 4437 12207 4471
rect 12541 4437 12575 4471
rect 13185 4437 13219 4471
rect 13921 4437 13955 4471
rect 1501 4233 1535 4267
rect 1685 4233 1719 4267
rect 1869 4233 1903 4267
rect 9781 4233 9815 4267
rect 10609 4233 10643 4267
rect 11529 4233 11563 4267
rect 12725 4233 12759 4267
rect 13093 4233 13127 4267
rect 14105 4233 14139 4267
rect 15577 4233 15611 4267
rect 3608 4165 3642 4199
rect 9045 4165 9079 4199
rect 9689 4165 9723 4199
rect 13553 4165 13587 4199
rect 14749 4165 14783 4199
rect 2982 4097 3016 4131
rect 3249 4097 3283 4131
rect 3341 4097 3375 4131
rect 4813 4097 4847 4131
rect 5080 4097 5114 4131
rect 6837 4097 6871 4131
rect 6929 4097 6963 4131
rect 7196 4097 7230 4131
rect 8953 4097 8987 4131
rect 10517 4097 10551 4131
rect 11345 4097 11379 4131
rect 11897 4097 11931 4131
rect 14289 4097 14323 4131
rect 14657 4097 14691 4131
rect 6561 4029 6595 4063
rect 9137 4029 9171 4063
rect 9597 4029 9631 4063
rect 10333 4029 10367 4063
rect 11989 4029 12023 4063
rect 12081 4029 12115 4063
rect 12449 4029 12483 4063
rect 12633 4029 12667 4063
rect 13645 4029 13679 4063
rect 13737 4029 13771 4063
rect 15209 4029 15243 4063
rect 8493 3961 8527 3995
rect 11161 3961 11195 3995
rect 13185 3961 13219 3995
rect 14473 3961 14507 3995
rect 15025 3961 15059 3995
rect 4721 3893 4755 3927
rect 6193 3893 6227 3927
rect 8309 3893 8343 3927
rect 8585 3893 8619 3927
rect 10149 3893 10183 3927
rect 10977 3893 11011 3927
rect 15393 3893 15427 3927
rect 1593 3689 1627 3723
rect 3249 3689 3283 3723
rect 6837 3689 6871 3723
rect 7665 3689 7699 3723
rect 13093 3689 13127 3723
rect 15393 3689 15427 3723
rect 15577 3689 15611 3723
rect 5181 3621 5215 3655
rect 5273 3621 5307 3655
rect 8493 3621 8527 3655
rect 8769 3621 8803 3655
rect 9689 3621 9723 3655
rect 1869 3553 1903 3587
rect 3801 3553 3835 3587
rect 5457 3553 5491 3587
rect 7021 3553 7055 3587
rect 7205 3553 7239 3587
rect 7941 3553 7975 3587
rect 8033 3553 8067 3587
rect 9137 3553 9171 3587
rect 10333 3553 10367 3587
rect 11161 3553 11195 3587
rect 12081 3553 12115 3587
rect 12909 3553 12943 3587
rect 13645 3553 13679 3587
rect 1777 3485 1811 3519
rect 3341 3485 3375 3519
rect 4068 3485 4102 3519
rect 5724 3485 5758 3519
rect 9321 3485 9355 3519
rect 10149 3485 10183 3519
rect 11805 3485 11839 3519
rect 12633 3485 12667 3519
rect 13461 3485 13495 3519
rect 13553 3485 13587 3519
rect 14105 3485 14139 3519
rect 14933 3485 14967 3519
rect 15301 3485 15335 3519
rect 2114 3417 2148 3451
rect 8125 3417 8159 3451
rect 11897 3417 11931 3451
rect 14381 3417 14415 3451
rect 3525 3349 3559 3383
rect 7297 3349 7331 3383
rect 9229 3349 9263 3383
rect 9781 3349 9815 3383
rect 10241 3349 10275 3383
rect 10609 3349 10643 3383
rect 10977 3349 11011 3383
rect 11069 3349 11103 3383
rect 11437 3349 11471 3383
rect 12265 3349 12299 3383
rect 12725 3349 12759 3383
rect 14749 3349 14783 3383
rect 15117 3349 15151 3383
rect 2237 3145 2271 3179
rect 2697 3145 2731 3179
rect 6377 3145 6411 3179
rect 7481 3145 7515 3179
rect 7573 3145 7607 3179
rect 7941 3145 7975 3179
rect 10609 3145 10643 3179
rect 11253 3145 11287 3179
rect 11529 3145 11563 3179
rect 12725 3145 12759 3179
rect 1593 3077 1627 3111
rect 5733 3077 5767 3111
rect 6745 3077 6779 3111
rect 8309 3077 8343 3111
rect 8953 3077 8987 3111
rect 9321 3077 9355 3111
rect 9413 3077 9447 3111
rect 10241 3077 10275 3111
rect 14933 3077 14967 3111
rect 1869 3009 1903 3043
rect 2329 3009 2363 3043
rect 2789 3009 2823 3043
rect 3045 3009 3079 3043
rect 4537 3009 4571 3043
rect 4905 3009 4939 3043
rect 4997 3009 5031 3043
rect 5825 3009 5859 3043
rect 8401 3009 8435 3043
rect 11161 3009 11195 3043
rect 11897 3009 11931 3043
rect 11989 3009 12023 3043
rect 13185 3009 13219 3043
rect 13737 3009 13771 3043
rect 14565 3009 14599 3043
rect 14657 3009 14691 3043
rect 15209 3009 15243 3043
rect 2053 2941 2087 2975
rect 4721 2941 4755 2975
rect 5549 2941 5583 2975
rect 6837 2941 6871 2975
rect 6929 2941 6963 2975
rect 7297 2941 7331 2975
rect 8125 2941 8159 2975
rect 9229 2941 9263 2975
rect 10057 2941 10091 2975
rect 10149 2941 10183 2975
rect 10977 2941 11011 2975
rect 12173 2941 12207 2975
rect 12449 2941 12483 2975
rect 12633 2941 12667 2975
rect 13369 2941 13403 2975
rect 14013 2941 14047 2975
rect 15485 2941 15519 2975
rect 4353 2873 4387 2907
rect 5365 2873 5399 2907
rect 6193 2873 6227 2907
rect 8769 2873 8803 2907
rect 4169 2805 4203 2839
rect 9781 2805 9815 2839
rect 13093 2805 13127 2839
rect 14381 2805 14415 2839
rect 4537 2601 4571 2635
rect 5365 2601 5399 2635
rect 9689 2601 9723 2635
rect 13921 2601 13955 2635
rect 15577 2601 15611 2635
rect 5457 2533 5491 2567
rect 12357 2533 12391 2567
rect 14197 2533 14231 2567
rect 1685 2465 1719 2499
rect 2145 2465 2179 2499
rect 2329 2465 2363 2499
rect 2973 2465 3007 2499
rect 3985 2465 4019 2499
rect 4077 2465 4111 2499
rect 4813 2465 4847 2499
rect 5917 2465 5951 2499
rect 6009 2465 6043 2499
rect 6469 2465 6503 2499
rect 6653 2465 6687 2499
rect 7389 2465 7423 2499
rect 7481 2465 7515 2499
rect 8217 2465 8251 2499
rect 9045 2465 9079 2499
rect 9229 2465 9263 2499
rect 9965 2465 9999 2499
rect 10057 2465 10091 2499
rect 11069 2465 11103 2499
rect 11161 2465 11195 2499
rect 12081 2465 12115 2499
rect 12909 2465 12943 2499
rect 13277 2465 13311 2499
rect 13461 2465 13495 2499
rect 14749 2465 14783 2499
rect 1869 2397 1903 2431
rect 3249 2397 3283 2431
rect 5825 2397 5859 2431
rect 6745 2397 6779 2431
rect 11897 2397 11931 2431
rect 12817 2397 12851 2431
rect 13553 2397 13587 2431
rect 14381 2397 14415 2431
rect 14473 2397 14507 2431
rect 15025 2397 15059 2431
rect 2421 2329 2455 2363
rect 4169 2329 4203 2363
rect 4997 2329 5031 2363
rect 8401 2329 8435 2363
rect 10149 2329 10183 2363
rect 11989 2329 12023 2363
rect 12725 2329 12759 2363
rect 15301 2329 15335 2363
rect 2789 2261 2823 2295
rect 3157 2261 3191 2295
rect 3617 2261 3651 2295
rect 4905 2261 4939 2295
rect 7113 2261 7147 2295
rect 7573 2261 7607 2295
rect 7941 2261 7975 2295
rect 8309 2261 8343 2295
rect 8769 2261 8803 2295
rect 9321 2261 9355 2295
rect 10517 2261 10551 2295
rect 10609 2261 10643 2295
rect 10977 2261 11011 2295
rect 11529 2261 11563 2295
<< metal1 >>
rect 4062 17960 4068 18012
rect 4120 18000 4126 18012
rect 6362 18000 6368 18012
rect 4120 17972 6368 18000
rect 4120 17960 4126 17972
rect 6362 17960 6368 17972
rect 6420 17960 6426 18012
rect 13906 17824 13912 17876
rect 13964 17864 13970 17876
rect 15470 17864 15476 17876
rect 13964 17836 15476 17864
rect 13964 17824 13970 17836
rect 15470 17824 15476 17836
rect 15528 17824 15534 17876
rect 1104 17434 16008 17456
rect 1104 17382 4698 17434
rect 4750 17382 4762 17434
rect 4814 17382 4826 17434
rect 4878 17382 4890 17434
rect 4942 17382 4954 17434
rect 5006 17382 8446 17434
rect 8498 17382 8510 17434
rect 8562 17382 8574 17434
rect 8626 17382 8638 17434
rect 8690 17382 8702 17434
rect 8754 17382 12194 17434
rect 12246 17382 12258 17434
rect 12310 17382 12322 17434
rect 12374 17382 12386 17434
rect 12438 17382 12450 17434
rect 12502 17382 16008 17434
rect 1104 17360 16008 17382
rect 934 17212 940 17264
rect 992 17252 998 17264
rect 2133 17255 2191 17261
rect 2133 17252 2145 17255
rect 992 17224 2145 17252
rect 992 17212 998 17224
rect 2133 17221 2145 17224
rect 2179 17221 2191 17255
rect 2133 17215 2191 17221
rect 2409 17187 2467 17193
rect 2409 17153 2421 17187
rect 2455 17184 2467 17187
rect 3142 17184 3148 17196
rect 2455 17156 3148 17184
rect 2455 17153 2467 17156
rect 2409 17147 2467 17153
rect 3142 17144 3148 17156
rect 3200 17144 3206 17196
rect 13078 17048 13084 17060
rect 8266 17020 13084 17048
rect 1946 16940 1952 16992
rect 2004 16980 2010 16992
rect 8266 16980 8294 17020
rect 13078 17008 13084 17020
rect 13136 17048 13142 17060
rect 13998 17048 14004 17060
rect 13136 17020 14004 17048
rect 13136 17008 13142 17020
rect 13998 17008 14004 17020
rect 14056 17008 14062 17060
rect 2004 16952 8294 16980
rect 2004 16940 2010 16952
rect 1104 16890 16008 16912
rect 1104 16838 2824 16890
rect 2876 16838 2888 16890
rect 2940 16838 2952 16890
rect 3004 16838 3016 16890
rect 3068 16838 3080 16890
rect 3132 16838 6572 16890
rect 6624 16838 6636 16890
rect 6688 16838 6700 16890
rect 6752 16838 6764 16890
rect 6816 16838 6828 16890
rect 6880 16838 10320 16890
rect 10372 16838 10384 16890
rect 10436 16838 10448 16890
rect 10500 16838 10512 16890
rect 10564 16838 10576 16890
rect 10628 16838 14068 16890
rect 14120 16838 14132 16890
rect 14184 16838 14196 16890
rect 14248 16838 14260 16890
rect 14312 16838 14324 16890
rect 14376 16838 16008 16890
rect 1104 16816 16008 16838
rect 1578 16736 1584 16788
rect 1636 16776 1642 16788
rect 9766 16776 9772 16788
rect 1636 16748 9772 16776
rect 1636 16736 1642 16748
rect 9766 16736 9772 16748
rect 9824 16736 9830 16788
rect 1762 16668 1768 16720
rect 1820 16708 1826 16720
rect 1820 16680 8340 16708
rect 1820 16668 1826 16680
rect 6178 16532 6184 16584
rect 6236 16572 6242 16584
rect 8202 16572 8208 16584
rect 6236 16544 8208 16572
rect 6236 16532 6242 16544
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 8312 16572 8340 16680
rect 10042 16572 10048 16584
rect 8312 16544 10048 16572
rect 10042 16532 10048 16544
rect 10100 16532 10106 16584
rect 2314 16396 2320 16448
rect 2372 16436 2378 16448
rect 7742 16436 7748 16448
rect 2372 16408 7748 16436
rect 2372 16396 2378 16408
rect 7742 16396 7748 16408
rect 7800 16396 7806 16448
rect 1104 16346 16008 16368
rect 1104 16294 4698 16346
rect 4750 16294 4762 16346
rect 4814 16294 4826 16346
rect 4878 16294 4890 16346
rect 4942 16294 4954 16346
rect 5006 16294 8446 16346
rect 8498 16294 8510 16346
rect 8562 16294 8574 16346
rect 8626 16294 8638 16346
rect 8690 16294 8702 16346
rect 8754 16294 12194 16346
rect 12246 16294 12258 16346
rect 12310 16294 12322 16346
rect 12374 16294 12386 16346
rect 12438 16294 12450 16346
rect 12502 16294 16008 16346
rect 1104 16272 16008 16294
rect 5350 16232 5356 16244
rect 5311 16204 5356 16232
rect 5350 16192 5356 16204
rect 5408 16192 5414 16244
rect 2038 16124 2044 16176
rect 2096 16164 2102 16176
rect 4893 16167 4951 16173
rect 4893 16164 4905 16167
rect 2096 16136 4905 16164
rect 2096 16124 2102 16136
rect 4893 16133 4905 16136
rect 4939 16133 4951 16167
rect 4893 16127 4951 16133
rect 5169 16099 5227 16105
rect 5169 16065 5181 16099
rect 5215 16096 5227 16099
rect 5368 16096 5396 16192
rect 5215 16068 5396 16096
rect 5215 16065 5227 16068
rect 5169 16059 5227 16065
rect 7834 16056 7840 16108
rect 7892 16096 7898 16108
rect 12894 16096 12900 16108
rect 7892 16068 12900 16096
rect 7892 16056 7898 16068
rect 12894 16056 12900 16068
rect 12952 16056 12958 16108
rect 2498 15988 2504 16040
rect 2556 16028 2562 16040
rect 5534 16028 5540 16040
rect 2556 16000 5540 16028
rect 2556 15988 2562 16000
rect 5534 15988 5540 16000
rect 5592 15988 5598 16040
rect 5810 15988 5816 16040
rect 5868 16028 5874 16040
rect 9398 16028 9404 16040
rect 5868 16000 9404 16028
rect 5868 15988 5874 16000
rect 9398 15988 9404 16000
rect 9456 15988 9462 16040
rect 5626 15920 5632 15972
rect 5684 15960 5690 15972
rect 10226 15960 10232 15972
rect 5684 15932 10232 15960
rect 5684 15920 5690 15932
rect 10226 15920 10232 15932
rect 10284 15960 10290 15972
rect 13814 15960 13820 15972
rect 10284 15932 13820 15960
rect 10284 15920 10290 15932
rect 13814 15920 13820 15932
rect 13872 15920 13878 15972
rect 1026 15852 1032 15904
rect 1084 15892 1090 15904
rect 1670 15892 1676 15904
rect 1084 15864 1676 15892
rect 1084 15852 1090 15864
rect 1670 15852 1676 15864
rect 1728 15852 1734 15904
rect 3694 15892 3700 15904
rect 3655 15864 3700 15892
rect 3694 15852 3700 15864
rect 3752 15852 3758 15904
rect 9398 15852 9404 15904
rect 9456 15892 9462 15904
rect 15102 15892 15108 15904
rect 9456 15864 15108 15892
rect 9456 15852 9462 15864
rect 15102 15852 15108 15864
rect 15160 15892 15166 15904
rect 15746 15892 15752 15904
rect 15160 15864 15752 15892
rect 15160 15852 15166 15864
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 1104 15802 16008 15824
rect 1104 15750 2824 15802
rect 2876 15750 2888 15802
rect 2940 15750 2952 15802
rect 3004 15750 3016 15802
rect 3068 15750 3080 15802
rect 3132 15750 6572 15802
rect 6624 15750 6636 15802
rect 6688 15750 6700 15802
rect 6752 15750 6764 15802
rect 6816 15750 6828 15802
rect 6880 15750 10320 15802
rect 10372 15750 10384 15802
rect 10436 15750 10448 15802
rect 10500 15750 10512 15802
rect 10564 15750 10576 15802
rect 10628 15750 14068 15802
rect 14120 15750 14132 15802
rect 14184 15750 14196 15802
rect 14248 15750 14260 15802
rect 14312 15750 14324 15802
rect 14376 15750 16008 15802
rect 1104 15728 16008 15750
rect 3234 15648 3240 15700
rect 3292 15688 3298 15700
rect 3421 15691 3479 15697
rect 3421 15688 3433 15691
rect 3292 15660 3433 15688
rect 3292 15648 3298 15660
rect 3421 15657 3433 15660
rect 3467 15657 3479 15691
rect 3421 15651 3479 15657
rect 3510 15648 3516 15700
rect 3568 15688 3574 15700
rect 4433 15691 4491 15697
rect 4433 15688 4445 15691
rect 3568 15660 4445 15688
rect 3568 15648 3574 15660
rect 4433 15657 4445 15660
rect 4479 15657 4491 15691
rect 4433 15651 4491 15657
rect 4985 15691 5043 15697
rect 4985 15657 4997 15691
rect 5031 15688 5043 15691
rect 5350 15688 5356 15700
rect 5031 15660 5356 15688
rect 5031 15657 5043 15660
rect 4985 15651 5043 15657
rect 5350 15648 5356 15660
rect 5408 15648 5414 15700
rect 7006 15688 7012 15700
rect 6967 15660 7012 15688
rect 7006 15648 7012 15660
rect 7064 15648 7070 15700
rect 7653 15691 7711 15697
rect 7653 15657 7665 15691
rect 7699 15688 7711 15691
rect 7742 15688 7748 15700
rect 7699 15660 7748 15688
rect 7699 15657 7711 15660
rect 7653 15651 7711 15657
rect 7742 15648 7748 15660
rect 7800 15648 7806 15700
rect 9950 15688 9956 15700
rect 7852 15660 9956 15688
rect 2406 15580 2412 15632
rect 2464 15620 2470 15632
rect 3602 15620 3608 15632
rect 2464 15592 3608 15620
rect 2464 15580 2470 15592
rect 3602 15580 3608 15592
rect 3660 15580 3666 15632
rect 5169 15623 5227 15629
rect 5169 15620 5181 15623
rect 3712 15592 5181 15620
rect 3050 15512 3056 15564
rect 3108 15552 3114 15564
rect 3712 15552 3740 15592
rect 5169 15589 5181 15592
rect 5215 15620 5227 15623
rect 7852 15620 7880 15660
rect 9950 15648 9956 15660
rect 10008 15688 10014 15700
rect 10870 15688 10876 15700
rect 10008 15660 10876 15688
rect 10008 15648 10014 15660
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 5215 15592 7880 15620
rect 5215 15589 5227 15592
rect 5169 15583 5227 15589
rect 9214 15580 9220 15632
rect 9272 15620 9278 15632
rect 11790 15620 11796 15632
rect 9272 15592 11796 15620
rect 9272 15580 9278 15592
rect 11790 15580 11796 15592
rect 11848 15620 11854 15632
rect 14550 15620 14556 15632
rect 11848 15592 14556 15620
rect 11848 15580 11854 15592
rect 14550 15580 14556 15592
rect 14608 15580 14614 15632
rect 3970 15552 3976 15564
rect 3108 15524 3740 15552
rect 3931 15524 3976 15552
rect 3108 15512 3114 15524
rect 3970 15512 3976 15524
rect 4028 15512 4034 15564
rect 5350 15552 5356 15564
rect 4264 15524 5356 15552
rect 4264 15493 4292 15524
rect 5350 15512 5356 15524
rect 5408 15512 5414 15564
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 7377 15555 7435 15561
rect 7377 15552 7389 15555
rect 5592 15524 7389 15552
rect 5592 15512 5598 15524
rect 7377 15521 7389 15524
rect 7423 15552 7435 15555
rect 7423 15524 9628 15552
rect 7423 15521 7435 15524
rect 7377 15515 7435 15521
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15453 3663 15487
rect 3605 15447 3663 15453
rect 4249 15487 4307 15493
rect 4249 15453 4261 15487
rect 4295 15453 4307 15487
rect 4249 15447 4307 15453
rect 3620 15416 3648 15447
rect 4338 15444 4344 15496
rect 4396 15484 4402 15496
rect 4617 15487 4675 15493
rect 4617 15484 4629 15487
rect 4396 15456 4629 15484
rect 4396 15444 4402 15456
rect 4617 15453 4629 15456
rect 4663 15484 4675 15487
rect 4801 15487 4859 15493
rect 4801 15484 4813 15487
rect 4663 15456 4813 15484
rect 4663 15453 4675 15456
rect 4617 15447 4675 15453
rect 4801 15453 4813 15456
rect 4847 15484 4859 15487
rect 5994 15484 6000 15496
rect 4847 15456 6000 15484
rect 4847 15453 4859 15456
rect 4801 15447 4859 15453
rect 5994 15444 6000 15456
rect 6052 15444 6058 15496
rect 6270 15444 6276 15496
rect 6328 15484 6334 15496
rect 6457 15487 6515 15493
rect 6457 15484 6469 15487
rect 6328 15456 6469 15484
rect 6328 15444 6334 15456
rect 6457 15453 6469 15456
rect 6503 15453 6515 15487
rect 6457 15447 6515 15453
rect 8018 15444 8024 15496
rect 8076 15484 8082 15496
rect 9030 15484 9036 15496
rect 8076 15456 9036 15484
rect 8076 15444 8082 15456
rect 9030 15444 9036 15456
rect 9088 15444 9094 15496
rect 9600 15484 9628 15524
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 15562 15552 15568 15564
rect 9732 15524 15568 15552
rect 9732 15512 9738 15524
rect 15562 15512 15568 15524
rect 15620 15512 15626 15564
rect 10686 15484 10692 15496
rect 9600 15456 10692 15484
rect 10686 15444 10692 15456
rect 10744 15444 10750 15496
rect 3694 15416 3700 15428
rect 3607 15388 3700 15416
rect 3694 15376 3700 15388
rect 3752 15416 3758 15428
rect 4430 15416 4436 15428
rect 3752 15388 4436 15416
rect 3752 15376 3758 15388
rect 4430 15376 4436 15388
rect 4488 15376 4494 15428
rect 4522 15376 4528 15428
rect 4580 15416 4586 15428
rect 7285 15419 7343 15425
rect 7285 15416 7297 15419
rect 4580 15388 7297 15416
rect 4580 15376 4586 15388
rect 7285 15385 7297 15388
rect 7331 15416 7343 15419
rect 10134 15416 10140 15428
rect 7331 15388 10140 15416
rect 7331 15385 7343 15388
rect 7285 15379 7343 15385
rect 10134 15376 10140 15388
rect 10192 15376 10198 15428
rect 3234 15308 3240 15360
rect 3292 15348 3298 15360
rect 4338 15348 4344 15360
rect 3292 15320 4344 15348
rect 3292 15308 3298 15320
rect 4338 15308 4344 15320
rect 4396 15308 4402 15360
rect 5534 15348 5540 15360
rect 5495 15320 5540 15348
rect 5534 15308 5540 15320
rect 5592 15308 5598 15360
rect 6178 15308 6184 15360
rect 6236 15348 6242 15360
rect 6273 15351 6331 15357
rect 6273 15348 6285 15351
rect 6236 15320 6285 15348
rect 6236 15308 6242 15320
rect 6273 15317 6285 15320
rect 6319 15317 6331 15351
rect 7742 15348 7748 15360
rect 7703 15320 7748 15348
rect 6273 15311 6331 15317
rect 7742 15308 7748 15320
rect 7800 15308 7806 15360
rect 8021 15351 8079 15357
rect 8021 15317 8033 15351
rect 8067 15348 8079 15351
rect 8110 15348 8116 15360
rect 8067 15320 8116 15348
rect 8067 15317 8079 15320
rect 8021 15311 8079 15317
rect 8110 15308 8116 15320
rect 8168 15308 8174 15360
rect 9766 15308 9772 15360
rect 9824 15348 9830 15360
rect 15194 15348 15200 15360
rect 9824 15320 15200 15348
rect 9824 15308 9830 15320
rect 15194 15308 15200 15320
rect 15252 15308 15258 15360
rect 1104 15258 16008 15280
rect 1104 15206 4698 15258
rect 4750 15206 4762 15258
rect 4814 15206 4826 15258
rect 4878 15206 4890 15258
rect 4942 15206 4954 15258
rect 5006 15206 8446 15258
rect 8498 15206 8510 15258
rect 8562 15206 8574 15258
rect 8626 15206 8638 15258
rect 8690 15206 8702 15258
rect 8754 15206 12194 15258
rect 12246 15206 12258 15258
rect 12310 15206 12322 15258
rect 12374 15206 12386 15258
rect 12438 15206 12450 15258
rect 12502 15206 16008 15258
rect 1104 15184 16008 15206
rect 3050 15144 3056 15156
rect 3011 15116 3056 15144
rect 3050 15104 3056 15116
rect 3108 15104 3114 15156
rect 3234 15144 3240 15156
rect 3195 15116 3240 15144
rect 3234 15104 3240 15116
rect 3292 15104 3298 15156
rect 3602 15144 3608 15156
rect 3563 15116 3608 15144
rect 3602 15104 3608 15116
rect 3660 15104 3666 15156
rect 4065 15147 4123 15153
rect 4065 15113 4077 15147
rect 4111 15113 4123 15147
rect 4065 15107 4123 15113
rect 4433 15147 4491 15153
rect 4433 15113 4445 15147
rect 4479 15144 4491 15147
rect 4522 15144 4528 15156
rect 4479 15116 4528 15144
rect 4479 15113 4491 15116
rect 4433 15107 4491 15113
rect 750 15036 756 15088
rect 808 15076 814 15088
rect 3252 15076 3280 15104
rect 808 15048 3280 15076
rect 808 15036 814 15048
rect 3326 15036 3332 15088
rect 3384 15076 3390 15088
rect 4080 15076 4108 15107
rect 4338 15076 4344 15088
rect 3384 15048 4108 15076
rect 4251 15048 4344 15076
rect 3384 15036 3390 15048
rect 3421 15011 3479 15017
rect 3421 14977 3433 15011
rect 3467 15008 3479 15011
rect 3694 15008 3700 15020
rect 3467 14980 3700 15008
rect 3467 14977 3479 14980
rect 3421 14971 3479 14977
rect 3694 14968 3700 14980
rect 3752 14968 3758 15020
rect 3786 14968 3792 15020
rect 3844 15008 3850 15020
rect 4264 15017 4292 15048
rect 4338 15036 4344 15048
rect 4396 15076 4402 15088
rect 4448 15076 4476 15107
rect 4522 15104 4528 15116
rect 4580 15104 4586 15156
rect 5077 15147 5135 15153
rect 5077 15113 5089 15147
rect 5123 15144 5135 15147
rect 5350 15144 5356 15156
rect 5123 15116 5356 15144
rect 5123 15113 5135 15116
rect 5077 15107 5135 15113
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 5997 15147 6055 15153
rect 5997 15144 6009 15147
rect 5776 15116 6009 15144
rect 5776 15104 5782 15116
rect 5997 15113 6009 15116
rect 6043 15113 6055 15147
rect 6362 15144 6368 15156
rect 6323 15116 6368 15144
rect 5997 15107 6055 15113
rect 6362 15104 6368 15116
rect 6420 15104 6426 15156
rect 7282 15104 7288 15156
rect 7340 15144 7346 15156
rect 7837 15147 7895 15153
rect 7837 15144 7849 15147
rect 7340 15116 7849 15144
rect 7340 15104 7346 15116
rect 7837 15113 7849 15116
rect 7883 15113 7895 15147
rect 7837 15107 7895 15113
rect 4396 15048 4476 15076
rect 4396 15036 4402 15048
rect 6086 15036 6092 15088
rect 6144 15076 6150 15088
rect 6917 15079 6975 15085
rect 6917 15076 6929 15079
rect 6144 15048 6929 15076
rect 6144 15036 6150 15048
rect 6917 15045 6929 15048
rect 6963 15045 6975 15079
rect 6917 15039 6975 15045
rect 4249 15011 4307 15017
rect 3844 14980 3889 15008
rect 3844 14968 3850 14980
rect 4249 14977 4261 15011
rect 4295 14977 4307 15011
rect 4617 15011 4675 15017
rect 4617 15008 4629 15011
rect 4249 14971 4307 14977
rect 4356 14980 4629 15008
rect 2869 14943 2927 14949
rect 2869 14940 2881 14943
rect 2746 14912 2881 14940
rect 2746 14816 2774 14912
rect 2869 14909 2881 14912
rect 2915 14940 2927 14943
rect 3804 14940 3832 14968
rect 4356 14940 4384 14980
rect 4617 14977 4629 14980
rect 4663 14977 4675 15011
rect 5166 15008 5172 15020
rect 5127 14980 5172 15008
rect 4617 14971 4675 14977
rect 5166 14968 5172 14980
rect 5224 14968 5230 15020
rect 5442 15008 5448 15020
rect 5403 14980 5448 15008
rect 5442 14968 5448 14980
rect 5500 14968 5506 15020
rect 6178 15008 6184 15020
rect 6091 14980 6184 15008
rect 6178 14968 6184 14980
rect 6236 15008 6242 15020
rect 7558 15008 7564 15020
rect 6236 14980 7564 15008
rect 6236 14968 6242 14980
rect 7558 14968 7564 14980
rect 7616 14968 7622 15020
rect 7653 15011 7711 15017
rect 7653 14977 7665 15011
rect 7699 15008 7711 15011
rect 7742 15008 7748 15020
rect 7699 14980 7748 15008
rect 7699 14977 7711 14980
rect 7653 14971 7711 14977
rect 7742 14968 7748 14980
rect 7800 14968 7806 15020
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 14977 8079 15011
rect 8021 14971 8079 14977
rect 2915 14912 4384 14940
rect 2915 14909 2927 14912
rect 2869 14903 2927 14909
rect 4430 14900 4436 14952
rect 4488 14940 4494 14952
rect 4801 14943 4859 14949
rect 4801 14940 4813 14943
rect 4488 14912 4813 14940
rect 4488 14900 4494 14912
rect 4801 14909 4813 14912
rect 4847 14909 4859 14943
rect 5350 14940 5356 14952
rect 4801 14903 4859 14909
rect 4908 14912 5356 14940
rect 3050 14832 3056 14884
rect 3108 14872 3114 14884
rect 3234 14872 3240 14884
rect 3108 14844 3240 14872
rect 3108 14832 3114 14844
rect 3234 14832 3240 14844
rect 3292 14832 3298 14884
rect 3970 14832 3976 14884
rect 4028 14872 4034 14884
rect 4908 14872 4936 14912
rect 5350 14900 5356 14912
rect 5408 14900 5414 14952
rect 5534 14900 5540 14952
rect 5592 14940 5598 14952
rect 5813 14943 5871 14949
rect 5813 14940 5825 14943
rect 5592 14912 5825 14940
rect 5592 14900 5598 14912
rect 5813 14909 5825 14912
rect 5859 14909 5871 14943
rect 7006 14940 7012 14952
rect 6967 14912 7012 14940
rect 5813 14903 5871 14909
rect 7006 14900 7012 14912
rect 7064 14900 7070 14952
rect 7098 14900 7104 14952
rect 7156 14940 7162 14952
rect 7156 14912 7201 14940
rect 7156 14900 7162 14912
rect 4028 14844 4936 14872
rect 5629 14875 5687 14881
rect 4028 14832 4034 14844
rect 5629 14841 5641 14875
rect 5675 14872 5687 14875
rect 6086 14872 6092 14884
rect 5675 14844 6092 14872
rect 5675 14841 5687 14844
rect 5629 14835 5687 14841
rect 6086 14832 6092 14844
rect 6144 14832 6150 14884
rect 7190 14832 7196 14884
rect 7248 14872 7254 14884
rect 7469 14875 7527 14881
rect 7469 14872 7481 14875
rect 7248 14844 7481 14872
rect 7248 14832 7254 14844
rect 7469 14841 7481 14844
rect 7515 14841 7527 14875
rect 8036 14872 8064 14971
rect 8478 14900 8484 14952
rect 8536 14940 8542 14952
rect 12802 14940 12808 14952
rect 8536 14912 12808 14940
rect 8536 14900 8542 14912
rect 12802 14900 12808 14912
rect 12860 14900 12866 14952
rect 8036 14844 8892 14872
rect 7469 14835 7527 14841
rect 8864 14816 8892 14844
rect 1118 14764 1124 14816
rect 1176 14804 1182 14816
rect 2593 14807 2651 14813
rect 2593 14804 2605 14807
rect 1176 14776 2605 14804
rect 1176 14764 1182 14776
rect 2593 14773 2605 14776
rect 2639 14773 2651 14807
rect 2593 14767 2651 14773
rect 2682 14764 2688 14816
rect 2740 14776 2774 14816
rect 2740 14764 2746 14776
rect 5350 14764 5356 14816
rect 5408 14804 5414 14816
rect 6549 14807 6607 14813
rect 6549 14804 6561 14807
rect 5408 14776 6561 14804
rect 5408 14764 5414 14776
rect 6549 14773 6561 14776
rect 6595 14773 6607 14807
rect 6549 14767 6607 14773
rect 7374 14764 7380 14816
rect 7432 14804 7438 14816
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 7432 14776 8217 14804
rect 7432 14764 7438 14776
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 8478 14804 8484 14816
rect 8439 14776 8484 14804
rect 8205 14767 8263 14773
rect 8478 14764 8484 14776
rect 8536 14764 8542 14816
rect 8662 14804 8668 14816
rect 8623 14776 8668 14804
rect 8662 14764 8668 14776
rect 8720 14764 8726 14816
rect 8846 14804 8852 14816
rect 8807 14776 8852 14804
rect 8846 14764 8852 14776
rect 8904 14764 8910 14816
rect 9674 14764 9680 14816
rect 9732 14804 9738 14816
rect 12066 14804 12072 14816
rect 9732 14776 12072 14804
rect 9732 14764 9738 14776
rect 12066 14764 12072 14776
rect 12124 14764 12130 14816
rect 1104 14714 16008 14736
rect 1104 14662 2824 14714
rect 2876 14662 2888 14714
rect 2940 14662 2952 14714
rect 3004 14662 3016 14714
rect 3068 14662 3080 14714
rect 3132 14662 6572 14714
rect 6624 14662 6636 14714
rect 6688 14662 6700 14714
rect 6752 14662 6764 14714
rect 6816 14662 6828 14714
rect 6880 14662 10320 14714
rect 10372 14662 10384 14714
rect 10436 14662 10448 14714
rect 10500 14662 10512 14714
rect 10564 14662 10576 14714
rect 10628 14662 14068 14714
rect 14120 14662 14132 14714
rect 14184 14662 14196 14714
rect 14248 14662 14260 14714
rect 14312 14662 14324 14714
rect 14376 14662 16008 14714
rect 1104 14640 16008 14662
rect 1210 14560 1216 14612
rect 1268 14600 1274 14612
rect 4522 14600 4528 14612
rect 1268 14572 4528 14600
rect 1268 14560 1274 14572
rect 4522 14560 4528 14572
rect 4580 14560 4586 14612
rect 4614 14560 4620 14612
rect 4672 14600 4678 14612
rect 5261 14603 5319 14609
rect 5261 14600 5273 14603
rect 4672 14572 5273 14600
rect 4672 14560 4678 14572
rect 5261 14569 5273 14572
rect 5307 14569 5319 14603
rect 7193 14603 7251 14609
rect 7193 14600 7205 14603
rect 5261 14563 5319 14569
rect 5368 14572 7205 14600
rect 842 14492 848 14544
rect 900 14532 906 14544
rect 2498 14532 2504 14544
rect 900 14504 2504 14532
rect 900 14492 906 14504
rect 2498 14492 2504 14504
rect 2556 14532 2562 14544
rect 2593 14535 2651 14541
rect 2593 14532 2605 14535
rect 2556 14504 2605 14532
rect 2556 14492 2562 14504
rect 2593 14501 2605 14504
rect 2639 14501 2651 14535
rect 3326 14532 3332 14544
rect 3287 14504 3332 14532
rect 2593 14495 2651 14501
rect 3326 14492 3332 14504
rect 3384 14492 3390 14544
rect 3602 14532 3608 14544
rect 3563 14504 3608 14532
rect 3602 14492 3608 14504
rect 3660 14492 3666 14544
rect 4154 14492 4160 14544
rect 4212 14532 4218 14544
rect 4893 14535 4951 14541
rect 4893 14532 4905 14535
rect 4212 14504 4905 14532
rect 4212 14492 4218 14504
rect 4893 14501 4905 14504
rect 4939 14501 4951 14535
rect 4893 14495 4951 14501
rect 1946 14464 1952 14476
rect 1907 14436 1952 14464
rect 1946 14424 1952 14436
rect 2004 14424 2010 14476
rect 2222 14464 2228 14476
rect 2183 14436 2228 14464
rect 2222 14424 2228 14436
rect 2280 14424 2286 14476
rect 2869 14467 2927 14473
rect 2869 14433 2881 14467
rect 2915 14464 2927 14467
rect 3053 14467 3111 14473
rect 3053 14464 3065 14467
rect 2915 14436 3065 14464
rect 2915 14433 2927 14436
rect 2869 14427 2927 14433
rect 3053 14433 3065 14436
rect 3099 14464 3111 14467
rect 3099 14436 4016 14464
rect 3099 14433 3111 14436
rect 3053 14427 3111 14433
rect 2501 14399 2559 14405
rect 2501 14365 2513 14399
rect 2547 14396 2559 14399
rect 3602 14396 3608 14408
rect 2547 14368 3608 14396
rect 2547 14365 2559 14368
rect 2501 14359 2559 14365
rect 3602 14356 3608 14368
rect 3660 14356 3666 14408
rect 3786 14396 3792 14408
rect 3747 14368 3792 14396
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 3988 14396 4016 14436
rect 4062 14424 4068 14476
rect 4120 14464 4126 14476
rect 5368 14464 5396 14572
rect 7193 14569 7205 14572
rect 7239 14569 7251 14603
rect 7193 14563 7251 14569
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 8113 14603 8171 14609
rect 8113 14600 8125 14603
rect 7708 14572 8125 14600
rect 7708 14560 7714 14572
rect 8113 14569 8125 14572
rect 8159 14569 8171 14603
rect 8113 14563 8171 14569
rect 8202 14560 8208 14612
rect 8260 14600 8266 14612
rect 8481 14603 8539 14609
rect 8481 14600 8493 14603
rect 8260 14572 8493 14600
rect 8260 14560 8266 14572
rect 8481 14569 8493 14572
rect 8527 14569 8539 14603
rect 8481 14563 8539 14569
rect 8846 14560 8852 14612
rect 8904 14600 8910 14612
rect 9769 14603 9827 14609
rect 9769 14600 9781 14603
rect 8904 14572 9781 14600
rect 8904 14560 8910 14572
rect 9769 14569 9781 14572
rect 9815 14600 9827 14603
rect 14642 14600 14648 14612
rect 9815 14572 14648 14600
rect 9815 14569 9827 14572
rect 9769 14563 9827 14569
rect 14642 14560 14648 14572
rect 14700 14560 14706 14612
rect 5442 14492 5448 14544
rect 5500 14492 5506 14544
rect 5718 14492 5724 14544
rect 5776 14532 5782 14544
rect 6365 14535 6423 14541
rect 6365 14532 6377 14535
rect 5776 14504 6377 14532
rect 5776 14492 5782 14504
rect 6365 14501 6377 14504
rect 6411 14501 6423 14535
rect 6365 14495 6423 14501
rect 7834 14492 7840 14544
rect 7892 14532 7898 14544
rect 9033 14535 9091 14541
rect 9033 14532 9045 14535
rect 7892 14504 9045 14532
rect 7892 14492 7898 14504
rect 9033 14501 9045 14504
rect 9079 14532 9091 14535
rect 9214 14532 9220 14544
rect 9079 14504 9220 14532
rect 9079 14501 9091 14504
rect 9033 14495 9091 14501
rect 9214 14492 9220 14504
rect 9272 14492 9278 14544
rect 9398 14492 9404 14544
rect 9456 14532 9462 14544
rect 12618 14532 12624 14544
rect 9456 14504 12624 14532
rect 9456 14492 9462 14504
rect 12618 14492 12624 14504
rect 12676 14492 12682 14544
rect 4120 14436 5396 14464
rect 5460 14464 5488 14492
rect 6086 14464 6092 14476
rect 5460 14436 6092 14464
rect 4120 14424 4126 14436
rect 6086 14424 6092 14436
rect 6144 14424 6150 14476
rect 6917 14467 6975 14473
rect 6917 14464 6929 14467
rect 6196 14436 6929 14464
rect 4338 14396 4344 14408
rect 3988 14368 4344 14396
rect 4338 14356 4344 14368
rect 4396 14356 4402 14408
rect 4525 14399 4583 14405
rect 4525 14365 4537 14399
rect 4571 14365 4583 14399
rect 4525 14359 4583 14365
rect 2038 14288 2044 14340
rect 2096 14328 2102 14340
rect 2682 14328 2688 14340
rect 2096 14300 2688 14328
rect 2096 14288 2102 14300
rect 2682 14288 2688 14300
rect 2740 14328 2746 14340
rect 3145 14331 3203 14337
rect 3145 14328 3157 14331
rect 2740 14300 3157 14328
rect 2740 14288 2746 14300
rect 3145 14297 3157 14300
rect 3191 14297 3203 14331
rect 3145 14291 3203 14297
rect 3326 14288 3332 14340
rect 3384 14328 3390 14340
rect 3510 14328 3516 14340
rect 3384 14300 3516 14328
rect 3384 14288 3390 14300
rect 3510 14288 3516 14300
rect 3568 14288 3574 14340
rect 3694 14288 3700 14340
rect 3752 14328 3758 14340
rect 3973 14331 4031 14337
rect 3973 14328 3985 14331
rect 3752 14300 3985 14328
rect 3752 14288 3758 14300
rect 3973 14297 3985 14300
rect 4019 14297 4031 14331
rect 3973 14291 4031 14297
rect 4246 14288 4252 14340
rect 4304 14328 4310 14340
rect 4540 14328 4568 14359
rect 4614 14356 4620 14408
rect 4672 14396 4678 14408
rect 5077 14399 5135 14405
rect 4672 14368 5028 14396
rect 4672 14356 4678 14368
rect 5000 14328 5028 14368
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5166 14396 5172 14408
rect 5123 14368 5172 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 5445 14399 5503 14405
rect 5445 14365 5457 14399
rect 5491 14396 5503 14399
rect 5534 14396 5540 14408
rect 5491 14368 5540 14396
rect 5491 14365 5503 14368
rect 5445 14359 5503 14365
rect 5460 14328 5488 14359
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 5902 14396 5908 14408
rect 5863 14368 5908 14396
rect 5902 14356 5908 14368
rect 5960 14356 5966 14408
rect 4304 14300 4384 14328
rect 4540 14300 4752 14328
rect 5000 14300 5488 14328
rect 4304 14288 4310 14300
rect 934 14220 940 14272
rect 992 14260 998 14272
rect 1673 14263 1731 14269
rect 1673 14260 1685 14263
rect 992 14232 1685 14260
rect 992 14220 998 14232
rect 1673 14229 1685 14232
rect 1719 14260 1731 14263
rect 4154 14260 4160 14272
rect 1719 14232 4160 14260
rect 1719 14229 1731 14232
rect 1673 14223 1731 14229
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 4356 14269 4384 14300
rect 4724 14269 4752 14300
rect 5626 14288 5632 14340
rect 5684 14328 5690 14340
rect 6196 14328 6224 14436
rect 6917 14433 6929 14436
rect 6963 14433 6975 14467
rect 6917 14427 6975 14433
rect 7466 14424 7472 14476
rect 7524 14464 7530 14476
rect 7745 14467 7803 14473
rect 7745 14464 7757 14467
rect 7524 14436 7757 14464
rect 7524 14424 7530 14436
rect 7745 14433 7757 14436
rect 7791 14433 7803 14467
rect 7745 14427 7803 14433
rect 8202 14424 8208 14476
rect 8260 14464 8266 14476
rect 9125 14467 9183 14473
rect 8260 14436 8616 14464
rect 8260 14424 8266 14436
rect 6822 14396 6828 14408
rect 6783 14368 6828 14396
rect 6822 14356 6828 14368
rect 6880 14356 6886 14408
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 7653 14399 7711 14405
rect 7653 14396 7665 14399
rect 7432 14368 7665 14396
rect 7432 14356 7438 14368
rect 7653 14365 7665 14368
rect 7699 14396 7711 14399
rect 7926 14396 7932 14408
rect 7699 14368 7932 14396
rect 7699 14365 7711 14368
rect 7653 14359 7711 14365
rect 7926 14356 7932 14368
rect 7984 14356 7990 14408
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 8478 14396 8484 14408
rect 8343 14368 8484 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 5684 14300 6224 14328
rect 6733 14331 6791 14337
rect 5684 14288 5690 14300
rect 6733 14297 6745 14331
rect 6779 14328 6791 14331
rect 7282 14328 7288 14340
rect 6779 14300 7288 14328
rect 6779 14297 6791 14300
rect 6733 14291 6791 14297
rect 7282 14288 7288 14300
rect 7340 14288 7346 14340
rect 7558 14328 7564 14340
rect 7519 14300 7564 14328
rect 7558 14288 7564 14300
rect 7616 14288 7622 14340
rect 8588 14328 8616 14436
rect 9125 14433 9137 14467
rect 9171 14464 9183 14467
rect 11698 14464 11704 14476
rect 9171 14436 11704 14464
rect 9171 14433 9183 14436
rect 9125 14427 9183 14433
rect 8665 14399 8723 14405
rect 8665 14365 8677 14399
rect 8711 14396 8723 14399
rect 9140 14396 9168 14427
rect 11698 14424 11704 14436
rect 11756 14424 11762 14476
rect 9582 14396 9588 14408
rect 8711 14368 9168 14396
rect 9495 14368 9588 14396
rect 8711 14365 8723 14368
rect 8665 14359 8723 14365
rect 9582 14356 9588 14368
rect 9640 14396 9646 14408
rect 11790 14396 11796 14408
rect 9640 14368 11796 14396
rect 9640 14356 9646 14368
rect 11790 14356 11796 14368
rect 11848 14356 11854 14408
rect 12986 14396 12992 14408
rect 12268 14368 12992 14396
rect 12268 14328 12296 14368
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 13630 14328 13636 14340
rect 8588 14300 12296 14328
rect 12406 14300 13636 14328
rect 4341 14263 4399 14269
rect 4341 14229 4353 14263
rect 4387 14229 4399 14263
rect 4341 14223 4399 14229
rect 4709 14263 4767 14269
rect 4709 14229 4721 14263
rect 4755 14260 4767 14263
rect 5166 14260 5172 14272
rect 4755 14232 5172 14260
rect 4755 14229 4767 14232
rect 4709 14223 4767 14229
rect 5166 14220 5172 14232
rect 5224 14220 5230 14272
rect 5534 14260 5540 14272
rect 5495 14232 5540 14260
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 5994 14220 6000 14272
rect 6052 14260 6058 14272
rect 6052 14232 6097 14260
rect 6052 14220 6058 14232
rect 6178 14220 6184 14272
rect 6236 14260 6242 14272
rect 9306 14260 9312 14272
rect 6236 14232 9312 14260
rect 6236 14220 6242 14232
rect 9306 14220 9312 14232
rect 9364 14220 9370 14272
rect 9398 14220 9404 14272
rect 9456 14260 9462 14272
rect 12406 14260 12434 14300
rect 13630 14288 13636 14300
rect 13688 14288 13694 14340
rect 9456 14232 12434 14260
rect 9456 14220 9462 14232
rect 1104 14170 16008 14192
rect 1104 14118 4698 14170
rect 4750 14118 4762 14170
rect 4814 14118 4826 14170
rect 4878 14118 4890 14170
rect 4942 14118 4954 14170
rect 5006 14118 8446 14170
rect 8498 14118 8510 14170
rect 8562 14118 8574 14170
rect 8626 14118 8638 14170
rect 8690 14118 8702 14170
rect 8754 14118 12194 14170
rect 12246 14118 12258 14170
rect 12310 14118 12322 14170
rect 12374 14118 12386 14170
rect 12438 14118 12450 14170
rect 12502 14118 16008 14170
rect 1104 14096 16008 14118
rect 1486 14056 1492 14068
rect 1447 14028 1492 14056
rect 1486 14016 1492 14028
rect 1544 14016 1550 14068
rect 1946 14016 1952 14068
rect 2004 14056 2010 14068
rect 3789 14059 3847 14065
rect 3789 14056 3801 14059
rect 2004 14028 3801 14056
rect 2004 14016 2010 14028
rect 3789 14025 3801 14028
rect 3835 14025 3847 14059
rect 3789 14019 3847 14025
rect 3878 14016 3884 14068
rect 3936 14056 3942 14068
rect 5905 14059 5963 14065
rect 5905 14056 5917 14059
rect 3936 14028 5917 14056
rect 3936 14016 3942 14028
rect 5905 14025 5917 14028
rect 5951 14025 5963 14059
rect 8849 14059 8907 14065
rect 5905 14019 5963 14025
rect 6288 14028 8800 14056
rect 1673 13991 1731 13997
rect 1673 13957 1685 13991
rect 1719 13988 1731 13991
rect 2130 13988 2136 14000
rect 1719 13960 2136 13988
rect 1719 13957 1731 13960
rect 1673 13951 1731 13957
rect 2130 13948 2136 13960
rect 2188 13948 2194 14000
rect 2777 13991 2835 13997
rect 2777 13957 2789 13991
rect 2823 13988 2835 13991
rect 3418 13988 3424 14000
rect 2823 13960 3424 13988
rect 2823 13957 2835 13960
rect 2777 13951 2835 13957
rect 3418 13948 3424 13960
rect 3476 13948 3482 14000
rect 3510 13948 3516 14000
rect 3568 13988 3574 14000
rect 3605 13991 3663 13997
rect 3605 13988 3617 13991
rect 3568 13960 3617 13988
rect 3568 13948 3574 13960
rect 3605 13957 3617 13960
rect 3651 13957 3663 13991
rect 4154 13988 4160 14000
rect 4115 13960 4160 13988
rect 3605 13951 3663 13957
rect 4154 13948 4160 13960
rect 4212 13948 4218 14000
rect 4249 13991 4307 13997
rect 4249 13957 4261 13991
rect 4295 13988 4307 13991
rect 5534 13988 5540 14000
rect 4295 13960 5540 13988
rect 4295 13957 4307 13960
rect 4249 13951 4307 13957
rect 5534 13948 5540 13960
rect 5592 13948 5598 14000
rect 6288 13988 6316 14028
rect 5736 13960 6316 13988
rect 1857 13923 1915 13929
rect 1857 13889 1869 13923
rect 1903 13920 1915 13923
rect 2038 13920 2044 13932
rect 1903 13892 2044 13920
rect 1903 13889 1915 13892
rect 1857 13883 1915 13889
rect 2038 13880 2044 13892
rect 2096 13880 2102 13932
rect 2148 13920 2176 13948
rect 2406 13920 2412 13932
rect 2148 13892 2268 13920
rect 2367 13892 2412 13920
rect 1394 13812 1400 13864
rect 1452 13852 1458 13864
rect 2133 13855 2191 13861
rect 2133 13852 2145 13855
rect 1452 13824 2145 13852
rect 1452 13812 1458 13824
rect 2133 13821 2145 13824
rect 2179 13821 2191 13855
rect 2133 13815 2191 13821
rect 1854 13744 1860 13796
rect 1912 13784 1918 13796
rect 2240 13784 2268 13892
rect 2406 13880 2412 13892
rect 2464 13880 2470 13932
rect 3050 13920 3056 13932
rect 3011 13892 3056 13920
rect 3050 13880 3056 13892
rect 3108 13880 3114 13932
rect 3234 13920 3240 13932
rect 3195 13892 3240 13920
rect 3234 13880 3240 13892
rect 3292 13880 3298 13932
rect 4985 13923 5043 13929
rect 3528 13892 4476 13920
rect 3528 13864 3556 13892
rect 3326 13812 3332 13864
rect 3384 13852 3390 13864
rect 3421 13855 3479 13861
rect 3421 13852 3433 13855
rect 3384 13824 3433 13852
rect 3384 13812 3390 13824
rect 3421 13821 3433 13824
rect 3467 13821 3479 13855
rect 3421 13815 3479 13821
rect 3510 13812 3516 13864
rect 3568 13812 3574 13864
rect 4338 13852 4344 13864
rect 4299 13824 4344 13852
rect 4338 13812 4344 13824
rect 4396 13812 4402 13864
rect 4448 13852 4476 13892
rect 4985 13889 4997 13923
rect 5031 13889 5043 13923
rect 4985 13883 5043 13889
rect 5077 13923 5135 13929
rect 5077 13889 5089 13923
rect 5123 13920 5135 13923
rect 5166 13920 5172 13932
rect 5123 13892 5172 13920
rect 5123 13889 5135 13892
rect 5077 13883 5135 13889
rect 5000 13852 5028 13883
rect 5166 13880 5172 13892
rect 5224 13880 5230 13932
rect 5442 13880 5448 13932
rect 5500 13920 5506 13932
rect 5736 13920 5764 13960
rect 6362 13948 6368 14000
rect 6420 13988 6426 14000
rect 6641 13991 6699 13997
rect 6641 13988 6653 13991
rect 6420 13960 6653 13988
rect 6420 13948 6426 13960
rect 6641 13957 6653 13960
rect 6687 13957 6699 13991
rect 6641 13951 6699 13957
rect 6730 13948 6736 14000
rect 6788 13988 6794 14000
rect 8202 13988 8208 14000
rect 6788 13960 8208 13988
rect 6788 13948 6794 13960
rect 8202 13948 8208 13960
rect 8260 13988 8266 14000
rect 8481 13991 8539 13997
rect 8481 13988 8493 13991
rect 8260 13960 8493 13988
rect 8260 13948 8266 13960
rect 8481 13957 8493 13960
rect 8527 13957 8539 13991
rect 8481 13951 8539 13957
rect 5500 13892 5764 13920
rect 5813 13923 5871 13929
rect 5500 13880 5506 13892
rect 5813 13889 5825 13923
rect 5859 13889 5871 13923
rect 5813 13883 5871 13889
rect 5261 13855 5319 13861
rect 5261 13852 5273 13855
rect 4448 13824 5028 13852
rect 5184 13824 5273 13852
rect 5184 13796 5212 13824
rect 5261 13821 5273 13824
rect 5307 13821 5319 13855
rect 5261 13815 5319 13821
rect 5534 13812 5540 13864
rect 5592 13852 5598 13864
rect 5828 13852 5856 13883
rect 5902 13880 5908 13932
rect 5960 13920 5966 13932
rect 7098 13920 7104 13932
rect 5960 13892 7104 13920
rect 5960 13880 5966 13892
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 7558 13880 7564 13932
rect 7616 13920 7622 13932
rect 8662 13920 8668 13932
rect 7616 13892 8668 13920
rect 7616 13880 7622 13892
rect 8662 13880 8668 13892
rect 8720 13880 8726 13932
rect 6086 13852 6092 13864
rect 5592 13824 5856 13852
rect 6047 13824 6092 13852
rect 5592 13812 5598 13824
rect 6086 13812 6092 13824
rect 6144 13812 6150 13864
rect 7006 13812 7012 13864
rect 7064 13852 7070 13864
rect 8205 13855 8263 13861
rect 8205 13852 8217 13855
rect 7064 13824 8217 13852
rect 7064 13812 7070 13824
rect 8205 13821 8217 13824
rect 8251 13821 8263 13855
rect 8772 13852 8800 14028
rect 8849 14025 8861 14059
rect 8895 14056 8907 14059
rect 9122 14056 9128 14068
rect 8895 14028 9128 14056
rect 8895 14025 8907 14028
rect 8849 14019 8907 14025
rect 9122 14016 9128 14028
rect 9180 14016 9186 14068
rect 9217 14059 9275 14065
rect 9217 14025 9229 14059
rect 9263 14025 9275 14059
rect 9217 14019 9275 14025
rect 8938 13948 8944 14000
rect 8996 13988 9002 14000
rect 9232 13988 9260 14019
rect 9398 14016 9404 14068
rect 9456 14056 9462 14068
rect 10045 14059 10103 14065
rect 10045 14056 10057 14059
rect 9456 14028 10057 14056
rect 9456 14016 9462 14028
rect 10045 14025 10057 14028
rect 10091 14025 10103 14059
rect 10045 14019 10103 14025
rect 9861 13991 9919 13997
rect 9861 13988 9873 13991
rect 8996 13960 9260 13988
rect 9324 13960 9873 13988
rect 8996 13948 9002 13960
rect 9033 13923 9091 13929
rect 9033 13889 9045 13923
rect 9079 13920 9091 13923
rect 9324 13920 9352 13960
rect 9861 13957 9873 13960
rect 9907 13988 9919 13991
rect 10226 13988 10232 14000
rect 9907 13960 10232 13988
rect 9907 13957 9919 13960
rect 9861 13951 9919 13957
rect 10226 13948 10232 13960
rect 10284 13948 10290 14000
rect 9079 13892 9352 13920
rect 9401 13923 9459 13929
rect 9079 13889 9091 13892
rect 9033 13883 9091 13889
rect 9401 13889 9413 13923
rect 9447 13889 9459 13923
rect 9582 13920 9588 13932
rect 9543 13892 9588 13920
rect 9401 13883 9459 13889
rect 9416 13852 9444 13883
rect 9582 13880 9588 13892
rect 9640 13880 9646 13932
rect 9677 13855 9735 13861
rect 9677 13852 9689 13855
rect 8772 13824 9352 13852
rect 9416 13824 9689 13852
rect 8205 13815 8263 13821
rect 1912 13756 2268 13784
rect 1912 13744 1918 13756
rect 2682 13744 2688 13796
rect 2740 13784 2746 13796
rect 4430 13784 4436 13796
rect 2740 13756 4436 13784
rect 2740 13744 2746 13756
rect 4430 13744 4436 13756
rect 4488 13744 4494 13796
rect 5166 13744 5172 13796
rect 5224 13744 5230 13796
rect 6638 13744 6644 13796
rect 6696 13744 6702 13796
rect 7190 13744 7196 13796
rect 7248 13784 7254 13796
rect 9122 13784 9128 13796
rect 7248 13756 9128 13784
rect 7248 13744 7254 13756
rect 9122 13744 9128 13756
rect 9180 13744 9186 13796
rect 9324 13784 9352 13824
rect 9677 13821 9689 13824
rect 9723 13852 9735 13855
rect 9766 13852 9772 13864
rect 9723 13824 9772 13852
rect 9723 13821 9735 13824
rect 9677 13815 9735 13821
rect 9766 13812 9772 13824
rect 9824 13812 9830 13864
rect 10042 13812 10048 13864
rect 10100 13852 10106 13864
rect 15470 13852 15476 13864
rect 10100 13824 15476 13852
rect 10100 13812 10106 13824
rect 15470 13812 15476 13824
rect 15528 13812 15534 13864
rect 9582 13784 9588 13796
rect 9324 13756 9588 13784
rect 9582 13744 9588 13756
rect 9640 13744 9646 13796
rect 10134 13744 10140 13796
rect 10192 13784 10198 13796
rect 11146 13784 11152 13796
rect 10192 13756 11152 13784
rect 10192 13744 10198 13756
rect 11146 13744 11152 13756
rect 11204 13744 11210 13796
rect 4522 13676 4528 13728
rect 4580 13716 4586 13728
rect 4617 13719 4675 13725
rect 4617 13716 4629 13719
rect 4580 13688 4629 13716
rect 4580 13676 4586 13688
rect 4617 13685 4629 13688
rect 4663 13685 4675 13719
rect 4617 13679 4675 13685
rect 4890 13676 4896 13728
rect 4948 13716 4954 13728
rect 5445 13719 5503 13725
rect 5445 13716 5457 13719
rect 4948 13688 5457 13716
rect 4948 13676 4954 13688
rect 5445 13685 5457 13688
rect 5491 13685 5503 13719
rect 5445 13679 5503 13685
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 6457 13719 6515 13725
rect 6457 13716 6469 13719
rect 6420 13688 6469 13716
rect 6420 13676 6426 13688
rect 6457 13685 6469 13688
rect 6503 13685 6515 13719
rect 6656 13716 6684 13744
rect 8938 13716 8944 13728
rect 6656 13688 8944 13716
rect 6457 13679 6515 13685
rect 8938 13676 8944 13688
rect 8996 13716 9002 13728
rect 13262 13716 13268 13728
rect 8996 13688 13268 13716
rect 8996 13676 9002 13688
rect 13262 13676 13268 13688
rect 13320 13676 13326 13728
rect 1104 13626 16008 13648
rect 1104 13574 2824 13626
rect 2876 13574 2888 13626
rect 2940 13574 2952 13626
rect 3004 13574 3016 13626
rect 3068 13574 3080 13626
rect 3132 13574 6572 13626
rect 6624 13574 6636 13626
rect 6688 13574 6700 13626
rect 6752 13574 6764 13626
rect 6816 13574 6828 13626
rect 6880 13574 10320 13626
rect 10372 13574 10384 13626
rect 10436 13574 10448 13626
rect 10500 13574 10512 13626
rect 10564 13574 10576 13626
rect 10628 13574 14068 13626
rect 14120 13574 14132 13626
rect 14184 13574 14196 13626
rect 14248 13574 14260 13626
rect 14312 13574 14324 13626
rect 14376 13574 16008 13626
rect 1104 13552 16008 13574
rect 2682 13512 2688 13524
rect 2643 13484 2688 13512
rect 2682 13472 2688 13484
rect 2740 13472 2746 13524
rect 3602 13472 3608 13524
rect 3660 13512 3666 13524
rect 3789 13515 3847 13521
rect 3789 13512 3801 13515
rect 3660 13484 3801 13512
rect 3660 13472 3666 13484
rect 3789 13481 3801 13484
rect 3835 13481 3847 13515
rect 3789 13475 3847 13481
rect 4430 13472 4436 13524
rect 4488 13512 4494 13524
rect 4801 13515 4859 13521
rect 4801 13512 4813 13515
rect 4488 13484 4813 13512
rect 4488 13472 4494 13484
rect 4801 13481 4813 13484
rect 4847 13512 4859 13515
rect 5994 13512 6000 13524
rect 4847 13484 6000 13512
rect 4847 13481 4859 13484
rect 4801 13475 4859 13481
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 6457 13515 6515 13521
rect 6457 13481 6469 13515
rect 6503 13512 6515 13515
rect 7098 13512 7104 13524
rect 6503 13484 7104 13512
rect 6503 13481 6515 13484
rect 6457 13475 6515 13481
rect 7098 13472 7104 13484
rect 7156 13472 7162 13524
rect 8294 13472 8300 13524
rect 8352 13512 8358 13524
rect 8573 13515 8631 13521
rect 8573 13512 8585 13515
rect 8352 13484 8585 13512
rect 8352 13472 8358 13484
rect 8573 13481 8585 13484
rect 8619 13481 8631 13515
rect 8573 13475 8631 13481
rect 9030 13472 9036 13524
rect 9088 13512 9094 13524
rect 9490 13512 9496 13524
rect 9088 13484 9133 13512
rect 9451 13484 9496 13512
rect 9088 13472 9094 13484
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 9582 13472 9588 13524
rect 9640 13512 9646 13524
rect 10042 13512 10048 13524
rect 9640 13484 10048 13512
rect 9640 13472 9646 13484
rect 10042 13472 10048 13484
rect 10100 13472 10106 13524
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 10505 13515 10563 13521
rect 10505 13512 10517 13515
rect 10192 13484 10517 13512
rect 10192 13472 10198 13484
rect 10505 13481 10517 13484
rect 10551 13481 10563 13515
rect 10686 13512 10692 13524
rect 10647 13484 10692 13512
rect 10505 13475 10563 13481
rect 10686 13472 10692 13484
rect 10744 13512 10750 13524
rect 11514 13512 11520 13524
rect 10744 13484 11520 13512
rect 10744 13472 10750 13484
rect 11514 13472 11520 13484
rect 11572 13472 11578 13524
rect 9214 13444 9220 13456
rect 1964 13416 4568 13444
rect 1670 13376 1676 13388
rect 1631 13348 1676 13376
rect 1670 13336 1676 13348
rect 1728 13336 1734 13388
rect 1964 13317 1992 13416
rect 3418 13336 3424 13388
rect 3476 13376 3482 13388
rect 3513 13379 3571 13385
rect 3513 13376 3525 13379
rect 3476 13348 3525 13376
rect 3476 13336 3482 13348
rect 3513 13345 3525 13348
rect 3559 13376 3571 13379
rect 3786 13376 3792 13388
rect 3559 13348 3792 13376
rect 3559 13345 3571 13348
rect 3513 13339 3571 13345
rect 3786 13336 3792 13348
rect 3844 13336 3850 13388
rect 4430 13376 4436 13388
rect 4391 13348 4436 13376
rect 4430 13336 4436 13348
rect 4488 13336 4494 13388
rect 4540 13376 4568 13416
rect 5736 13416 9220 13444
rect 4890 13376 4896 13388
rect 4540 13348 4896 13376
rect 4890 13336 4896 13348
rect 4948 13336 4954 13388
rect 5258 13336 5264 13388
rect 5316 13376 5322 13388
rect 5445 13379 5503 13385
rect 5445 13376 5457 13379
rect 5316 13348 5457 13376
rect 5316 13336 5322 13348
rect 5445 13345 5457 13348
rect 5491 13345 5503 13379
rect 5445 13339 5503 13345
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13277 2007 13311
rect 1949 13271 2007 13277
rect 2501 13311 2559 13317
rect 2501 13277 2513 13311
rect 2547 13308 2559 13311
rect 3234 13308 3240 13320
rect 2547 13280 3240 13308
rect 2547 13277 2559 13280
rect 2501 13271 2559 13277
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 3329 13311 3387 13317
rect 3329 13277 3341 13311
rect 3375 13308 3387 13311
rect 5736 13308 5764 13416
rect 9214 13404 9220 13416
rect 9272 13404 9278 13456
rect 9950 13404 9956 13456
rect 10008 13444 10014 13456
rect 10229 13447 10287 13453
rect 10229 13444 10241 13447
rect 10008 13416 10241 13444
rect 10008 13404 10014 13416
rect 10229 13413 10241 13416
rect 10275 13413 10287 13447
rect 10229 13407 10287 13413
rect 5905 13379 5963 13385
rect 5905 13345 5917 13379
rect 5951 13376 5963 13379
rect 6546 13376 6552 13388
rect 5951 13348 6552 13376
rect 5951 13345 5963 13348
rect 5905 13339 5963 13345
rect 6546 13336 6552 13348
rect 6604 13336 6610 13388
rect 6733 13379 6791 13385
rect 6733 13345 6745 13379
rect 6779 13376 6791 13379
rect 7374 13376 7380 13388
rect 6779 13348 7380 13376
rect 6779 13345 6791 13348
rect 6733 13339 6791 13345
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 7558 13376 7564 13388
rect 7519 13348 7564 13376
rect 7558 13336 7564 13348
rect 7616 13336 7622 13388
rect 7834 13376 7840 13388
rect 7760 13348 7840 13376
rect 3375 13280 5764 13308
rect 3375 13277 3387 13280
rect 3329 13271 3387 13277
rect 5810 13268 5816 13320
rect 5868 13308 5874 13320
rect 6089 13311 6147 13317
rect 6089 13308 6101 13311
rect 5868 13280 6101 13308
rect 5868 13268 5874 13280
rect 6089 13277 6101 13280
rect 6135 13277 6147 13311
rect 6914 13308 6920 13320
rect 6875 13280 6920 13308
rect 6089 13271 6147 13277
rect 6914 13268 6920 13280
rect 6972 13268 6978 13320
rect 7760 13317 7788 13348
rect 7834 13336 7840 13348
rect 7892 13336 7898 13388
rect 7926 13336 7932 13388
rect 7984 13376 7990 13388
rect 8294 13376 8300 13388
rect 7984 13348 8300 13376
rect 7984 13336 7990 13348
rect 8294 13336 8300 13348
rect 8352 13336 8358 13388
rect 11330 13376 11336 13388
rect 8680 13348 11336 13376
rect 7745 13311 7803 13317
rect 7745 13277 7757 13311
rect 7791 13277 7803 13311
rect 7745 13271 7803 13277
rect 2222 13240 2228 13252
rect 2183 13212 2228 13240
rect 2222 13200 2228 13212
rect 2280 13200 2286 13252
rect 4249 13243 4307 13249
rect 4249 13209 4261 13243
rect 4295 13240 4307 13243
rect 5353 13243 5411 13249
rect 4295 13212 4936 13240
rect 4295 13209 4307 13212
rect 4249 13203 4307 13209
rect 2682 13132 2688 13184
rect 2740 13172 2746 13184
rect 2869 13175 2927 13181
rect 2869 13172 2881 13175
rect 2740 13144 2881 13172
rect 2740 13132 2746 13144
rect 2869 13141 2881 13144
rect 2915 13141 2927 13175
rect 2869 13135 2927 13141
rect 3237 13175 3295 13181
rect 3237 13141 3249 13175
rect 3283 13172 3295 13175
rect 3326 13172 3332 13184
rect 3283 13144 3332 13172
rect 3283 13141 3295 13144
rect 3237 13135 3295 13141
rect 3326 13132 3332 13144
rect 3384 13132 3390 13184
rect 4157 13175 4215 13181
rect 4157 13141 4169 13175
rect 4203 13172 4215 13175
rect 4614 13172 4620 13184
rect 4203 13144 4620 13172
rect 4203 13141 4215 13144
rect 4157 13135 4215 13141
rect 4614 13132 4620 13144
rect 4672 13132 4678 13184
rect 4908 13181 4936 13212
rect 5353 13209 5365 13243
rect 5399 13240 5411 13243
rect 6730 13240 6736 13252
rect 5399 13212 6736 13240
rect 5399 13209 5411 13212
rect 5353 13203 5411 13209
rect 6730 13200 6736 13212
rect 6788 13200 6794 13252
rect 6825 13243 6883 13249
rect 6825 13209 6837 13243
rect 6871 13240 6883 13243
rect 7834 13240 7840 13252
rect 6871 13212 7840 13240
rect 6871 13209 6883 13212
rect 6825 13203 6883 13209
rect 7834 13200 7840 13212
rect 7892 13200 7898 13252
rect 7926 13200 7932 13252
rect 7984 13240 7990 13252
rect 8205 13243 8263 13249
rect 8205 13240 8217 13243
rect 7984 13212 8217 13240
rect 7984 13200 7990 13212
rect 8205 13209 8217 13212
rect 8251 13209 8263 13243
rect 8205 13203 8263 13209
rect 4893 13175 4951 13181
rect 4893 13141 4905 13175
rect 4939 13141 4951 13175
rect 4893 13135 4951 13141
rect 5261 13175 5319 13181
rect 5261 13141 5273 13175
rect 5307 13172 5319 13175
rect 5442 13172 5448 13184
rect 5307 13144 5448 13172
rect 5307 13141 5319 13144
rect 5261 13135 5319 13141
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 5997 13175 6055 13181
rect 5997 13141 6009 13175
rect 6043 13172 6055 13175
rect 7098 13172 7104 13184
rect 6043 13144 7104 13172
rect 6043 13141 6055 13144
rect 5997 13135 6055 13141
rect 7098 13132 7104 13144
rect 7156 13132 7162 13184
rect 7190 13132 7196 13184
rect 7248 13172 7254 13184
rect 7285 13175 7343 13181
rect 7285 13172 7297 13175
rect 7248 13144 7297 13172
rect 7248 13132 7254 13144
rect 7285 13141 7297 13144
rect 7331 13141 7343 13175
rect 7285 13135 7343 13141
rect 7653 13175 7711 13181
rect 7653 13141 7665 13175
rect 7699 13172 7711 13175
rect 7742 13172 7748 13184
rect 7699 13144 7748 13172
rect 7699 13141 7711 13144
rect 7653 13135 7711 13141
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 8113 13175 8171 13181
rect 8113 13141 8125 13175
rect 8159 13172 8171 13175
rect 8680 13172 8708 13348
rect 11330 13336 11336 13348
rect 11388 13336 11394 13388
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13277 8815 13311
rect 8757 13271 8815 13277
rect 9217 13311 9275 13317
rect 9217 13277 9229 13311
rect 9263 13308 9275 13311
rect 9398 13308 9404 13320
rect 9263 13280 9404 13308
rect 9263 13277 9275 13280
rect 9217 13271 9275 13277
rect 8772 13240 8800 13271
rect 9398 13268 9404 13280
rect 9456 13268 9462 13320
rect 9677 13311 9735 13317
rect 9677 13277 9689 13311
rect 9723 13308 9735 13311
rect 10045 13311 10103 13317
rect 10045 13308 10057 13311
rect 9723 13280 10057 13308
rect 9723 13277 9735 13280
rect 9677 13271 9735 13277
rect 10045 13277 10057 13280
rect 10091 13308 10103 13311
rect 10778 13308 10784 13320
rect 10091 13280 10784 13308
rect 10091 13277 10103 13280
rect 10045 13271 10103 13277
rect 10778 13268 10784 13280
rect 10836 13268 10842 13320
rect 10870 13268 10876 13320
rect 10928 13308 10934 13320
rect 10928 13280 10973 13308
rect 10928 13268 10934 13280
rect 10413 13243 10471 13249
rect 10413 13240 10425 13243
rect 8772 13212 10425 13240
rect 10413 13209 10425 13212
rect 10459 13240 10471 13243
rect 11238 13240 11244 13252
rect 10459 13212 11244 13240
rect 10459 13209 10471 13212
rect 10413 13203 10471 13209
rect 11238 13200 11244 13212
rect 11296 13200 11302 13252
rect 11606 13200 11612 13252
rect 11664 13240 11670 13252
rect 14826 13240 14832 13252
rect 11664 13212 14832 13240
rect 11664 13200 11670 13212
rect 14826 13200 14832 13212
rect 14884 13200 14890 13252
rect 8159 13144 8708 13172
rect 8159 13141 8171 13144
rect 8113 13135 8171 13141
rect 9582 13132 9588 13184
rect 9640 13172 9646 13184
rect 9769 13175 9827 13181
rect 9769 13172 9781 13175
rect 9640 13144 9781 13172
rect 9640 13132 9646 13144
rect 9769 13141 9781 13144
rect 9815 13172 9827 13175
rect 10594 13172 10600 13184
rect 9815 13144 10600 13172
rect 9815 13141 9827 13144
rect 9769 13135 9827 13141
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 10686 13132 10692 13184
rect 10744 13172 10750 13184
rect 13170 13172 13176 13184
rect 10744 13144 13176 13172
rect 10744 13132 10750 13144
rect 13170 13132 13176 13144
rect 13228 13132 13234 13184
rect 1104 13082 16008 13104
rect 1104 13030 4698 13082
rect 4750 13030 4762 13082
rect 4814 13030 4826 13082
rect 4878 13030 4890 13082
rect 4942 13030 4954 13082
rect 5006 13030 8446 13082
rect 8498 13030 8510 13082
rect 8562 13030 8574 13082
rect 8626 13030 8638 13082
rect 8690 13030 8702 13082
rect 8754 13030 12194 13082
rect 12246 13030 12258 13082
rect 12310 13030 12322 13082
rect 12374 13030 12386 13082
rect 12438 13030 12450 13082
rect 12502 13030 16008 13082
rect 1104 13008 16008 13030
rect 1673 12971 1731 12977
rect 1673 12937 1685 12971
rect 1719 12968 1731 12971
rect 1762 12968 1768 12980
rect 1719 12940 1768 12968
rect 1719 12937 1731 12940
rect 1673 12931 1731 12937
rect 1762 12928 1768 12940
rect 1820 12928 1826 12980
rect 2130 12968 2136 12980
rect 2091 12940 2136 12968
rect 2130 12928 2136 12940
rect 2188 12928 2194 12980
rect 2314 12968 2320 12980
rect 2275 12940 2320 12968
rect 2314 12928 2320 12940
rect 2372 12928 2378 12980
rect 2958 12928 2964 12980
rect 3016 12968 3022 12980
rect 3053 12971 3111 12977
rect 3053 12968 3065 12971
rect 3016 12940 3065 12968
rect 3016 12928 3022 12940
rect 3053 12937 3065 12940
rect 3099 12968 3111 12971
rect 3786 12968 3792 12980
rect 3099 12940 3792 12968
rect 3099 12937 3111 12940
rect 3053 12931 3111 12937
rect 3786 12928 3792 12940
rect 3844 12928 3850 12980
rect 4614 12968 4620 12980
rect 4575 12940 4620 12968
rect 4614 12928 4620 12940
rect 4672 12928 4678 12980
rect 5721 12971 5779 12977
rect 5721 12937 5733 12971
rect 5767 12968 5779 12971
rect 5994 12968 6000 12980
rect 5767 12940 6000 12968
rect 5767 12937 5779 12940
rect 5721 12931 5779 12937
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 6454 12928 6460 12980
rect 6512 12968 6518 12980
rect 6549 12971 6607 12977
rect 6549 12968 6561 12971
rect 6512 12940 6561 12968
rect 6512 12928 6518 12940
rect 6549 12937 6561 12940
rect 6595 12937 6607 12971
rect 6549 12931 6607 12937
rect 6730 12928 6736 12980
rect 6788 12968 6794 12980
rect 8481 12971 8539 12977
rect 8481 12968 8493 12971
rect 6788 12940 8493 12968
rect 6788 12928 6794 12940
rect 8481 12937 8493 12940
rect 8527 12937 8539 12971
rect 8481 12931 8539 12937
rect 9214 12928 9220 12980
rect 9272 12968 9278 12980
rect 9309 12971 9367 12977
rect 9309 12968 9321 12971
rect 9272 12940 9321 12968
rect 9272 12928 9278 12940
rect 9309 12937 9321 12940
rect 9355 12937 9367 12971
rect 9309 12931 9367 12937
rect 9582 12928 9588 12980
rect 9640 12968 9646 12980
rect 9677 12971 9735 12977
rect 9677 12968 9689 12971
rect 9640 12940 9689 12968
rect 9640 12928 9646 12940
rect 9677 12937 9689 12940
rect 9723 12937 9735 12971
rect 11606 12968 11612 12980
rect 9677 12931 9735 12937
rect 9784 12940 11612 12968
rect 2332 12900 2360 12928
rect 7006 12900 7012 12912
rect 1596 12872 2360 12900
rect 4356 12872 7012 12900
rect 1596 12773 1624 12872
rect 1762 12832 1768 12844
rect 1723 12804 1768 12832
rect 1762 12792 1768 12804
rect 1820 12792 1826 12844
rect 4356 12841 4384 12872
rect 7006 12860 7012 12872
rect 7064 12860 7070 12912
rect 9784 12909 9812 12940
rect 11606 12928 11612 12940
rect 11664 12928 11670 12980
rect 11790 12928 11796 12980
rect 11848 12968 11854 12980
rect 15838 12968 15844 12980
rect 11848 12940 15844 12968
rect 11848 12928 11854 12940
rect 15838 12928 15844 12940
rect 15896 12928 15902 12980
rect 7285 12903 7343 12909
rect 7285 12869 7297 12903
rect 7331 12900 7343 12903
rect 9769 12903 9827 12909
rect 7331 12872 9720 12900
rect 7331 12869 7343 12872
rect 7285 12863 7343 12869
rect 4341 12835 4399 12841
rect 4341 12801 4353 12835
rect 4387 12801 4399 12835
rect 4982 12832 4988 12844
rect 4943 12804 4988 12832
rect 4341 12795 4399 12801
rect 4982 12792 4988 12804
rect 5040 12792 5046 12844
rect 5077 12835 5135 12841
rect 5077 12801 5089 12835
rect 5123 12832 5135 12835
rect 5442 12832 5448 12844
rect 5123 12804 5448 12832
rect 5123 12801 5135 12804
rect 5077 12795 5135 12801
rect 5442 12792 5448 12804
rect 5500 12792 5506 12844
rect 5813 12835 5871 12841
rect 5813 12801 5825 12835
rect 5859 12832 5871 12835
rect 5902 12832 5908 12844
rect 5859 12804 5908 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 1581 12767 1639 12773
rect 1581 12733 1593 12767
rect 1627 12733 1639 12767
rect 5258 12764 5264 12776
rect 5219 12736 5264 12764
rect 1581 12727 1639 12733
rect 5258 12724 5264 12736
rect 5316 12724 5322 12776
rect 5629 12767 5687 12773
rect 5629 12733 5641 12767
rect 5675 12764 5687 12767
rect 5718 12764 5724 12776
rect 5675 12736 5724 12764
rect 5675 12733 5687 12736
rect 5629 12727 5687 12733
rect 5718 12724 5724 12736
rect 5776 12724 5782 12776
rect 4246 12656 4252 12708
rect 4304 12696 4310 12708
rect 5166 12696 5172 12708
rect 4304 12668 5172 12696
rect 4304 12656 4310 12668
rect 5166 12656 5172 12668
rect 5224 12656 5230 12708
rect 2498 12628 2504 12640
rect 2411 12600 2504 12628
rect 2498 12588 2504 12600
rect 2556 12628 2562 12640
rect 4525 12631 4583 12637
rect 4525 12628 4537 12631
rect 2556 12600 4537 12628
rect 2556 12588 2562 12600
rect 4525 12597 4537 12600
rect 4571 12628 4583 12631
rect 5828 12628 5856 12795
rect 5902 12792 5908 12804
rect 5960 12792 5966 12844
rect 6362 12792 6368 12844
rect 6420 12832 6426 12844
rect 6733 12835 6791 12841
rect 6733 12832 6745 12835
rect 6420 12804 6745 12832
rect 6420 12792 6426 12804
rect 6733 12801 6745 12804
rect 6779 12801 6791 12835
rect 6733 12795 6791 12801
rect 7193 12835 7251 12841
rect 7193 12801 7205 12835
rect 7239 12832 7251 12835
rect 8018 12832 8024 12844
rect 7239 12804 7880 12832
rect 7979 12804 8024 12832
rect 7239 12801 7251 12804
rect 7193 12795 7251 12801
rect 7466 12764 7472 12776
rect 5920 12736 7472 12764
rect 5920 12708 5948 12736
rect 7466 12724 7472 12736
rect 7524 12724 7530 12776
rect 7742 12764 7748 12776
rect 7703 12736 7748 12764
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 5902 12656 5908 12708
rect 5960 12656 5966 12708
rect 6181 12699 6239 12705
rect 6181 12665 6193 12699
rect 6227 12696 6239 12699
rect 7190 12696 7196 12708
rect 6227 12668 7196 12696
rect 6227 12665 6239 12668
rect 6181 12659 6239 12665
rect 7190 12656 7196 12668
rect 7248 12656 7254 12708
rect 4571 12600 5856 12628
rect 4571 12597 4583 12600
rect 4525 12591 4583 12597
rect 6270 12588 6276 12640
rect 6328 12628 6334 12640
rect 6825 12631 6883 12637
rect 6825 12628 6837 12631
rect 6328 12600 6837 12628
rect 6328 12588 6334 12600
rect 6825 12597 6837 12600
rect 6871 12597 6883 12631
rect 7852 12628 7880 12804
rect 8018 12792 8024 12804
rect 8076 12792 8082 12844
rect 8294 12792 8300 12844
rect 8352 12832 8358 12844
rect 8849 12835 8907 12841
rect 8352 12804 8708 12832
rect 8352 12792 8358 12804
rect 7929 12767 7987 12773
rect 7929 12733 7941 12767
rect 7975 12764 7987 12767
rect 8202 12764 8208 12776
rect 7975 12736 8208 12764
rect 7975 12733 7987 12736
rect 7929 12727 7987 12733
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 8294 12656 8300 12708
rect 8352 12696 8358 12708
rect 8389 12699 8447 12705
rect 8389 12696 8401 12699
rect 8352 12668 8401 12696
rect 8352 12656 8358 12668
rect 8389 12665 8401 12668
rect 8435 12665 8447 12699
rect 8680 12696 8708 12804
rect 8849 12801 8861 12835
rect 8895 12832 8907 12835
rect 9490 12832 9496 12844
rect 8895 12804 9496 12832
rect 8895 12801 8907 12804
rect 8849 12795 8907 12801
rect 9490 12792 9496 12804
rect 9548 12792 9554 12844
rect 9692 12832 9720 12872
rect 9769 12869 9781 12903
rect 9815 12869 9827 12903
rect 9769 12863 9827 12869
rect 9858 12860 9864 12912
rect 9916 12900 9922 12912
rect 10226 12900 10232 12912
rect 9916 12872 10232 12900
rect 9916 12860 9922 12872
rect 10226 12860 10232 12872
rect 10284 12860 10290 12912
rect 10594 12900 10600 12912
rect 10555 12872 10600 12900
rect 10594 12860 10600 12872
rect 10652 12860 10658 12912
rect 10873 12903 10931 12909
rect 10873 12900 10885 12903
rect 10695 12872 10885 12900
rect 10695 12832 10723 12872
rect 10873 12869 10885 12872
rect 10919 12900 10931 12903
rect 16206 12900 16212 12912
rect 10919 12872 16212 12900
rect 10919 12869 10931 12872
rect 10873 12863 10931 12869
rect 16206 12860 16212 12872
rect 16264 12860 16270 12912
rect 9692 12804 10723 12832
rect 10781 12835 10839 12841
rect 10781 12801 10793 12835
rect 10827 12832 10839 12835
rect 11146 12832 11152 12844
rect 10827 12804 11152 12832
rect 10827 12801 10839 12804
rect 10781 12795 10839 12801
rect 11146 12792 11152 12804
rect 11204 12832 11210 12844
rect 11204 12804 12020 12832
rect 11204 12792 11210 12804
rect 8754 12724 8760 12776
rect 8812 12764 8818 12776
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 8812 12736 8953 12764
rect 8812 12724 8818 12736
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 9030 12724 9036 12776
rect 9088 12764 9094 12776
rect 9858 12764 9864 12776
rect 9088 12736 9133 12764
rect 9819 12736 9864 12764
rect 9088 12724 9094 12736
rect 9858 12724 9864 12736
rect 9916 12724 9922 12776
rect 10686 12764 10692 12776
rect 10520 12736 10692 12764
rect 9214 12696 9220 12708
rect 8680 12668 9220 12696
rect 8389 12659 8447 12665
rect 9214 12656 9220 12668
rect 9272 12696 9278 12708
rect 10137 12699 10195 12705
rect 10137 12696 10149 12699
rect 9272 12668 10149 12696
rect 9272 12656 9278 12668
rect 10137 12665 10149 12668
rect 10183 12696 10195 12699
rect 10520 12696 10548 12736
rect 10686 12724 10692 12736
rect 10744 12724 10750 12776
rect 10962 12724 10968 12776
rect 11020 12764 11026 12776
rect 11057 12767 11115 12773
rect 11057 12764 11069 12767
rect 11020 12736 11069 12764
rect 11020 12724 11026 12736
rect 11057 12733 11069 12736
rect 11103 12733 11115 12767
rect 11057 12727 11115 12733
rect 10183 12668 10548 12696
rect 11333 12699 11391 12705
rect 10183 12665 10195 12668
rect 10137 12659 10195 12665
rect 11333 12665 11345 12699
rect 11379 12696 11391 12699
rect 11514 12696 11520 12708
rect 11379 12668 11520 12696
rect 11379 12665 11391 12668
rect 11333 12659 11391 12665
rect 11514 12656 11520 12668
rect 11572 12656 11578 12708
rect 11609 12699 11667 12705
rect 11609 12665 11621 12699
rect 11655 12696 11667 12699
rect 11698 12696 11704 12708
rect 11655 12668 11704 12696
rect 11655 12665 11667 12668
rect 11609 12659 11667 12665
rect 11698 12656 11704 12668
rect 11756 12656 11762 12708
rect 11790 12656 11796 12708
rect 11848 12696 11854 12708
rect 11992 12705 12020 12804
rect 11977 12699 12035 12705
rect 11848 12668 11893 12696
rect 11848 12656 11854 12668
rect 11977 12665 11989 12699
rect 12023 12696 12035 12699
rect 12526 12696 12532 12708
rect 12023 12668 12532 12696
rect 12023 12665 12035 12668
rect 11977 12659 12035 12665
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 9582 12628 9588 12640
rect 7852 12600 9588 12628
rect 6825 12591 6883 12597
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 9766 12588 9772 12640
rect 9824 12628 9830 12640
rect 10321 12631 10379 12637
rect 10321 12628 10333 12631
rect 9824 12600 10333 12628
rect 9824 12588 9830 12600
rect 10321 12597 10333 12600
rect 10367 12597 10379 12631
rect 10321 12591 10379 12597
rect 10686 12588 10692 12640
rect 10744 12628 10750 12640
rect 12342 12628 12348 12640
rect 10744 12600 12348 12628
rect 10744 12588 10750 12600
rect 12342 12588 12348 12600
rect 12400 12588 12406 12640
rect 1104 12538 16008 12560
rect 1104 12486 2824 12538
rect 2876 12486 2888 12538
rect 2940 12486 2952 12538
rect 3004 12486 3016 12538
rect 3068 12486 3080 12538
rect 3132 12486 6572 12538
rect 6624 12486 6636 12538
rect 6688 12486 6700 12538
rect 6752 12486 6764 12538
rect 6816 12486 6828 12538
rect 6880 12486 10320 12538
rect 10372 12486 10384 12538
rect 10436 12486 10448 12538
rect 10500 12486 10512 12538
rect 10564 12486 10576 12538
rect 10628 12486 14068 12538
rect 14120 12486 14132 12538
rect 14184 12486 14196 12538
rect 14248 12486 14260 12538
rect 14312 12486 14324 12538
rect 14376 12486 16008 12538
rect 1104 12464 16008 12486
rect 2869 12427 2927 12433
rect 2869 12393 2881 12427
rect 2915 12424 2927 12427
rect 3234 12424 3240 12436
rect 2915 12396 3240 12424
rect 2915 12393 2927 12396
rect 2869 12387 2927 12393
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 5074 12384 5080 12436
rect 5132 12424 5138 12436
rect 5261 12427 5319 12433
rect 5261 12424 5273 12427
rect 5132 12396 5273 12424
rect 5132 12384 5138 12396
rect 5261 12393 5273 12396
rect 5307 12393 5319 12427
rect 5261 12387 5319 12393
rect 5368 12396 6960 12424
rect 2774 12316 2780 12368
rect 2832 12356 2838 12368
rect 5368 12356 5396 12396
rect 2832 12328 5396 12356
rect 5537 12359 5595 12365
rect 2832 12316 2838 12328
rect 5537 12325 5549 12359
rect 5583 12356 5595 12359
rect 5626 12356 5632 12368
rect 5583 12328 5632 12356
rect 5583 12325 5595 12328
rect 5537 12319 5595 12325
rect 5626 12316 5632 12328
rect 5684 12316 5690 12368
rect 1578 12248 1584 12300
rect 1636 12288 1642 12300
rect 1673 12291 1731 12297
rect 1673 12288 1685 12291
rect 1636 12260 1685 12288
rect 1636 12248 1642 12260
rect 1673 12257 1685 12260
rect 1719 12257 1731 12291
rect 2222 12288 2228 12300
rect 2183 12260 2228 12288
rect 1673 12251 1731 12257
rect 2222 12248 2228 12260
rect 2280 12248 2286 12300
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12288 2375 12291
rect 2682 12288 2688 12300
rect 2363 12260 2688 12288
rect 2363 12257 2375 12260
rect 2317 12251 2375 12257
rect 2682 12248 2688 12260
rect 2740 12248 2746 12300
rect 3050 12248 3056 12300
rect 3108 12288 3114 12300
rect 3329 12291 3387 12297
rect 3329 12288 3341 12291
rect 3108 12260 3341 12288
rect 3108 12248 3114 12260
rect 3329 12257 3341 12260
rect 3375 12257 3387 12291
rect 3329 12251 3387 12257
rect 3418 12248 3424 12300
rect 3476 12288 3482 12300
rect 3970 12288 3976 12300
rect 3476 12260 3521 12288
rect 3620 12260 3976 12288
rect 3476 12248 3482 12260
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12189 2007 12223
rect 1949 12183 2007 12189
rect 2409 12223 2467 12229
rect 2409 12189 2421 12223
rect 2455 12220 2467 12223
rect 3620 12220 3648 12260
rect 3970 12248 3976 12260
rect 4028 12248 4034 12300
rect 6932 12288 6960 12396
rect 7190 12384 7196 12436
rect 7248 12424 7254 12436
rect 7248 12396 7972 12424
rect 7248 12384 7254 12396
rect 7944 12356 7972 12396
rect 8018 12384 8024 12436
rect 8076 12424 8082 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 8076 12396 8585 12424
rect 8076 12384 8082 12396
rect 8573 12393 8585 12396
rect 8619 12393 8631 12427
rect 9398 12424 9404 12436
rect 8573 12387 8631 12393
rect 8680 12396 9404 12424
rect 8680 12356 8708 12396
rect 9398 12384 9404 12396
rect 9456 12384 9462 12436
rect 9490 12384 9496 12436
rect 9548 12424 9554 12436
rect 9769 12427 9827 12433
rect 9769 12424 9781 12427
rect 9548 12396 9781 12424
rect 9548 12384 9554 12396
rect 9769 12393 9781 12396
rect 9815 12393 9827 12427
rect 9769 12387 9827 12393
rect 11425 12427 11483 12433
rect 11425 12393 11437 12427
rect 11471 12424 11483 12427
rect 11790 12424 11796 12436
rect 11471 12396 11796 12424
rect 11471 12393 11483 12396
rect 11425 12387 11483 12393
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 11974 12424 11980 12436
rect 11935 12396 11980 12424
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 12434 12424 12440 12436
rect 12268 12396 12440 12424
rect 7944 12328 8708 12356
rect 8938 12316 8944 12368
rect 8996 12356 9002 12368
rect 10686 12356 10692 12368
rect 8996 12328 10692 12356
rect 8996 12316 9002 12328
rect 10686 12316 10692 12328
rect 10744 12356 10750 12368
rect 10781 12359 10839 12365
rect 10781 12356 10793 12359
rect 10744 12328 10793 12356
rect 10744 12316 10750 12328
rect 10781 12325 10793 12328
rect 10827 12325 10839 12359
rect 10781 12319 10839 12325
rect 10870 12316 10876 12368
rect 10928 12356 10934 12368
rect 10928 12328 11284 12356
rect 10928 12316 10934 12328
rect 9493 12291 9551 12297
rect 9493 12288 9505 12291
rect 5368 12260 5948 12288
rect 6932 12260 7144 12288
rect 3786 12220 3792 12232
rect 2455 12192 3648 12220
rect 3747 12192 3792 12220
rect 2455 12189 2467 12192
rect 2409 12183 2467 12189
rect 1964 12152 1992 12183
rect 3786 12180 3792 12192
rect 3844 12180 3850 12232
rect 4522 12220 4528 12232
rect 3896 12192 4528 12220
rect 3896 12152 3924 12192
rect 4522 12180 4528 12192
rect 4580 12180 4586 12232
rect 4617 12223 4675 12229
rect 4617 12189 4629 12223
rect 4663 12220 4675 12223
rect 5074 12220 5080 12232
rect 4663 12192 5080 12220
rect 4663 12189 4675 12192
rect 4617 12183 4675 12189
rect 5074 12180 5080 12192
rect 5132 12180 5138 12232
rect 1964 12124 3924 12152
rect 658 12044 664 12096
rect 716 12084 722 12096
rect 1118 12084 1124 12096
rect 716 12056 1124 12084
rect 716 12044 722 12056
rect 1118 12044 1124 12056
rect 1176 12044 1182 12096
rect 2777 12087 2835 12093
rect 2777 12053 2789 12087
rect 2823 12084 2835 12087
rect 3142 12084 3148 12096
rect 2823 12056 3148 12084
rect 2823 12053 2835 12056
rect 2777 12047 2835 12053
rect 3142 12044 3148 12056
rect 3200 12044 3206 12096
rect 3237 12087 3295 12093
rect 3237 12053 3249 12087
rect 3283 12084 3295 12087
rect 3602 12084 3608 12096
rect 3283 12056 3608 12084
rect 3283 12053 3295 12056
rect 3237 12047 3295 12053
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 5077 12087 5135 12093
rect 5077 12053 5089 12087
rect 5123 12084 5135 12087
rect 5368 12084 5396 12260
rect 5445 12223 5503 12229
rect 5445 12189 5457 12223
rect 5491 12189 5503 12223
rect 5920 12220 5948 12260
rect 6270 12220 6276 12232
rect 5920 12192 6276 12220
rect 5445 12183 5503 12189
rect 5123 12056 5396 12084
rect 5460 12084 5488 12183
rect 6270 12180 6276 12192
rect 6328 12180 6334 12232
rect 6650 12223 6708 12229
rect 6650 12189 6662 12223
rect 6696 12189 6708 12223
rect 6650 12183 6708 12189
rect 5626 12112 5632 12164
rect 5684 12152 5690 12164
rect 6546 12152 6552 12164
rect 5684 12124 6552 12152
rect 5684 12112 5690 12124
rect 6546 12112 6552 12124
rect 6604 12112 6610 12164
rect 6656 12152 6684 12183
rect 6822 12180 6828 12232
rect 6880 12220 6886 12232
rect 6917 12223 6975 12229
rect 6917 12220 6929 12223
rect 6880 12192 6929 12220
rect 6880 12180 6886 12192
rect 6917 12189 6929 12192
rect 6963 12220 6975 12223
rect 7009 12223 7067 12229
rect 7009 12220 7021 12223
rect 6963 12192 7021 12220
rect 6963 12189 6975 12192
rect 6917 12183 6975 12189
rect 7009 12189 7021 12192
rect 7055 12189 7067 12223
rect 7116 12220 7144 12260
rect 8036 12260 9505 12288
rect 7265 12223 7323 12229
rect 7265 12220 7277 12223
rect 7116 12192 7277 12220
rect 7009 12183 7067 12189
rect 7265 12189 7277 12192
rect 7311 12189 7323 12223
rect 7265 12183 7323 12189
rect 7558 12180 7564 12232
rect 7616 12220 7622 12232
rect 8036 12220 8064 12260
rect 9493 12257 9505 12260
rect 9539 12257 9551 12291
rect 9493 12251 9551 12257
rect 9674 12248 9680 12300
rect 9732 12248 9738 12300
rect 9858 12248 9864 12300
rect 9916 12288 9922 12300
rect 10321 12291 10379 12297
rect 10321 12288 10333 12291
rect 9916 12260 10333 12288
rect 9916 12248 9922 12260
rect 10321 12257 10333 12260
rect 10367 12257 10379 12291
rect 11146 12288 11152 12300
rect 10321 12251 10379 12257
rect 10612 12260 11152 12288
rect 7616 12192 8064 12220
rect 7616 12180 7622 12192
rect 8110 12180 8116 12232
rect 8168 12220 8174 12232
rect 8757 12223 8815 12229
rect 8757 12220 8769 12223
rect 8168 12192 8769 12220
rect 8168 12180 8174 12192
rect 8757 12189 8769 12192
rect 8803 12189 8815 12223
rect 8757 12183 8815 12189
rect 6730 12152 6736 12164
rect 6656 12124 6736 12152
rect 6730 12112 6736 12124
rect 6788 12112 6794 12164
rect 8772 12152 8800 12183
rect 9214 12180 9220 12232
rect 9272 12220 9278 12232
rect 9309 12223 9367 12229
rect 9309 12220 9321 12223
rect 9272 12192 9321 12220
rect 9272 12180 9278 12192
rect 9309 12189 9321 12192
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9398 12180 9404 12232
rect 9456 12220 9462 12232
rect 9456 12192 9501 12220
rect 9456 12180 9462 12192
rect 9692 12152 9720 12248
rect 10042 12180 10048 12232
rect 10100 12220 10106 12232
rect 10612 12229 10640 12260
rect 11146 12248 11152 12260
rect 11204 12248 11210 12300
rect 11256 12297 11284 12328
rect 11606 12316 11612 12368
rect 11664 12356 11670 12368
rect 12268 12365 12296 12396
rect 12434 12384 12440 12396
rect 12492 12384 12498 12436
rect 12897 12427 12955 12433
rect 12897 12393 12909 12427
rect 12943 12424 12955 12427
rect 13538 12424 13544 12436
rect 12943 12396 13544 12424
rect 12943 12393 12955 12396
rect 12897 12387 12955 12393
rect 11701 12359 11759 12365
rect 11701 12356 11713 12359
rect 11664 12328 11713 12356
rect 11664 12316 11670 12328
rect 11701 12325 11713 12328
rect 11747 12356 11759 12359
rect 12253 12359 12311 12365
rect 12253 12356 12265 12359
rect 11747 12328 12265 12356
rect 11747 12325 11759 12328
rect 11701 12319 11759 12325
rect 12253 12325 12265 12328
rect 12299 12325 12311 12359
rect 12253 12319 12311 12325
rect 12342 12316 12348 12368
rect 12400 12356 12406 12368
rect 12912 12356 12940 12387
rect 13538 12384 13544 12396
rect 13596 12384 13602 12436
rect 13814 12384 13820 12436
rect 13872 12424 13878 12436
rect 14277 12427 14335 12433
rect 14277 12424 14289 12427
rect 13872 12396 14289 12424
rect 13872 12384 13878 12396
rect 14277 12393 14289 12396
rect 14323 12393 14335 12427
rect 14277 12387 14335 12393
rect 12400 12328 12940 12356
rect 12400 12316 12406 12328
rect 13446 12316 13452 12368
rect 13504 12356 13510 12368
rect 16942 12356 16948 12368
rect 13504 12328 16948 12356
rect 13504 12316 13510 12328
rect 16942 12316 16948 12328
rect 17000 12316 17006 12368
rect 11241 12291 11299 12297
rect 11241 12257 11253 12291
rect 11287 12288 11299 12291
rect 11974 12288 11980 12300
rect 11287 12260 11980 12288
rect 11287 12257 11299 12260
rect 11241 12251 11299 12257
rect 11974 12248 11980 12260
rect 12032 12248 12038 12300
rect 12526 12288 12532 12300
rect 12439 12260 12532 12288
rect 12526 12248 12532 12260
rect 12584 12288 12590 12300
rect 14090 12288 14096 12300
rect 12584 12260 14096 12288
rect 12584 12248 12590 12260
rect 14090 12248 14096 12260
rect 14148 12248 14154 12300
rect 14458 12288 14464 12300
rect 14419 12260 14464 12288
rect 14458 12248 14464 12260
rect 14516 12248 14522 12300
rect 10229 12223 10287 12229
rect 10229 12220 10241 12223
rect 10100 12192 10241 12220
rect 10100 12180 10106 12192
rect 10229 12189 10241 12192
rect 10275 12220 10287 12223
rect 10597 12223 10655 12229
rect 10597 12220 10609 12223
rect 10275 12192 10609 12220
rect 10275 12189 10287 12192
rect 10229 12183 10287 12189
rect 10597 12189 10609 12192
rect 10643 12189 10655 12223
rect 13262 12220 13268 12232
rect 10597 12183 10655 12189
rect 10980 12192 13268 12220
rect 9858 12152 9864 12164
rect 6840 12124 8616 12152
rect 8772 12124 9260 12152
rect 9692 12124 9864 12152
rect 5718 12084 5724 12096
rect 5460 12056 5724 12084
rect 5123 12053 5135 12056
rect 5077 12047 5135 12053
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 5994 12044 6000 12096
rect 6052 12084 6058 12096
rect 6840 12084 6868 12124
rect 6052 12056 6868 12084
rect 6052 12044 6058 12056
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 8202 12084 8208 12096
rect 6972 12056 8208 12084
rect 6972 12044 6978 12056
rect 8202 12044 8208 12056
rect 8260 12084 8266 12096
rect 8389 12087 8447 12093
rect 8389 12084 8401 12087
rect 8260 12056 8401 12084
rect 8260 12044 8266 12056
rect 8389 12053 8401 12056
rect 8435 12053 8447 12087
rect 8588 12084 8616 12124
rect 9232 12096 9260 12124
rect 9858 12112 9864 12124
rect 9916 12112 9922 12164
rect 10137 12155 10195 12161
rect 10137 12121 10149 12155
rect 10183 12152 10195 12155
rect 10870 12152 10876 12164
rect 10183 12124 10876 12152
rect 10183 12121 10195 12124
rect 10137 12115 10195 12121
rect 10870 12112 10876 12124
rect 10928 12112 10934 12164
rect 8941 12087 8999 12093
rect 8941 12084 8953 12087
rect 8588 12056 8953 12084
rect 8389 12047 8447 12053
rect 8941 12053 8953 12056
rect 8987 12053 8999 12087
rect 8941 12047 8999 12053
rect 9214 12044 9220 12096
rect 9272 12044 9278 12096
rect 9582 12044 9588 12096
rect 9640 12084 9646 12096
rect 10980 12093 11008 12192
rect 13262 12180 13268 12192
rect 13320 12180 13326 12232
rect 11514 12112 11520 12164
rect 11572 12152 11578 12164
rect 11609 12155 11667 12161
rect 11609 12152 11621 12155
rect 11572 12124 11621 12152
rect 11572 12112 11578 12124
rect 11609 12121 11621 12124
rect 11655 12152 11667 12155
rect 13354 12152 13360 12164
rect 11655 12124 13360 12152
rect 11655 12121 11667 12124
rect 11609 12115 11667 12121
rect 13354 12112 13360 12124
rect 13412 12112 13418 12164
rect 14550 12152 14556 12164
rect 14108 12124 14556 12152
rect 10965 12087 11023 12093
rect 10965 12084 10977 12087
rect 9640 12056 10977 12084
rect 9640 12044 9646 12056
rect 10965 12053 10977 12056
rect 11011 12053 11023 12087
rect 10965 12047 11023 12053
rect 11790 12044 11796 12096
rect 11848 12084 11854 12096
rect 12069 12087 12127 12093
rect 12069 12084 12081 12087
rect 11848 12056 12081 12084
rect 11848 12044 11854 12056
rect 12069 12053 12081 12056
rect 12115 12053 12127 12087
rect 12618 12084 12624 12096
rect 12579 12056 12624 12084
rect 12069 12047 12127 12053
rect 12618 12044 12624 12056
rect 12676 12044 12682 12096
rect 13446 12084 13452 12096
rect 13407 12056 13452 12084
rect 13446 12044 13452 12056
rect 13504 12044 13510 12096
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 14108 12093 14136 12124
rect 14550 12112 14556 12124
rect 14608 12112 14614 12164
rect 14921 12155 14979 12161
rect 14921 12121 14933 12155
rect 14967 12152 14979 12155
rect 16482 12152 16488 12164
rect 14967 12124 16488 12152
rect 14967 12121 14979 12124
rect 14921 12115 14979 12121
rect 16482 12112 16488 12124
rect 16540 12112 16546 12164
rect 14093 12087 14151 12093
rect 14093 12084 14105 12087
rect 14056 12056 14105 12084
rect 14056 12044 14062 12056
rect 14093 12053 14105 12056
rect 14139 12053 14151 12087
rect 14093 12047 14151 12053
rect 14182 12044 14188 12096
rect 14240 12084 14246 12096
rect 15289 12087 15347 12093
rect 15289 12084 15301 12087
rect 14240 12056 15301 12084
rect 14240 12044 14246 12056
rect 15289 12053 15301 12056
rect 15335 12084 15347 12087
rect 16666 12084 16672 12096
rect 15335 12056 16672 12084
rect 15335 12053 15347 12056
rect 15289 12047 15347 12053
rect 16666 12044 16672 12056
rect 16724 12044 16730 12096
rect 1104 11994 16008 12016
rect 1104 11942 4698 11994
rect 4750 11942 4762 11994
rect 4814 11942 4826 11994
rect 4878 11942 4890 11994
rect 4942 11942 4954 11994
rect 5006 11942 8446 11994
rect 8498 11942 8510 11994
rect 8562 11942 8574 11994
rect 8626 11942 8638 11994
rect 8690 11942 8702 11994
rect 8754 11942 12194 11994
rect 12246 11942 12258 11994
rect 12310 11942 12322 11994
rect 12374 11942 12386 11994
rect 12438 11942 12450 11994
rect 12502 11942 16008 11994
rect 1104 11920 16008 11942
rect 1118 11840 1124 11892
rect 1176 11880 1182 11892
rect 1302 11880 1308 11892
rect 1176 11852 1308 11880
rect 1176 11840 1182 11852
rect 1302 11840 1308 11852
rect 1360 11840 1366 11892
rect 1578 11840 1584 11892
rect 1636 11880 1642 11892
rect 1765 11883 1823 11889
rect 1765 11880 1777 11883
rect 1636 11852 1777 11880
rect 1636 11840 1642 11852
rect 1765 11849 1777 11852
rect 1811 11849 1823 11883
rect 1765 11843 1823 11849
rect 2225 11883 2283 11889
rect 2225 11849 2237 11883
rect 2271 11880 2283 11883
rect 2406 11880 2412 11892
rect 2271 11852 2412 11880
rect 2271 11849 2283 11852
rect 2225 11843 2283 11849
rect 2406 11840 2412 11852
rect 2464 11840 2470 11892
rect 2682 11880 2688 11892
rect 2643 11852 2688 11880
rect 2682 11840 2688 11852
rect 2740 11840 2746 11892
rect 3050 11880 3056 11892
rect 3011 11852 3056 11880
rect 3050 11840 3056 11852
rect 3108 11840 3114 11892
rect 3878 11880 3884 11892
rect 3839 11852 3884 11880
rect 3878 11840 3884 11852
rect 3936 11840 3942 11892
rect 4338 11840 4344 11892
rect 4396 11840 4402 11892
rect 4709 11883 4767 11889
rect 4709 11849 4721 11883
rect 4755 11880 4767 11883
rect 5718 11880 5724 11892
rect 4755 11852 5724 11880
rect 4755 11849 4767 11852
rect 4709 11843 4767 11849
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 6270 11840 6276 11892
rect 6328 11880 6334 11892
rect 6328 11852 8993 11880
rect 6328 11840 6334 11852
rect 2590 11772 2596 11824
rect 2648 11812 2654 11824
rect 3421 11815 3479 11821
rect 3421 11812 3433 11815
rect 2648 11784 3433 11812
rect 2648 11772 2654 11784
rect 3421 11781 3433 11784
rect 3467 11781 3479 11815
rect 3421 11775 3479 11781
rect 3513 11815 3571 11821
rect 3513 11781 3525 11815
rect 3559 11812 3571 11815
rect 4062 11812 4068 11824
rect 3559 11784 4068 11812
rect 3559 11781 3571 11784
rect 3513 11775 3571 11781
rect 4062 11772 4068 11784
rect 4120 11772 4126 11824
rect 4356 11812 4384 11840
rect 4356 11784 5212 11812
rect 1854 11744 1860 11756
rect 1815 11716 1860 11744
rect 1854 11704 1860 11716
rect 1912 11704 1918 11756
rect 3970 11704 3976 11756
rect 4028 11744 4034 11756
rect 4249 11747 4307 11753
rect 4249 11744 4261 11747
rect 4028 11716 4261 11744
rect 4028 11704 4034 11716
rect 4249 11713 4261 11716
rect 4295 11713 4307 11747
rect 4249 11707 4307 11713
rect 4341 11747 4399 11753
rect 4341 11713 4353 11747
rect 4387 11744 4399 11747
rect 4614 11744 4620 11756
rect 4387 11716 4620 11744
rect 4387 11713 4399 11716
rect 4341 11707 4399 11713
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 5057 11747 5115 11753
rect 5057 11744 5069 11747
rect 4724 11716 5069 11744
rect 1578 11676 1584 11688
rect 1539 11648 1584 11676
rect 1578 11636 1584 11648
rect 1636 11636 1642 11688
rect 2501 11679 2559 11685
rect 2501 11645 2513 11679
rect 2547 11645 2559 11679
rect 2501 11639 2559 11645
rect 2516 11608 2544 11639
rect 2590 11636 2596 11688
rect 2648 11676 2654 11688
rect 3329 11679 3387 11685
rect 2648 11648 2693 11676
rect 2648 11636 2654 11648
rect 3329 11645 3341 11679
rect 3375 11676 3387 11679
rect 3602 11676 3608 11688
rect 3375 11648 3608 11676
rect 3375 11645 3387 11648
rect 3329 11639 3387 11645
rect 3602 11636 3608 11648
rect 3660 11636 3666 11688
rect 4062 11636 4068 11688
rect 4120 11676 4126 11688
rect 4157 11679 4215 11685
rect 4157 11676 4169 11679
rect 4120 11648 4169 11676
rect 4120 11636 4126 11648
rect 4157 11645 4169 11648
rect 4203 11645 4215 11679
rect 4157 11639 4215 11645
rect 3620 11608 3648 11636
rect 4522 11608 4528 11620
rect 2516 11580 2774 11608
rect 3620 11580 4528 11608
rect 2746 11540 2774 11580
rect 4522 11568 4528 11580
rect 4580 11608 4586 11620
rect 4724 11608 4752 11716
rect 5057 11713 5069 11716
rect 5103 11713 5115 11747
rect 5184 11744 5212 11784
rect 6730 11772 6736 11824
rect 6788 11812 6794 11824
rect 6788 11784 7420 11812
rect 6788 11772 6794 11784
rect 6621 11747 6679 11753
rect 6621 11744 6633 11747
rect 5184 11716 6633 11744
rect 5057 11707 5115 11713
rect 6621 11713 6633 11716
rect 6667 11713 6679 11747
rect 6621 11707 6679 11713
rect 4801 11679 4859 11685
rect 4801 11645 4813 11679
rect 4847 11645 4859 11679
rect 6362 11676 6368 11688
rect 6323 11648 6368 11676
rect 4801 11639 4859 11645
rect 4580 11580 4752 11608
rect 4580 11568 4586 11580
rect 4154 11540 4160 11552
rect 2746 11512 4160 11540
rect 4154 11500 4160 11512
rect 4212 11540 4218 11552
rect 4706 11540 4712 11552
rect 4212 11512 4712 11540
rect 4212 11500 4218 11512
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 4816 11540 4844 11639
rect 6362 11636 6368 11648
rect 6420 11636 6426 11688
rect 7392 11676 7420 11784
rect 8110 11772 8116 11824
rect 8168 11812 8174 11824
rect 8297 11815 8355 11821
rect 8297 11812 8309 11815
rect 8168 11784 8309 11812
rect 8168 11772 8174 11784
rect 8297 11781 8309 11784
rect 8343 11781 8355 11815
rect 8965 11812 8993 11852
rect 9030 11840 9036 11892
rect 9088 11880 9094 11892
rect 10042 11880 10048 11892
rect 9088 11852 9133 11880
rect 9692 11852 10048 11880
rect 9088 11840 9094 11852
rect 9692 11812 9720 11852
rect 10042 11840 10048 11852
rect 10100 11840 10106 11892
rect 10410 11840 10416 11892
rect 10468 11880 10474 11892
rect 11514 11880 11520 11892
rect 10468 11852 11520 11880
rect 10468 11840 10474 11852
rect 11514 11840 11520 11852
rect 11572 11840 11578 11892
rect 12529 11883 12587 11889
rect 12529 11849 12541 11883
rect 12575 11880 12587 11883
rect 12894 11880 12900 11892
rect 12575 11852 12900 11880
rect 12575 11849 12587 11852
rect 12529 11843 12587 11849
rect 12894 11840 12900 11852
rect 12952 11880 12958 11892
rect 13906 11880 13912 11892
rect 12952 11852 13912 11880
rect 12952 11840 12958 11852
rect 13906 11840 13912 11852
rect 13964 11840 13970 11892
rect 14550 11880 14556 11892
rect 14511 11852 14556 11880
rect 14550 11840 14556 11852
rect 14608 11840 14614 11892
rect 14734 11840 14740 11892
rect 14792 11880 14798 11892
rect 14829 11883 14887 11889
rect 14829 11880 14841 11883
rect 14792 11852 14841 11880
rect 14792 11840 14798 11852
rect 14829 11849 14841 11852
rect 14875 11849 14887 11883
rect 14829 11843 14887 11849
rect 10689 11815 10747 11821
rect 10689 11812 10701 11815
rect 8965 11784 9720 11812
rect 9784 11784 10701 11812
rect 8297 11775 8355 11781
rect 8205 11747 8263 11753
rect 8205 11713 8217 11747
rect 8251 11744 8263 11747
rect 8662 11744 8668 11756
rect 8251 11716 8668 11744
rect 8251 11713 8263 11716
rect 8205 11707 8263 11713
rect 8662 11704 8668 11716
rect 8720 11704 8726 11756
rect 8846 11704 8852 11756
rect 8904 11744 8910 11756
rect 8941 11747 8999 11753
rect 8941 11744 8953 11747
rect 8904 11716 8953 11744
rect 8904 11704 8910 11716
rect 8941 11713 8953 11716
rect 8987 11713 8999 11747
rect 8941 11707 8999 11713
rect 8294 11676 8300 11688
rect 7392 11648 8300 11676
rect 8294 11636 8300 11648
rect 8352 11676 8358 11688
rect 8389 11679 8447 11685
rect 8389 11676 8401 11679
rect 8352 11648 8401 11676
rect 8352 11636 8358 11648
rect 8389 11645 8401 11648
rect 8435 11645 8447 11679
rect 8757 11679 8815 11685
rect 8757 11676 8769 11679
rect 8389 11639 8447 11645
rect 8680 11648 8769 11676
rect 6086 11568 6092 11620
rect 6144 11608 6150 11620
rect 6181 11611 6239 11617
rect 6181 11608 6193 11611
rect 6144 11580 6193 11608
rect 6144 11568 6150 11580
rect 6181 11577 6193 11580
rect 6227 11608 6239 11611
rect 6270 11608 6276 11620
rect 6227 11580 6276 11608
rect 6227 11577 6239 11580
rect 6181 11571 6239 11577
rect 6270 11568 6276 11580
rect 6328 11568 6334 11620
rect 7837 11611 7895 11617
rect 7837 11608 7849 11611
rect 7300 11580 7849 11608
rect 5166 11540 5172 11552
rect 4816 11512 5172 11540
rect 5166 11500 5172 11512
rect 5224 11500 5230 11552
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 7300 11540 7328 11580
rect 7837 11577 7849 11580
rect 7883 11577 7895 11611
rect 7837 11571 7895 11577
rect 5500 11512 7328 11540
rect 5500 11500 5506 11512
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 7524 11512 7757 11540
rect 7524 11500 7530 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 7745 11503 7803 11509
rect 8202 11500 8208 11552
rect 8260 11540 8266 11552
rect 8680 11540 8708 11648
rect 8757 11645 8769 11648
rect 8803 11645 8815 11679
rect 8956 11676 8984 11707
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 9784 11744 9812 11784
rect 10689 11781 10701 11784
rect 10735 11781 10747 11815
rect 10689 11775 10747 11781
rect 10781 11815 10839 11821
rect 10781 11781 10793 11815
rect 10827 11812 10839 11815
rect 11790 11812 11796 11824
rect 10827 11784 11796 11812
rect 10827 11781 10839 11784
rect 10781 11775 10839 11781
rect 11790 11772 11796 11784
rect 11848 11772 11854 11824
rect 11885 11815 11943 11821
rect 11885 11781 11897 11815
rect 11931 11812 11943 11815
rect 11974 11812 11980 11824
rect 11931 11784 11980 11812
rect 11931 11781 11943 11784
rect 11885 11775 11943 11781
rect 11974 11772 11980 11784
rect 12032 11812 12038 11824
rect 12032 11784 12204 11812
rect 12032 11772 12038 11784
rect 9640 11716 9812 11744
rect 9861 11747 9919 11753
rect 9640 11704 9646 11716
rect 9861 11713 9873 11747
rect 9907 11713 9919 11747
rect 9861 11707 9919 11713
rect 8956 11648 9628 11676
rect 8757 11639 8815 11645
rect 8938 11568 8944 11620
rect 8996 11608 9002 11620
rect 9493 11611 9551 11617
rect 9493 11608 9505 11611
rect 8996 11580 9505 11608
rect 8996 11568 9002 11580
rect 9493 11577 9505 11580
rect 9539 11577 9551 11611
rect 9600 11608 9628 11648
rect 9674 11636 9680 11688
rect 9732 11676 9738 11688
rect 9876 11676 9904 11707
rect 10594 11704 10600 11756
rect 10652 11704 10658 11756
rect 11146 11744 11152 11756
rect 11107 11716 11152 11744
rect 11146 11704 11152 11716
rect 11204 11704 11210 11756
rect 11238 11704 11244 11756
rect 11296 11744 11302 11756
rect 12069 11747 12127 11753
rect 12069 11744 12081 11747
rect 11296 11716 12081 11744
rect 11296 11704 11302 11716
rect 9732 11648 9904 11676
rect 9953 11679 10011 11685
rect 9732 11636 9738 11648
rect 9953 11645 9965 11679
rect 9999 11645 10011 11679
rect 9953 11639 10011 11645
rect 10137 11679 10195 11685
rect 10137 11645 10149 11679
rect 10183 11676 10195 11679
rect 10226 11676 10232 11688
rect 10183 11648 10232 11676
rect 10183 11645 10195 11648
rect 10137 11639 10195 11645
rect 9766 11608 9772 11620
rect 9600 11580 9772 11608
rect 9493 11571 9551 11577
rect 9766 11568 9772 11580
rect 9824 11568 9830 11620
rect 9858 11568 9864 11620
rect 9916 11568 9922 11620
rect 9968 11608 9996 11639
rect 10226 11636 10232 11648
rect 10284 11676 10290 11688
rect 10410 11676 10416 11688
rect 10284 11648 10416 11676
rect 10284 11636 10290 11648
rect 10410 11636 10416 11648
rect 10468 11636 10474 11688
rect 10612 11676 10640 11704
rect 11532 11688 11560 11716
rect 12069 11713 12081 11716
rect 12115 11713 12127 11747
rect 12176 11744 12204 11784
rect 12434 11772 12440 11824
rect 12492 11812 12498 11824
rect 13078 11812 13084 11824
rect 12492 11784 13084 11812
rect 12492 11772 12498 11784
rect 13078 11772 13084 11784
rect 13136 11812 13142 11824
rect 13173 11815 13231 11821
rect 13173 11812 13185 11815
rect 13136 11784 13185 11812
rect 13136 11772 13142 11784
rect 13173 11781 13185 11784
rect 13219 11781 13231 11815
rect 15381 11815 15439 11821
rect 15381 11812 15393 11815
rect 13173 11775 13231 11781
rect 13280 11784 15393 11812
rect 13280 11744 13308 11784
rect 15381 11781 15393 11784
rect 15427 11812 15439 11815
rect 16206 11812 16212 11824
rect 15427 11784 16212 11812
rect 15427 11781 15439 11784
rect 15381 11775 15439 11781
rect 16206 11772 16212 11784
rect 16264 11772 16270 11824
rect 12176 11716 13308 11744
rect 12069 11707 12127 11713
rect 13354 11704 13360 11756
rect 13412 11744 13418 11756
rect 14737 11747 14795 11753
rect 14737 11744 14749 11747
rect 13412 11716 14749 11744
rect 13412 11704 13418 11716
rect 14737 11713 14749 11716
rect 14783 11744 14795 11747
rect 16298 11744 16304 11756
rect 14783 11716 16304 11744
rect 14783 11713 14795 11716
rect 14737 11707 14795 11713
rect 16298 11704 16304 11716
rect 16356 11704 16362 11756
rect 10873 11679 10931 11685
rect 10873 11676 10885 11679
rect 10612 11648 10885 11676
rect 10873 11645 10885 11648
rect 10919 11645 10931 11679
rect 10873 11639 10931 11645
rect 11514 11636 11520 11688
rect 11572 11636 11578 11688
rect 11793 11679 11851 11685
rect 11793 11645 11805 11679
rect 11839 11676 11851 11679
rect 11974 11676 11980 11688
rect 11839 11648 11980 11676
rect 11839 11645 11851 11648
rect 11793 11639 11851 11645
rect 11808 11608 11836 11639
rect 11974 11636 11980 11648
rect 12032 11636 12038 11688
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11645 12311 11679
rect 12253 11639 12311 11645
rect 12268 11608 12296 11639
rect 12342 11636 12348 11688
rect 12400 11676 12406 11688
rect 12526 11676 12532 11688
rect 12400 11648 12532 11676
rect 12400 11636 12406 11648
rect 12526 11636 12532 11648
rect 12584 11676 12590 11688
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 12584 11648 12633 11676
rect 12584 11636 12590 11648
rect 12621 11645 12633 11648
rect 12667 11676 12679 11679
rect 13817 11679 13875 11685
rect 12667 11648 13768 11676
rect 12667 11645 12679 11648
rect 12621 11639 12679 11645
rect 9968 11580 11836 11608
rect 11900 11580 12296 11608
rect 13740 11608 13768 11648
rect 13817 11645 13829 11679
rect 13863 11676 13875 11679
rect 13906 11676 13912 11688
rect 13863 11648 13912 11676
rect 13863 11645 13875 11648
rect 13817 11639 13875 11645
rect 13906 11636 13912 11648
rect 13964 11636 13970 11688
rect 15013 11679 15071 11685
rect 15013 11676 15025 11679
rect 14016 11648 15025 11676
rect 14016 11617 14044 11648
rect 15013 11645 15025 11648
rect 15059 11676 15071 11679
rect 15102 11676 15108 11688
rect 15059 11648 15108 11676
rect 15059 11645 15071 11648
rect 15013 11639 15071 11645
rect 15102 11636 15108 11648
rect 15160 11636 15166 11688
rect 15378 11636 15384 11688
rect 15436 11676 15442 11688
rect 15930 11676 15936 11688
rect 15436 11648 15936 11676
rect 15436 11636 15442 11648
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 14001 11611 14059 11617
rect 14001 11608 14013 11611
rect 13740 11580 14013 11608
rect 9398 11540 9404 11552
rect 8260 11512 8708 11540
rect 9359 11512 9404 11540
rect 8260 11500 8266 11512
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 9876 11540 9904 11568
rect 10888 11552 10916 11580
rect 10321 11543 10379 11549
rect 10321 11540 10333 11543
rect 9876 11512 10333 11540
rect 10321 11509 10333 11512
rect 10367 11509 10379 11543
rect 10321 11503 10379 11509
rect 10870 11500 10876 11552
rect 10928 11500 10934 11552
rect 11238 11500 11244 11552
rect 11296 11540 11302 11552
rect 11900 11540 11928 11580
rect 14001 11577 14013 11580
rect 14047 11577 14059 11611
rect 14001 11571 14059 11577
rect 14090 11568 14096 11620
rect 14148 11568 14154 11620
rect 14274 11568 14280 11620
rect 14332 11608 14338 11620
rect 14369 11611 14427 11617
rect 14369 11608 14381 11611
rect 14332 11580 14381 11608
rect 14332 11568 14338 11580
rect 14369 11577 14381 11580
rect 14415 11608 14427 11611
rect 16022 11608 16028 11620
rect 14415 11580 16028 11608
rect 14415 11577 14427 11580
rect 14369 11571 14427 11577
rect 16022 11568 16028 11580
rect 16080 11568 16086 11620
rect 11296 11512 11928 11540
rect 11296 11500 11302 11512
rect 12250 11500 12256 11552
rect 12308 11540 12314 11552
rect 12805 11543 12863 11549
rect 12805 11540 12817 11543
rect 12308 11512 12817 11540
rect 12308 11500 12314 11512
rect 12805 11509 12817 11512
rect 12851 11509 12863 11543
rect 13078 11540 13084 11552
rect 13039 11512 13084 11540
rect 12805 11503 12863 11509
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13354 11540 13360 11552
rect 13315 11512 13360 11540
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 13633 11543 13691 11549
rect 13633 11509 13645 11543
rect 13679 11540 13691 11543
rect 14108 11540 14136 11568
rect 14185 11543 14243 11549
rect 14185 11540 14197 11543
rect 13679 11512 14197 11540
rect 13679 11509 13691 11512
rect 13633 11503 13691 11509
rect 14185 11509 14197 11512
rect 14231 11540 14243 11543
rect 15010 11540 15016 11552
rect 14231 11512 15016 11540
rect 14231 11509 14243 11512
rect 14185 11503 14243 11509
rect 15010 11500 15016 11512
rect 15068 11500 15074 11552
rect 15289 11543 15347 11549
rect 15289 11509 15301 11543
rect 15335 11540 15347 11543
rect 15378 11540 15384 11552
rect 15335 11512 15384 11540
rect 15335 11509 15347 11512
rect 15289 11503 15347 11509
rect 15378 11500 15384 11512
rect 15436 11500 15442 11552
rect 15562 11540 15568 11552
rect 15523 11512 15568 11540
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 1104 11450 16008 11472
rect 1104 11398 2824 11450
rect 2876 11398 2888 11450
rect 2940 11398 2952 11450
rect 3004 11398 3016 11450
rect 3068 11398 3080 11450
rect 3132 11398 6572 11450
rect 6624 11398 6636 11450
rect 6688 11398 6700 11450
rect 6752 11398 6764 11450
rect 6816 11398 6828 11450
rect 6880 11398 10320 11450
rect 10372 11398 10384 11450
rect 10436 11398 10448 11450
rect 10500 11398 10512 11450
rect 10564 11398 10576 11450
rect 10628 11398 14068 11450
rect 14120 11398 14132 11450
rect 14184 11398 14196 11450
rect 14248 11398 14260 11450
rect 14312 11398 14324 11450
rect 14376 11398 16008 11450
rect 1104 11376 16008 11398
rect 3510 11336 3516 11348
rect 2884 11308 3516 11336
rect 2777 11271 2835 11277
rect 2777 11237 2789 11271
rect 2823 11268 2835 11271
rect 2884 11268 2912 11308
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 4154 11296 4160 11348
rect 4212 11336 4218 11348
rect 4338 11336 4344 11348
rect 4212 11308 4344 11336
rect 4212 11296 4218 11308
rect 4338 11296 4344 11308
rect 4396 11296 4402 11348
rect 4614 11336 4620 11348
rect 4575 11308 4620 11336
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 5442 11336 5448 11348
rect 4724 11308 5448 11336
rect 4724 11268 4752 11308
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 7190 11336 7196 11348
rect 6380 11308 7196 11336
rect 2823 11240 2912 11268
rect 2985 11240 4752 11268
rect 2823 11237 2835 11240
rect 2777 11231 2835 11237
rect 1670 11200 1676 11212
rect 1631 11172 1676 11200
rect 1670 11160 1676 11172
rect 1728 11160 1734 11212
rect 2222 11200 2228 11212
rect 2183 11172 2228 11200
rect 2222 11160 2228 11172
rect 2280 11160 2286 11212
rect 1946 11132 1952 11144
rect 1907 11104 1952 11132
rect 1946 11092 1952 11104
rect 2004 11092 2010 11144
rect 2409 11135 2467 11141
rect 2409 11101 2421 11135
rect 2455 11132 2467 11135
rect 2985 11132 3013 11240
rect 6086 11228 6092 11280
rect 6144 11268 6150 11280
rect 6181 11271 6239 11277
rect 6181 11268 6193 11271
rect 6144 11240 6193 11268
rect 6144 11228 6150 11240
rect 6181 11237 6193 11240
rect 6227 11268 6239 11271
rect 6380 11268 6408 11308
rect 7190 11296 7196 11308
rect 7248 11296 7254 11348
rect 7282 11296 7288 11348
rect 7340 11336 7346 11348
rect 7653 11339 7711 11345
rect 7653 11336 7665 11339
rect 7340 11308 7665 11336
rect 7340 11296 7346 11308
rect 7653 11305 7665 11308
rect 7699 11305 7711 11339
rect 7653 11299 7711 11305
rect 8941 11339 8999 11345
rect 8941 11305 8953 11339
rect 8987 11336 8999 11339
rect 9030 11336 9036 11348
rect 8987 11308 9036 11336
rect 8987 11305 8999 11308
rect 8941 11299 8999 11305
rect 9030 11296 9036 11308
rect 9088 11296 9094 11348
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 9364 11308 9812 11336
rect 9364 11296 9370 11308
rect 9784 11277 9812 11308
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10597 11339 10655 11345
rect 10597 11336 10609 11339
rect 10192 11308 10609 11336
rect 10192 11296 10198 11308
rect 10597 11305 10609 11308
rect 10643 11305 10655 11339
rect 11974 11336 11980 11348
rect 10597 11299 10655 11305
rect 10695 11308 11980 11336
rect 9769 11271 9827 11277
rect 6227 11240 6408 11268
rect 8220 11240 9536 11268
rect 6227 11237 6239 11240
rect 6181 11231 6239 11237
rect 3326 11200 3332 11212
rect 3287 11172 3332 11200
rect 3326 11160 3332 11172
rect 3384 11160 3390 11212
rect 3513 11203 3571 11209
rect 3513 11169 3525 11203
rect 3559 11200 3571 11203
rect 3786 11200 3792 11212
rect 3559 11172 3792 11200
rect 3559 11169 3571 11172
rect 3513 11163 3571 11169
rect 3786 11160 3792 11172
rect 3844 11160 3850 11212
rect 4062 11200 4068 11212
rect 4023 11172 4068 11200
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4157 11203 4215 11209
rect 4157 11169 4169 11203
rect 4203 11200 4215 11203
rect 5074 11200 5080 11212
rect 4203 11172 5080 11200
rect 4203 11169 4215 11172
rect 4157 11163 4215 11169
rect 4172 11132 4200 11163
rect 5074 11160 5080 11172
rect 5132 11160 5138 11212
rect 7926 11160 7932 11212
rect 7984 11200 7990 11212
rect 8220 11209 8248 11240
rect 8205 11203 8263 11209
rect 8205 11200 8217 11203
rect 7984 11172 8217 11200
rect 7984 11160 7990 11172
rect 8205 11169 8217 11172
rect 8251 11169 8263 11203
rect 8205 11163 8263 11169
rect 8665 11203 8723 11209
rect 8665 11169 8677 11203
rect 8711 11200 8723 11203
rect 8846 11200 8852 11212
rect 8711 11172 8852 11200
rect 8711 11169 8723 11172
rect 8665 11163 8723 11169
rect 8846 11160 8852 11172
rect 8904 11160 8910 11212
rect 9508 11209 9536 11240
rect 9769 11237 9781 11271
rect 9815 11237 9827 11271
rect 10695 11268 10723 11308
rect 11974 11296 11980 11308
rect 12032 11336 12038 11348
rect 12434 11336 12440 11348
rect 12032 11308 12440 11336
rect 12032 11296 12038 11308
rect 12434 11296 12440 11308
rect 12492 11296 12498 11348
rect 12710 11336 12716 11348
rect 12671 11308 12716 11336
rect 12710 11296 12716 11308
rect 12768 11296 12774 11348
rect 12894 11336 12900 11348
rect 12855 11308 12900 11336
rect 12894 11296 12900 11308
rect 12952 11296 12958 11348
rect 12986 11296 12992 11348
rect 13044 11336 13050 11348
rect 13173 11339 13231 11345
rect 13173 11336 13185 11339
rect 13044 11308 13185 11336
rect 13044 11296 13050 11308
rect 13173 11305 13185 11308
rect 13219 11305 13231 11339
rect 13173 11299 13231 11305
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 14277 11339 14335 11345
rect 14277 11336 14289 11339
rect 13596 11308 14289 11336
rect 13596 11296 13602 11308
rect 14277 11305 14289 11308
rect 14323 11305 14335 11339
rect 14550 11336 14556 11348
rect 14511 11308 14556 11336
rect 14277 11299 14335 11305
rect 14550 11296 14556 11308
rect 14608 11296 14614 11348
rect 15378 11336 15384 11348
rect 14844 11308 15384 11336
rect 9769 11231 9827 11237
rect 10244 11240 10723 11268
rect 11072 11240 11284 11268
rect 9401 11203 9459 11209
rect 9401 11169 9413 11203
rect 9447 11169 9459 11203
rect 9401 11163 9459 11169
rect 9493 11203 9551 11209
rect 9493 11169 9505 11203
rect 9539 11169 9551 11203
rect 10244 11200 10272 11240
rect 9493 11163 9551 11169
rect 9784 11172 10272 11200
rect 5994 11132 6000 11144
rect 2455 11104 3013 11132
rect 3068 11104 4200 11132
rect 4448 11104 6000 11132
rect 2455 11101 2467 11104
rect 2409 11095 2467 11101
rect 2314 11064 2320 11076
rect 2275 11036 2320 11064
rect 2314 11024 2320 11036
rect 2372 11024 2378 11076
rect 3068 11064 3096 11104
rect 2424 11036 3096 11064
rect 3237 11067 3295 11073
rect 1578 10956 1584 11008
rect 1636 10996 1642 11008
rect 2424 10996 2452 11036
rect 3237 11033 3249 11067
rect 3283 11064 3295 11067
rect 4448 11064 4476 11104
rect 5994 11092 6000 11104
rect 6052 11092 6058 11144
rect 6089 11135 6147 11141
rect 6089 11101 6101 11135
rect 6135 11132 6147 11135
rect 6362 11132 6368 11144
rect 6135 11104 6368 11132
rect 6135 11101 6147 11104
rect 6089 11095 6147 11101
rect 6362 11092 6368 11104
rect 6420 11132 6426 11144
rect 7561 11135 7619 11141
rect 7561 11132 7573 11135
rect 6420 11104 7573 11132
rect 6420 11092 6426 11104
rect 7561 11101 7573 11104
rect 7607 11101 7619 11135
rect 7561 11095 7619 11101
rect 7742 11092 7748 11144
rect 7800 11092 7806 11144
rect 7834 11092 7840 11144
rect 7892 11132 7898 11144
rect 8018 11132 8024 11144
rect 7892 11104 8024 11132
rect 7892 11092 7898 11104
rect 8018 11092 8024 11104
rect 8076 11092 8082 11144
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 9214 11132 9220 11144
rect 8444 11104 9220 11132
rect 8444 11092 8450 11104
rect 9214 11092 9220 11104
rect 9272 11092 9278 11144
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9416 11132 9444 11163
rect 9784 11132 9812 11172
rect 10318 11160 10324 11212
rect 10376 11200 10382 11212
rect 11072 11200 11100 11240
rect 10376 11172 10421 11200
rect 10520 11172 11100 11200
rect 11149 11203 11207 11209
rect 10376 11160 10382 11172
rect 9416 11104 9812 11132
rect 9309 11095 9367 11101
rect 3283 11036 4476 11064
rect 3283 11033 3295 11036
rect 3237 11027 3295 11033
rect 4522 11024 4528 11076
rect 4580 11064 4586 11076
rect 4580 11036 4752 11064
rect 4580 11024 4586 11036
rect 1636 10968 2452 10996
rect 1636 10956 1642 10968
rect 2590 10956 2596 11008
rect 2648 10996 2654 11008
rect 2869 10999 2927 11005
rect 2869 10996 2881 10999
rect 2648 10968 2881 10996
rect 2648 10956 2654 10968
rect 2869 10965 2881 10968
rect 2915 10965 2927 10999
rect 2869 10959 2927 10965
rect 4246 10956 4252 11008
rect 4304 10996 4310 11008
rect 4724 11005 4752 11036
rect 4890 11024 4896 11076
rect 4948 11064 4954 11076
rect 5442 11064 5448 11076
rect 4948 11036 5448 11064
rect 4948 11024 4954 11036
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 5810 11024 5816 11076
rect 5868 11073 5874 11076
rect 5868 11064 5880 11073
rect 7316 11067 7374 11073
rect 5868 11036 5913 11064
rect 5868 11027 5880 11036
rect 7316 11033 7328 11067
rect 7362 11064 7374 11067
rect 7650 11064 7656 11076
rect 7362 11036 7656 11064
rect 7362 11033 7374 11036
rect 7316 11027 7374 11033
rect 5868 11024 5874 11027
rect 7650 11024 7656 11036
rect 7708 11024 7714 11076
rect 7760 11064 7788 11092
rect 9030 11064 9036 11076
rect 7760 11036 9036 11064
rect 9030 11024 9036 11036
rect 9088 11024 9094 11076
rect 9324 11064 9352 11095
rect 9858 11092 9864 11144
rect 9916 11132 9922 11144
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 9916 11104 10149 11132
rect 9916 11092 9922 11104
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 10137 11095 10195 11101
rect 10229 11135 10287 11141
rect 10229 11101 10241 11135
rect 10275 11132 10287 11135
rect 10520 11132 10548 11172
rect 11149 11169 11161 11203
rect 11195 11169 11207 11203
rect 11256 11200 11284 11240
rect 11514 11228 11520 11280
rect 11572 11268 11578 11280
rect 11572 11240 12112 11268
rect 11572 11228 11578 11240
rect 11606 11200 11612 11212
rect 11256 11172 11612 11200
rect 11149 11163 11207 11169
rect 10275 11104 10548 11132
rect 10275 11101 10287 11104
rect 10229 11095 10287 11101
rect 10594 11092 10600 11144
rect 10652 11132 10658 11144
rect 11164 11132 11192 11163
rect 11606 11160 11612 11172
rect 11664 11160 11670 11212
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 11808 11172 11989 11200
rect 11808 11132 11836 11172
rect 11977 11169 11989 11172
rect 12023 11169 12035 11203
rect 12084 11200 12112 11240
rect 12158 11228 12164 11280
rect 12216 11268 12222 11280
rect 12216 11240 14044 11268
rect 12216 11228 12222 11240
rect 14016 11212 14044 11240
rect 14366 11228 14372 11280
rect 14424 11268 14430 11280
rect 14844 11268 14872 11308
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 15473 11339 15531 11345
rect 15473 11305 15485 11339
rect 15519 11336 15531 11339
rect 15562 11336 15568 11348
rect 15519 11308 15568 11336
rect 15519 11305 15531 11308
rect 15473 11299 15531 11305
rect 15562 11296 15568 11308
rect 15620 11336 15626 11348
rect 15838 11336 15844 11348
rect 15620 11308 15844 11336
rect 15620 11296 15626 11308
rect 15838 11296 15844 11308
rect 15896 11296 15902 11348
rect 14424 11240 14872 11268
rect 14921 11271 14979 11277
rect 14424 11228 14430 11240
rect 14921 11237 14933 11271
rect 14967 11268 14979 11271
rect 16574 11268 16580 11280
rect 14967 11240 16580 11268
rect 14967 11237 14979 11240
rect 14921 11231 14979 11237
rect 13446 11200 13452 11212
rect 12084 11172 12480 11200
rect 11977 11163 12035 11169
rect 10652 11104 11192 11132
rect 11256 11104 11836 11132
rect 11885 11135 11943 11141
rect 10652 11092 10658 11104
rect 9950 11064 9956 11076
rect 9324 11036 9956 11064
rect 9950 11024 9956 11036
rect 10008 11064 10014 11076
rect 10502 11064 10508 11076
rect 10008 11036 10508 11064
rect 10008 11024 10014 11036
rect 10502 11024 10508 11036
rect 10560 11024 10566 11076
rect 10962 11064 10968 11076
rect 10923 11036 10968 11064
rect 10962 11024 10968 11036
rect 11020 11024 11026 11076
rect 11057 11067 11115 11073
rect 11057 11033 11069 11067
rect 11103 11064 11115 11067
rect 11146 11064 11152 11076
rect 11103 11036 11152 11064
rect 11103 11033 11115 11036
rect 11057 11027 11115 11033
rect 11146 11024 11152 11036
rect 11204 11024 11210 11076
rect 4709 10999 4767 11005
rect 4304 10968 4349 10996
rect 4304 10956 4310 10968
rect 4709 10965 4721 10999
rect 4755 10965 4767 10999
rect 4709 10959 4767 10965
rect 6822 10956 6828 11008
rect 6880 10996 6886 11008
rect 7466 10996 7472 11008
rect 6880 10968 7472 10996
rect 6880 10956 6886 10968
rect 7466 10956 7472 10968
rect 7524 10956 7530 11008
rect 7742 10956 7748 11008
rect 7800 10996 7806 11008
rect 8021 10999 8079 11005
rect 8021 10996 8033 10999
rect 7800 10968 8033 10996
rect 7800 10956 7806 10968
rect 8021 10965 8033 10968
rect 8067 10965 8079 10999
rect 8021 10959 8079 10965
rect 8113 10999 8171 11005
rect 8113 10965 8125 10999
rect 8159 10996 8171 10999
rect 10134 10996 10140 11008
rect 8159 10968 10140 10996
rect 8159 10965 8171 10968
rect 8113 10959 8171 10965
rect 10134 10956 10140 10968
rect 10192 10956 10198 11008
rect 10318 10956 10324 11008
rect 10376 10996 10382 11008
rect 11256 10996 11284 11104
rect 11885 11101 11897 11135
rect 11931 11132 11943 11135
rect 12342 11132 12348 11144
rect 11931 11104 12348 11132
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 11606 11024 11612 11076
rect 11664 11064 11670 11076
rect 12250 11064 12256 11076
rect 11664 11036 12256 11064
rect 11664 11024 11670 11036
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 12452 11064 12480 11172
rect 13096 11172 13452 11200
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 13096 11132 13124 11172
rect 13446 11160 13452 11172
rect 13504 11200 13510 11212
rect 13725 11203 13783 11209
rect 13725 11200 13737 11203
rect 13504 11172 13737 11200
rect 13504 11160 13510 11172
rect 13725 11169 13737 11172
rect 13771 11169 13783 11203
rect 13725 11163 13783 11169
rect 13998 11160 14004 11212
rect 14056 11200 14062 11212
rect 14936 11200 14964 11231
rect 16574 11228 16580 11240
rect 16632 11228 16638 11280
rect 14056 11172 14964 11200
rect 14056 11160 14062 11172
rect 12860 11104 13124 11132
rect 12860 11092 12866 11104
rect 13170 11092 13176 11144
rect 13228 11132 13234 11144
rect 13357 11135 13415 11141
rect 13357 11132 13369 11135
rect 13228 11104 13369 11132
rect 13228 11092 13234 11104
rect 13357 11101 13369 11104
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 13556 11104 13860 11132
rect 13556 11064 13584 11104
rect 12452 11036 13584 11064
rect 11422 10996 11428 11008
rect 10376 10968 11284 10996
rect 11383 10968 11428 10996
rect 10376 10956 10382 10968
rect 11422 10956 11428 10968
rect 11480 10956 11486 11008
rect 11698 10956 11704 11008
rect 11756 10996 11762 11008
rect 11793 10999 11851 11005
rect 11793 10996 11805 10999
rect 11756 10968 11805 10996
rect 11756 10956 11762 10968
rect 11793 10965 11805 10968
rect 11839 10996 11851 10999
rect 12894 10996 12900 11008
rect 11839 10968 12900 10996
rect 11839 10965 11851 10968
rect 11793 10959 11851 10965
rect 12894 10956 12900 10968
rect 12952 10996 12958 11008
rect 12989 10999 13047 11005
rect 12989 10996 13001 10999
rect 12952 10968 13001 10996
rect 12952 10956 12958 10968
rect 12989 10965 13001 10968
rect 13035 10965 13047 10999
rect 12989 10959 13047 10965
rect 13354 10956 13360 11008
rect 13412 10996 13418 11008
rect 13541 10999 13599 11005
rect 13541 10996 13553 10999
rect 13412 10968 13553 10996
rect 13412 10956 13418 10968
rect 13541 10965 13553 10968
rect 13587 10996 13599 10999
rect 13630 10996 13636 11008
rect 13587 10968 13636 10996
rect 13587 10965 13599 10968
rect 13541 10959 13599 10965
rect 13630 10956 13636 10968
rect 13688 10956 13694 11008
rect 13832 10996 13860 11104
rect 13906 11092 13912 11144
rect 13964 11132 13970 11144
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 13964 11104 14197 11132
rect 13964 11092 13970 11104
rect 14185 11101 14197 11104
rect 14231 11132 14243 11135
rect 14642 11132 14648 11144
rect 14231 11104 14648 11132
rect 14231 11101 14243 11104
rect 14185 11095 14243 11101
rect 14642 11092 14648 11104
rect 14700 11092 14706 11144
rect 14918 11092 14924 11144
rect 14976 11132 14982 11144
rect 15378 11132 15384 11144
rect 14976 11104 15384 11132
rect 14976 11092 14982 11104
rect 15378 11092 15384 11104
rect 15436 11092 15442 11144
rect 14090 11024 14096 11076
rect 14148 11064 14154 11076
rect 15013 11067 15071 11073
rect 15013 11064 15025 11067
rect 14148 11036 15025 11064
rect 14148 11024 14154 11036
rect 15013 11033 15025 11036
rect 15059 11033 15071 11067
rect 15562 11064 15568 11076
rect 15523 11036 15568 11064
rect 15013 11027 15071 11033
rect 15562 11024 15568 11036
rect 15620 11064 15626 11076
rect 15746 11064 15752 11076
rect 15620 11036 15752 11064
rect 15620 11024 15626 11036
rect 15746 11024 15752 11036
rect 15804 11024 15810 11076
rect 14182 10996 14188 11008
rect 13832 10968 14188 10996
rect 14182 10956 14188 10968
rect 14240 10956 14246 11008
rect 14734 10996 14740 11008
rect 14695 10968 14740 10996
rect 14734 10956 14740 10968
rect 14792 10956 14798 11008
rect 15102 10956 15108 11008
rect 15160 10996 15166 11008
rect 15197 10999 15255 11005
rect 15197 10996 15209 10999
rect 15160 10968 15209 10996
rect 15160 10956 15166 10968
rect 15197 10965 15209 10968
rect 15243 10965 15255 10999
rect 15197 10959 15255 10965
rect 1104 10906 16008 10928
rect 1104 10854 4698 10906
rect 4750 10854 4762 10906
rect 4814 10854 4826 10906
rect 4878 10854 4890 10906
rect 4942 10854 4954 10906
rect 5006 10854 8446 10906
rect 8498 10854 8510 10906
rect 8562 10854 8574 10906
rect 8626 10854 8638 10906
rect 8690 10854 8702 10906
rect 8754 10854 12194 10906
rect 12246 10854 12258 10906
rect 12310 10854 12322 10906
rect 12374 10854 12386 10906
rect 12438 10854 12450 10906
rect 12502 10854 16008 10906
rect 1104 10832 16008 10854
rect 1578 10792 1584 10804
rect 1539 10764 1584 10792
rect 1578 10752 1584 10764
rect 1636 10752 1642 10804
rect 1949 10795 2007 10801
rect 1949 10761 1961 10795
rect 1995 10792 2007 10795
rect 2130 10792 2136 10804
rect 1995 10764 2136 10792
rect 1995 10761 2007 10764
rect 1949 10755 2007 10761
rect 2130 10752 2136 10764
rect 2188 10752 2194 10804
rect 2409 10795 2467 10801
rect 2409 10761 2421 10795
rect 2455 10792 2467 10795
rect 3326 10792 3332 10804
rect 2455 10764 3332 10792
rect 2455 10761 2467 10764
rect 2409 10755 2467 10761
rect 3326 10752 3332 10764
rect 3384 10752 3390 10804
rect 5626 10792 5632 10804
rect 3436 10764 5632 10792
rect 2774 10684 2780 10736
rect 2832 10724 2838 10736
rect 2832 10696 2877 10724
rect 2832 10684 2838 10696
rect 3050 10684 3056 10736
rect 3108 10724 3114 10736
rect 3436 10724 3464 10764
rect 5626 10752 5632 10764
rect 5684 10752 5690 10804
rect 6914 10792 6920 10804
rect 5951 10764 6920 10792
rect 5166 10724 5172 10736
rect 3108 10696 3464 10724
rect 3528 10696 5172 10724
rect 3108 10684 3114 10696
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 2498 10656 2504 10668
rect 2087 10628 2504 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 2498 10616 2504 10628
rect 2556 10616 2562 10668
rect 2869 10659 2927 10665
rect 2869 10625 2881 10659
rect 2915 10656 2927 10659
rect 3329 10659 3387 10665
rect 2915 10628 3188 10656
rect 2915 10625 2927 10628
rect 2869 10619 2927 10625
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10557 1915 10591
rect 2682 10588 2688 10600
rect 2643 10560 2688 10588
rect 1857 10551 1915 10557
rect 1872 10520 1900 10551
rect 2682 10548 2688 10560
rect 2740 10548 2746 10600
rect 3050 10520 3056 10532
rect 1872 10492 3056 10520
rect 3050 10480 3056 10492
rect 3108 10480 3114 10532
rect 3160 10452 3188 10628
rect 3329 10625 3341 10659
rect 3375 10656 3387 10659
rect 3528 10656 3556 10696
rect 5166 10684 5172 10696
rect 5224 10684 5230 10736
rect 5258 10684 5264 10736
rect 5316 10684 5322 10736
rect 5951 10733 5979 10764
rect 6914 10752 6920 10764
rect 6972 10752 6978 10804
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 7064 10764 7144 10792
rect 7064 10752 7070 10764
rect 5936 10727 5994 10733
rect 5936 10693 5948 10727
rect 5982 10693 5994 10727
rect 7116 10724 7144 10764
rect 9122 10752 9128 10804
rect 9180 10792 9186 10804
rect 9677 10795 9735 10801
rect 9677 10792 9689 10795
rect 9180 10764 9689 10792
rect 9180 10752 9186 10764
rect 9677 10761 9689 10764
rect 9723 10761 9735 10795
rect 9677 10755 9735 10761
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10873 10795 10931 10801
rect 10873 10792 10885 10795
rect 10100 10764 10885 10792
rect 10100 10752 10106 10764
rect 10873 10761 10885 10764
rect 10919 10761 10931 10795
rect 10873 10755 10931 10761
rect 10962 10752 10968 10804
rect 11020 10792 11026 10804
rect 11514 10792 11520 10804
rect 11020 10764 11065 10792
rect 11475 10764 11520 10792
rect 11020 10752 11026 10764
rect 11514 10752 11520 10764
rect 11572 10752 11578 10804
rect 11882 10752 11888 10804
rect 11940 10792 11946 10804
rect 11977 10795 12035 10801
rect 11977 10792 11989 10795
rect 11940 10764 11989 10792
rect 11940 10752 11946 10764
rect 11977 10761 11989 10764
rect 12023 10761 12035 10795
rect 11977 10755 12035 10761
rect 12713 10795 12771 10801
rect 12713 10761 12725 10795
rect 12759 10792 12771 10795
rect 12986 10792 12992 10804
rect 12759 10764 12992 10792
rect 12759 10761 12771 10764
rect 12713 10755 12771 10761
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 13170 10752 13176 10804
rect 13228 10792 13234 10804
rect 13998 10792 14004 10804
rect 13228 10764 13860 10792
rect 13959 10764 14004 10792
rect 13228 10752 13234 10764
rect 7837 10727 7895 10733
rect 7837 10724 7849 10727
rect 5936 10687 5994 10693
rect 6104 10696 7052 10724
rect 7116 10696 7849 10724
rect 3375 10628 3556 10656
rect 3596 10659 3654 10665
rect 3375 10625 3387 10628
rect 3329 10619 3387 10625
rect 3596 10625 3608 10659
rect 3642 10656 3654 10659
rect 3878 10656 3884 10668
rect 3642 10628 3884 10656
rect 3642 10625 3654 10628
rect 3596 10619 3654 10625
rect 3878 10616 3884 10628
rect 3936 10616 3942 10668
rect 4798 10616 4804 10668
rect 4856 10656 4862 10668
rect 5276 10656 5304 10684
rect 6104 10656 6132 10696
rect 6638 10665 6644 10668
rect 6632 10656 6644 10665
rect 4856 10628 6132 10656
rect 6599 10628 6644 10656
rect 4856 10616 4862 10628
rect 6632 10619 6644 10628
rect 6638 10616 6644 10619
rect 6696 10616 6702 10668
rect 7024 10656 7052 10696
rect 7837 10693 7849 10696
rect 7883 10693 7895 10727
rect 8938 10724 8944 10736
rect 7837 10687 7895 10693
rect 7944 10696 8944 10724
rect 7944 10656 7972 10696
rect 8938 10684 8944 10696
rect 8996 10684 9002 10736
rect 10980 10724 11008 10752
rect 13354 10724 13360 10736
rect 9048 10696 11008 10724
rect 11900 10696 13360 10724
rect 7024 10628 7972 10656
rect 8110 10616 8116 10668
rect 8168 10656 8174 10668
rect 9048 10656 9076 10696
rect 8168 10628 9076 10656
rect 10045 10659 10103 10665
rect 8168 10616 8174 10628
rect 10045 10625 10057 10659
rect 10091 10656 10103 10659
rect 10870 10656 10876 10668
rect 10091 10628 10876 10656
rect 10091 10625 10103 10628
rect 10045 10619 10103 10625
rect 10870 10616 10876 10628
rect 10928 10656 10934 10668
rect 11146 10656 11152 10668
rect 10928 10628 11152 10656
rect 10928 10616 10934 10628
rect 11146 10616 11152 10628
rect 11204 10616 11210 10668
rect 11900 10665 11928 10696
rect 13354 10684 13360 10696
rect 13412 10724 13418 10736
rect 13725 10727 13783 10733
rect 13725 10724 13737 10727
rect 13412 10696 13737 10724
rect 13412 10684 13418 10696
rect 13725 10693 13737 10696
rect 13771 10693 13783 10727
rect 13832 10724 13860 10764
rect 13998 10752 14004 10764
rect 14056 10752 14062 10804
rect 14090 10752 14096 10804
rect 14148 10792 14154 10804
rect 14148 10764 14193 10792
rect 14148 10752 14154 10764
rect 14274 10752 14280 10804
rect 14332 10792 14338 10804
rect 15102 10792 15108 10804
rect 14332 10764 15108 10792
rect 14332 10752 14338 10764
rect 15102 10752 15108 10764
rect 15160 10792 15166 10804
rect 15289 10795 15347 10801
rect 15289 10792 15301 10795
rect 15160 10764 15301 10792
rect 15160 10752 15166 10764
rect 15289 10761 15301 10764
rect 15335 10761 15347 10795
rect 15289 10755 15347 10761
rect 15473 10795 15531 10801
rect 15473 10761 15485 10795
rect 15519 10792 15531 10795
rect 16206 10792 16212 10804
rect 15519 10764 16212 10792
rect 15519 10761 15531 10764
rect 15473 10755 15531 10761
rect 16206 10752 16212 10764
rect 16264 10752 16270 10804
rect 14366 10724 14372 10736
rect 13832 10696 14372 10724
rect 13725 10687 13783 10693
rect 14366 10684 14372 10696
rect 14424 10724 14430 10736
rect 14829 10727 14887 10733
rect 14829 10724 14841 10727
rect 14424 10696 14841 10724
rect 14424 10684 14430 10696
rect 14829 10693 14841 10696
rect 14875 10693 14887 10727
rect 14829 10687 14887 10693
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 12434 10616 12440 10668
rect 12492 10656 12498 10668
rect 13162 10659 13220 10665
rect 12492 10628 13032 10656
rect 12492 10616 12498 10628
rect 6181 10591 6239 10597
rect 6181 10557 6193 10591
rect 6227 10588 6239 10591
rect 6362 10588 6368 10600
rect 6227 10560 6368 10588
rect 6227 10557 6239 10560
rect 6181 10551 6239 10557
rect 6362 10548 6368 10560
rect 6420 10548 6426 10600
rect 7834 10588 7840 10600
rect 7392 10560 7840 10588
rect 3237 10523 3295 10529
rect 3237 10489 3249 10523
rect 3283 10520 3295 10523
rect 3326 10520 3332 10532
rect 3283 10492 3332 10520
rect 3283 10489 3295 10492
rect 3237 10483 3295 10489
rect 3326 10480 3332 10492
rect 3384 10480 3390 10532
rect 4264 10492 5028 10520
rect 4264 10452 4292 10492
rect 3160 10424 4292 10452
rect 4338 10412 4344 10464
rect 4396 10452 4402 10464
rect 4614 10452 4620 10464
rect 4396 10424 4620 10452
rect 4396 10412 4402 10424
rect 4614 10412 4620 10424
rect 4672 10452 4678 10464
rect 4709 10455 4767 10461
rect 4709 10452 4721 10455
rect 4672 10424 4721 10452
rect 4672 10412 4678 10424
rect 4709 10421 4721 10424
rect 4755 10421 4767 10455
rect 4709 10415 4767 10421
rect 4798 10412 4804 10464
rect 4856 10452 4862 10464
rect 5000 10452 5028 10492
rect 7392 10452 7420 10560
rect 7834 10548 7840 10560
rect 7892 10548 7898 10600
rect 7926 10548 7932 10600
rect 7984 10588 7990 10600
rect 9306 10588 9312 10600
rect 7984 10560 9312 10588
rect 7984 10548 7990 10560
rect 9306 10548 9312 10560
rect 9364 10548 9370 10600
rect 9493 10591 9551 10597
rect 9493 10557 9505 10591
rect 9539 10588 9551 10591
rect 10134 10588 10140 10600
rect 9539 10560 9720 10588
rect 10095 10560 10140 10588
rect 9539 10557 9551 10560
rect 9493 10551 9551 10557
rect 7650 10480 7656 10532
rect 7708 10520 7714 10532
rect 9692 10520 9720 10560
rect 10134 10548 10140 10560
rect 10192 10548 10198 10600
rect 10229 10591 10287 10597
rect 10229 10557 10241 10591
rect 10275 10557 10287 10591
rect 10229 10551 10287 10557
rect 9950 10520 9956 10532
rect 7708 10492 9628 10520
rect 9692 10492 9956 10520
rect 7708 10480 7714 10492
rect 4856 10424 4901 10452
rect 5000 10424 7420 10452
rect 7745 10455 7803 10461
rect 4856 10412 4862 10424
rect 7745 10421 7757 10455
rect 7791 10452 7803 10455
rect 8386 10452 8392 10464
rect 7791 10424 8392 10452
rect 7791 10421 7803 10424
rect 7745 10415 7803 10421
rect 8386 10412 8392 10424
rect 8444 10412 8450 10464
rect 9600 10452 9628 10492
rect 9950 10480 9956 10492
rect 10008 10480 10014 10532
rect 10244 10520 10272 10551
rect 10318 10548 10324 10600
rect 10376 10588 10382 10600
rect 11057 10591 11115 10597
rect 11057 10588 11069 10591
rect 10376 10560 11069 10588
rect 10376 10548 10382 10560
rect 11057 10557 11069 10560
rect 11103 10557 11115 10591
rect 11057 10551 11115 10557
rect 11698 10548 11704 10600
rect 11756 10588 11762 10600
rect 12069 10591 12127 10597
rect 12069 10588 12081 10591
rect 11756 10560 12081 10588
rect 11756 10548 11762 10560
rect 12069 10557 12081 10560
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 12342 10548 12348 10600
rect 12400 10588 12406 10600
rect 13004 10597 13032 10628
rect 13162 10625 13174 10659
rect 13208 10656 13220 10659
rect 13446 10656 13452 10668
rect 13208 10628 13452 10656
rect 13208 10625 13220 10628
rect 13162 10619 13220 10625
rect 13446 10616 13452 10628
rect 13504 10656 13510 10668
rect 14461 10659 14519 10665
rect 14461 10656 14473 10659
rect 13504 10628 14473 10656
rect 13504 10616 13510 10628
rect 14461 10625 14473 10628
rect 14507 10625 14519 10659
rect 14461 10619 14519 10625
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12400 10560 12817 10588
rect 12400 10548 12406 10560
rect 12805 10557 12817 10560
rect 12851 10557 12863 10591
rect 12805 10551 12863 10557
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10557 13047 10591
rect 12989 10551 13047 10557
rect 13357 10591 13415 10597
rect 13357 10557 13369 10591
rect 13403 10557 13415 10591
rect 13357 10551 13415 10557
rect 11882 10520 11888 10532
rect 10060 10492 11888 10520
rect 10060 10452 10088 10492
rect 11882 10480 11888 10492
rect 11940 10480 11946 10532
rect 13372 10520 13400 10551
rect 14090 10548 14096 10600
rect 14148 10588 14154 10600
rect 14550 10588 14556 10600
rect 14148 10560 14556 10588
rect 14148 10548 14154 10560
rect 14550 10548 14556 10560
rect 14608 10588 14614 10600
rect 15013 10591 15071 10597
rect 15013 10588 15025 10591
rect 14608 10560 15025 10588
rect 14608 10548 14614 10560
rect 15013 10557 15025 10560
rect 15059 10557 15071 10591
rect 15013 10551 15071 10557
rect 13446 10520 13452 10532
rect 13372 10492 13452 10520
rect 13446 10480 13452 10492
rect 13504 10480 13510 10532
rect 14182 10480 14188 10532
rect 14240 10520 14246 10532
rect 15565 10523 15623 10529
rect 15565 10520 15577 10523
rect 14240 10492 15577 10520
rect 14240 10480 14246 10492
rect 15565 10489 15577 10492
rect 15611 10520 15623 10523
rect 16574 10520 16580 10532
rect 15611 10492 16580 10520
rect 15611 10489 15623 10492
rect 15565 10483 15623 10489
rect 16574 10480 16580 10492
rect 16632 10480 16638 10532
rect 9600 10424 10088 10452
rect 10134 10412 10140 10464
rect 10192 10452 10198 10464
rect 10505 10455 10563 10461
rect 10505 10452 10517 10455
rect 10192 10424 10517 10452
rect 10192 10412 10198 10424
rect 10505 10421 10517 10424
rect 10551 10421 10563 10455
rect 10505 10415 10563 10421
rect 10686 10412 10692 10464
rect 10744 10452 10750 10464
rect 11514 10452 11520 10464
rect 10744 10424 11520 10452
rect 10744 10412 10750 10424
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 11974 10412 11980 10464
rect 12032 10452 12038 10464
rect 12345 10455 12403 10461
rect 12345 10452 12357 10455
rect 12032 10424 12357 10452
rect 12032 10412 12038 10424
rect 12345 10421 12357 10424
rect 12391 10421 12403 10455
rect 12345 10415 12403 10421
rect 12710 10412 12716 10464
rect 12768 10452 12774 10464
rect 13630 10452 13636 10464
rect 12768 10424 13636 10452
rect 12768 10412 12774 10424
rect 13630 10412 13636 10424
rect 13688 10412 13694 10464
rect 14734 10452 14740 10464
rect 14695 10424 14740 10452
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 1104 10362 16008 10384
rect 1104 10310 2824 10362
rect 2876 10310 2888 10362
rect 2940 10310 2952 10362
rect 3004 10310 3016 10362
rect 3068 10310 3080 10362
rect 3132 10310 6572 10362
rect 6624 10310 6636 10362
rect 6688 10310 6700 10362
rect 6752 10310 6764 10362
rect 6816 10310 6828 10362
rect 6880 10310 10320 10362
rect 10372 10310 10384 10362
rect 10436 10310 10448 10362
rect 10500 10310 10512 10362
rect 10564 10310 10576 10362
rect 10628 10310 14068 10362
rect 14120 10310 14132 10362
rect 14184 10310 14196 10362
rect 14248 10310 14260 10362
rect 14312 10310 14324 10362
rect 14376 10310 16008 10362
rect 1104 10288 16008 10310
rect 6914 10248 6920 10260
rect 1596 10220 6920 10248
rect 1596 10121 1624 10220
rect 6914 10208 6920 10220
rect 6972 10208 6978 10260
rect 8110 10208 8116 10260
rect 8168 10248 8174 10260
rect 8168 10220 9996 10248
rect 8168 10208 8174 10220
rect 2130 10180 2136 10192
rect 2091 10152 2136 10180
rect 2130 10140 2136 10152
rect 2188 10140 2194 10192
rect 3605 10183 3663 10189
rect 3605 10149 3617 10183
rect 3651 10180 3663 10183
rect 4154 10180 4160 10192
rect 3651 10152 4160 10180
rect 3651 10149 3663 10152
rect 3605 10143 3663 10149
rect 4154 10140 4160 10152
rect 4212 10140 4218 10192
rect 5442 10140 5448 10192
rect 5500 10180 5506 10192
rect 7377 10183 7435 10189
rect 7377 10180 7389 10183
rect 5500 10152 7389 10180
rect 5500 10140 5506 10152
rect 7377 10149 7389 10152
rect 7423 10149 7435 10183
rect 7377 10143 7435 10149
rect 1581 10115 1639 10121
rect 1581 10081 1593 10115
rect 1627 10081 1639 10115
rect 1581 10075 1639 10081
rect 1673 10115 1731 10121
rect 1673 10081 1685 10115
rect 1719 10112 1731 10115
rect 1946 10112 1952 10124
rect 1719 10084 1952 10112
rect 1719 10081 1731 10084
rect 1673 10075 1731 10081
rect 1578 9936 1584 9988
rect 1636 9976 1642 9988
rect 1688 9976 1716 10075
rect 1946 10072 1952 10084
rect 2004 10072 2010 10124
rect 5166 10112 5172 10124
rect 5127 10084 5172 10112
rect 5166 10072 5172 10084
rect 5224 10072 5230 10124
rect 7285 10115 7343 10121
rect 7285 10081 7297 10115
rect 7331 10112 7343 10115
rect 7742 10112 7748 10124
rect 7331 10084 7748 10112
rect 7331 10081 7343 10084
rect 7285 10075 7343 10081
rect 7742 10072 7748 10084
rect 7800 10072 7806 10124
rect 8757 10115 8815 10121
rect 8757 10081 8769 10115
rect 8803 10081 8815 10115
rect 8757 10075 8815 10081
rect 2222 10044 2228 10056
rect 2183 10016 2228 10044
rect 2222 10004 2228 10016
rect 2280 10004 2286 10056
rect 3234 10044 3240 10056
rect 2424 10016 3240 10044
rect 2424 9976 2452 10016
rect 3234 10004 3240 10016
rect 3292 10004 3298 10056
rect 4338 10044 4344 10056
rect 3344 10016 4344 10044
rect 1636 9948 1716 9976
rect 1780 9948 2452 9976
rect 2492 9979 2550 9985
rect 1636 9936 1642 9948
rect 1780 9920 1808 9948
rect 2492 9945 2504 9979
rect 2538 9976 2550 9979
rect 2590 9976 2596 9988
rect 2538 9948 2596 9976
rect 2538 9945 2550 9948
rect 2492 9939 2550 9945
rect 2590 9936 2596 9948
rect 2648 9936 2654 9988
rect 2774 9936 2780 9988
rect 2832 9976 2838 9988
rect 3344 9976 3372 10016
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 4614 10004 4620 10056
rect 4672 10044 4678 10056
rect 6730 10044 6736 10056
rect 4672 10016 6736 10044
rect 4672 10004 4678 10016
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 7374 10004 7380 10056
rect 7432 10044 7438 10056
rect 8772 10044 8800 10075
rect 8846 10072 8852 10124
rect 8904 10112 8910 10124
rect 9968 10112 9996 10220
rect 10134 10208 10140 10260
rect 10192 10248 10198 10260
rect 10321 10251 10379 10257
rect 10321 10248 10333 10251
rect 10192 10220 10333 10248
rect 10192 10208 10198 10220
rect 10321 10217 10333 10220
rect 10367 10217 10379 10251
rect 11238 10248 11244 10260
rect 11199 10220 11244 10248
rect 10321 10211 10379 10217
rect 11238 10208 11244 10220
rect 11296 10208 11302 10260
rect 12710 10248 12716 10260
rect 11900 10220 12716 10248
rect 10042 10140 10048 10192
rect 10100 10180 10106 10192
rect 10413 10183 10471 10189
rect 10413 10180 10425 10183
rect 10100 10152 10425 10180
rect 10100 10140 10106 10152
rect 10413 10149 10425 10152
rect 10459 10149 10471 10183
rect 11900 10180 11928 10220
rect 12710 10208 12716 10220
rect 12768 10248 12774 10260
rect 12768 10220 13400 10248
rect 12768 10208 12774 10220
rect 10413 10143 10471 10149
rect 10704 10152 11928 10180
rect 10704 10112 10732 10152
rect 11974 10140 11980 10192
rect 12032 10180 12038 10192
rect 13372 10180 13400 10220
rect 13814 10208 13820 10260
rect 13872 10248 13878 10260
rect 14277 10251 14335 10257
rect 14277 10248 14289 10251
rect 13872 10220 14289 10248
rect 13872 10208 13878 10220
rect 14277 10217 14289 10220
rect 14323 10217 14335 10251
rect 15654 10248 15660 10260
rect 15615 10220 15660 10248
rect 14277 10211 14335 10217
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 12032 10152 12756 10180
rect 13372 10152 13492 10180
rect 12032 10140 12038 10152
rect 8904 10084 9076 10112
rect 9968 10084 10732 10112
rect 8904 10072 8910 10084
rect 8938 10044 8944 10056
rect 7432 10016 8616 10044
rect 8772 10016 8944 10044
rect 7432 10004 7438 10016
rect 2832 9948 3372 9976
rect 2832 9936 2838 9948
rect 3418 9936 3424 9988
rect 3476 9936 3482 9988
rect 4522 9936 4528 9988
rect 4580 9976 4586 9988
rect 4902 9979 4960 9985
rect 4902 9976 4914 9979
rect 4580 9948 4914 9976
rect 4580 9936 4586 9948
rect 4902 9945 4914 9948
rect 4948 9945 4960 9979
rect 4902 9939 4960 9945
rect 5261 9979 5319 9985
rect 5261 9945 5273 9979
rect 5307 9976 5319 9979
rect 5810 9976 5816 9988
rect 5307 9948 5816 9976
rect 5307 9945 5319 9948
rect 5261 9939 5319 9945
rect 5810 9936 5816 9948
rect 5868 9936 5874 9988
rect 5902 9936 5908 9988
rect 5960 9976 5966 9988
rect 5960 9948 8294 9976
rect 5960 9936 5966 9948
rect 1762 9908 1768 9920
rect 1723 9880 1768 9908
rect 1762 9868 1768 9880
rect 1820 9868 1826 9920
rect 2038 9868 2044 9920
rect 2096 9908 2102 9920
rect 3234 9908 3240 9920
rect 2096 9880 3240 9908
rect 2096 9868 2102 9880
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 3436 9908 3464 9936
rect 3789 9911 3847 9917
rect 3789 9908 3801 9911
rect 3436 9880 3801 9908
rect 3789 9877 3801 9880
rect 3835 9908 3847 9911
rect 3878 9908 3884 9920
rect 3835 9880 3884 9908
rect 3835 9877 3847 9880
rect 3789 9871 3847 9877
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 4614 9908 4620 9920
rect 4120 9880 4620 9908
rect 4120 9868 4126 9880
rect 4614 9868 4620 9880
rect 4672 9868 4678 9920
rect 6362 9868 6368 9920
rect 6420 9908 6426 9920
rect 6549 9911 6607 9917
rect 6549 9908 6561 9911
rect 6420 9880 6561 9908
rect 6420 9868 6426 9880
rect 6549 9877 6561 9880
rect 6595 9877 6607 9911
rect 8266 9908 8294 9948
rect 8386 9936 8392 9988
rect 8444 9976 8450 9988
rect 8490 9979 8548 9985
rect 8490 9976 8502 9979
rect 8444 9948 8502 9976
rect 8444 9936 8450 9948
rect 8490 9945 8502 9948
rect 8536 9945 8548 9979
rect 8588 9976 8616 10016
rect 8938 10004 8944 10016
rect 8996 10004 9002 10056
rect 9048 10044 9076 10084
rect 10778 10072 10784 10124
rect 10836 10112 10842 10124
rect 10873 10115 10931 10121
rect 10873 10112 10885 10115
rect 10836 10084 10885 10112
rect 10836 10072 10842 10084
rect 10873 10081 10885 10084
rect 10919 10081 10931 10115
rect 10873 10075 10931 10081
rect 10965 10115 11023 10121
rect 10965 10081 10977 10115
rect 11011 10112 11023 10115
rect 11698 10112 11704 10124
rect 11011 10084 11704 10112
rect 11011 10081 11023 10084
rect 10965 10075 11023 10081
rect 9048 10016 10548 10044
rect 9186 9979 9244 9985
rect 9186 9976 9198 9979
rect 8588 9948 9198 9976
rect 8490 9939 8548 9945
rect 9186 9945 9198 9948
rect 9232 9945 9244 9979
rect 10520 9976 10548 10016
rect 10594 10004 10600 10056
rect 10652 10044 10658 10056
rect 10980 10044 11008 10075
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 11882 10112 11888 10124
rect 11843 10084 11888 10112
rect 11882 10072 11888 10084
rect 11940 10112 11946 10124
rect 12618 10112 12624 10124
rect 11940 10084 12624 10112
rect 11940 10072 11946 10084
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 12728 10112 12756 10152
rect 13078 10112 13084 10124
rect 12728 10084 13084 10112
rect 13078 10072 13084 10084
rect 13136 10112 13142 10124
rect 13464 10121 13492 10152
rect 14182 10140 14188 10192
rect 14240 10180 14246 10192
rect 14461 10183 14519 10189
rect 14461 10180 14473 10183
rect 14240 10152 14473 10180
rect 14240 10140 14246 10152
rect 14461 10149 14473 10152
rect 14507 10180 14519 10183
rect 15197 10183 15255 10189
rect 15197 10180 15209 10183
rect 14507 10152 15209 10180
rect 14507 10149 14519 10152
rect 14461 10143 14519 10149
rect 15197 10149 15209 10152
rect 15243 10149 15255 10183
rect 15197 10143 15255 10149
rect 13449 10115 13507 10121
rect 13136 10084 13400 10112
rect 13136 10072 13142 10084
rect 12437 10047 12495 10053
rect 12437 10044 12449 10047
rect 10652 10016 11008 10044
rect 11072 10016 12449 10044
rect 10652 10004 10658 10016
rect 11072 9976 11100 10016
rect 12437 10013 12449 10016
rect 12483 10013 12495 10047
rect 12437 10007 12495 10013
rect 13170 10004 13176 10056
rect 13228 10044 13234 10056
rect 13265 10047 13323 10053
rect 13265 10044 13277 10047
rect 13228 10016 13277 10044
rect 13228 10004 13234 10016
rect 13265 10013 13277 10016
rect 13311 10013 13323 10047
rect 13372 10044 13400 10084
rect 13449 10081 13461 10115
rect 13495 10081 13507 10115
rect 13449 10075 13507 10081
rect 13630 10072 13636 10124
rect 13688 10112 13694 10124
rect 15013 10115 15071 10121
rect 15013 10112 15025 10115
rect 13688 10084 15025 10112
rect 13688 10072 13694 10084
rect 15013 10081 15025 10084
rect 15059 10081 15071 10115
rect 15013 10075 15071 10081
rect 13725 10047 13783 10053
rect 13725 10044 13737 10047
rect 13372 10016 13737 10044
rect 13265 10007 13323 10013
rect 13725 10013 13737 10016
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 13814 10004 13820 10056
rect 13872 10044 13878 10056
rect 14645 10047 14703 10053
rect 14645 10044 14657 10047
rect 13872 10016 14657 10044
rect 13872 10004 13878 10016
rect 14645 10013 14657 10016
rect 14691 10013 14703 10047
rect 14645 10007 14703 10013
rect 10520 9948 11100 9976
rect 11609 9979 11667 9985
rect 9186 9939 9244 9945
rect 11609 9945 11621 9979
rect 11655 9976 11667 9979
rect 11655 9948 12940 9976
rect 11655 9945 11667 9948
rect 11609 9939 11667 9945
rect 10594 9908 10600 9920
rect 8266 9880 10600 9908
rect 6549 9871 6607 9877
rect 10594 9868 10600 9880
rect 10652 9868 10658 9920
rect 10781 9911 10839 9917
rect 10781 9877 10793 9911
rect 10827 9908 10839 9911
rect 11146 9908 11152 9920
rect 10827 9880 11152 9908
rect 10827 9877 10839 9880
rect 10781 9871 10839 9877
rect 11146 9868 11152 9880
rect 11204 9868 11210 9920
rect 11698 9908 11704 9920
rect 11659 9880 11704 9908
rect 11698 9868 11704 9880
rect 11756 9868 11762 9920
rect 12066 9908 12072 9920
rect 12027 9880 12072 9908
rect 12066 9868 12072 9880
rect 12124 9868 12130 9920
rect 12529 9911 12587 9917
rect 12529 9877 12541 9911
rect 12575 9908 12587 9911
rect 12802 9908 12808 9920
rect 12575 9880 12808 9908
rect 12575 9877 12587 9880
rect 12529 9871 12587 9877
rect 12802 9868 12808 9880
rect 12860 9868 12866 9920
rect 12912 9917 12940 9948
rect 12897 9911 12955 9917
rect 12897 9877 12909 9911
rect 12943 9877 12955 9911
rect 13188 9908 13216 10004
rect 13354 9976 13360 9988
rect 13315 9948 13360 9976
rect 13354 9936 13360 9948
rect 13412 9936 13418 9988
rect 14550 9936 14556 9988
rect 14608 9976 14614 9988
rect 15381 9979 15439 9985
rect 15381 9976 15393 9979
rect 14608 9948 15393 9976
rect 14608 9936 14614 9948
rect 15381 9945 15393 9948
rect 15427 9945 15439 9979
rect 15381 9939 15439 9945
rect 13630 9908 13636 9920
rect 13188 9880 13636 9908
rect 12897 9871 12955 9877
rect 13630 9868 13636 9880
rect 13688 9868 13694 9920
rect 14090 9908 14096 9920
rect 14051 9880 14096 9908
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 14182 9868 14188 9920
rect 14240 9908 14246 9920
rect 14829 9911 14887 9917
rect 14829 9908 14841 9911
rect 14240 9880 14841 9908
rect 14240 9868 14246 9880
rect 14829 9877 14841 9880
rect 14875 9877 14887 9911
rect 14829 9871 14887 9877
rect 1104 9818 16008 9840
rect 1104 9766 4698 9818
rect 4750 9766 4762 9818
rect 4814 9766 4826 9818
rect 4878 9766 4890 9818
rect 4942 9766 4954 9818
rect 5006 9766 8446 9818
rect 8498 9766 8510 9818
rect 8562 9766 8574 9818
rect 8626 9766 8638 9818
rect 8690 9766 8702 9818
rect 8754 9766 12194 9818
rect 12246 9766 12258 9818
rect 12310 9766 12322 9818
rect 12374 9766 12386 9818
rect 12438 9766 12450 9818
rect 12502 9766 16008 9818
rect 1104 9744 16008 9766
rect 2498 9664 2504 9716
rect 2556 9704 2562 9716
rect 4338 9704 4344 9716
rect 2556 9676 4344 9704
rect 2556 9664 2562 9676
rect 4338 9664 4344 9676
rect 4396 9664 4402 9716
rect 4709 9707 4767 9713
rect 4709 9673 4721 9707
rect 4755 9704 4767 9707
rect 6181 9707 6239 9713
rect 4755 9676 6132 9704
rect 4755 9673 4767 9676
rect 4709 9667 4767 9673
rect 1765 9639 1823 9645
rect 1765 9605 1777 9639
rect 1811 9636 1823 9639
rect 5166 9636 5172 9648
rect 1811 9608 3188 9636
rect 1811 9605 1823 9608
rect 1765 9599 1823 9605
rect 1489 9571 1547 9577
rect 1489 9537 1501 9571
rect 1535 9568 1547 9571
rect 2682 9568 2688 9580
rect 1535 9540 2688 9568
rect 1535 9537 1547 9540
rect 1489 9531 1547 9537
rect 2682 9528 2688 9540
rect 2740 9528 2746 9580
rect 2958 9568 2964 9580
rect 3016 9577 3022 9580
rect 2928 9540 2964 9568
rect 2958 9528 2964 9540
rect 3016 9531 3028 9577
rect 3016 9528 3022 9531
rect 3160 9500 3188 9608
rect 3344 9608 5172 9636
rect 3344 9577 3372 9608
rect 3237 9571 3295 9577
rect 3237 9537 3249 9571
rect 3283 9568 3295 9571
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 3283 9540 3341 9568
rect 3283 9537 3295 9540
rect 3237 9531 3295 9537
rect 3329 9537 3341 9540
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 3418 9528 3424 9580
rect 3476 9568 3482 9580
rect 3585 9571 3643 9577
rect 3585 9568 3597 9571
rect 3476 9540 3597 9568
rect 3476 9528 3482 9540
rect 3585 9537 3597 9540
rect 3631 9537 3643 9571
rect 3585 9531 3643 9537
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4430 9568 4436 9580
rect 4212 9540 4436 9568
rect 4212 9528 4218 9540
rect 4430 9528 4436 9540
rect 4488 9568 4494 9580
rect 4816 9577 4844 9608
rect 5166 9596 5172 9608
rect 5224 9596 5230 9648
rect 6104 9636 6132 9676
rect 6181 9673 6193 9707
rect 6227 9704 6239 9707
rect 6227 9676 6675 9704
rect 6227 9673 6239 9676
rect 6181 9667 6239 9673
rect 6454 9636 6460 9648
rect 6104 9608 6460 9636
rect 6454 9596 6460 9608
rect 6512 9596 6518 9648
rect 4801 9571 4859 9577
rect 4488 9540 4752 9568
rect 4488 9528 4494 9540
rect 4724 9500 4752 9540
rect 4801 9537 4813 9571
rect 4847 9537 4859 9571
rect 5057 9571 5115 9577
rect 5057 9568 5069 9571
rect 4801 9531 4859 9537
rect 4908 9540 5069 9568
rect 4908 9500 4936 9540
rect 5057 9537 5069 9540
rect 5103 9537 5115 9571
rect 6362 9568 6368 9580
rect 6323 9540 6368 9568
rect 5057 9531 5115 9537
rect 6362 9528 6368 9540
rect 6420 9528 6426 9580
rect 6647 9577 6675 9676
rect 6914 9664 6920 9716
rect 6972 9704 6978 9716
rect 7837 9707 7895 9713
rect 7837 9704 7849 9707
rect 6972 9676 7849 9704
rect 6972 9664 6978 9676
rect 7837 9673 7849 9676
rect 7883 9673 7895 9707
rect 7837 9667 7895 9673
rect 7926 9664 7932 9716
rect 7984 9704 7990 9716
rect 9030 9704 9036 9716
rect 7984 9676 9036 9704
rect 7984 9664 7990 9676
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 9858 9664 9864 9716
rect 9916 9704 9922 9716
rect 11422 9704 11428 9716
rect 9916 9676 11428 9704
rect 9916 9664 9922 9676
rect 11422 9664 11428 9676
rect 11480 9664 11486 9716
rect 11808 9676 12388 9704
rect 6730 9596 6736 9648
rect 6788 9636 6794 9648
rect 7374 9636 7380 9648
rect 6788 9608 7380 9636
rect 6788 9596 6794 9608
rect 7374 9596 7380 9608
rect 7432 9596 7438 9648
rect 7742 9596 7748 9648
rect 7800 9636 7806 9648
rect 9576 9639 9634 9645
rect 9576 9636 9588 9639
rect 7800 9608 9588 9636
rect 7800 9596 7806 9608
rect 9576 9605 9588 9608
rect 9622 9636 9634 9639
rect 11057 9639 11115 9645
rect 9622 9608 11008 9636
rect 9622 9605 9634 9608
rect 9576 9599 9634 9605
rect 6632 9571 6690 9577
rect 6632 9537 6644 9571
rect 6678 9568 6690 9571
rect 8202 9568 8208 9580
rect 6678 9540 8208 9568
rect 6678 9537 6690 9540
rect 6632 9531 6690 9537
rect 8202 9528 8208 9540
rect 8260 9528 8266 9580
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 8950 9571 9008 9577
rect 8950 9568 8962 9571
rect 8720 9540 8962 9568
rect 8720 9528 8726 9540
rect 8950 9537 8962 9540
rect 8996 9537 9008 9571
rect 8950 9531 9008 9537
rect 9122 9528 9128 9580
rect 9180 9568 9186 9580
rect 9217 9571 9275 9577
rect 9217 9568 9229 9571
rect 9180 9540 9229 9568
rect 9180 9528 9186 9540
rect 9217 9537 9229 9540
rect 9263 9568 9275 9571
rect 9309 9571 9367 9577
rect 9309 9568 9321 9571
rect 9263 9540 9321 9568
rect 9263 9537 9275 9540
rect 9217 9531 9275 9537
rect 9309 9537 9321 9540
rect 9355 9537 9367 9571
rect 9309 9531 9367 9537
rect 9950 9528 9956 9580
rect 10008 9568 10014 9580
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 10008 9540 10793 9568
rect 10008 9528 10014 9540
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 10980 9568 11008 9608
rect 11057 9605 11069 9639
rect 11103 9636 11115 9639
rect 11808 9636 11836 9676
rect 11103 9608 11836 9636
rect 11885 9639 11943 9645
rect 11103 9605 11115 9608
rect 11057 9599 11115 9605
rect 11885 9605 11897 9639
rect 11931 9605 11943 9639
rect 11885 9599 11943 9605
rect 10980 9540 11192 9568
rect 10781 9531 10839 9537
rect 3160 9472 3280 9500
rect 4724 9472 4936 9500
rect 1670 9392 1676 9444
rect 1728 9432 1734 9444
rect 1854 9432 1860 9444
rect 1728 9404 1860 9432
rect 1728 9392 1734 9404
rect 1854 9392 1860 9404
rect 1912 9392 1918 9444
rect 3252 9364 3280 9472
rect 10594 9460 10600 9512
rect 10652 9500 10658 9512
rect 11164 9500 11192 9540
rect 11422 9528 11428 9580
rect 11480 9568 11486 9580
rect 11900 9568 11928 9599
rect 11480 9540 11928 9568
rect 12360 9568 12388 9676
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 12713 9707 12771 9713
rect 12713 9704 12725 9707
rect 12584 9676 12725 9704
rect 12584 9664 12590 9676
rect 12713 9673 12725 9676
rect 12759 9704 12771 9707
rect 13354 9704 13360 9716
rect 12759 9676 13360 9704
rect 12759 9673 12771 9676
rect 12713 9667 12771 9673
rect 13354 9664 13360 9676
rect 13412 9704 13418 9716
rect 14182 9704 14188 9716
rect 13412 9676 14188 9704
rect 13412 9664 13418 9676
rect 14182 9664 14188 9676
rect 14240 9664 14246 9716
rect 14369 9707 14427 9713
rect 14369 9673 14381 9707
rect 14415 9704 14427 9707
rect 14734 9704 14740 9716
rect 14415 9676 14740 9704
rect 14415 9673 14427 9676
rect 14369 9667 14427 9673
rect 14734 9664 14740 9676
rect 14792 9664 14798 9716
rect 14826 9664 14832 9716
rect 14884 9704 14890 9716
rect 14884 9676 14929 9704
rect 14884 9664 14890 9676
rect 15102 9664 15108 9716
rect 15160 9704 15166 9716
rect 15289 9707 15347 9713
rect 15289 9704 15301 9707
rect 15160 9676 15301 9704
rect 15160 9664 15166 9676
rect 15289 9673 15301 9676
rect 15335 9673 15347 9707
rect 15289 9667 15347 9673
rect 12434 9596 12440 9648
rect 12492 9636 12498 9648
rect 13541 9639 13599 9645
rect 13541 9636 13553 9639
rect 12492 9608 13553 9636
rect 12492 9596 12498 9608
rect 13541 9605 13553 9608
rect 13587 9605 13599 9639
rect 13541 9599 13599 9605
rect 13740 9608 15424 9636
rect 12526 9568 12532 9580
rect 12360 9540 12532 9568
rect 11480 9528 11486 9540
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 12805 9571 12863 9577
rect 12805 9537 12817 9571
rect 12851 9568 12863 9571
rect 12986 9568 12992 9580
rect 12851 9540 12992 9568
rect 12851 9537 12863 9540
rect 12805 9531 12863 9537
rect 12986 9528 12992 9540
rect 13044 9568 13050 9580
rect 13446 9568 13452 9580
rect 13044 9540 13452 9568
rect 13044 9528 13050 9540
rect 13446 9528 13452 9540
rect 13504 9528 13510 9580
rect 10652 9472 11100 9500
rect 11164 9472 11652 9500
rect 10652 9460 10658 9472
rect 7650 9392 7656 9444
rect 7708 9432 7714 9444
rect 7745 9435 7803 9441
rect 7745 9432 7757 9435
rect 7708 9404 7757 9432
rect 7708 9392 7714 9404
rect 7745 9401 7757 9404
rect 7791 9401 7803 9435
rect 10778 9432 10784 9444
rect 7745 9395 7803 9401
rect 10244 9404 10784 9432
rect 4246 9364 4252 9376
rect 3252 9336 4252 9364
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 4430 9324 4436 9376
rect 4488 9364 4494 9376
rect 5442 9364 5448 9376
rect 4488 9336 5448 9364
rect 4488 9324 4494 9336
rect 5442 9324 5448 9336
rect 5500 9324 5506 9376
rect 5810 9324 5816 9376
rect 5868 9364 5874 9376
rect 7098 9364 7104 9376
rect 5868 9336 7104 9364
rect 5868 9324 5874 9336
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 8938 9324 8944 9376
rect 8996 9364 9002 9376
rect 9674 9364 9680 9376
rect 8996 9336 9680 9364
rect 8996 9324 9002 9336
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 9950 9324 9956 9376
rect 10008 9364 10014 9376
rect 10244 9364 10272 9404
rect 10778 9392 10784 9404
rect 10836 9392 10842 9444
rect 10686 9364 10692 9376
rect 10008 9336 10272 9364
rect 10647 9336 10692 9364
rect 10008 9324 10014 9336
rect 10686 9324 10692 9336
rect 10744 9324 10750 9376
rect 11072 9364 11100 9472
rect 11517 9367 11575 9373
rect 11517 9364 11529 9367
rect 11072 9336 11529 9364
rect 11517 9333 11529 9336
rect 11563 9333 11575 9367
rect 11624 9364 11652 9472
rect 11882 9460 11888 9512
rect 11940 9500 11946 9512
rect 11977 9503 12035 9509
rect 11977 9500 11989 9503
rect 11940 9472 11989 9500
rect 11940 9460 11946 9472
rect 11977 9469 11989 9472
rect 12023 9469 12035 9503
rect 11977 9463 12035 9469
rect 12066 9460 12072 9512
rect 12124 9500 12130 9512
rect 12894 9500 12900 9512
rect 12124 9472 12169 9500
rect 12855 9472 12900 9500
rect 12124 9460 12130 9472
rect 12894 9460 12900 9472
rect 12952 9460 12958 9512
rect 13078 9460 13084 9512
rect 13136 9500 13142 9512
rect 13633 9503 13691 9509
rect 13633 9500 13645 9503
rect 13136 9472 13645 9500
rect 13136 9460 13142 9472
rect 13633 9469 13645 9472
rect 13679 9469 13691 9503
rect 13633 9463 13691 9469
rect 11790 9392 11796 9444
rect 11848 9432 11854 9444
rect 12345 9435 12403 9441
rect 12345 9432 12357 9435
rect 11848 9404 12357 9432
rect 11848 9392 11854 9404
rect 12345 9401 12357 9404
rect 12391 9401 12403 9435
rect 13740 9432 13768 9608
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9568 14519 9571
rect 14642 9568 14648 9580
rect 14507 9540 14648 9568
rect 14507 9537 14519 9540
rect 14461 9531 14519 9537
rect 14642 9528 14648 9540
rect 14700 9528 14706 9580
rect 14826 9528 14832 9580
rect 14884 9568 14890 9580
rect 15197 9571 15255 9577
rect 15197 9568 15209 9571
rect 14884 9540 15209 9568
rect 14884 9528 14890 9540
rect 15197 9537 15209 9540
rect 15243 9537 15255 9571
rect 15197 9531 15255 9537
rect 13817 9503 13875 9509
rect 13817 9469 13829 9503
rect 13863 9469 13875 9503
rect 14550 9500 14556 9512
rect 14511 9472 14556 9500
rect 13817 9463 13875 9469
rect 12345 9395 12403 9401
rect 12452 9404 13768 9432
rect 12452 9364 12480 9404
rect 13170 9364 13176 9376
rect 11624 9336 12480 9364
rect 13131 9336 13176 9364
rect 11517 9327 11575 9333
rect 13170 9324 13176 9336
rect 13228 9324 13234 9376
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 13832 9364 13860 9463
rect 14550 9460 14556 9472
rect 14608 9460 14614 9512
rect 15396 9509 15424 9608
rect 15381 9503 15439 9509
rect 15381 9469 15393 9503
rect 15427 9469 15439 9503
rect 15381 9463 15439 9469
rect 14458 9392 14464 9444
rect 14516 9432 14522 9444
rect 14826 9432 14832 9444
rect 14516 9404 14832 9432
rect 14516 9392 14522 9404
rect 14826 9392 14832 9404
rect 14884 9392 14890 9444
rect 13780 9336 13860 9364
rect 14001 9367 14059 9373
rect 13780 9324 13786 9336
rect 14001 9333 14013 9367
rect 14047 9364 14059 9367
rect 15286 9364 15292 9376
rect 14047 9336 15292 9364
rect 14047 9333 14059 9336
rect 14001 9327 14059 9333
rect 15286 9324 15292 9336
rect 15344 9324 15350 9376
rect 1104 9274 16008 9296
rect 1104 9222 2824 9274
rect 2876 9222 2888 9274
rect 2940 9222 2952 9274
rect 3004 9222 3016 9274
rect 3068 9222 3080 9274
rect 3132 9222 6572 9274
rect 6624 9222 6636 9274
rect 6688 9222 6700 9274
rect 6752 9222 6764 9274
rect 6816 9222 6828 9274
rect 6880 9222 10320 9274
rect 10372 9222 10384 9274
rect 10436 9222 10448 9274
rect 10500 9222 10512 9274
rect 10564 9222 10576 9274
rect 10628 9222 14068 9274
rect 14120 9222 14132 9274
rect 14184 9222 14196 9274
rect 14248 9222 14260 9274
rect 14312 9222 14324 9274
rect 14376 9222 16008 9274
rect 1104 9200 16008 9222
rect 3510 9160 3516 9172
rect 1596 9132 3516 9160
rect 1596 9033 1624 9132
rect 3510 9120 3516 9132
rect 3568 9120 3574 9172
rect 3786 9120 3792 9172
rect 3844 9160 3850 9172
rect 4246 9160 4252 9172
rect 3844 9132 4252 9160
rect 3844 9120 3850 9132
rect 4246 9120 4252 9132
rect 4304 9120 4310 9172
rect 4614 9120 4620 9172
rect 4672 9160 4678 9172
rect 6914 9160 6920 9172
rect 4672 9132 6920 9160
rect 4672 9120 4678 9132
rect 6914 9120 6920 9132
rect 6972 9120 6978 9172
rect 8941 9163 8999 9169
rect 8941 9129 8953 9163
rect 8987 9160 8999 9163
rect 9030 9160 9036 9172
rect 8987 9132 9036 9160
rect 8987 9129 8999 9132
rect 8941 9123 8999 9129
rect 9030 9120 9036 9132
rect 9088 9120 9094 9172
rect 9398 9120 9404 9172
rect 9456 9160 9462 9172
rect 10413 9163 10471 9169
rect 10413 9160 10425 9163
rect 9456 9132 10425 9160
rect 9456 9120 9462 9132
rect 10413 9129 10425 9132
rect 10459 9129 10471 9163
rect 11238 9160 11244 9172
rect 11199 9132 11244 9160
rect 10413 9123 10471 9129
rect 11238 9120 11244 9132
rect 11296 9120 11302 9172
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 12069 9163 12127 9169
rect 12069 9160 12081 9163
rect 11756 9132 12081 9160
rect 11756 9120 11762 9132
rect 12069 9129 12081 9132
rect 12115 9129 12127 9163
rect 14550 9160 14556 9172
rect 12069 9123 12127 9129
rect 12176 9132 14556 9160
rect 2130 9092 2136 9104
rect 2091 9064 2136 9092
rect 2130 9052 2136 9064
rect 2188 9052 2194 9104
rect 3605 9095 3663 9101
rect 3605 9061 3617 9095
rect 3651 9092 3663 9095
rect 3878 9092 3884 9104
rect 3651 9064 3884 9092
rect 3651 9061 3663 9064
rect 3605 9055 3663 9061
rect 3878 9052 3884 9064
rect 3936 9052 3942 9104
rect 5902 9092 5908 9104
rect 5863 9064 5908 9092
rect 5902 9052 5908 9064
rect 5960 9052 5966 9104
rect 6178 9052 6184 9104
rect 6236 9052 6242 9104
rect 10686 9052 10692 9104
rect 10744 9092 10750 9104
rect 12176 9092 12204 9132
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 14921 9163 14979 9169
rect 14921 9129 14933 9163
rect 14967 9160 14979 9163
rect 15470 9160 15476 9172
rect 14967 9132 15476 9160
rect 14967 9129 14979 9132
rect 14921 9123 14979 9129
rect 15470 9120 15476 9132
rect 15528 9120 15534 9172
rect 12894 9092 12900 9104
rect 10744 9064 12204 9092
rect 12855 9064 12900 9092
rect 10744 9052 10750 9064
rect 12894 9052 12900 9064
rect 12952 9052 12958 9104
rect 13630 9052 13636 9104
rect 13688 9092 13694 9104
rect 14093 9095 14151 9101
rect 13688 9064 13768 9092
rect 13688 9052 13694 9064
rect 1581 9027 1639 9033
rect 1581 8993 1593 9027
rect 1627 8993 1639 9027
rect 1581 8987 1639 8993
rect 1670 8984 1676 9036
rect 1728 9024 1734 9036
rect 2222 9024 2228 9036
rect 1728 8996 1773 9024
rect 2183 8996 2228 9024
rect 1728 8984 1734 8996
rect 2222 8984 2228 8996
rect 2280 8984 2286 9036
rect 3970 9024 3976 9036
rect 3931 8996 3976 9024
rect 3970 8984 3976 8996
rect 4028 8984 4034 9036
rect 6196 9024 6224 9052
rect 5727 8996 6224 9024
rect 1118 8916 1124 8968
rect 1176 8956 1182 8968
rect 2481 8959 2539 8965
rect 2481 8956 2493 8959
rect 1176 8928 2493 8956
rect 1176 8916 1182 8928
rect 2481 8925 2493 8928
rect 2527 8925 2539 8959
rect 2481 8919 2539 8925
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8925 3847 8959
rect 5534 8956 5540 8968
rect 5592 8965 5598 8968
rect 3789 8919 3847 8925
rect 3988 8928 5212 8956
rect 5504 8928 5540 8956
rect 3142 8848 3148 8900
rect 3200 8888 3206 8900
rect 3804 8888 3832 8919
rect 3200 8860 3832 8888
rect 3200 8848 3206 8860
rect 1765 8823 1823 8829
rect 1765 8789 1777 8823
rect 1811 8820 1823 8823
rect 3988 8820 4016 8928
rect 1811 8792 4016 8820
rect 1811 8789 1823 8792
rect 1765 8783 1823 8789
rect 4246 8780 4252 8832
rect 4304 8820 4310 8832
rect 4433 8823 4491 8829
rect 4433 8820 4445 8823
rect 4304 8792 4445 8820
rect 4304 8780 4310 8792
rect 4433 8789 4445 8792
rect 4479 8820 4491 8823
rect 5074 8820 5080 8832
rect 4479 8792 5080 8820
rect 4479 8789 4491 8792
rect 4433 8783 4491 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 5184 8820 5212 8928
rect 5534 8916 5540 8928
rect 5592 8919 5604 8965
rect 5727 8956 5755 8996
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 10965 9027 11023 9033
rect 10965 9024 10977 9027
rect 8444 8996 9260 9024
rect 8444 8984 8450 8996
rect 5644 8928 5755 8956
rect 5813 8959 5871 8965
rect 5592 8916 5598 8919
rect 5644 8820 5672 8928
rect 5813 8925 5825 8959
rect 5859 8956 5871 8959
rect 6178 8956 6184 8968
rect 5859 8928 6184 8956
rect 5859 8925 5871 8928
rect 5813 8919 5871 8925
rect 6178 8916 6184 8928
rect 6236 8956 6242 8968
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 6236 8928 7297 8956
rect 6236 8916 6242 8928
rect 7285 8925 7297 8928
rect 7331 8956 7343 8959
rect 7377 8959 7435 8965
rect 7377 8956 7389 8959
rect 7331 8928 7389 8956
rect 7331 8925 7343 8928
rect 7285 8919 7343 8925
rect 7377 8925 7389 8928
rect 7423 8956 7435 8959
rect 9122 8956 9128 8968
rect 7423 8928 9128 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 9232 8956 9260 8996
rect 10244 8996 10977 9024
rect 9490 8956 9496 8968
rect 9232 8928 9496 8956
rect 9490 8916 9496 8928
rect 9548 8956 9554 8968
rect 10244 8956 10272 8996
rect 10965 8993 10977 8996
rect 11011 8993 11023 9027
rect 11882 9024 11888 9036
rect 11843 8996 11888 9024
rect 10965 8987 11023 8993
rect 11882 8984 11888 8996
rect 11940 8984 11946 9036
rect 12710 9024 12716 9036
rect 12671 8996 12716 9024
rect 12710 8984 12716 8996
rect 12768 8984 12774 9036
rect 13262 8984 13268 9036
rect 13320 9024 13326 9036
rect 13357 9027 13415 9033
rect 13357 9024 13369 9027
rect 13320 8996 13369 9024
rect 13320 8984 13326 8996
rect 13357 8993 13369 8996
rect 13403 8993 13415 9027
rect 13357 8987 13415 8993
rect 13541 9027 13599 9033
rect 13541 8993 13553 9027
rect 13587 9024 13599 9027
rect 13740 9024 13768 9064
rect 14093 9061 14105 9095
rect 14139 9092 14151 9095
rect 14458 9092 14464 9104
rect 14139 9064 14464 9092
rect 14139 9061 14151 9064
rect 14093 9055 14151 9061
rect 14458 9052 14464 9064
rect 14516 9052 14522 9104
rect 14568 9092 14596 9120
rect 14568 9064 14688 9092
rect 14550 9024 14556 9036
rect 13587 8996 13676 9024
rect 13740 8996 14556 9024
rect 13587 8993 13599 8996
rect 13541 8987 13599 8993
rect 9548 8928 10272 8956
rect 10321 8959 10379 8965
rect 9548 8916 9554 8928
rect 10321 8925 10333 8959
rect 10367 8956 10379 8959
rect 10502 8956 10508 8968
rect 10367 8928 10508 8956
rect 10367 8925 10379 8928
rect 10321 8919 10379 8925
rect 10502 8916 10508 8928
rect 10560 8916 10566 8968
rect 10778 8916 10784 8968
rect 10836 8956 10842 8968
rect 10873 8959 10931 8965
rect 10873 8956 10885 8959
rect 10836 8928 10885 8956
rect 10836 8916 10842 8928
rect 10873 8925 10885 8928
rect 10919 8925 10931 8959
rect 10873 8919 10931 8925
rect 11054 8916 11060 8968
rect 11112 8956 11118 8968
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 11112 8928 11621 8956
rect 11112 8916 11118 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 11790 8916 11796 8968
rect 11848 8956 11854 8968
rect 12066 8956 12072 8968
rect 11848 8928 12072 8956
rect 11848 8916 11854 8928
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 12158 8916 12164 8968
rect 12216 8956 12222 8968
rect 12437 8959 12495 8965
rect 12437 8956 12449 8959
rect 12216 8928 12449 8956
rect 12216 8916 12222 8928
rect 12437 8925 12449 8928
rect 12483 8956 12495 8959
rect 12802 8956 12808 8968
rect 12483 8928 12808 8956
rect 12483 8925 12495 8928
rect 12437 8919 12495 8925
rect 12802 8916 12808 8928
rect 12860 8916 12866 8968
rect 13648 8956 13676 8996
rect 14550 8984 14556 8996
rect 14608 8984 14614 9036
rect 14660 9033 14688 9064
rect 14826 9052 14832 9104
rect 14884 9092 14890 9104
rect 15286 9092 15292 9104
rect 14884 9064 15292 9092
rect 14884 9052 14890 9064
rect 15286 9052 15292 9064
rect 15344 9052 15350 9104
rect 16114 9092 16120 9104
rect 15396 9064 16120 9092
rect 15396 9033 15424 9064
rect 16114 9052 16120 9064
rect 16172 9092 16178 9104
rect 16574 9092 16580 9104
rect 16172 9064 16580 9092
rect 16172 9052 16178 9064
rect 16574 9052 16580 9064
rect 16632 9052 16638 9104
rect 14645 9027 14703 9033
rect 14645 8993 14657 9027
rect 14691 8993 14703 9027
rect 14645 8987 14703 8993
rect 15381 9027 15439 9033
rect 15381 8993 15393 9027
rect 15427 8993 15439 9027
rect 15381 8987 15439 8993
rect 15473 9027 15531 9033
rect 15473 8993 15485 9027
rect 15519 8993 15531 9027
rect 15473 8987 15531 8993
rect 15488 8956 15516 8987
rect 13648 8928 15516 8956
rect 7006 8848 7012 8900
rect 7064 8897 7070 8900
rect 7064 8888 7076 8897
rect 7064 8860 7109 8888
rect 7064 8851 7076 8860
rect 7064 8848 7070 8851
rect 7190 8848 7196 8900
rect 7248 8888 7254 8900
rect 7622 8891 7680 8897
rect 7622 8888 7634 8891
rect 7248 8860 7634 8888
rect 7248 8848 7254 8860
rect 7622 8857 7634 8860
rect 7668 8857 7680 8891
rect 7622 8851 7680 8857
rect 8220 8860 8984 8888
rect 5184 8792 5672 8820
rect 5718 8780 5724 8832
rect 5776 8820 5782 8832
rect 8220 8820 8248 8860
rect 5776 8792 8248 8820
rect 8757 8823 8815 8829
rect 5776 8780 5782 8792
rect 8757 8789 8769 8823
rect 8803 8820 8815 8823
rect 8846 8820 8852 8832
rect 8803 8792 8852 8820
rect 8803 8789 8815 8792
rect 8757 8783 8815 8789
rect 8846 8780 8852 8792
rect 8904 8780 8910 8832
rect 8956 8820 8984 8860
rect 9674 8848 9680 8900
rect 9732 8888 9738 8900
rect 10076 8891 10134 8897
rect 10076 8888 10088 8891
rect 9732 8860 10088 8888
rect 9732 8848 9738 8860
rect 10076 8857 10088 8860
rect 10122 8888 10134 8891
rect 10226 8888 10232 8900
rect 10122 8860 10232 8888
rect 10122 8857 10134 8860
rect 10076 8851 10134 8857
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 11701 8891 11759 8897
rect 11701 8888 11713 8891
rect 10428 8860 11713 8888
rect 10428 8820 10456 8860
rect 11701 8857 11713 8860
rect 11747 8857 11759 8891
rect 11701 8851 11759 8857
rect 12529 8891 12587 8897
rect 12529 8857 12541 8891
rect 12575 8888 12587 8891
rect 13078 8888 13084 8900
rect 12575 8860 13084 8888
rect 12575 8857 12587 8860
rect 12529 8851 12587 8857
rect 13078 8848 13084 8860
rect 13136 8848 13142 8900
rect 13265 8891 13323 8897
rect 13265 8857 13277 8891
rect 13311 8888 13323 8891
rect 13538 8888 13544 8900
rect 13311 8860 13544 8888
rect 13311 8857 13323 8860
rect 13265 8851 13323 8857
rect 13538 8848 13544 8860
rect 13596 8848 13602 8900
rect 10778 8820 10784 8832
rect 8956 8792 10456 8820
rect 10739 8792 10784 8820
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 11238 8780 11244 8832
rect 11296 8820 11302 8832
rect 13648 8820 13676 8928
rect 14461 8891 14519 8897
rect 14461 8857 14473 8891
rect 14507 8888 14519 8891
rect 15654 8888 15660 8900
rect 14507 8860 15660 8888
rect 14507 8857 14519 8860
rect 14461 8851 14519 8857
rect 15654 8848 15660 8860
rect 15712 8848 15718 8900
rect 11296 8792 13676 8820
rect 13725 8823 13783 8829
rect 11296 8780 11302 8792
rect 13725 8789 13737 8823
rect 13771 8820 13783 8823
rect 13814 8820 13820 8832
rect 13771 8792 13820 8820
rect 13771 8789 13783 8792
rect 13725 8783 13783 8789
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 15289 8823 15347 8829
rect 15289 8789 15301 8823
rect 15335 8820 15347 8823
rect 16206 8820 16212 8832
rect 15335 8792 16212 8820
rect 15335 8789 15347 8792
rect 15289 8783 15347 8789
rect 16206 8780 16212 8792
rect 16264 8820 16270 8832
rect 16390 8820 16396 8832
rect 16264 8792 16396 8820
rect 16264 8780 16270 8792
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 1104 8730 16008 8752
rect 1104 8678 4698 8730
rect 4750 8678 4762 8730
rect 4814 8678 4826 8730
rect 4878 8678 4890 8730
rect 4942 8678 4954 8730
rect 5006 8678 8446 8730
rect 8498 8678 8510 8730
rect 8562 8678 8574 8730
rect 8626 8678 8638 8730
rect 8690 8678 8702 8730
rect 8754 8678 12194 8730
rect 12246 8678 12258 8730
rect 12310 8678 12322 8730
rect 12374 8678 12386 8730
rect 12438 8678 12450 8730
rect 12502 8678 16008 8730
rect 1104 8656 16008 8678
rect 1857 8619 1915 8625
rect 1857 8585 1869 8619
rect 1903 8616 1915 8619
rect 2406 8616 2412 8628
rect 1903 8588 2412 8616
rect 1903 8585 1915 8588
rect 1857 8579 1915 8585
rect 2406 8576 2412 8588
rect 2464 8576 2470 8628
rect 3326 8616 3332 8628
rect 3160 8588 3332 8616
rect 2992 8551 3050 8557
rect 2992 8517 3004 8551
rect 3038 8548 3050 8551
rect 3160 8548 3188 8588
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 4801 8619 4859 8625
rect 4801 8585 4813 8619
rect 4847 8616 4859 8619
rect 5994 8616 6000 8628
rect 4847 8588 6000 8616
rect 4847 8585 4859 8588
rect 4801 8579 4859 8585
rect 3038 8520 3188 8548
rect 3252 8520 4752 8548
rect 3038 8517 3050 8520
rect 2992 8511 3050 8517
rect 1765 8483 1823 8489
rect 1765 8449 1777 8483
rect 1811 8480 1823 8483
rect 1946 8480 1952 8492
rect 1811 8452 1952 8480
rect 1811 8449 1823 8452
rect 1765 8443 1823 8449
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 3252 8489 3280 8520
rect 4724 8492 4752 8520
rect 3237 8483 3295 8489
rect 3237 8449 3249 8483
rect 3283 8449 3295 8483
rect 4154 8480 4160 8492
rect 3237 8443 3295 8449
rect 3344 8452 4160 8480
rect 1394 8304 1400 8356
rect 1452 8344 1458 8356
rect 3344 8353 3372 8452
rect 4154 8440 4160 8452
rect 4212 8440 4218 8492
rect 4430 8480 4436 8492
rect 4488 8489 4494 8492
rect 4400 8452 4436 8480
rect 4430 8440 4436 8452
rect 4488 8443 4500 8489
rect 4488 8440 4494 8443
rect 4706 8440 4712 8492
rect 4764 8480 4770 8492
rect 4764 8452 4809 8480
rect 4764 8440 4770 8452
rect 1581 8347 1639 8353
rect 1581 8344 1593 8347
rect 1452 8316 1593 8344
rect 1452 8304 1458 8316
rect 1581 8313 1593 8316
rect 1627 8313 1639 8347
rect 1581 8307 1639 8313
rect 3329 8347 3387 8353
rect 3329 8313 3341 8347
rect 3375 8313 3387 8347
rect 3329 8307 3387 8313
rect 2590 8236 2596 8288
rect 2648 8276 2654 8288
rect 3418 8276 3424 8288
rect 2648 8248 3424 8276
rect 2648 8236 2654 8248
rect 3418 8236 3424 8248
rect 3476 8276 3482 8288
rect 4908 8276 4936 8588
rect 5994 8576 6000 8588
rect 6052 8576 6058 8628
rect 7742 8616 7748 8628
rect 7703 8588 7748 8616
rect 7742 8576 7748 8588
rect 7800 8576 7806 8628
rect 9122 8616 9128 8628
rect 9083 8588 9128 8616
rect 9122 8576 9128 8588
rect 9180 8576 9186 8628
rect 11238 8616 11244 8628
rect 9600 8588 11244 8616
rect 5810 8508 5816 8560
rect 5868 8548 5874 8560
rect 6610 8551 6668 8557
rect 6610 8548 6622 8551
rect 5868 8520 6622 8548
rect 5868 8508 5874 8520
rect 6610 8517 6622 8520
rect 6656 8517 6668 8551
rect 6610 8511 6668 8517
rect 7006 8508 7012 8560
rect 7064 8548 7070 8560
rect 9600 8548 9628 8588
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 11514 8616 11520 8628
rect 11475 8588 11520 8616
rect 11514 8576 11520 8588
rect 11572 8576 11578 8628
rect 11790 8576 11796 8628
rect 11848 8616 11854 8628
rect 11977 8619 12035 8625
rect 11977 8616 11989 8619
rect 11848 8588 11989 8616
rect 11848 8576 11854 8588
rect 11977 8585 11989 8588
rect 12023 8585 12035 8619
rect 12345 8619 12403 8625
rect 12345 8616 12357 8619
rect 11977 8579 12035 8585
rect 12176 8588 12357 8616
rect 12176 8560 12204 8588
rect 12345 8585 12357 8588
rect 12391 8585 12403 8619
rect 13170 8616 13176 8628
rect 13131 8588 13176 8616
rect 12345 8579 12403 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13541 8619 13599 8625
rect 13541 8585 13553 8619
rect 13587 8616 13599 8619
rect 13906 8616 13912 8628
rect 13587 8588 13912 8616
rect 13587 8585 13599 8588
rect 13541 8579 13599 8585
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 14458 8576 14464 8628
rect 14516 8616 14522 8628
rect 14734 8616 14740 8628
rect 14516 8588 14740 8616
rect 14516 8576 14522 8588
rect 14734 8576 14740 8588
rect 14792 8576 14798 8628
rect 15194 8616 15200 8628
rect 15155 8588 15200 8616
rect 15194 8576 15200 8588
rect 15252 8576 15258 8628
rect 15289 8619 15347 8625
rect 15289 8585 15301 8619
rect 15335 8616 15347 8619
rect 15562 8616 15568 8628
rect 15335 8588 15568 8616
rect 15335 8585 15347 8588
rect 15289 8579 15347 8585
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 10226 8548 10232 8560
rect 7064 8520 9628 8548
rect 9692 8520 10232 8548
rect 7064 8508 7070 8520
rect 5442 8440 5448 8492
rect 5500 8480 5506 8492
rect 5914 8483 5972 8489
rect 5914 8480 5926 8483
rect 5500 8452 5926 8480
rect 5500 8440 5506 8452
rect 5914 8449 5926 8452
rect 5960 8449 5972 8483
rect 5914 8443 5972 8449
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7834 8480 7840 8492
rect 7156 8452 7840 8480
rect 7156 8440 7162 8452
rect 7834 8440 7840 8452
rect 7892 8440 7898 8492
rect 9692 8489 9720 8520
rect 10226 8508 10232 8520
rect 10284 8508 10290 8560
rect 10410 8508 10416 8560
rect 10468 8548 10474 8560
rect 11149 8551 11207 8557
rect 11149 8548 11161 8551
rect 10468 8520 11161 8548
rect 10468 8508 10474 8520
rect 11149 8517 11161 8520
rect 11195 8548 11207 8551
rect 11698 8548 11704 8560
rect 11195 8520 11704 8548
rect 11195 8517 11207 8520
rect 11149 8511 11207 8517
rect 11698 8508 11704 8520
rect 11756 8508 11762 8560
rect 12158 8508 12164 8560
rect 12216 8508 12222 8560
rect 12986 8548 12992 8560
rect 12360 8520 12992 8548
rect 12360 8492 12388 8520
rect 12986 8508 12992 8520
rect 13044 8508 13050 8560
rect 13354 8508 13360 8560
rect 13412 8548 13418 8560
rect 13633 8551 13691 8557
rect 13633 8548 13645 8551
rect 13412 8520 13645 8548
rect 13412 8508 13418 8520
rect 13633 8517 13645 8520
rect 13679 8517 13691 8551
rect 13633 8511 13691 8517
rect 9677 8483 9735 8489
rect 9677 8449 9689 8483
rect 9723 8449 9735 8483
rect 9933 8483 9991 8489
rect 9933 8480 9945 8483
rect 9677 8443 9735 8449
rect 9784 8452 9945 8480
rect 6178 8412 6184 8424
rect 6139 8384 6184 8412
rect 6178 8372 6184 8384
rect 6236 8412 6242 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 6236 8384 6377 8412
rect 6236 8372 6242 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 7374 8372 7380 8424
rect 7432 8412 7438 8424
rect 9784 8412 9812 8452
rect 9933 8449 9945 8452
rect 9979 8449 9991 8483
rect 9933 8443 9991 8449
rect 11606 8440 11612 8492
rect 11664 8480 11670 8492
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11664 8452 11897 8480
rect 11664 8440 11670 8452
rect 11885 8449 11897 8452
rect 11931 8480 11943 8483
rect 12250 8480 12256 8492
rect 11931 8452 12256 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 12342 8440 12348 8492
rect 12400 8440 12406 8492
rect 12710 8480 12716 8492
rect 12671 8452 12716 8480
rect 12710 8440 12716 8452
rect 12768 8440 12774 8492
rect 12805 8483 12863 8489
rect 12805 8449 12817 8483
rect 12851 8480 12863 8483
rect 13170 8480 13176 8492
rect 12851 8452 13176 8480
rect 12851 8449 12863 8452
rect 12805 8443 12863 8449
rect 13170 8440 13176 8452
rect 13228 8440 13234 8492
rect 14369 8483 14427 8489
rect 14369 8480 14381 8483
rect 13648 8452 14381 8480
rect 13648 8424 13676 8452
rect 14369 8449 14381 8452
rect 14415 8449 14427 8483
rect 14369 8443 14427 8449
rect 14550 8440 14556 8492
rect 14608 8480 14614 8492
rect 14826 8480 14832 8492
rect 14608 8452 14832 8480
rect 14608 8440 14614 8452
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 7432 8384 9812 8412
rect 7432 8372 7438 8384
rect 10686 8372 10692 8424
rect 10744 8412 10750 8424
rect 11790 8412 11796 8424
rect 10744 8384 11796 8412
rect 10744 8372 10750 8384
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 12161 8415 12219 8421
rect 12161 8381 12173 8415
rect 12207 8381 12219 8415
rect 12161 8375 12219 8381
rect 12176 8344 12204 8375
rect 12618 8372 12624 8424
rect 12676 8412 12682 8424
rect 12897 8415 12955 8421
rect 12897 8412 12909 8415
rect 12676 8384 12909 8412
rect 12676 8372 12682 8384
rect 12897 8381 12909 8384
rect 12943 8381 12955 8415
rect 12897 8375 12955 8381
rect 12986 8372 12992 8424
rect 13044 8412 13050 8424
rect 13538 8412 13544 8424
rect 13044 8384 13544 8412
rect 13044 8372 13050 8384
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 13630 8372 13636 8424
rect 13688 8372 13694 8424
rect 13817 8415 13875 8421
rect 13817 8381 13829 8415
rect 13863 8412 13875 8415
rect 13863 8384 13952 8412
rect 13863 8381 13875 8384
rect 13817 8375 13875 8381
rect 13924 8344 13952 8384
rect 13998 8372 14004 8424
rect 14056 8412 14062 8424
rect 14461 8415 14519 8421
rect 14461 8412 14473 8415
rect 14056 8384 14473 8412
rect 14056 8372 14062 8384
rect 14461 8381 14473 8384
rect 14507 8381 14519 8415
rect 14461 8375 14519 8381
rect 14645 8415 14703 8421
rect 14645 8381 14657 8415
rect 14691 8381 14703 8415
rect 14645 8375 14703 8381
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8412 15531 8415
rect 15654 8412 15660 8424
rect 15519 8384 15660 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 7300 8316 9674 8344
rect 3476 8248 4936 8276
rect 3476 8236 3482 8248
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 7300 8276 7328 8316
rect 5500 8248 7328 8276
rect 9646 8276 9674 8316
rect 10888 8316 13952 8344
rect 10888 8276 10916 8316
rect 14550 8304 14556 8356
rect 14608 8344 14614 8356
rect 14660 8344 14688 8375
rect 15654 8372 15660 8384
rect 15712 8372 15718 8424
rect 14608 8316 14688 8344
rect 14608 8304 14614 8316
rect 11054 8276 11060 8288
rect 9646 8248 10916 8276
rect 11015 8248 11060 8276
rect 5500 8236 5506 8248
rect 11054 8236 11060 8248
rect 11112 8236 11118 8288
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 12526 8276 12532 8288
rect 11756 8248 12532 8276
rect 11756 8236 11762 8248
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 12894 8236 12900 8288
rect 12952 8276 12958 8288
rect 14001 8279 14059 8285
rect 14001 8276 14013 8279
rect 12952 8248 14013 8276
rect 12952 8236 12958 8248
rect 14001 8245 14013 8248
rect 14047 8245 14059 8279
rect 14001 8239 14059 8245
rect 14829 8279 14887 8285
rect 14829 8245 14841 8279
rect 14875 8276 14887 8279
rect 16758 8276 16764 8288
rect 14875 8248 16764 8276
rect 14875 8245 14887 8248
rect 14829 8239 14887 8245
rect 16758 8236 16764 8248
rect 16816 8236 16822 8288
rect 1104 8186 16008 8208
rect 1104 8134 2824 8186
rect 2876 8134 2888 8186
rect 2940 8134 2952 8186
rect 3004 8134 3016 8186
rect 3068 8134 3080 8186
rect 3132 8134 6572 8186
rect 6624 8134 6636 8186
rect 6688 8134 6700 8186
rect 6752 8134 6764 8186
rect 6816 8134 6828 8186
rect 6880 8134 10320 8186
rect 10372 8134 10384 8186
rect 10436 8134 10448 8186
rect 10500 8134 10512 8186
rect 10564 8134 10576 8186
rect 10628 8134 14068 8186
rect 14120 8134 14132 8186
rect 14184 8134 14196 8186
rect 14248 8134 14260 8186
rect 14312 8134 14324 8186
rect 14376 8134 16008 8186
rect 1104 8112 16008 8134
rect 1854 8072 1860 8084
rect 1767 8044 1860 8072
rect 1854 8032 1860 8044
rect 1912 8072 1918 8084
rect 2222 8072 2228 8084
rect 1912 8044 2228 8072
rect 1912 8032 1918 8044
rect 2222 8032 2228 8044
rect 2280 8032 2286 8084
rect 4706 8032 4712 8084
rect 4764 8072 4770 8084
rect 4801 8075 4859 8081
rect 4801 8072 4813 8075
rect 4764 8044 4813 8072
rect 4764 8032 4770 8044
rect 4801 8041 4813 8044
rect 4847 8072 4859 8075
rect 5166 8072 5172 8084
rect 4847 8044 5172 8072
rect 4847 8041 4859 8044
rect 4801 8035 4859 8041
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 5776 8044 8953 8072
rect 5776 8032 5782 8044
rect 8941 8041 8953 8044
rect 8987 8072 8999 8075
rect 10686 8072 10692 8084
rect 8987 8044 10692 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 10686 8032 10692 8044
rect 10744 8032 10750 8084
rect 10778 8032 10784 8084
rect 10836 8072 10842 8084
rect 10836 8044 11928 8072
rect 10836 8032 10842 8044
rect 4433 8007 4491 8013
rect 4433 7973 4445 8007
rect 4479 8004 4491 8007
rect 11900 8004 11928 8044
rect 12250 8032 12256 8084
rect 12308 8072 12314 8084
rect 12308 8044 12572 8072
rect 12308 8032 12314 8044
rect 12544 8004 12572 8044
rect 13354 8032 13360 8084
rect 13412 8072 13418 8084
rect 16114 8072 16120 8084
rect 13412 8044 16120 8072
rect 13412 8032 13418 8044
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 13998 8004 14004 8016
rect 4479 7976 8800 8004
rect 11900 7976 12480 8004
rect 12544 7976 14004 8004
rect 4479 7973 4491 7976
rect 4433 7967 4491 7973
rect 2130 7896 2136 7948
rect 2188 7936 2194 7948
rect 5166 7936 5172 7948
rect 2188 7908 5172 7936
rect 2188 7896 2194 7908
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 8481 7939 8539 7945
rect 8481 7936 8493 7939
rect 5684 7908 8493 7936
rect 5684 7896 5690 7908
rect 8481 7905 8493 7908
rect 8527 7905 8539 7939
rect 8481 7899 8539 7905
rect 3602 7868 3608 7880
rect 3563 7840 3608 7868
rect 3602 7828 3608 7840
rect 3660 7828 3666 7880
rect 3694 7828 3700 7880
rect 3752 7868 3758 7880
rect 3973 7871 4031 7877
rect 3973 7868 3985 7871
rect 3752 7840 3985 7868
rect 3752 7828 3758 7840
rect 3973 7837 3985 7840
rect 4019 7837 4031 7871
rect 3973 7831 4031 7837
rect 4062 7828 4068 7880
rect 4120 7868 4126 7880
rect 4249 7871 4307 7877
rect 4249 7868 4261 7871
rect 4120 7840 4261 7868
rect 4120 7828 4126 7840
rect 4249 7837 4261 7840
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 5350 7828 5356 7880
rect 5408 7868 5414 7880
rect 6365 7871 6423 7877
rect 6365 7868 6377 7871
rect 5408 7840 6377 7868
rect 5408 7828 5414 7840
rect 6365 7837 6377 7840
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 6454 7828 6460 7880
rect 6512 7868 6518 7880
rect 6512 7840 7788 7868
rect 6512 7828 6518 7840
rect 3145 7803 3203 7809
rect 3145 7769 3157 7803
rect 3191 7800 3203 7803
rect 6273 7803 6331 7809
rect 3191 7772 5672 7800
rect 3191 7769 3203 7772
rect 3145 7763 3203 7769
rect 5644 7744 5672 7772
rect 6273 7769 6285 7803
rect 6319 7769 6331 7803
rect 7760 7800 7788 7840
rect 7834 7828 7840 7880
rect 7892 7868 7898 7880
rect 8772 7877 8800 7976
rect 12158 7936 12164 7948
rect 11716 7908 12164 7936
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7892 7840 7941 7868
rect 7892 7828 7898 7840
rect 7929 7837 7941 7840
rect 7975 7837 7987 7871
rect 7929 7831 7987 7837
rect 8757 7871 8815 7877
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 9306 7868 9312 7880
rect 8803 7840 9312 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 9306 7828 9312 7840
rect 9364 7828 9370 7880
rect 9766 7828 9772 7880
rect 9824 7868 9830 7880
rect 10226 7868 10232 7880
rect 9824 7840 10232 7868
rect 9824 7828 9830 7840
rect 10226 7828 10232 7840
rect 10284 7868 10290 7880
rect 10321 7871 10379 7877
rect 10321 7868 10333 7871
rect 10284 7840 10333 7868
rect 10284 7828 10290 7840
rect 10321 7837 10333 7840
rect 10367 7868 10379 7871
rect 10413 7871 10471 7877
rect 10413 7868 10425 7871
rect 10367 7840 10425 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 10413 7837 10425 7840
rect 10459 7837 10471 7871
rect 11716 7868 11744 7908
rect 12158 7896 12164 7908
rect 12216 7896 12222 7948
rect 12342 7936 12348 7948
rect 12303 7908 12348 7936
rect 12342 7896 12348 7908
rect 12400 7896 12406 7948
rect 12452 7945 12480 7976
rect 13998 7964 14004 7976
rect 14056 7964 14062 8016
rect 14093 8007 14151 8013
rect 14093 7973 14105 8007
rect 14139 8004 14151 8007
rect 15378 8004 15384 8016
rect 14139 7976 15384 8004
rect 14139 7973 14151 7976
rect 14093 7967 14151 7973
rect 15378 7964 15384 7976
rect 15436 7964 15442 8016
rect 12437 7939 12495 7945
rect 12437 7905 12449 7939
rect 12483 7905 12495 7939
rect 12437 7899 12495 7905
rect 12897 7939 12955 7945
rect 12897 7905 12909 7939
rect 12943 7905 12955 7939
rect 12897 7899 12955 7905
rect 10413 7831 10471 7837
rect 10612 7840 11744 7868
rect 9030 7800 9036 7812
rect 7760 7772 9036 7800
rect 6273 7763 6331 7769
rect 3418 7732 3424 7744
rect 3379 7704 3424 7732
rect 3418 7692 3424 7704
rect 3476 7692 3482 7744
rect 5626 7692 5632 7744
rect 5684 7732 5690 7744
rect 6288 7732 6316 7763
rect 9030 7760 9036 7772
rect 9088 7760 9094 7812
rect 9398 7760 9404 7812
rect 9456 7800 9462 7812
rect 10054 7803 10112 7809
rect 10054 7800 10066 7803
rect 9456 7772 10066 7800
rect 9456 7760 9462 7772
rect 10054 7769 10066 7772
rect 10100 7800 10112 7803
rect 10612 7800 10640 7840
rect 11790 7828 11796 7880
rect 11848 7868 11854 7880
rect 12912 7868 12940 7899
rect 13538 7896 13544 7948
rect 13596 7936 13602 7948
rect 13817 7939 13875 7945
rect 13817 7936 13829 7939
rect 13596 7908 13829 7936
rect 13596 7896 13602 7908
rect 13817 7905 13829 7908
rect 13863 7905 13875 7939
rect 13817 7899 13875 7905
rect 14737 7939 14795 7945
rect 14737 7905 14749 7939
rect 14783 7936 14795 7939
rect 15102 7936 15108 7948
rect 14783 7908 15108 7936
rect 14783 7905 14795 7908
rect 14737 7899 14795 7905
rect 15102 7896 15108 7908
rect 15160 7896 15166 7948
rect 15470 7936 15476 7948
rect 15431 7908 15476 7936
rect 15470 7896 15476 7908
rect 15528 7896 15534 7948
rect 13998 7868 14004 7880
rect 11848 7840 14004 7868
rect 11848 7828 11854 7840
rect 13998 7828 14004 7840
rect 14056 7868 14062 7880
rect 15654 7868 15660 7880
rect 14056 7840 15660 7868
rect 14056 7828 14062 7840
rect 15654 7828 15660 7840
rect 15712 7828 15718 7880
rect 10686 7809 10692 7812
rect 10100 7772 10640 7800
rect 10100 7769 10112 7772
rect 10054 7763 10112 7769
rect 10680 7763 10692 7809
rect 10744 7800 10750 7812
rect 12253 7803 12311 7809
rect 12253 7800 12265 7803
rect 10744 7772 10780 7800
rect 11072 7772 12265 7800
rect 10686 7760 10692 7763
rect 10744 7760 10750 7772
rect 7834 7732 7840 7744
rect 5684 7704 7840 7732
rect 5684 7692 5690 7704
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 7926 7692 7932 7744
rect 7984 7732 7990 7744
rect 11072 7732 11100 7772
rect 12253 7769 12265 7772
rect 12299 7769 12311 7803
rect 12253 7763 12311 7769
rect 12618 7760 12624 7812
rect 12676 7800 12682 7812
rect 13722 7800 13728 7812
rect 12676 7772 13728 7800
rect 12676 7760 12682 7772
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 13814 7760 13820 7812
rect 13872 7800 13878 7812
rect 14090 7800 14096 7812
rect 13872 7772 14096 7800
rect 13872 7760 13878 7772
rect 14090 7760 14096 7772
rect 14148 7760 14154 7812
rect 14553 7803 14611 7809
rect 14553 7769 14565 7803
rect 14599 7800 14611 7803
rect 14642 7800 14648 7812
rect 14599 7772 14648 7800
rect 14599 7769 14611 7772
rect 14553 7763 14611 7769
rect 14642 7760 14648 7772
rect 14700 7800 14706 7812
rect 15102 7800 15108 7812
rect 14700 7772 15108 7800
rect 14700 7760 14706 7772
rect 15102 7760 15108 7772
rect 15160 7760 15166 7812
rect 15194 7760 15200 7812
rect 15252 7800 15258 7812
rect 15381 7803 15439 7809
rect 15381 7800 15393 7803
rect 15252 7772 15393 7800
rect 15252 7760 15258 7772
rect 15381 7769 15393 7772
rect 15427 7800 15439 7803
rect 16114 7800 16120 7812
rect 15427 7772 16120 7800
rect 15427 7769 15439 7772
rect 15381 7763 15439 7769
rect 16114 7760 16120 7772
rect 16172 7760 16178 7812
rect 7984 7704 11100 7732
rect 7984 7692 7990 7704
rect 11238 7692 11244 7744
rect 11296 7732 11302 7744
rect 11790 7732 11796 7744
rect 11296 7704 11796 7732
rect 11296 7692 11302 7704
rect 11790 7692 11796 7704
rect 11848 7692 11854 7744
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 12986 7732 12992 7744
rect 11940 7704 11985 7732
rect 12947 7704 12992 7732
rect 11940 7692 11946 7704
rect 12986 7692 12992 7704
rect 13044 7692 13050 7744
rect 13081 7735 13139 7741
rect 13081 7701 13093 7735
rect 13127 7732 13139 7735
rect 13262 7732 13268 7744
rect 13127 7704 13268 7732
rect 13127 7701 13139 7704
rect 13081 7695 13139 7701
rect 13262 7692 13268 7704
rect 13320 7692 13326 7744
rect 13446 7732 13452 7744
rect 13407 7704 13452 7732
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13541 7735 13599 7741
rect 13541 7701 13553 7735
rect 13587 7732 13599 7735
rect 13906 7732 13912 7744
rect 13587 7704 13912 7732
rect 13587 7701 13599 7704
rect 13541 7695 13599 7701
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 14458 7732 14464 7744
rect 14419 7704 14464 7732
rect 14458 7692 14464 7704
rect 14516 7692 14522 7744
rect 14734 7692 14740 7744
rect 14792 7732 14798 7744
rect 14921 7735 14979 7741
rect 14921 7732 14933 7735
rect 14792 7704 14933 7732
rect 14792 7692 14798 7704
rect 14921 7701 14933 7704
rect 14967 7701 14979 7735
rect 15286 7732 15292 7744
rect 15199 7704 15292 7732
rect 14921 7695 14979 7701
rect 15286 7692 15292 7704
rect 15344 7732 15350 7744
rect 15654 7732 15660 7744
rect 15344 7704 15660 7732
rect 15344 7692 15350 7704
rect 15654 7692 15660 7704
rect 15712 7692 15718 7744
rect 1104 7642 16008 7664
rect 1104 7590 4698 7642
rect 4750 7590 4762 7642
rect 4814 7590 4826 7642
rect 4878 7590 4890 7642
rect 4942 7590 4954 7642
rect 5006 7590 8446 7642
rect 8498 7590 8510 7642
rect 8562 7590 8574 7642
rect 8626 7590 8638 7642
rect 8690 7590 8702 7642
rect 8754 7590 12194 7642
rect 12246 7590 12258 7642
rect 12310 7590 12322 7642
rect 12374 7590 12386 7642
rect 12438 7590 12450 7642
rect 12502 7590 16008 7642
rect 1104 7568 16008 7590
rect 2130 7488 2136 7540
rect 2188 7528 2194 7540
rect 3329 7531 3387 7537
rect 3329 7528 3341 7531
rect 2188 7500 3341 7528
rect 2188 7488 2194 7500
rect 3329 7497 3341 7500
rect 3375 7497 3387 7531
rect 3329 7491 3387 7497
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 4801 7531 4859 7537
rect 4801 7528 4813 7531
rect 4580 7500 4813 7528
rect 4580 7488 4586 7500
rect 4801 7497 4813 7500
rect 4847 7497 4859 7531
rect 4801 7491 4859 7497
rect 5074 7488 5080 7540
rect 5132 7528 5138 7540
rect 8018 7528 8024 7540
rect 5132 7500 8024 7528
rect 5132 7488 5138 7500
rect 4154 7420 4160 7472
rect 4212 7460 4218 7472
rect 4212 7432 4752 7460
rect 4212 7420 4218 7432
rect 1486 7392 1492 7404
rect 1447 7364 1492 7392
rect 1486 7352 1492 7364
rect 1544 7352 1550 7404
rect 1854 7392 1860 7404
rect 1815 7364 1860 7392
rect 1854 7352 1860 7364
rect 1912 7352 1918 7404
rect 2124 7395 2182 7401
rect 2124 7361 2136 7395
rect 2170 7392 2182 7395
rect 2498 7392 2504 7404
rect 2170 7364 2504 7392
rect 2170 7361 2182 7364
rect 2124 7355 2182 7361
rect 2498 7352 2504 7364
rect 2556 7352 2562 7404
rect 4453 7395 4511 7401
rect 4453 7361 4465 7395
rect 4499 7392 4511 7395
rect 4614 7392 4620 7404
rect 4499 7364 4620 7392
rect 4499 7361 4511 7364
rect 4453 7355 4511 7361
rect 4614 7352 4620 7364
rect 4672 7352 4678 7404
rect 4724 7401 4752 7432
rect 5166 7420 5172 7472
rect 5224 7460 5230 7472
rect 5951 7469 5979 7500
rect 8018 7488 8024 7500
rect 8076 7528 8082 7540
rect 8076 7500 9444 7528
rect 8076 7488 8082 7500
rect 5936 7463 5994 7469
rect 5224 7432 5865 7460
rect 5224 7420 5230 7432
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 5442 7392 5448 7404
rect 4709 7355 4767 7361
rect 4816 7364 5448 7392
rect 4632 7324 4660 7352
rect 4816 7324 4844 7364
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 5837 7392 5865 7432
rect 5936 7429 5948 7463
rect 5982 7429 5994 7463
rect 9416 7460 9444 7500
rect 10042 7488 10048 7540
rect 10100 7528 10106 7540
rect 10962 7528 10968 7540
rect 10100 7500 10968 7528
rect 10100 7488 10106 7500
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11146 7528 11152 7540
rect 11107 7500 11152 7528
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 12345 7531 12403 7537
rect 12345 7528 12357 7531
rect 11808 7500 12357 7528
rect 11238 7460 11244 7472
rect 5936 7423 5994 7429
rect 6840 7432 8064 7460
rect 9416 7432 11244 7460
rect 6840 7392 6868 7432
rect 8036 7404 8064 7432
rect 11238 7420 11244 7432
rect 11296 7420 11302 7472
rect 5837 7364 6868 7392
rect 6914 7352 6920 7404
rect 6972 7392 6978 7404
rect 7478 7395 7536 7401
rect 7478 7392 7490 7395
rect 6972 7364 7490 7392
rect 6972 7352 6978 7364
rect 7478 7361 7490 7364
rect 7524 7361 7536 7395
rect 7478 7355 7536 7361
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 7892 7364 7937 7392
rect 7892 7352 7898 7364
rect 8018 7352 8024 7404
rect 8076 7352 8082 7404
rect 9030 7352 9036 7404
rect 9088 7392 9094 7404
rect 9490 7392 9496 7404
rect 9088 7364 9496 7392
rect 9088 7352 9094 7364
rect 9490 7352 9496 7364
rect 9548 7352 9554 7404
rect 9585 7395 9643 7401
rect 9585 7361 9597 7395
rect 9631 7392 9643 7395
rect 9677 7395 9735 7401
rect 9677 7392 9689 7395
rect 9631 7364 9689 7392
rect 9631 7361 9643 7364
rect 9585 7355 9643 7361
rect 9677 7361 9689 7364
rect 9723 7392 9735 7395
rect 9766 7392 9772 7404
rect 9723 7364 9772 7392
rect 9723 7361 9735 7364
rect 9677 7355 9735 7361
rect 6178 7324 6184 7336
rect 4632 7296 4844 7324
rect 6139 7296 6184 7324
rect 6178 7284 6184 7296
rect 6236 7284 6242 7336
rect 7745 7327 7803 7333
rect 7745 7293 7757 7327
rect 7791 7324 7803 7327
rect 9306 7324 9312 7336
rect 7791 7296 9312 7324
rect 7791 7293 7803 7296
rect 7745 7287 7803 7293
rect 9306 7284 9312 7296
rect 9364 7324 9370 7336
rect 9600 7324 9628 7355
rect 9766 7352 9772 7364
rect 9824 7352 9830 7404
rect 9950 7401 9956 7404
rect 9944 7355 9956 7401
rect 10008 7392 10014 7404
rect 10008 7364 10044 7392
rect 9950 7352 9956 7355
rect 10008 7352 10014 7364
rect 11146 7352 11152 7404
rect 11204 7392 11210 7404
rect 11808 7392 11836 7500
rect 12345 7497 12357 7500
rect 12391 7497 12403 7531
rect 12345 7491 12403 7497
rect 13262 7488 13268 7540
rect 13320 7528 13326 7540
rect 13541 7531 13599 7537
rect 13541 7528 13553 7531
rect 13320 7500 13553 7528
rect 13320 7488 13326 7500
rect 13541 7497 13553 7500
rect 13587 7528 13599 7531
rect 13722 7528 13728 7540
rect 13587 7500 13728 7528
rect 13587 7497 13599 7500
rect 13541 7491 13599 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 14369 7531 14427 7537
rect 14369 7497 14381 7531
rect 14415 7528 14427 7531
rect 14918 7528 14924 7540
rect 14415 7500 14924 7528
rect 14415 7497 14427 7500
rect 14369 7491 14427 7497
rect 14918 7488 14924 7500
rect 14976 7488 14982 7540
rect 15028 7500 15424 7528
rect 11885 7463 11943 7469
rect 11885 7429 11897 7463
rect 11931 7460 11943 7463
rect 12250 7460 12256 7472
rect 11931 7432 12256 7460
rect 11931 7429 11943 7432
rect 11885 7423 11943 7429
rect 12250 7420 12256 7432
rect 12308 7420 12314 7472
rect 12805 7463 12863 7469
rect 12805 7429 12817 7463
rect 12851 7429 12863 7463
rect 12805 7423 12863 7429
rect 11974 7392 11980 7404
rect 11204 7364 11836 7392
rect 11935 7364 11980 7392
rect 11204 7352 11210 7364
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 12434 7352 12440 7404
rect 12492 7392 12498 7404
rect 12710 7392 12716 7404
rect 12492 7364 12716 7392
rect 12492 7352 12498 7364
rect 12710 7352 12716 7364
rect 12768 7352 12774 7404
rect 12820 7392 12848 7423
rect 12986 7420 12992 7472
rect 13044 7460 13050 7472
rect 15028 7460 15056 7500
rect 15194 7460 15200 7472
rect 13044 7432 15056 7460
rect 15155 7432 15200 7460
rect 13044 7420 13050 7432
rect 15194 7420 15200 7432
rect 15252 7420 15258 7472
rect 13449 7395 13507 7401
rect 12820 7364 13400 7392
rect 9364 7296 9628 7324
rect 9364 7284 9370 7296
rect 10686 7284 10692 7336
rect 10744 7324 10750 7336
rect 10962 7324 10968 7336
rect 10744 7296 10968 7324
rect 10744 7284 10750 7296
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11238 7284 11244 7336
rect 11296 7324 11302 7336
rect 12161 7327 12219 7333
rect 12161 7324 12173 7327
rect 11296 7296 11652 7324
rect 11296 7284 11302 7296
rect 3050 7216 3056 7268
rect 3108 7256 3114 7268
rect 3237 7259 3295 7265
rect 3237 7256 3249 7259
rect 3108 7228 3249 7256
rect 3108 7216 3114 7228
rect 3237 7225 3249 7228
rect 3283 7225 3295 7259
rect 8202 7256 8208 7268
rect 3237 7219 3295 7225
rect 7760 7228 8208 7256
rect 1673 7191 1731 7197
rect 1673 7157 1685 7191
rect 1719 7188 1731 7191
rect 2222 7188 2228 7200
rect 1719 7160 2228 7188
rect 1719 7157 1731 7160
rect 1673 7151 1731 7157
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 3326 7148 3332 7200
rect 3384 7188 3390 7200
rect 6365 7191 6423 7197
rect 6365 7188 6377 7191
rect 3384 7160 6377 7188
rect 3384 7148 3390 7160
rect 6365 7157 6377 7160
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 6454 7148 6460 7200
rect 6512 7188 6518 7200
rect 7760 7188 7788 7228
rect 8202 7216 8208 7228
rect 8260 7256 8266 7268
rect 9398 7256 9404 7268
rect 8260 7228 9404 7256
rect 8260 7216 8266 7228
rect 9398 7216 9404 7228
rect 9456 7216 9462 7268
rect 11514 7256 11520 7268
rect 11475 7228 11520 7256
rect 11514 7216 11520 7228
rect 11572 7216 11578 7268
rect 11624 7256 11652 7296
rect 11992 7296 12173 7324
rect 11992 7256 12020 7296
rect 12161 7293 12173 7296
rect 12207 7293 12219 7327
rect 12897 7327 12955 7333
rect 12897 7324 12909 7327
rect 12161 7287 12219 7293
rect 12268 7296 12909 7324
rect 12268 7256 12296 7296
rect 12897 7293 12909 7296
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 13265 7327 13323 7333
rect 13265 7293 13277 7327
rect 13311 7293 13323 7327
rect 13372 7324 13400 7364
rect 13449 7361 13461 7395
rect 13495 7392 13507 7395
rect 13538 7392 13544 7404
rect 13495 7364 13544 7392
rect 13495 7361 13507 7364
rect 13449 7355 13507 7361
rect 13538 7352 13544 7364
rect 13596 7392 13602 7404
rect 14366 7392 14372 7404
rect 13596 7364 14372 7392
rect 13596 7352 13602 7364
rect 14366 7352 14372 7364
rect 14424 7352 14430 7404
rect 14461 7395 14519 7401
rect 14461 7361 14473 7395
rect 14507 7392 14519 7395
rect 14550 7392 14556 7404
rect 14507 7364 14556 7392
rect 14507 7361 14519 7364
rect 14461 7355 14519 7361
rect 14550 7352 14556 7364
rect 14608 7392 14614 7404
rect 15010 7392 15016 7404
rect 14608 7364 15016 7392
rect 14608 7352 14614 7364
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 13722 7324 13728 7336
rect 13372 7296 13728 7324
rect 13265 7287 13323 7293
rect 11624 7228 12020 7256
rect 12176 7228 12296 7256
rect 6512 7160 7788 7188
rect 6512 7148 6518 7160
rect 7834 7148 7840 7200
rect 7892 7188 7898 7200
rect 10686 7188 10692 7200
rect 7892 7160 10692 7188
rect 7892 7148 7898 7160
rect 10686 7148 10692 7160
rect 10744 7148 10750 7200
rect 11054 7188 11060 7200
rect 11015 7160 11060 7188
rect 11054 7148 11060 7160
rect 11112 7148 11118 7200
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 12176 7188 12204 7228
rect 12342 7216 12348 7268
rect 12400 7256 12406 7268
rect 12618 7256 12624 7268
rect 12400 7228 12624 7256
rect 12400 7216 12406 7228
rect 12618 7216 12624 7228
rect 12676 7216 12682 7268
rect 12710 7216 12716 7268
rect 12768 7256 12774 7268
rect 13280 7256 13308 7287
rect 13722 7284 13728 7296
rect 13780 7284 13786 7336
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 13832 7296 14657 7324
rect 12768 7228 13308 7256
rect 12768 7216 12774 7228
rect 11204 7160 12204 7188
rect 11204 7148 11210 7160
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 12802 7188 12808 7200
rect 12584 7160 12808 7188
rect 12584 7148 12590 7160
rect 12802 7148 12808 7160
rect 12860 7188 12866 7200
rect 13832 7188 13860 7296
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 15286 7324 15292 7336
rect 15247 7296 15292 7324
rect 14645 7287 14703 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 15396 7333 15424 7500
rect 15381 7327 15439 7333
rect 15381 7293 15393 7327
rect 15427 7293 15439 7327
rect 15381 7287 15439 7293
rect 13998 7256 14004 7268
rect 13959 7228 14004 7256
rect 13998 7216 14004 7228
rect 14056 7216 14062 7268
rect 15194 7256 15200 7268
rect 14660 7228 15200 7256
rect 12860 7160 13860 7188
rect 13909 7191 13967 7197
rect 12860 7148 12866 7160
rect 13909 7157 13921 7191
rect 13955 7188 13967 7191
rect 14660 7188 14688 7228
rect 15194 7216 15200 7228
rect 15252 7216 15258 7268
rect 13955 7160 14688 7188
rect 14829 7191 14887 7197
rect 13955 7157 13967 7160
rect 13909 7151 13967 7157
rect 14829 7157 14841 7191
rect 14875 7188 14887 7191
rect 15010 7188 15016 7200
rect 14875 7160 15016 7188
rect 14875 7157 14887 7160
rect 14829 7151 14887 7157
rect 15010 7148 15016 7160
rect 15068 7148 15074 7200
rect 1104 7098 16008 7120
rect 1104 7046 2824 7098
rect 2876 7046 2888 7098
rect 2940 7046 2952 7098
rect 3004 7046 3016 7098
rect 3068 7046 3080 7098
rect 3132 7046 6572 7098
rect 6624 7046 6636 7098
rect 6688 7046 6700 7098
rect 6752 7046 6764 7098
rect 6816 7046 6828 7098
rect 6880 7046 10320 7098
rect 10372 7046 10384 7098
rect 10436 7046 10448 7098
rect 10500 7046 10512 7098
rect 10564 7046 10576 7098
rect 10628 7046 14068 7098
rect 14120 7046 14132 7098
rect 14184 7046 14196 7098
rect 14248 7046 14260 7098
rect 14312 7046 14324 7098
rect 14376 7046 16008 7098
rect 1104 7024 16008 7046
rect 3878 6944 3884 6996
rect 3936 6984 3942 6996
rect 7098 6984 7104 6996
rect 3936 6956 7104 6984
rect 3936 6944 3942 6956
rect 7098 6944 7104 6956
rect 7156 6944 7162 6996
rect 7650 6944 7656 6996
rect 7708 6984 7714 6996
rect 9674 6984 9680 6996
rect 7708 6956 9680 6984
rect 7708 6944 7714 6956
rect 9674 6944 9680 6956
rect 9732 6944 9738 6996
rect 9950 6944 9956 6996
rect 10008 6984 10014 6996
rect 10778 6984 10784 6996
rect 10008 6956 10784 6984
rect 10008 6944 10014 6956
rect 10778 6944 10784 6956
rect 10836 6944 10842 6996
rect 11146 6944 11152 6996
rect 11204 6984 11210 6996
rect 11882 6984 11888 6996
rect 11204 6956 11888 6984
rect 11204 6944 11210 6956
rect 11882 6944 11888 6956
rect 11940 6944 11946 6996
rect 12069 6987 12127 6993
rect 12069 6984 12081 6987
rect 11992 6956 12081 6984
rect 5905 6919 5963 6925
rect 5905 6885 5917 6919
rect 5951 6916 5963 6919
rect 6270 6916 6276 6928
rect 5951 6888 6276 6916
rect 5951 6885 5963 6888
rect 5905 6879 5963 6885
rect 6270 6876 6276 6888
rect 6328 6876 6334 6928
rect 10962 6876 10968 6928
rect 11020 6916 11026 6928
rect 11241 6919 11299 6925
rect 11241 6916 11253 6919
rect 11020 6888 11253 6916
rect 11020 6876 11026 6888
rect 11241 6885 11253 6888
rect 11287 6885 11299 6919
rect 11241 6879 11299 6885
rect 11330 6876 11336 6928
rect 11388 6916 11394 6928
rect 11992 6916 12020 6956
rect 12069 6953 12081 6956
rect 12115 6953 12127 6987
rect 12069 6947 12127 6953
rect 12158 6944 12164 6996
rect 12216 6984 12222 6996
rect 12216 6956 13492 6984
rect 12216 6944 12222 6956
rect 11388 6888 12020 6916
rect 11388 6876 11394 6888
rect 12250 6876 12256 6928
rect 12308 6916 12314 6928
rect 13262 6916 13268 6928
rect 12308 6888 13268 6916
rect 12308 6876 12314 6888
rect 13262 6876 13268 6888
rect 13320 6876 13326 6928
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6848 1639 6851
rect 2590 6848 2596 6860
rect 1627 6820 2596 6848
rect 1627 6817 1639 6820
rect 1581 6811 1639 6817
rect 2590 6808 2596 6820
rect 2648 6808 2654 6860
rect 3970 6848 3976 6860
rect 3931 6820 3976 6848
rect 3970 6808 3976 6820
rect 4028 6808 4034 6860
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6848 5871 6851
rect 6178 6848 6184 6860
rect 5859 6820 6184 6848
rect 5859 6817 5871 6820
rect 5813 6811 5871 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 8757 6851 8815 6857
rect 8757 6817 8769 6851
rect 8803 6848 8815 6851
rect 9306 6848 9312 6860
rect 8803 6820 9312 6848
rect 8803 6817 8815 6820
rect 8757 6811 8815 6817
rect 9306 6808 9312 6820
rect 9364 6808 9370 6860
rect 10597 6851 10655 6857
rect 10244 6820 10548 6848
rect 10244 6792 10272 6820
rect 842 6740 848 6792
rect 900 6780 906 6792
rect 1486 6780 1492 6792
rect 900 6752 1492 6780
rect 900 6740 906 6752
rect 1486 6740 1492 6752
rect 1544 6780 1550 6792
rect 1765 6783 1823 6789
rect 1765 6780 1777 6783
rect 1544 6752 1777 6780
rect 1544 6740 1550 6752
rect 1765 6749 1777 6752
rect 1811 6749 1823 6783
rect 3510 6780 3516 6792
rect 1765 6743 1823 6749
rect 2746 6752 3516 6780
rect 2746 6712 2774 6752
rect 3510 6740 3516 6752
rect 3568 6740 3574 6792
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6780 3663 6783
rect 4154 6780 4160 6792
rect 3651 6752 4160 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 5166 6780 5172 6792
rect 4295 6752 5172 6780
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 7285 6783 7343 6789
rect 5460 6752 7236 6780
rect 2148 6684 2774 6712
rect 3360 6715 3418 6721
rect 1670 6644 1676 6656
rect 1631 6616 1676 6644
rect 1670 6604 1676 6616
rect 1728 6604 1734 6656
rect 2148 6653 2176 6684
rect 3360 6681 3372 6715
rect 3406 6712 3418 6715
rect 5460 6712 5488 6752
rect 3406 6684 5488 6712
rect 5546 6715 5604 6721
rect 3406 6681 3418 6684
rect 3360 6675 3418 6681
rect 5546 6681 5558 6715
rect 5592 6681 5604 6715
rect 5546 6675 5604 6681
rect 2133 6647 2191 6653
rect 2133 6613 2145 6647
rect 2179 6613 2191 6647
rect 2133 6607 2191 6613
rect 2225 6647 2283 6653
rect 2225 6613 2237 6647
rect 2271 6644 2283 6647
rect 2406 6644 2412 6656
rect 2271 6616 2412 6644
rect 2271 6613 2283 6616
rect 2225 6607 2283 6613
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 4430 6644 4436 6656
rect 4391 6616 4436 6644
rect 4430 6604 4436 6616
rect 4488 6604 4494 6656
rect 5258 6604 5264 6656
rect 5316 6644 5322 6656
rect 5442 6644 5448 6656
rect 5316 6616 5448 6644
rect 5316 6604 5322 6616
rect 5442 6604 5448 6616
rect 5500 6644 5506 6656
rect 5552 6644 5580 6675
rect 7006 6672 7012 6724
rect 7064 6721 7070 6724
rect 7064 6712 7076 6721
rect 7064 6684 7109 6712
rect 7064 6675 7076 6684
rect 7064 6672 7070 6675
rect 5500 6616 5580 6644
rect 7208 6644 7236 6752
rect 7285 6749 7297 6783
rect 7331 6780 7343 6783
rect 7742 6780 7748 6792
rect 7331 6752 7748 6780
rect 7331 6749 7343 6752
rect 7285 6743 7343 6749
rect 7742 6740 7748 6752
rect 7800 6740 7806 6792
rect 8110 6740 8116 6792
rect 8168 6780 8174 6792
rect 8168 6752 9987 6780
rect 8168 6740 8174 6752
rect 8512 6715 8570 6721
rect 8512 6681 8524 6715
rect 8558 6712 8570 6715
rect 9858 6712 9864 6724
rect 8558 6684 9864 6712
rect 8558 6681 8570 6684
rect 8512 6675 8570 6681
rect 9858 6672 9864 6684
rect 9916 6672 9922 6724
rect 7377 6647 7435 6653
rect 7377 6644 7389 6647
rect 7208 6616 7389 6644
rect 5500 6604 5506 6616
rect 7377 6613 7389 6616
rect 7423 6644 7435 6647
rect 7834 6644 7840 6656
rect 7423 6616 7840 6644
rect 7423 6613 7435 6616
rect 7377 6607 7435 6613
rect 7834 6604 7840 6616
rect 7892 6604 7898 6656
rect 7926 6604 7932 6656
rect 7984 6644 7990 6656
rect 8941 6647 8999 6653
rect 8941 6644 8953 6647
rect 7984 6616 8953 6644
rect 7984 6604 7990 6616
rect 8941 6613 8953 6616
rect 8987 6613 8999 6647
rect 8941 6607 8999 6613
rect 9122 6604 9128 6656
rect 9180 6644 9186 6656
rect 9398 6644 9404 6656
rect 9180 6616 9404 6644
rect 9180 6604 9186 6616
rect 9398 6604 9404 6616
rect 9456 6604 9462 6656
rect 9490 6604 9496 6656
rect 9548 6644 9554 6656
rect 9766 6644 9772 6656
rect 9548 6616 9772 6644
rect 9548 6604 9554 6616
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 9959 6644 9987 6752
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10318 6740 10324 6792
rect 10376 6780 10382 6792
rect 10520 6780 10548 6820
rect 10597 6817 10609 6851
rect 10643 6848 10655 6851
rect 10686 6848 10692 6860
rect 10643 6820 10692 6848
rect 10643 6817 10655 6820
rect 10597 6811 10655 6817
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 11514 6808 11520 6860
rect 11572 6848 11578 6860
rect 11790 6848 11796 6860
rect 11572 6820 11796 6848
rect 11572 6808 11578 6820
rect 11790 6808 11796 6820
rect 11848 6808 11854 6860
rect 11882 6808 11888 6860
rect 11940 6848 11946 6860
rect 12621 6851 12679 6857
rect 12621 6848 12633 6851
rect 11940 6820 12633 6848
rect 11940 6808 11946 6820
rect 12621 6817 12633 6820
rect 12667 6817 12679 6851
rect 12621 6811 12679 6817
rect 12710 6808 12716 6860
rect 12768 6848 12774 6860
rect 12894 6848 12900 6860
rect 12768 6820 12900 6848
rect 12768 6808 12774 6820
rect 12894 6808 12900 6820
rect 12952 6808 12958 6860
rect 13354 6848 13360 6860
rect 13315 6820 13360 6848
rect 13354 6808 13360 6820
rect 13412 6808 13418 6860
rect 13464 6857 13492 6956
rect 13630 6944 13636 6996
rect 13688 6944 13694 6996
rect 13722 6944 13728 6996
rect 13780 6984 13786 6996
rect 13780 6956 14320 6984
rect 13780 6944 13786 6956
rect 13449 6851 13507 6857
rect 13449 6817 13461 6851
rect 13495 6817 13507 6851
rect 13648 6848 13676 6944
rect 14292 6928 14320 6956
rect 15562 6944 15568 6996
rect 15620 6944 15626 6996
rect 14274 6876 14280 6928
rect 14332 6876 14338 6928
rect 13909 6851 13967 6857
rect 13909 6848 13921 6851
rect 13648 6820 13921 6848
rect 13449 6811 13507 6817
rect 13909 6817 13921 6820
rect 13955 6817 13967 6851
rect 14642 6848 14648 6860
rect 14603 6820 14648 6848
rect 13909 6811 13967 6817
rect 14642 6808 14648 6820
rect 14700 6808 14706 6860
rect 15194 6808 15200 6860
rect 15252 6848 15258 6860
rect 15580 6857 15608 6944
rect 15381 6851 15439 6857
rect 15381 6848 15393 6851
rect 15252 6820 15393 6848
rect 15252 6808 15258 6820
rect 15381 6817 15393 6820
rect 15427 6817 15439 6851
rect 15381 6811 15439 6817
rect 15565 6851 15623 6857
rect 15565 6817 15577 6851
rect 15611 6817 15623 6851
rect 15565 6811 15623 6817
rect 10376 6752 10421 6780
rect 10520 6752 11100 6780
rect 10376 6740 10382 6752
rect 10076 6715 10134 6721
rect 10076 6681 10088 6715
rect 10122 6712 10134 6715
rect 10410 6712 10416 6724
rect 10122 6684 10416 6712
rect 10122 6681 10134 6684
rect 10076 6675 10134 6681
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 10781 6715 10839 6721
rect 10781 6681 10793 6715
rect 10827 6712 10839 6715
rect 10962 6712 10968 6724
rect 10827 6684 10968 6712
rect 10827 6681 10839 6684
rect 10781 6675 10839 6681
rect 10962 6672 10968 6684
rect 11020 6672 11026 6724
rect 11072 6712 11100 6752
rect 11606 6740 11612 6792
rect 11664 6780 11670 6792
rect 11664 6752 11709 6780
rect 11664 6740 11670 6752
rect 12434 6740 12440 6792
rect 12492 6780 12498 6792
rect 13265 6783 13323 6789
rect 12492 6752 12537 6780
rect 12492 6740 12498 6752
rect 13265 6749 13277 6783
rect 13311 6749 13323 6783
rect 13265 6743 13323 6749
rect 12529 6715 12587 6721
rect 11072 6684 11928 6712
rect 10594 6644 10600 6656
rect 9959 6616 10600 6644
rect 10594 6604 10600 6616
rect 10652 6644 10658 6656
rect 10689 6647 10747 6653
rect 10689 6644 10701 6647
rect 10652 6616 10701 6644
rect 10652 6604 10658 6616
rect 10689 6613 10701 6616
rect 10735 6613 10747 6647
rect 10689 6607 10747 6613
rect 10870 6604 10876 6656
rect 10928 6644 10934 6656
rect 11149 6647 11207 6653
rect 11149 6644 11161 6647
rect 10928 6616 11161 6644
rect 10928 6604 10934 6616
rect 11149 6613 11161 6616
rect 11195 6613 11207 6647
rect 11149 6607 11207 6613
rect 11701 6647 11759 6653
rect 11701 6613 11713 6647
rect 11747 6644 11759 6647
rect 11790 6644 11796 6656
rect 11747 6616 11796 6644
rect 11747 6613 11759 6616
rect 11701 6607 11759 6613
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 11900 6644 11928 6684
rect 12529 6681 12541 6715
rect 12575 6712 12587 6715
rect 13078 6712 13084 6724
rect 12575 6684 13084 6712
rect 12575 6681 12587 6684
rect 12529 6675 12587 6681
rect 13078 6672 13084 6684
rect 13136 6672 13142 6724
rect 13280 6712 13308 6743
rect 13722 6740 13728 6792
rect 13780 6780 13786 6792
rect 14550 6780 14556 6792
rect 13780 6752 14556 6780
rect 13780 6740 13786 6752
rect 14550 6740 14556 6752
rect 14608 6740 14614 6792
rect 14826 6712 14832 6724
rect 13280 6684 14832 6712
rect 14826 6672 14832 6684
rect 14884 6672 14890 6724
rect 12897 6647 12955 6653
rect 12897 6644 12909 6647
rect 11900 6616 12909 6644
rect 12897 6613 12909 6616
rect 12943 6613 12955 6647
rect 12897 6607 12955 6613
rect 13538 6604 13544 6656
rect 13596 6644 13602 6656
rect 13906 6644 13912 6656
rect 13596 6616 13912 6644
rect 13596 6604 13602 6616
rect 13906 6604 13912 6616
rect 13964 6604 13970 6656
rect 14090 6644 14096 6656
rect 14051 6616 14096 6644
rect 14090 6604 14096 6616
rect 14148 6604 14154 6656
rect 14182 6604 14188 6656
rect 14240 6644 14246 6656
rect 14461 6647 14519 6653
rect 14461 6644 14473 6647
rect 14240 6616 14473 6644
rect 14240 6604 14246 6616
rect 14461 6613 14473 6616
rect 14507 6613 14519 6647
rect 14461 6607 14519 6613
rect 14550 6604 14556 6656
rect 14608 6644 14614 6656
rect 14918 6644 14924 6656
rect 14608 6616 14653 6644
rect 14879 6616 14924 6644
rect 14608 6604 14614 6616
rect 14918 6604 14924 6616
rect 14976 6604 14982 6656
rect 15102 6604 15108 6656
rect 15160 6644 15166 6656
rect 15289 6647 15347 6653
rect 15289 6644 15301 6647
rect 15160 6616 15301 6644
rect 15160 6604 15166 6616
rect 15289 6613 15301 6616
rect 15335 6613 15347 6647
rect 15289 6607 15347 6613
rect 1104 6554 16008 6576
rect 1104 6502 4698 6554
rect 4750 6502 4762 6554
rect 4814 6502 4826 6554
rect 4878 6502 4890 6554
rect 4942 6502 4954 6554
rect 5006 6502 8446 6554
rect 8498 6502 8510 6554
rect 8562 6502 8574 6554
rect 8626 6502 8638 6554
rect 8690 6502 8702 6554
rect 8754 6502 12194 6554
rect 12246 6502 12258 6554
rect 12310 6502 12322 6554
rect 12374 6502 12386 6554
rect 12438 6502 12450 6554
rect 12502 6502 16008 6554
rect 1104 6480 16008 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 3602 6440 3608 6452
rect 1627 6412 3608 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 3602 6400 3608 6412
rect 3660 6400 3666 6452
rect 4614 6400 4620 6452
rect 4672 6440 4678 6452
rect 4709 6443 4767 6449
rect 4709 6440 4721 6443
rect 4672 6412 4721 6440
rect 4672 6400 4678 6412
rect 4709 6409 4721 6412
rect 4755 6409 4767 6443
rect 4709 6403 4767 6409
rect 6086 6400 6092 6452
rect 6144 6440 6150 6452
rect 7745 6443 7803 6449
rect 7745 6440 7757 6443
rect 6144 6412 7757 6440
rect 6144 6400 6150 6412
rect 7745 6409 7757 6412
rect 7791 6440 7803 6443
rect 8110 6440 8116 6452
rect 7791 6412 8116 6440
rect 7791 6409 7803 6412
rect 7745 6403 7803 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 8294 6400 8300 6452
rect 8352 6440 8358 6452
rect 10778 6440 10784 6452
rect 8352 6412 10784 6440
rect 8352 6400 8358 6412
rect 10778 6400 10784 6412
rect 10836 6400 10842 6452
rect 12621 6443 12679 6449
rect 12176 6412 12572 6440
rect 12176 6384 12204 6412
rect 2222 6372 2228 6384
rect 1872 6344 2228 6372
rect 1872 6316 1900 6344
rect 2222 6332 2228 6344
rect 2280 6372 2286 6384
rect 2280 6344 2774 6372
rect 2280 6332 2286 6344
rect 1762 6304 1768 6316
rect 1723 6276 1768 6304
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 1854 6264 1860 6316
rect 1912 6304 1918 6316
rect 2130 6313 2136 6316
rect 2124 6304 2136 6313
rect 1912 6276 1957 6304
rect 2091 6276 2136 6304
rect 1912 6264 1918 6276
rect 2124 6267 2136 6276
rect 2130 6264 2136 6267
rect 2188 6264 2194 6316
rect 2746 6304 2774 6344
rect 4154 6332 4160 6384
rect 4212 6372 4218 6384
rect 4212 6344 6408 6372
rect 4212 6332 4218 6344
rect 4816 6316 4844 6344
rect 3329 6307 3387 6313
rect 3329 6304 3341 6307
rect 2746 6276 3341 6304
rect 3329 6273 3341 6276
rect 3375 6273 3387 6307
rect 3329 6267 3387 6273
rect 3596 6307 3654 6313
rect 3596 6273 3608 6307
rect 3642 6304 3654 6307
rect 4522 6304 4528 6316
rect 3642 6276 4528 6304
rect 3642 6273 3654 6276
rect 3596 6267 3654 6273
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 4798 6304 4804 6316
rect 4711 6276 4804 6304
rect 4798 6264 4804 6276
rect 4856 6264 4862 6316
rect 5068 6307 5126 6313
rect 5068 6304 5080 6307
rect 4917 6276 5080 6304
rect 4917 6236 4945 6276
rect 5068 6273 5080 6276
rect 5114 6304 5126 6307
rect 5350 6304 5356 6316
rect 5114 6276 5356 6304
rect 5114 6273 5126 6276
rect 5068 6267 5126 6273
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 6380 6313 6408 6344
rect 7190 6332 7196 6384
rect 7248 6372 7254 6384
rect 7248 6344 9352 6372
rect 7248 6332 7254 6344
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6304 6423 6307
rect 6454 6304 6460 6316
rect 6411 6276 6460 6304
rect 6411 6273 6423 6276
rect 6365 6267 6423 6273
rect 6454 6264 6460 6276
rect 6512 6264 6518 6316
rect 6632 6307 6690 6313
rect 6632 6273 6644 6307
rect 6678 6304 6690 6307
rect 7006 6304 7012 6316
rect 6678 6276 7012 6304
rect 6678 6273 6690 6276
rect 6632 6267 6690 6273
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 7742 6264 7748 6316
rect 7800 6304 7806 6316
rect 7837 6307 7895 6313
rect 7837 6304 7849 6307
rect 7800 6276 7849 6304
rect 7800 6264 7806 6276
rect 7837 6273 7849 6276
rect 7883 6273 7895 6307
rect 7837 6267 7895 6273
rect 8104 6307 8162 6313
rect 8104 6273 8116 6307
rect 8150 6304 8162 6307
rect 8478 6304 8484 6316
rect 8150 6276 8484 6304
rect 8150 6273 8162 6276
rect 8104 6267 8162 6273
rect 8478 6264 8484 6276
rect 8536 6264 8542 6316
rect 9324 6304 9352 6344
rect 9398 6332 9404 6384
rect 9456 6372 9462 6384
rect 9554 6375 9612 6381
rect 9554 6372 9566 6375
rect 9456 6344 9566 6372
rect 9456 6332 9462 6344
rect 9554 6341 9566 6344
rect 9600 6341 9612 6375
rect 9674 6372 9680 6384
rect 9554 6335 9612 6341
rect 9646 6332 9680 6372
rect 9732 6332 9738 6384
rect 10134 6332 10140 6384
rect 10192 6372 10198 6384
rect 11514 6372 11520 6384
rect 10192 6344 11520 6372
rect 10192 6332 10198 6344
rect 11514 6332 11520 6344
rect 11572 6332 11578 6384
rect 12158 6332 12164 6384
rect 12216 6332 12222 6384
rect 9646 6304 9674 6332
rect 9324 6276 9674 6304
rect 9858 6264 9864 6316
rect 9916 6304 9922 6316
rect 11241 6307 11299 6313
rect 9916 6276 11192 6304
rect 9916 6264 9922 6276
rect 11164 6248 11192 6276
rect 11241 6273 11253 6307
rect 11287 6304 11299 6307
rect 11606 6304 11612 6316
rect 11287 6276 11612 6304
rect 11287 6273 11299 6276
rect 11241 6267 11299 6273
rect 11606 6264 11612 6276
rect 11664 6264 11670 6316
rect 11698 6264 11704 6316
rect 11756 6304 11762 6316
rect 11885 6307 11943 6313
rect 11885 6304 11897 6307
rect 11756 6276 11897 6304
rect 11756 6264 11762 6276
rect 11885 6273 11897 6276
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 11977 6307 12035 6313
rect 11977 6273 11989 6307
rect 12023 6304 12035 6307
rect 12544 6304 12572 6412
rect 12621 6409 12633 6443
rect 12667 6409 12679 6443
rect 12621 6403 12679 6409
rect 12713 6443 12771 6449
rect 12713 6409 12725 6443
rect 12759 6440 12771 6443
rect 13081 6443 13139 6449
rect 12759 6412 13032 6440
rect 12759 6409 12771 6412
rect 12713 6403 12771 6409
rect 12636 6372 12664 6403
rect 12894 6372 12900 6384
rect 12636 6344 12900 6372
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 13004 6372 13032 6412
rect 13081 6409 13093 6443
rect 13127 6440 13139 6443
rect 13538 6440 13544 6452
rect 13127 6412 13400 6440
rect 13499 6412 13544 6440
rect 13127 6409 13139 6412
rect 13081 6403 13139 6409
rect 13262 6372 13268 6384
rect 13004 6344 13268 6372
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 13372 6372 13400 6412
rect 13538 6400 13544 6412
rect 13596 6400 13602 6452
rect 13998 6440 14004 6452
rect 13959 6412 14004 6440
rect 13998 6400 14004 6412
rect 14056 6400 14062 6452
rect 14090 6400 14096 6452
rect 14148 6440 14154 6452
rect 14642 6440 14648 6452
rect 14148 6412 14648 6440
rect 14148 6400 14154 6412
rect 14642 6400 14648 6412
rect 14700 6400 14706 6452
rect 13633 6375 13691 6381
rect 13633 6372 13645 6375
rect 13372 6344 13645 6372
rect 13633 6341 13645 6344
rect 13679 6341 13691 6375
rect 14918 6372 14924 6384
rect 13633 6335 13691 6341
rect 13786 6344 14924 6372
rect 13786 6304 13814 6344
rect 14918 6332 14924 6344
rect 14976 6332 14982 6384
rect 12023 6276 12204 6304
rect 12544 6276 13814 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 9306 6236 9312 6248
rect 4816 6208 4945 6236
rect 9267 6208 9312 6236
rect 4816 6168 4844 6208
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 10778 6196 10784 6248
rect 10836 6236 10842 6248
rect 10965 6239 11023 6245
rect 10965 6236 10977 6239
rect 10836 6208 10977 6236
rect 10836 6196 10842 6208
rect 10965 6205 10977 6208
rect 11011 6205 11023 6239
rect 10965 6199 11023 6205
rect 11146 6196 11152 6248
rect 11204 6236 11210 6248
rect 12066 6236 12072 6248
rect 11204 6208 12072 6236
rect 11204 6196 11210 6208
rect 12066 6196 12072 6208
rect 12124 6196 12130 6248
rect 12176 6236 12204 6276
rect 13906 6264 13912 6316
rect 13964 6304 13970 6316
rect 14369 6307 14427 6313
rect 14369 6304 14381 6307
rect 13964 6276 14381 6304
rect 13964 6264 13970 6276
rect 14369 6273 14381 6276
rect 14415 6273 14427 6307
rect 16022 6304 16028 6316
rect 14369 6267 14427 6273
rect 14568 6276 16028 6304
rect 12250 6236 12256 6248
rect 12176 6208 12256 6236
rect 12250 6196 12256 6208
rect 12308 6196 12314 6248
rect 12529 6239 12587 6245
rect 12529 6205 12541 6239
rect 12575 6236 12587 6239
rect 12802 6236 12808 6248
rect 12575 6208 12808 6236
rect 12575 6205 12587 6208
rect 12529 6199 12587 6205
rect 12802 6196 12808 6208
rect 12860 6196 12866 6248
rect 12894 6196 12900 6248
rect 12952 6236 12958 6248
rect 13078 6236 13084 6248
rect 12952 6208 13084 6236
rect 12952 6196 12958 6208
rect 13078 6196 13084 6208
rect 13136 6196 13142 6248
rect 13814 6236 13820 6248
rect 13775 6208 13820 6236
rect 13814 6196 13820 6208
rect 13872 6196 13878 6248
rect 14458 6236 14464 6248
rect 14419 6208 14464 6236
rect 14458 6196 14464 6208
rect 14516 6196 14522 6248
rect 14568 6245 14596 6276
rect 16022 6264 16028 6276
rect 16080 6264 16086 6316
rect 14553 6239 14611 6245
rect 14553 6205 14565 6239
rect 14599 6205 14611 6239
rect 14826 6236 14832 6248
rect 14787 6208 14832 6236
rect 14553 6199 14611 6205
rect 14826 6196 14832 6208
rect 14884 6196 14890 6248
rect 4356 6140 4844 6168
rect 3237 6103 3295 6109
rect 3237 6069 3249 6103
rect 3283 6100 3295 6103
rect 4356 6100 4384 6140
rect 9030 6128 9036 6180
rect 9088 6168 9094 6180
rect 9217 6171 9275 6177
rect 9217 6168 9229 6171
rect 9088 6140 9229 6168
rect 9088 6128 9094 6140
rect 9217 6137 9229 6140
rect 9263 6137 9275 6171
rect 11517 6171 11575 6177
rect 11517 6168 11529 6171
rect 9217 6131 9275 6137
rect 10244 6140 11529 6168
rect 3283 6072 4384 6100
rect 3283 6069 3295 6072
rect 3237 6063 3295 6069
rect 4522 6060 4528 6112
rect 4580 6100 4586 6112
rect 5902 6100 5908 6112
rect 4580 6072 5908 6100
rect 4580 6060 4586 6072
rect 5902 6060 5908 6072
rect 5960 6060 5966 6112
rect 6178 6100 6184 6112
rect 6091 6072 6184 6100
rect 6178 6060 6184 6072
rect 6236 6100 6242 6112
rect 7098 6100 7104 6112
rect 6236 6072 7104 6100
rect 6236 6060 6242 6072
rect 7098 6060 7104 6072
rect 7156 6060 7162 6112
rect 7558 6060 7564 6112
rect 7616 6100 7622 6112
rect 9122 6100 9128 6112
rect 7616 6072 9128 6100
rect 7616 6060 7622 6072
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 9306 6060 9312 6112
rect 9364 6100 9370 6112
rect 10244 6100 10272 6140
rect 11517 6137 11529 6140
rect 11563 6137 11575 6171
rect 11517 6131 11575 6137
rect 11606 6128 11612 6180
rect 11664 6168 11670 6180
rect 14182 6168 14188 6180
rect 11664 6140 14188 6168
rect 11664 6128 11670 6140
rect 14182 6128 14188 6140
rect 14240 6128 14246 6180
rect 14274 6128 14280 6180
rect 14332 6168 14338 6180
rect 14642 6168 14648 6180
rect 14332 6140 14648 6168
rect 14332 6128 14338 6140
rect 14642 6128 14648 6140
rect 14700 6168 14706 6180
rect 15289 6171 15347 6177
rect 15289 6168 15301 6171
rect 14700 6140 15301 6168
rect 14700 6128 14706 6140
rect 15289 6137 15301 6140
rect 15335 6137 15347 6171
rect 15289 6131 15347 6137
rect 15565 6171 15623 6177
rect 15565 6137 15577 6171
rect 15611 6168 15623 6171
rect 15654 6168 15660 6180
rect 15611 6140 15660 6168
rect 15611 6137 15623 6140
rect 15565 6131 15623 6137
rect 15654 6128 15660 6140
rect 15712 6168 15718 6180
rect 16022 6168 16028 6180
rect 15712 6140 16028 6168
rect 15712 6128 15718 6140
rect 16022 6128 16028 6140
rect 16080 6128 16086 6180
rect 9364 6072 10272 6100
rect 10689 6103 10747 6109
rect 9364 6060 9370 6072
rect 10689 6069 10701 6103
rect 10735 6100 10747 6103
rect 10778 6100 10784 6112
rect 10735 6072 10784 6100
rect 10735 6069 10747 6072
rect 10689 6063 10747 6069
rect 10778 6060 10784 6072
rect 10836 6060 10842 6112
rect 10962 6060 10968 6112
rect 11020 6100 11026 6112
rect 11422 6100 11428 6112
rect 11020 6072 11428 6100
rect 11020 6060 11026 6072
rect 11422 6060 11428 6072
rect 11480 6100 11486 6112
rect 12894 6100 12900 6112
rect 11480 6072 12900 6100
rect 11480 6060 11486 6072
rect 12894 6060 12900 6072
rect 12952 6060 12958 6112
rect 13170 6100 13176 6112
rect 13131 6072 13176 6100
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 14918 6100 14924 6112
rect 13872 6072 14924 6100
rect 13872 6060 13878 6072
rect 14918 6060 14924 6072
rect 14976 6060 14982 6112
rect 15197 6103 15255 6109
rect 15197 6069 15209 6103
rect 15243 6100 15255 6103
rect 15930 6100 15936 6112
rect 15243 6072 15936 6100
rect 15243 6069 15255 6072
rect 15197 6063 15255 6069
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 1104 6010 16008 6032
rect 1104 5958 2824 6010
rect 2876 5958 2888 6010
rect 2940 5958 2952 6010
rect 3004 5958 3016 6010
rect 3068 5958 3080 6010
rect 3132 5958 6572 6010
rect 6624 5958 6636 6010
rect 6688 5958 6700 6010
rect 6752 5958 6764 6010
rect 6816 5958 6828 6010
rect 6880 5958 10320 6010
rect 10372 5958 10384 6010
rect 10436 5958 10448 6010
rect 10500 5958 10512 6010
rect 10564 5958 10576 6010
rect 10628 5958 14068 6010
rect 14120 5958 14132 6010
rect 14184 5958 14196 6010
rect 14248 5958 14260 6010
rect 14312 5958 14324 6010
rect 14376 5958 16008 6010
rect 1104 5936 16008 5958
rect 1946 5856 1952 5908
rect 2004 5896 2010 5908
rect 2130 5896 2136 5908
rect 2004 5868 2136 5896
rect 2004 5856 2010 5868
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 3421 5899 3479 5905
rect 3421 5865 3433 5899
rect 3467 5896 3479 5899
rect 4154 5896 4160 5908
rect 3467 5868 4160 5896
rect 3467 5865 3479 5868
rect 3421 5859 3479 5865
rect 4154 5856 4160 5868
rect 4212 5856 4218 5908
rect 5169 5899 5227 5905
rect 5169 5865 5181 5899
rect 5215 5896 5227 5899
rect 7374 5896 7380 5908
rect 5215 5868 7380 5896
rect 5215 5865 5227 5868
rect 5169 5859 5227 5865
rect 7374 5856 7380 5868
rect 7432 5856 7438 5908
rect 7466 5856 7472 5908
rect 7524 5896 7530 5908
rect 7834 5896 7840 5908
rect 7524 5868 7840 5896
rect 7524 5856 7530 5868
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 10505 5899 10563 5905
rect 8588 5868 10456 5896
rect 3786 5788 3792 5840
rect 3844 5788 3850 5840
rect 8478 5828 8484 5840
rect 8439 5800 8484 5828
rect 8478 5788 8484 5800
rect 8536 5788 8542 5840
rect 3804 5760 3832 5788
rect 3620 5732 3832 5760
rect 3620 5701 3648 5732
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5661 3663 5695
rect 3605 5655 3663 5661
rect 3789 5695 3847 5701
rect 3789 5661 3801 5695
rect 3835 5692 3847 5695
rect 4798 5692 4804 5704
rect 3835 5664 4804 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5692 5319 5695
rect 5626 5692 5632 5704
rect 5307 5664 5632 5692
rect 5307 5661 5319 5664
rect 5261 5655 5319 5661
rect 3145 5627 3203 5633
rect 3145 5593 3157 5627
rect 3191 5593 3203 5627
rect 3145 5587 3203 5593
rect 4056 5627 4114 5633
rect 4056 5593 4068 5627
rect 4102 5624 4114 5627
rect 5074 5624 5080 5636
rect 4102 5596 5080 5624
rect 4102 5593 4114 5596
rect 4056 5587 4114 5593
rect 1854 5556 1860 5568
rect 1815 5528 1860 5556
rect 1854 5516 1860 5528
rect 1912 5516 1918 5568
rect 3160 5556 3188 5587
rect 5074 5584 5080 5596
rect 5132 5584 5138 5636
rect 5258 5556 5264 5568
rect 3160 5528 5264 5556
rect 5258 5516 5264 5528
rect 5316 5556 5322 5568
rect 5368 5556 5396 5664
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 7101 5695 7159 5701
rect 7101 5661 7113 5695
rect 7147 5692 7159 5695
rect 7742 5692 7748 5704
rect 7147 5664 7748 5692
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 8588 5692 8616 5868
rect 9950 5828 9956 5840
rect 9876 5800 9956 5828
rect 8938 5720 8944 5772
rect 8996 5760 9002 5772
rect 9033 5763 9091 5769
rect 9033 5760 9045 5763
rect 8996 5732 9045 5760
rect 8996 5720 9002 5732
rect 9033 5729 9045 5732
rect 9079 5729 9091 5763
rect 9214 5760 9220 5772
rect 9175 5732 9220 5760
rect 9033 5723 9091 5729
rect 9214 5720 9220 5732
rect 9272 5720 9278 5772
rect 9876 5769 9904 5800
rect 9950 5788 9956 5800
rect 10008 5788 10014 5840
rect 10134 5788 10140 5840
rect 10192 5788 10198 5840
rect 10428 5828 10456 5868
rect 10505 5865 10517 5899
rect 10551 5896 10563 5899
rect 10551 5868 11652 5896
rect 10551 5865 10563 5868
rect 10505 5859 10563 5865
rect 10428 5800 11560 5828
rect 9861 5763 9919 5769
rect 9861 5729 9873 5763
rect 9907 5729 9919 5763
rect 10152 5760 10180 5788
rect 10689 5763 10747 5769
rect 10689 5760 10701 5763
rect 10152 5732 10701 5760
rect 9861 5723 9919 5729
rect 10689 5729 10701 5732
rect 10735 5729 10747 5763
rect 10689 5723 10747 5729
rect 10873 5763 10931 5769
rect 10873 5729 10885 5763
rect 10919 5760 10931 5763
rect 11054 5760 11060 5772
rect 10919 5732 11060 5760
rect 10919 5729 10931 5732
rect 10873 5723 10931 5729
rect 11054 5720 11060 5732
rect 11112 5720 11118 5772
rect 11532 5769 11560 5800
rect 11517 5763 11575 5769
rect 11517 5729 11529 5763
rect 11563 5729 11575 5763
rect 11624 5760 11652 5868
rect 11790 5856 11796 5908
rect 11848 5896 11854 5908
rect 12434 5896 12440 5908
rect 11848 5868 12440 5896
rect 11848 5856 11854 5868
rect 12434 5856 12440 5868
rect 12492 5856 12498 5908
rect 12894 5856 12900 5908
rect 12952 5896 12958 5908
rect 14737 5899 14795 5905
rect 12952 5868 14228 5896
rect 12952 5856 12958 5868
rect 11698 5788 11704 5840
rect 11756 5828 11762 5840
rect 12158 5828 12164 5840
rect 11756 5800 12164 5828
rect 11756 5788 11762 5800
rect 12158 5788 12164 5800
rect 12216 5788 12222 5840
rect 12618 5828 12624 5840
rect 12544 5800 12624 5828
rect 12544 5760 12572 5800
rect 12618 5788 12624 5800
rect 12676 5788 12682 5840
rect 12802 5788 12808 5840
rect 12860 5828 12866 5840
rect 12860 5800 13124 5828
rect 12860 5788 12866 5800
rect 12710 5760 12716 5772
rect 11624 5732 12572 5760
rect 12636 5732 12716 5760
rect 11517 5723 11575 5729
rect 8404 5664 8616 5692
rect 6454 5584 6460 5636
rect 6512 5624 6518 5636
rect 7368 5627 7426 5633
rect 7368 5624 7380 5627
rect 6512 5596 7380 5624
rect 6512 5584 6518 5596
rect 7368 5593 7380 5596
rect 7414 5624 7426 5627
rect 8404 5624 8432 5664
rect 8662 5652 8668 5704
rect 8720 5692 8726 5704
rect 8757 5695 8815 5701
rect 8757 5692 8769 5695
rect 8720 5664 8769 5692
rect 8720 5652 8726 5664
rect 8757 5661 8769 5664
rect 8803 5661 8815 5695
rect 8757 5655 8815 5661
rect 10137 5695 10195 5701
rect 10137 5661 10149 5695
rect 10183 5692 10195 5695
rect 10962 5692 10968 5704
rect 10183 5664 10968 5692
rect 10183 5661 10195 5664
rect 10137 5655 10195 5661
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 11606 5652 11612 5704
rect 11664 5692 11670 5704
rect 11793 5695 11851 5701
rect 11793 5692 11805 5695
rect 11664 5664 11805 5692
rect 11664 5652 11670 5664
rect 11793 5661 11805 5664
rect 11839 5661 11851 5695
rect 11793 5655 11851 5661
rect 12526 5652 12532 5704
rect 12584 5652 12590 5704
rect 12636 5701 12664 5732
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 12894 5720 12900 5772
rect 12952 5760 12958 5772
rect 13096 5760 13124 5800
rect 13262 5788 13268 5840
rect 13320 5828 13326 5840
rect 13998 5828 14004 5840
rect 13320 5800 14004 5828
rect 13320 5788 13326 5800
rect 13998 5788 14004 5800
rect 14056 5788 14062 5840
rect 13633 5763 13691 5769
rect 13633 5760 13645 5763
rect 12952 5732 12997 5760
rect 13096 5732 13645 5760
rect 12952 5720 12958 5732
rect 13633 5729 13645 5732
rect 13679 5729 13691 5763
rect 13633 5723 13691 5729
rect 12621 5695 12679 5701
rect 12621 5661 12633 5695
rect 12667 5661 12679 5695
rect 13538 5692 13544 5704
rect 13499 5664 13544 5692
rect 12621 5655 12679 5661
rect 13538 5652 13544 5664
rect 13596 5652 13602 5704
rect 7414 5596 8432 5624
rect 7414 5593 7426 5596
rect 7368 5587 7426 5593
rect 8570 5584 8576 5636
rect 8628 5624 8634 5636
rect 12066 5624 12072 5636
rect 8628 5596 12072 5624
rect 8628 5584 8634 5596
rect 12066 5584 12072 5596
rect 12124 5584 12130 5636
rect 12544 5624 12572 5652
rect 14090 5624 14096 5636
rect 12544 5596 14096 5624
rect 14090 5584 14096 5596
rect 14148 5584 14154 5636
rect 14200 5624 14228 5868
rect 14737 5865 14749 5899
rect 14783 5896 14795 5899
rect 14918 5896 14924 5908
rect 14783 5868 14924 5896
rect 14783 5865 14795 5868
rect 14737 5859 14795 5865
rect 14918 5856 14924 5868
rect 14976 5856 14982 5908
rect 15473 5899 15531 5905
rect 15473 5865 15485 5899
rect 15519 5896 15531 5899
rect 16574 5896 16580 5908
rect 15519 5868 16580 5896
rect 15519 5865 15531 5868
rect 15473 5859 15531 5865
rect 16574 5856 16580 5868
rect 16632 5856 16638 5908
rect 14826 5828 14832 5840
rect 14787 5800 14832 5828
rect 14826 5788 14832 5800
rect 14884 5788 14890 5840
rect 15289 5831 15347 5837
rect 15289 5797 15301 5831
rect 15335 5828 15347 5831
rect 16298 5828 16304 5840
rect 15335 5800 16304 5828
rect 15335 5797 15347 5800
rect 15289 5791 15347 5797
rect 16298 5788 16304 5800
rect 16356 5788 16362 5840
rect 14369 5763 14427 5769
rect 14369 5729 14381 5763
rect 14415 5760 14427 5763
rect 15746 5760 15752 5772
rect 14415 5732 15752 5760
rect 14415 5729 14427 5732
rect 14369 5723 14427 5729
rect 15746 5720 15752 5732
rect 15804 5720 15810 5772
rect 14553 5695 14611 5701
rect 14553 5661 14565 5695
rect 14599 5692 14611 5695
rect 15838 5692 15844 5704
rect 14599 5664 15844 5692
rect 14599 5661 14611 5664
rect 14553 5655 14611 5661
rect 15838 5652 15844 5664
rect 15896 5652 15902 5704
rect 14826 5624 14832 5636
rect 14200 5596 14832 5624
rect 14826 5584 14832 5596
rect 14884 5624 14890 5636
rect 15013 5627 15071 5633
rect 15013 5624 15025 5627
rect 14884 5596 15025 5624
rect 14884 5584 14890 5596
rect 15013 5593 15025 5596
rect 15059 5593 15071 5627
rect 15013 5587 15071 5593
rect 15657 5627 15715 5633
rect 15657 5593 15669 5627
rect 15703 5624 15715 5627
rect 15746 5624 15752 5636
rect 15703 5596 15752 5624
rect 15703 5593 15715 5596
rect 15657 5587 15715 5593
rect 15746 5584 15752 5596
rect 15804 5624 15810 5636
rect 16022 5624 16028 5636
rect 15804 5596 16028 5624
rect 15804 5584 15810 5596
rect 16022 5584 16028 5596
rect 16080 5584 16086 5636
rect 6546 5556 6552 5568
rect 5316 5528 5396 5556
rect 6507 5528 6552 5556
rect 5316 5516 5322 5528
rect 6546 5516 6552 5528
rect 6604 5516 6610 5568
rect 8202 5516 8208 5568
rect 8260 5556 8266 5568
rect 8588 5556 8616 5584
rect 8260 5528 8616 5556
rect 8260 5516 8266 5528
rect 9122 5516 9128 5568
rect 9180 5556 9186 5568
rect 9309 5559 9367 5565
rect 9309 5556 9321 5559
rect 9180 5528 9321 5556
rect 9180 5516 9186 5528
rect 9309 5525 9321 5528
rect 9355 5525 9367 5559
rect 9674 5556 9680 5568
rect 9635 5528 9680 5556
rect 9309 5519 9367 5525
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 9766 5516 9772 5568
rect 9824 5556 9830 5568
rect 10045 5559 10103 5565
rect 10045 5556 10057 5559
rect 9824 5528 10057 5556
rect 9824 5516 9830 5528
rect 10045 5525 10057 5528
rect 10091 5525 10103 5559
rect 10045 5519 10103 5525
rect 10502 5516 10508 5568
rect 10560 5556 10566 5568
rect 10778 5556 10784 5568
rect 10560 5528 10784 5556
rect 10560 5516 10566 5528
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 10965 5559 11023 5565
rect 10965 5525 10977 5559
rect 11011 5556 11023 5559
rect 11238 5556 11244 5568
rect 11011 5528 11244 5556
rect 11011 5525 11023 5528
rect 10965 5519 11023 5525
rect 11238 5516 11244 5528
rect 11296 5516 11302 5568
rect 11333 5559 11391 5565
rect 11333 5525 11345 5559
rect 11379 5556 11391 5559
rect 11422 5556 11428 5568
rect 11379 5528 11428 5556
rect 11379 5525 11391 5528
rect 11333 5519 11391 5525
rect 11422 5516 11428 5528
rect 11480 5516 11486 5568
rect 11514 5516 11520 5568
rect 11572 5556 11578 5568
rect 11701 5559 11759 5565
rect 11701 5556 11713 5559
rect 11572 5528 11713 5556
rect 11572 5516 11578 5528
rect 11701 5525 11713 5528
rect 11747 5556 11759 5559
rect 11790 5556 11796 5568
rect 11747 5528 11796 5556
rect 11747 5525 11759 5528
rect 11701 5519 11759 5525
rect 11790 5516 11796 5528
rect 11848 5516 11854 5568
rect 11974 5516 11980 5568
rect 12032 5556 12038 5568
rect 12161 5559 12219 5565
rect 12161 5556 12173 5559
rect 12032 5528 12173 5556
rect 12032 5516 12038 5528
rect 12161 5525 12173 5528
rect 12207 5525 12219 5559
rect 12161 5519 12219 5525
rect 12253 5559 12311 5565
rect 12253 5525 12265 5559
rect 12299 5556 12311 5559
rect 12526 5556 12532 5568
rect 12299 5528 12532 5556
rect 12299 5525 12311 5528
rect 12253 5519 12311 5525
rect 12526 5516 12532 5528
rect 12584 5516 12590 5568
rect 12618 5516 12624 5568
rect 12676 5556 12682 5568
rect 12713 5559 12771 5565
rect 12713 5556 12725 5559
rect 12676 5528 12725 5556
rect 12676 5516 12682 5528
rect 12713 5525 12725 5528
rect 12759 5525 12771 5559
rect 12713 5519 12771 5525
rect 12986 5516 12992 5568
rect 13044 5556 13050 5568
rect 13081 5559 13139 5565
rect 13081 5556 13093 5559
rect 13044 5528 13093 5556
rect 13044 5516 13050 5528
rect 13081 5525 13093 5528
rect 13127 5525 13139 5559
rect 13081 5519 13139 5525
rect 13449 5559 13507 5565
rect 13449 5525 13461 5559
rect 13495 5556 13507 5559
rect 16758 5556 16764 5568
rect 13495 5528 16764 5556
rect 13495 5525 13507 5528
rect 13449 5519 13507 5525
rect 16758 5516 16764 5528
rect 16816 5516 16822 5568
rect 1104 5466 16008 5488
rect 1104 5414 4698 5466
rect 4750 5414 4762 5466
rect 4814 5414 4826 5466
rect 4878 5414 4890 5466
rect 4942 5414 4954 5466
rect 5006 5414 8446 5466
rect 8498 5414 8510 5466
rect 8562 5414 8574 5466
rect 8626 5414 8638 5466
rect 8690 5414 8702 5466
rect 8754 5414 12194 5466
rect 12246 5414 12258 5466
rect 12310 5414 12322 5466
rect 12374 5414 12386 5466
rect 12438 5414 12450 5466
rect 12502 5414 16008 5466
rect 1104 5392 16008 5414
rect 1670 5312 1676 5364
rect 1728 5352 1734 5364
rect 1765 5355 1823 5361
rect 1765 5352 1777 5355
rect 1728 5324 1777 5352
rect 1728 5312 1734 5324
rect 1765 5321 1777 5324
rect 1811 5321 1823 5355
rect 2130 5352 2136 5364
rect 2091 5324 2136 5352
rect 1765 5315 1823 5321
rect 2130 5312 2136 5324
rect 2188 5312 2194 5364
rect 4338 5352 4344 5364
rect 2746 5324 4200 5352
rect 4299 5324 4344 5352
rect 2746 5284 2774 5324
rect 1596 5256 2774 5284
rect 1596 5157 1624 5256
rect 3786 5244 3792 5296
rect 3844 5284 3850 5296
rect 3881 5287 3939 5293
rect 3881 5284 3893 5287
rect 3844 5256 3893 5284
rect 3844 5244 3850 5256
rect 3881 5253 3893 5256
rect 3927 5253 3939 5287
rect 4172 5284 4200 5324
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 4801 5355 4859 5361
rect 4801 5321 4813 5355
rect 4847 5352 4859 5355
rect 5074 5352 5080 5364
rect 4847 5324 5080 5352
rect 4847 5321 4859 5324
rect 4801 5315 4859 5321
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 8018 5312 8024 5364
rect 8076 5352 8082 5364
rect 8938 5352 8944 5364
rect 8076 5324 8944 5352
rect 8076 5312 8082 5324
rect 8938 5312 8944 5324
rect 8996 5352 9002 5364
rect 10505 5355 10563 5361
rect 10505 5352 10517 5355
rect 8996 5324 10517 5352
rect 8996 5312 9002 5324
rect 10505 5321 10517 5324
rect 10551 5321 10563 5355
rect 10505 5315 10563 5321
rect 10594 5312 10600 5364
rect 10652 5352 10658 5364
rect 11057 5355 11115 5361
rect 11057 5352 11069 5355
rect 10652 5324 10697 5352
rect 10796 5324 11069 5352
rect 10652 5312 10658 5324
rect 5442 5284 5448 5296
rect 4172 5256 5448 5284
rect 3881 5247 3939 5253
rect 5442 5244 5448 5256
rect 5500 5244 5506 5296
rect 5914 5287 5972 5293
rect 5914 5253 5926 5287
rect 5960 5284 5972 5287
rect 6086 5284 6092 5296
rect 5960 5256 6092 5284
rect 5960 5253 5972 5256
rect 5914 5247 5972 5253
rect 6086 5244 6092 5256
rect 6144 5244 6150 5296
rect 6270 5244 6276 5296
rect 6328 5284 6334 5296
rect 7190 5284 7196 5296
rect 6328 5256 7196 5284
rect 6328 5244 6334 5256
rect 7190 5244 7196 5256
rect 7248 5244 7254 5296
rect 7500 5287 7558 5293
rect 7500 5253 7512 5287
rect 7546 5284 7558 5287
rect 7650 5284 7656 5296
rect 7546 5256 7656 5284
rect 7546 5253 7558 5256
rect 7500 5247 7558 5253
rect 7650 5244 7656 5256
rect 7708 5244 7714 5296
rect 8846 5284 8852 5296
rect 7944 5256 8852 5284
rect 2222 5216 2228 5228
rect 2183 5188 2228 5216
rect 2222 5176 2228 5188
rect 2280 5176 2286 5228
rect 2314 5176 2320 5228
rect 2372 5216 2378 5228
rect 2481 5219 2539 5225
rect 2481 5216 2493 5219
rect 2372 5188 2493 5216
rect 2372 5176 2378 5188
rect 2481 5185 2493 5188
rect 2527 5185 2539 5219
rect 2481 5179 2539 5185
rect 3234 5176 3240 5228
rect 3292 5216 3298 5228
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 3292 5188 4261 5216
rect 3292 5176 3298 5188
rect 4249 5185 4261 5188
rect 4295 5216 4307 5219
rect 5166 5216 5172 5228
rect 4295 5188 5172 5216
rect 4295 5185 4307 5188
rect 4249 5179 4307 5185
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 7742 5216 7748 5228
rect 7703 5188 7748 5216
rect 7742 5176 7748 5188
rect 7800 5216 7806 5228
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 7800 5188 7849 5216
rect 7800 5176 7806 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 1581 5151 1639 5157
rect 1581 5117 1593 5151
rect 1627 5117 1639 5151
rect 1581 5111 1639 5117
rect 1673 5151 1731 5157
rect 1673 5117 1685 5151
rect 1719 5117 1731 5151
rect 1673 5111 1731 5117
rect 4157 5151 4215 5157
rect 4157 5117 4169 5151
rect 4203 5148 4215 5151
rect 4430 5148 4436 5160
rect 4203 5120 4436 5148
rect 4203 5117 4215 5120
rect 4157 5111 4215 5117
rect 1302 5040 1308 5092
rect 1360 5080 1366 5092
rect 1688 5080 1716 5111
rect 4264 5092 4292 5120
rect 4430 5108 4436 5120
rect 4488 5108 4494 5160
rect 6181 5151 6239 5157
rect 6181 5117 6193 5151
rect 6227 5148 6239 5151
rect 6546 5148 6552 5160
rect 6227 5120 6552 5148
rect 6227 5117 6239 5120
rect 6181 5111 6239 5117
rect 1360 5052 1716 5080
rect 1360 5040 1366 5052
rect 4246 5040 4252 5092
rect 4304 5040 4310 5092
rect 5074 5080 5080 5092
rect 4540 5052 5080 5080
rect 3605 5015 3663 5021
rect 3605 4981 3617 5015
rect 3651 5012 3663 5015
rect 4540 5012 4568 5052
rect 5074 5040 5080 5052
rect 5132 5040 5138 5092
rect 3651 4984 4568 5012
rect 3651 4981 3663 4984
rect 3605 4975 3663 4981
rect 4614 4972 4620 5024
rect 4672 5012 4678 5024
rect 4709 5015 4767 5021
rect 4709 5012 4721 5015
rect 4672 4984 4721 5012
rect 4672 4972 4678 4984
rect 4709 4981 4721 4984
rect 4755 4981 4767 5015
rect 4709 4975 4767 4981
rect 4798 4972 4804 5024
rect 4856 5012 4862 5024
rect 5442 5012 5448 5024
rect 4856 4984 5448 5012
rect 4856 4972 4862 4984
rect 5442 4972 5448 4984
rect 5500 5012 5506 5024
rect 6196 5012 6224 5111
rect 6546 5108 6552 5120
rect 6604 5108 6610 5160
rect 7944 5148 7972 5256
rect 8846 5244 8852 5256
rect 8904 5244 8910 5296
rect 9677 5287 9735 5293
rect 9677 5253 9689 5287
rect 9723 5284 9735 5287
rect 10318 5284 10324 5296
rect 9723 5256 10324 5284
rect 9723 5253 9735 5256
rect 9677 5247 9735 5253
rect 10318 5244 10324 5256
rect 10376 5244 10382 5296
rect 10410 5244 10416 5296
rect 10468 5284 10474 5296
rect 10796 5284 10824 5324
rect 11057 5321 11069 5324
rect 11103 5321 11115 5355
rect 11517 5355 11575 5361
rect 11517 5352 11529 5355
rect 11057 5315 11115 5321
rect 11164 5324 11529 5352
rect 10468 5256 10824 5284
rect 10468 5244 10474 5256
rect 8110 5225 8116 5228
rect 8104 5216 8116 5225
rect 8071 5188 8116 5216
rect 8104 5179 8116 5188
rect 8168 5216 8174 5228
rect 10502 5216 10508 5228
rect 8168 5188 10508 5216
rect 8110 5176 8116 5179
rect 8168 5176 8174 5188
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 11054 5176 11060 5228
rect 11112 5216 11118 5228
rect 11164 5216 11192 5324
rect 11517 5321 11529 5324
rect 11563 5321 11575 5355
rect 11974 5352 11980 5364
rect 11935 5324 11980 5352
rect 11517 5315 11575 5321
rect 11974 5312 11980 5324
rect 12032 5312 12038 5364
rect 12894 5352 12900 5364
rect 12636 5324 12900 5352
rect 11790 5244 11796 5296
rect 11848 5284 11854 5296
rect 12526 5284 12532 5296
rect 11848 5256 12532 5284
rect 11848 5244 11854 5256
rect 12526 5244 12532 5256
rect 12584 5244 12590 5296
rect 12636 5293 12664 5324
rect 12894 5312 12900 5324
rect 12952 5312 12958 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 13004 5324 13461 5352
rect 12621 5287 12679 5293
rect 12621 5253 12633 5287
rect 12667 5253 12679 5287
rect 12621 5247 12679 5253
rect 11112 5188 11192 5216
rect 11241 5219 11299 5225
rect 11112 5176 11118 5188
rect 11241 5185 11253 5219
rect 11287 5216 11299 5219
rect 11606 5216 11612 5228
rect 11287 5188 11612 5216
rect 11287 5185 11299 5188
rect 11241 5179 11299 5185
rect 11606 5176 11612 5188
rect 11664 5176 11670 5228
rect 11885 5219 11943 5225
rect 11885 5185 11897 5219
rect 11931 5216 11943 5219
rect 11931 5188 12020 5216
rect 11931 5185 11943 5188
rect 11885 5179 11943 5185
rect 7760 5120 7972 5148
rect 6362 5080 6368 5092
rect 6323 5052 6368 5080
rect 6362 5040 6368 5052
rect 6420 5040 6426 5092
rect 5500 4984 6224 5012
rect 5500 4972 5506 4984
rect 6270 4972 6276 5024
rect 6328 5012 6334 5024
rect 7760 5012 7788 5120
rect 9214 5108 9220 5160
rect 9272 5148 9278 5160
rect 9769 5151 9827 5157
rect 9769 5148 9781 5151
rect 9272 5120 9781 5148
rect 9272 5108 9278 5120
rect 9769 5117 9781 5120
rect 9815 5117 9827 5151
rect 9769 5111 9827 5117
rect 9309 5083 9367 5089
rect 9309 5080 9321 5083
rect 8772 5052 9321 5080
rect 6328 4984 7788 5012
rect 6328 4972 6334 4984
rect 7834 4972 7840 5024
rect 7892 5012 7898 5024
rect 8772 5012 8800 5052
rect 9309 5049 9321 5052
rect 9355 5049 9367 5083
rect 9784 5080 9812 5111
rect 9858 5108 9864 5160
rect 9916 5148 9922 5160
rect 9916 5120 9961 5148
rect 9916 5108 9922 5120
rect 10226 5108 10232 5160
rect 10284 5148 10290 5160
rect 10689 5151 10747 5157
rect 10689 5148 10701 5151
rect 10284 5120 10701 5148
rect 10284 5108 10290 5120
rect 10689 5117 10701 5120
rect 10735 5117 10747 5151
rect 10689 5111 10747 5117
rect 11992 5092 12020 5188
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12713 5219 12771 5225
rect 12308 5188 12572 5216
rect 12308 5176 12314 5188
rect 12158 5148 12164 5160
rect 12119 5120 12164 5148
rect 12158 5108 12164 5120
rect 12216 5108 12222 5160
rect 12437 5151 12495 5157
rect 12437 5117 12449 5151
rect 12483 5117 12495 5151
rect 12544 5148 12572 5188
rect 12713 5185 12725 5219
rect 12759 5216 12771 5219
rect 12802 5216 12808 5228
rect 12759 5188 12808 5216
rect 12759 5185 12771 5188
rect 12713 5179 12771 5185
rect 12802 5176 12808 5188
rect 12860 5176 12866 5228
rect 13004 5216 13032 5324
rect 13449 5321 13461 5324
rect 13495 5321 13507 5355
rect 13449 5315 13507 5321
rect 13541 5355 13599 5361
rect 13541 5321 13553 5355
rect 13587 5352 13599 5355
rect 13722 5352 13728 5364
rect 13587 5324 13728 5352
rect 13587 5321 13599 5324
rect 13541 5315 13599 5321
rect 13078 5244 13084 5296
rect 13136 5284 13142 5296
rect 13556 5284 13584 5315
rect 13722 5312 13728 5324
rect 13780 5312 13786 5364
rect 13909 5355 13967 5361
rect 13909 5321 13921 5355
rect 13955 5352 13967 5355
rect 15286 5352 15292 5364
rect 13955 5324 15292 5352
rect 13955 5321 13967 5324
rect 13909 5315 13967 5321
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 15381 5355 15439 5361
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 15470 5352 15476 5364
rect 15427 5324 15476 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 15470 5312 15476 5324
rect 15528 5312 15534 5364
rect 13998 5284 14004 5296
rect 13136 5256 13584 5284
rect 13959 5256 14004 5284
rect 13136 5244 13142 5256
rect 13998 5244 14004 5256
rect 14056 5244 14062 5296
rect 14461 5287 14519 5293
rect 14461 5284 14473 5287
rect 14108 5256 14473 5284
rect 13630 5216 13636 5228
rect 12912 5188 13032 5216
rect 13372 5188 13636 5216
rect 12912 5148 12940 5188
rect 13372 5157 13400 5188
rect 13630 5176 13636 5188
rect 13688 5176 13694 5228
rect 13722 5176 13728 5228
rect 13780 5216 13786 5228
rect 14016 5216 14044 5244
rect 13780 5188 14044 5216
rect 13780 5176 13786 5188
rect 12544 5120 12940 5148
rect 13357 5151 13415 5157
rect 12437 5111 12495 5117
rect 13357 5117 13369 5151
rect 13403 5117 13415 5151
rect 14108 5148 14136 5256
rect 14461 5253 14473 5256
rect 14507 5284 14519 5287
rect 14642 5284 14648 5296
rect 14507 5256 14648 5284
rect 14507 5253 14519 5256
rect 14461 5247 14519 5253
rect 14642 5244 14648 5256
rect 14700 5244 14706 5296
rect 15197 5287 15255 5293
rect 15197 5253 15209 5287
rect 15243 5284 15255 5287
rect 15562 5284 15568 5296
rect 15243 5256 15568 5284
rect 15243 5253 15255 5256
rect 15197 5247 15255 5253
rect 15562 5244 15568 5256
rect 15620 5244 15626 5296
rect 14274 5216 14280 5228
rect 14235 5188 14280 5216
rect 14274 5176 14280 5188
rect 14332 5216 14338 5228
rect 14826 5216 14832 5228
rect 14332 5188 14832 5216
rect 14332 5176 14338 5188
rect 14826 5176 14832 5188
rect 14884 5176 14890 5228
rect 16114 5216 16120 5228
rect 14936 5188 16120 5216
rect 13357 5111 13415 5117
rect 13464 5120 14136 5148
rect 9784 5052 10272 5080
rect 9309 5043 9367 5049
rect 9214 5012 9220 5024
rect 7892 4984 8800 5012
rect 9175 4984 9220 5012
rect 7892 4972 7898 4984
rect 9214 4972 9220 4984
rect 9272 4972 9278 5024
rect 9582 4972 9588 5024
rect 9640 5012 9646 5024
rect 10137 5015 10195 5021
rect 10137 5012 10149 5015
rect 9640 4984 10149 5012
rect 9640 4972 9646 4984
rect 10137 4981 10149 4984
rect 10183 4981 10195 5015
rect 10244 5012 10272 5052
rect 11974 5040 11980 5092
rect 12032 5040 12038 5092
rect 12342 5080 12348 5092
rect 12176 5052 12348 5080
rect 12176 5012 12204 5052
rect 12342 5040 12348 5052
rect 12400 5040 12406 5092
rect 10244 4984 12204 5012
rect 10137 4975 10195 4981
rect 12250 4972 12256 5024
rect 12308 5012 12314 5024
rect 12452 5012 12480 5111
rect 13464 5080 13492 5120
rect 14182 5108 14188 5160
rect 14240 5148 14246 5160
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 14240 5120 14565 5148
rect 14240 5108 14246 5120
rect 14553 5117 14565 5120
rect 14599 5148 14611 5151
rect 14936 5148 14964 5188
rect 16114 5176 16120 5188
rect 16172 5176 16178 5228
rect 14599 5120 14964 5148
rect 15013 5151 15071 5157
rect 14599 5117 14611 5120
rect 14553 5111 14611 5117
rect 15013 5117 15025 5151
rect 15059 5148 15071 5151
rect 15470 5148 15476 5160
rect 15059 5120 15476 5148
rect 15059 5117 15071 5120
rect 15013 5111 15071 5117
rect 15470 5108 15476 5120
rect 15528 5108 15534 5160
rect 12636 5052 13492 5080
rect 12308 4984 12480 5012
rect 12308 4972 12314 4984
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 12636 5012 12664 5052
rect 14274 5040 14280 5092
rect 14332 5080 14338 5092
rect 14737 5083 14795 5089
rect 14737 5080 14749 5083
rect 14332 5052 14749 5080
rect 14332 5040 14338 5052
rect 14737 5049 14749 5052
rect 14783 5080 14795 5083
rect 15286 5080 15292 5092
rect 14783 5052 15292 5080
rect 14783 5049 14795 5052
rect 14737 5043 14795 5049
rect 15286 5040 15292 5052
rect 15344 5040 15350 5092
rect 12584 4984 12664 5012
rect 13081 5015 13139 5021
rect 12584 4972 12590 4984
rect 13081 4981 13093 5015
rect 13127 5012 13139 5015
rect 13354 5012 13360 5024
rect 13127 4984 13360 5012
rect 13127 4981 13139 4984
rect 13081 4975 13139 4981
rect 13354 4972 13360 4984
rect 13412 4972 13418 5024
rect 13814 4972 13820 5024
rect 13872 5012 13878 5024
rect 14642 5012 14648 5024
rect 13872 4984 14648 5012
rect 13872 4972 13878 4984
rect 14642 4972 14648 4984
rect 14700 4972 14706 5024
rect 15562 5012 15568 5024
rect 15523 4984 15568 5012
rect 15562 4972 15568 4984
rect 15620 5012 15626 5024
rect 16390 5012 16396 5024
rect 15620 4984 16396 5012
rect 15620 4972 15626 4984
rect 16390 4972 16396 4984
rect 16448 4972 16454 5024
rect 1104 4922 16008 4944
rect 1104 4870 2824 4922
rect 2876 4870 2888 4922
rect 2940 4870 2952 4922
rect 3004 4870 3016 4922
rect 3068 4870 3080 4922
rect 3132 4870 6572 4922
rect 6624 4870 6636 4922
rect 6688 4870 6700 4922
rect 6752 4870 6764 4922
rect 6816 4870 6828 4922
rect 6880 4870 10320 4922
rect 10372 4870 10384 4922
rect 10436 4870 10448 4922
rect 10500 4870 10512 4922
rect 10564 4870 10576 4922
rect 10628 4870 14068 4922
rect 14120 4870 14132 4922
rect 14184 4870 14196 4922
rect 14248 4870 14260 4922
rect 14312 4870 14324 4922
rect 14376 4870 16008 4922
rect 1104 4848 16008 4870
rect 2222 4808 2228 4820
rect 1872 4780 2228 4808
rect 1578 4672 1584 4684
rect 1539 4644 1584 4672
rect 1578 4632 1584 4644
rect 1636 4632 1642 4684
rect 1872 4681 1900 4780
rect 2222 4768 2228 4780
rect 2280 4768 2286 4820
rect 4430 4768 4436 4820
rect 4488 4808 4494 4820
rect 5169 4811 5227 4817
rect 4488 4780 5120 4808
rect 4488 4768 4494 4780
rect 5092 4740 5120 4780
rect 5169 4777 5181 4811
rect 5215 4808 5227 4811
rect 8110 4808 8116 4820
rect 5215 4780 8116 4808
rect 5215 4777 5227 4780
rect 5169 4771 5227 4777
rect 8110 4768 8116 4780
rect 8168 4768 8174 4820
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 8662 4808 8668 4820
rect 8260 4780 8668 4808
rect 8260 4768 8266 4780
rect 8662 4768 8668 4780
rect 8720 4768 8726 4820
rect 8757 4811 8815 4817
rect 8757 4777 8769 4811
rect 8803 4808 8815 4811
rect 9122 4808 9128 4820
rect 8803 4780 9128 4808
rect 8803 4777 8815 4780
rect 8757 4771 8815 4777
rect 9122 4768 9128 4780
rect 9180 4768 9186 4820
rect 9858 4768 9864 4820
rect 9916 4808 9922 4820
rect 9916 4780 10723 4808
rect 9916 4768 9922 4780
rect 7006 4740 7012 4752
rect 5092 4712 7012 4740
rect 7006 4700 7012 4712
rect 7064 4740 7070 4752
rect 7101 4743 7159 4749
rect 7101 4740 7113 4743
rect 7064 4712 7113 4740
rect 7064 4700 7070 4712
rect 7101 4709 7113 4712
rect 7147 4709 7159 4743
rect 7101 4703 7159 4709
rect 8478 4700 8484 4752
rect 8536 4740 8542 4752
rect 10695 4740 10723 4780
rect 10778 4768 10784 4820
rect 10836 4808 10842 4820
rect 11146 4808 11152 4820
rect 10836 4780 11152 4808
rect 10836 4768 10842 4780
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 11606 4768 11612 4820
rect 11664 4808 11670 4820
rect 12434 4808 12440 4820
rect 11664 4780 12440 4808
rect 11664 4768 11670 4780
rect 12434 4768 12440 4780
rect 12492 4768 12498 4820
rect 12989 4811 13047 4817
rect 12989 4777 13001 4811
rect 13035 4808 13047 4811
rect 14642 4808 14648 4820
rect 13035 4780 14648 4808
rect 13035 4777 13047 4780
rect 12989 4771 13047 4777
rect 14642 4768 14648 4780
rect 14700 4768 14706 4820
rect 14826 4808 14832 4820
rect 14787 4780 14832 4808
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 14918 4768 14924 4820
rect 14976 4808 14982 4820
rect 15102 4808 15108 4820
rect 14976 4780 15108 4808
rect 14976 4768 14982 4780
rect 15102 4768 15108 4780
rect 15160 4768 15166 4820
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 15565 4811 15623 4817
rect 15565 4808 15577 4811
rect 15344 4780 15577 4808
rect 15344 4768 15350 4780
rect 15565 4777 15577 4780
rect 15611 4777 15623 4811
rect 15565 4771 15623 4777
rect 8536 4712 10640 4740
rect 10695 4712 11376 4740
rect 8536 4700 8542 4712
rect 1857 4675 1915 4681
rect 1857 4641 1869 4675
rect 1903 4641 1915 4675
rect 1857 4635 1915 4641
rect 5166 4632 5172 4684
rect 5224 4672 5230 4684
rect 7282 4672 7288 4684
rect 5224 4644 7288 4672
rect 5224 4632 5230 4644
rect 7282 4632 7288 4644
rect 7340 4632 7346 4684
rect 8846 4632 8852 4684
rect 8904 4672 8910 4684
rect 9033 4675 9091 4681
rect 9033 4672 9045 4675
rect 8904 4644 9045 4672
rect 8904 4632 8910 4644
rect 9033 4641 9045 4644
rect 9079 4641 9091 4675
rect 9861 4675 9919 4681
rect 9861 4672 9873 4675
rect 9033 4635 9091 4641
rect 9232 4644 9873 4672
rect 1762 4564 1768 4616
rect 1820 4564 1826 4616
rect 2124 4607 2182 4613
rect 2124 4573 2136 4607
rect 2170 4604 2182 4607
rect 2406 4604 2412 4616
rect 2170 4576 2412 4604
rect 2170 4573 2182 4576
rect 2124 4567 2182 4573
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 3510 4564 3516 4616
rect 3568 4604 3574 4616
rect 3605 4607 3663 4613
rect 3605 4604 3617 4607
rect 3568 4576 3617 4604
rect 3568 4564 3574 4576
rect 3605 4573 3617 4576
rect 3651 4573 3663 4607
rect 3605 4567 3663 4573
rect 3789 4607 3847 4613
rect 3789 4573 3801 4607
rect 3835 4604 3847 4607
rect 4798 4604 4804 4616
rect 3835 4576 4804 4604
rect 3835 4573 3847 4576
rect 3789 4567 3847 4573
rect 4798 4564 4804 4576
rect 4856 4564 4862 4616
rect 5092 4576 6040 4604
rect 1780 4536 1808 4564
rect 4056 4539 4114 4545
rect 1780 4508 4016 4536
rect 750 4428 756 4480
rect 808 4468 814 4480
rect 1762 4468 1768 4480
rect 808 4440 1768 4468
rect 808 4428 814 4440
rect 1762 4428 1768 4440
rect 1820 4428 1826 4480
rect 3234 4468 3240 4480
rect 3195 4440 3240 4468
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 3421 4471 3479 4477
rect 3421 4437 3433 4471
rect 3467 4468 3479 4471
rect 3786 4468 3792 4480
rect 3467 4440 3792 4468
rect 3467 4437 3479 4440
rect 3421 4431 3479 4437
rect 3786 4428 3792 4440
rect 3844 4428 3850 4480
rect 3988 4468 4016 4508
rect 4056 4505 4068 4539
rect 4102 4536 4114 4539
rect 5092 4536 5120 4576
rect 5258 4536 5264 4548
rect 4102 4508 5120 4536
rect 5219 4508 5264 4536
rect 4102 4505 4114 4508
rect 4056 4499 4114 4505
rect 5258 4496 5264 4508
rect 5316 4496 5322 4548
rect 6012 4536 6040 4576
rect 6086 4564 6092 4616
rect 6144 4604 6150 4616
rect 6730 4604 6736 4616
rect 6144 4576 6736 4604
rect 6144 4564 6150 4576
rect 6730 4564 6736 4576
rect 6788 4564 6794 4616
rect 6914 4564 6920 4616
rect 6972 4604 6978 4616
rect 7009 4607 7067 4613
rect 7009 4604 7021 4607
rect 6972 4576 7021 4604
rect 6972 4564 6978 4576
rect 7009 4573 7021 4576
rect 7055 4604 7067 4607
rect 7742 4604 7748 4616
rect 7055 4576 7748 4604
rect 7055 4573 7067 4576
rect 7009 4567 7067 4573
rect 7742 4564 7748 4576
rect 7800 4604 7806 4616
rect 8481 4607 8539 4613
rect 8481 4604 8493 4607
rect 7800 4576 8493 4604
rect 7800 4564 7806 4576
rect 8481 4573 8493 4576
rect 8527 4573 8539 4607
rect 8481 4567 8539 4573
rect 8662 4564 8668 4616
rect 8720 4604 8726 4616
rect 9232 4604 9260 4644
rect 9861 4641 9873 4644
rect 9907 4641 9919 4675
rect 9861 4635 9919 4641
rect 10045 4675 10103 4681
rect 10045 4641 10057 4675
rect 10091 4672 10103 4675
rect 10318 4672 10324 4684
rect 10091 4644 10324 4672
rect 10091 4641 10103 4644
rect 10045 4635 10103 4641
rect 8720 4576 9260 4604
rect 9309 4607 9367 4613
rect 8720 4564 8726 4576
rect 9309 4573 9321 4607
rect 9355 4604 9367 4607
rect 9398 4604 9404 4616
rect 9355 4576 9404 4604
rect 9355 4573 9367 4576
rect 9309 4567 9367 4573
rect 9398 4564 9404 4576
rect 9456 4564 9462 4616
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 10137 4607 10195 4613
rect 10137 4604 10149 4607
rect 9732 4576 10149 4604
rect 9732 4564 9738 4576
rect 10137 4573 10149 4576
rect 10183 4573 10195 4607
rect 10137 4567 10195 4573
rect 6362 4536 6368 4548
rect 6012 4508 6368 4536
rect 6362 4496 6368 4508
rect 6420 4536 6426 4548
rect 8110 4536 8116 4548
rect 6420 4508 8116 4536
rect 6420 4496 6426 4508
rect 8110 4496 8116 4508
rect 8168 4496 8174 4548
rect 8202 4496 8208 4548
rect 8260 4545 8266 4548
rect 8260 4536 8272 4545
rect 10244 4536 10272 4644
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 10502 4604 10508 4616
rect 8260 4508 8305 4536
rect 9048 4508 10272 4536
rect 10336 4576 10508 4604
rect 8260 4499 8272 4508
rect 8260 4496 8266 4499
rect 6086 4468 6092 4480
rect 3988 4440 6092 4468
rect 6086 4428 6092 4440
rect 6144 4428 6150 4480
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 9048 4468 9076 4508
rect 9214 4468 9220 4480
rect 7064 4440 9076 4468
rect 9175 4440 9220 4468
rect 7064 4428 7070 4440
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 9306 4428 9312 4480
rect 9364 4468 9370 4480
rect 9582 4468 9588 4480
rect 9364 4440 9588 4468
rect 9364 4428 9370 4440
rect 9582 4428 9588 4440
rect 9640 4428 9646 4480
rect 9677 4471 9735 4477
rect 9677 4437 9689 4471
rect 9723 4468 9735 4471
rect 10336 4468 10364 4576
rect 10502 4564 10508 4576
rect 10560 4564 10566 4616
rect 10410 4496 10416 4548
rect 10468 4536 10474 4548
rect 10468 4508 10548 4536
rect 10468 4496 10474 4508
rect 10520 4477 10548 4508
rect 9723 4440 10364 4468
rect 10505 4471 10563 4477
rect 9723 4437 9735 4440
rect 9677 4431 9735 4437
rect 10505 4437 10517 4471
rect 10551 4437 10563 4471
rect 10612 4468 10640 4712
rect 10778 4672 10784 4684
rect 10739 4644 10784 4672
rect 10778 4632 10784 4644
rect 10836 4632 10842 4684
rect 10873 4675 10931 4681
rect 10873 4641 10885 4675
rect 10919 4672 10931 4675
rect 11238 4672 11244 4684
rect 10919 4644 11244 4672
rect 10919 4641 10931 4644
rect 10873 4635 10931 4641
rect 11238 4632 11244 4644
rect 11296 4632 11302 4684
rect 10962 4604 10968 4616
rect 10923 4576 10968 4604
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 11348 4604 11376 4712
rect 11422 4700 11428 4752
rect 11480 4740 11486 4752
rect 13541 4743 13599 4749
rect 11480 4712 13032 4740
rect 11480 4700 11486 4712
rect 13004 4684 13032 4712
rect 13541 4709 13553 4743
rect 13587 4740 13599 4743
rect 13630 4740 13636 4752
rect 13587 4712 13636 4740
rect 13587 4709 13599 4712
rect 13541 4703 13599 4709
rect 13630 4700 13636 4712
rect 13688 4700 13694 4752
rect 14185 4743 14243 4749
rect 14185 4709 14197 4743
rect 14231 4740 14243 4743
rect 15470 4740 15476 4752
rect 14231 4712 15476 4740
rect 14231 4709 14243 4712
rect 14185 4703 14243 4709
rect 15470 4700 15476 4712
rect 15528 4700 15534 4752
rect 11517 4675 11575 4681
rect 11517 4641 11529 4675
rect 11563 4641 11575 4675
rect 11701 4675 11759 4681
rect 11701 4672 11713 4675
rect 11517 4635 11575 4641
rect 11624 4644 11713 4672
rect 11532 4604 11560 4635
rect 11624 4616 11652 4644
rect 11701 4641 11713 4644
rect 11747 4641 11759 4675
rect 11882 4672 11888 4684
rect 11701 4635 11759 4641
rect 11808 4644 11888 4672
rect 11348 4576 11560 4604
rect 11606 4564 11612 4616
rect 11664 4564 11670 4616
rect 11808 4536 11836 4644
rect 11882 4632 11888 4644
rect 11940 4632 11946 4684
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 11992 4644 12357 4672
rect 11348 4508 11836 4536
rect 11238 4468 11244 4480
rect 10612 4440 11244 4468
rect 10505 4431 10563 4437
rect 11238 4428 11244 4440
rect 11296 4428 11302 4480
rect 11348 4477 11376 4508
rect 11333 4471 11391 4477
rect 11333 4437 11345 4471
rect 11379 4437 11391 4471
rect 11333 4431 11391 4437
rect 11698 4428 11704 4480
rect 11756 4468 11762 4480
rect 11793 4471 11851 4477
rect 11793 4468 11805 4471
rect 11756 4440 11805 4468
rect 11756 4428 11762 4440
rect 11793 4437 11805 4440
rect 11839 4437 11851 4471
rect 11793 4431 11851 4437
rect 11882 4428 11888 4480
rect 11940 4468 11946 4480
rect 11992 4468 12020 4644
rect 12345 4641 12357 4644
rect 12391 4641 12403 4675
rect 12345 4635 12403 4641
rect 12986 4632 12992 4684
rect 13044 4632 13050 4684
rect 14918 4672 14924 4684
rect 13096 4644 14924 4672
rect 12066 4564 12072 4616
rect 12124 4564 12130 4616
rect 12621 4607 12679 4613
rect 12621 4573 12633 4607
rect 12667 4604 12679 4607
rect 13096 4604 13124 4644
rect 14918 4632 14924 4644
rect 14976 4632 14982 4684
rect 15197 4675 15255 4681
rect 15197 4641 15209 4675
rect 15243 4672 15255 4675
rect 15654 4672 15660 4684
rect 15243 4644 15660 4672
rect 15243 4641 15255 4644
rect 15197 4635 15255 4641
rect 15396 4616 15424 4644
rect 15654 4632 15660 4644
rect 15712 4632 15718 4684
rect 12667 4576 13124 4604
rect 12667 4573 12679 4576
rect 12621 4567 12679 4573
rect 13262 4564 13268 4616
rect 13320 4604 13326 4616
rect 13357 4607 13415 4613
rect 13357 4604 13369 4607
rect 13320 4576 13369 4604
rect 13320 4564 13326 4576
rect 13357 4573 13369 4576
rect 13403 4573 13415 4607
rect 13357 4567 13415 4573
rect 13725 4607 13783 4613
rect 13725 4573 13737 4607
rect 13771 4604 13783 4607
rect 14182 4604 14188 4616
rect 13771 4576 14188 4604
rect 13771 4573 13783 4576
rect 13725 4567 13783 4573
rect 14182 4564 14188 4576
rect 14240 4564 14246 4616
rect 14369 4607 14427 4613
rect 14369 4573 14381 4607
rect 14415 4604 14427 4607
rect 15102 4604 15108 4616
rect 14415 4576 15108 4604
rect 14415 4573 14427 4576
rect 14369 4567 14427 4573
rect 15102 4564 15108 4576
rect 15160 4564 15166 4616
rect 15378 4564 15384 4616
rect 15436 4564 15442 4616
rect 12084 4536 12112 4564
rect 14461 4539 14519 4545
rect 14461 4536 14473 4539
rect 12084 4508 14473 4536
rect 14461 4505 14473 4508
rect 14507 4505 14519 4539
rect 15286 4536 15292 4548
rect 15247 4508 15292 4536
rect 14461 4499 14519 4505
rect 15286 4496 15292 4508
rect 15344 4496 15350 4548
rect 11940 4440 12020 4468
rect 11940 4428 11946 4440
rect 12066 4428 12072 4480
rect 12124 4468 12130 4480
rect 12161 4471 12219 4477
rect 12161 4468 12173 4471
rect 12124 4440 12173 4468
rect 12124 4428 12130 4440
rect 12161 4437 12173 4440
rect 12207 4437 12219 4471
rect 12526 4468 12532 4480
rect 12439 4440 12532 4468
rect 12161 4431 12219 4437
rect 12526 4428 12532 4440
rect 12584 4468 12590 4480
rect 13078 4468 13084 4480
rect 12584 4440 13084 4468
rect 12584 4428 12590 4440
rect 13078 4428 13084 4440
rect 13136 4428 13142 4480
rect 13173 4471 13231 4477
rect 13173 4437 13185 4471
rect 13219 4468 13231 4471
rect 13262 4468 13268 4480
rect 13219 4440 13268 4468
rect 13219 4437 13231 4440
rect 13173 4431 13231 4437
rect 13262 4428 13268 4440
rect 13320 4428 13326 4480
rect 13909 4471 13967 4477
rect 13909 4437 13921 4471
rect 13955 4468 13967 4471
rect 15746 4468 15752 4480
rect 13955 4440 15752 4468
rect 13955 4437 13967 4440
rect 13909 4431 13967 4437
rect 15746 4428 15752 4440
rect 15804 4468 15810 4480
rect 16482 4468 16488 4480
rect 15804 4440 16488 4468
rect 15804 4428 15810 4440
rect 16482 4428 16488 4440
rect 16540 4428 16546 4480
rect 1104 4378 16008 4400
rect 1104 4326 4698 4378
rect 4750 4326 4762 4378
rect 4814 4326 4826 4378
rect 4878 4326 4890 4378
rect 4942 4326 4954 4378
rect 5006 4326 8446 4378
rect 8498 4326 8510 4378
rect 8562 4326 8574 4378
rect 8626 4326 8638 4378
rect 8690 4326 8702 4378
rect 8754 4326 12194 4378
rect 12246 4326 12258 4378
rect 12310 4326 12322 4378
rect 12374 4326 12386 4378
rect 12438 4326 12450 4378
rect 12502 4326 16008 4378
rect 1104 4304 16008 4326
rect 1118 4224 1124 4276
rect 1176 4264 1182 4276
rect 1489 4267 1547 4273
rect 1489 4264 1501 4267
rect 1176 4236 1501 4264
rect 1176 4224 1182 4236
rect 1489 4233 1501 4236
rect 1535 4233 1547 4267
rect 1670 4264 1676 4276
rect 1631 4236 1676 4264
rect 1489 4227 1547 4233
rect 1504 4196 1532 4227
rect 1670 4224 1676 4236
rect 1728 4224 1734 4276
rect 1857 4267 1915 4273
rect 1857 4233 1869 4267
rect 1903 4264 1915 4267
rect 2038 4264 2044 4276
rect 1903 4236 2044 4264
rect 1903 4233 1915 4236
rect 1857 4227 1915 4233
rect 2038 4224 2044 4236
rect 2096 4264 2102 4276
rect 2314 4264 2320 4276
rect 2096 4236 2320 4264
rect 2096 4224 2102 4236
rect 2314 4224 2320 4236
rect 2372 4224 2378 4276
rect 2682 4224 2688 4276
rect 2740 4264 2746 4276
rect 3234 4264 3240 4276
rect 2740 4236 3240 4264
rect 2740 4224 2746 4236
rect 3234 4224 3240 4236
rect 3292 4224 3298 4276
rect 3878 4224 3884 4276
rect 3936 4264 3942 4276
rect 4430 4264 4436 4276
rect 3936 4236 4436 4264
rect 3936 4224 3942 4236
rect 4430 4224 4436 4236
rect 4488 4224 4494 4276
rect 8846 4264 8852 4276
rect 5561 4236 8852 4264
rect 2406 4196 2412 4208
rect 1504 4168 2412 4196
rect 2406 4156 2412 4168
rect 2464 4156 2470 4208
rect 3596 4199 3654 4205
rect 2884 4168 3188 4196
rect 1854 4088 1860 4140
rect 1912 4128 1918 4140
rect 2884 4128 2912 4168
rect 1912 4100 2912 4128
rect 1912 4088 1918 4100
rect 2958 4088 2964 4140
rect 3016 4137 3022 4140
rect 3016 4128 3028 4137
rect 3160 4128 3188 4168
rect 3596 4165 3608 4199
rect 3642 4196 3654 4199
rect 5561 4196 5589 4236
rect 8846 4224 8852 4236
rect 8904 4224 8910 4276
rect 9769 4267 9827 4273
rect 9769 4264 9781 4267
rect 8956 4236 9781 4264
rect 7742 4196 7748 4208
rect 3642 4168 5589 4196
rect 7576 4168 7748 4196
rect 3642 4165 3654 4168
rect 3596 4159 3654 4165
rect 5074 4137 5080 4140
rect 3237 4131 3295 4137
rect 3237 4128 3249 4131
rect 3016 4100 3061 4128
rect 3160 4100 3249 4128
rect 3016 4091 3028 4100
rect 3237 4097 3249 4100
rect 3283 4128 3295 4131
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 3283 4100 3341 4128
rect 3283 4097 3295 4100
rect 3237 4091 3295 4097
rect 3329 4097 3341 4100
rect 3375 4128 3387 4131
rect 4801 4131 4859 4137
rect 4801 4128 4813 4131
rect 3375 4100 4813 4128
rect 3375 4097 3387 4100
rect 3329 4091 3387 4097
rect 4801 4097 4813 4100
rect 4847 4097 4859 4131
rect 5068 4128 5080 4137
rect 4987 4100 5080 4128
rect 4801 4091 4859 4097
rect 5068 4091 5080 4100
rect 5132 4128 5138 4140
rect 6270 4128 6276 4140
rect 5132 4100 6276 4128
rect 3016 4088 3022 4091
rect 5074 4088 5080 4091
rect 5132 4088 5138 4100
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 6822 4128 6828 4140
rect 6783 4100 6828 4128
rect 6822 4088 6828 4100
rect 6880 4088 6886 4140
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 7184 4131 7242 4137
rect 6972 4100 7017 4128
rect 6972 4088 6978 4100
rect 7184 4097 7196 4131
rect 7230 4128 7242 4131
rect 7576 4128 7604 4168
rect 7742 4156 7748 4168
rect 7800 4156 7806 4208
rect 8018 4156 8024 4208
rect 8076 4196 8082 4208
rect 8956 4196 8984 4236
rect 9769 4233 9781 4236
rect 9815 4233 9827 4267
rect 9769 4227 9827 4233
rect 10502 4224 10508 4276
rect 10560 4264 10566 4276
rect 10597 4267 10655 4273
rect 10597 4264 10609 4267
rect 10560 4236 10609 4264
rect 10560 4224 10566 4236
rect 10597 4233 10609 4236
rect 10643 4233 10655 4267
rect 11517 4267 11575 4273
rect 11517 4264 11529 4267
rect 10597 4227 10655 4233
rect 11164 4236 11529 4264
rect 11164 4208 11192 4236
rect 11517 4233 11529 4236
rect 11563 4233 11575 4267
rect 11517 4227 11575 4233
rect 12618 4224 12624 4276
rect 12676 4264 12682 4276
rect 12713 4267 12771 4273
rect 12713 4264 12725 4267
rect 12676 4236 12725 4264
rect 12676 4224 12682 4236
rect 12713 4233 12725 4236
rect 12759 4233 12771 4267
rect 13078 4264 13084 4276
rect 13039 4236 13084 4264
rect 12713 4227 12771 4233
rect 8076 4168 8984 4196
rect 9033 4199 9091 4205
rect 8076 4156 8082 4168
rect 9033 4165 9045 4199
rect 9079 4196 9091 4199
rect 9398 4196 9404 4208
rect 9079 4168 9404 4196
rect 9079 4165 9091 4168
rect 9033 4159 9091 4165
rect 7230 4100 7604 4128
rect 7230 4097 7242 4100
rect 7184 4091 7242 4097
rect 7650 4088 7656 4140
rect 7708 4128 7714 4140
rect 7708 4100 7972 4128
rect 7708 4088 7714 4100
rect 6546 4060 6552 4072
rect 6507 4032 6552 4060
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 7944 3992 7972 4100
rect 8386 4088 8392 4140
rect 8444 4128 8450 4140
rect 8444 4100 8616 4128
rect 8444 4088 8450 4100
rect 8294 4020 8300 4072
rect 8352 4060 8358 4072
rect 8588 4060 8616 4100
rect 8754 4088 8760 4140
rect 8812 4128 8818 4140
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 8812 4100 8953 4128
rect 8812 4088 8818 4100
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 8941 4091 8999 4097
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 8352 4032 8524 4060
rect 8588 4032 9137 4060
rect 8352 4020 8358 4032
rect 8496 4001 8524 4032
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 8481 3995 8539 4001
rect 6104 3964 6914 3992
rect 7944 3964 8340 3992
rect 1762 3884 1768 3936
rect 1820 3924 1826 3936
rect 3510 3924 3516 3936
rect 1820 3896 3516 3924
rect 1820 3884 1826 3896
rect 3510 3884 3516 3896
rect 3568 3884 3574 3936
rect 4709 3927 4767 3933
rect 4709 3893 4721 3927
rect 4755 3924 4767 3927
rect 6104 3924 6132 3964
rect 4755 3896 6132 3924
rect 6181 3927 6239 3933
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 6181 3893 6193 3927
rect 6227 3924 6239 3927
rect 6270 3924 6276 3936
rect 6227 3896 6276 3924
rect 6227 3893 6239 3896
rect 6181 3887 6239 3893
rect 6270 3884 6276 3896
rect 6328 3884 6334 3936
rect 6886 3924 6914 3964
rect 8202 3924 8208 3936
rect 6886 3896 8208 3924
rect 8202 3884 8208 3896
rect 8260 3884 8266 3936
rect 8312 3933 8340 3964
rect 8481 3961 8493 3995
rect 8527 3992 8539 3995
rect 9232 3992 9260 4168
rect 9398 4156 9404 4168
rect 9456 4156 9462 4208
rect 9677 4199 9735 4205
rect 9677 4165 9689 4199
rect 9723 4196 9735 4199
rect 10318 4196 10324 4208
rect 9723 4168 10324 4196
rect 9723 4165 9735 4168
rect 9677 4159 9735 4165
rect 10318 4156 10324 4168
rect 10376 4156 10382 4208
rect 11054 4196 11060 4208
rect 10520 4168 11060 4196
rect 10134 4128 10140 4140
rect 9600 4100 10140 4128
rect 9600 4072 9628 4100
rect 10134 4088 10140 4100
rect 10192 4128 10198 4140
rect 10520 4137 10548 4168
rect 11054 4156 11060 4168
rect 11112 4156 11118 4208
rect 11146 4156 11152 4208
rect 11204 4156 11210 4208
rect 11238 4156 11244 4208
rect 11296 4196 11302 4208
rect 12728 4196 12756 4227
rect 13078 4224 13084 4236
rect 13136 4224 13142 4276
rect 14090 4264 14096 4276
rect 13347 4236 13676 4264
rect 14051 4236 14096 4264
rect 13347 4196 13375 4236
rect 13538 4196 13544 4208
rect 11296 4168 12664 4196
rect 12728 4168 13375 4196
rect 13499 4168 13544 4196
rect 11296 4156 11302 4168
rect 10505 4131 10563 4137
rect 10192 4100 10456 4128
rect 10192 4088 10198 4100
rect 9582 4060 9588 4072
rect 9543 4032 9588 4060
rect 9582 4020 9588 4032
rect 9640 4020 9646 4072
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 10321 4063 10379 4069
rect 10321 4060 10333 4063
rect 10008 4032 10333 4060
rect 10008 4020 10014 4032
rect 10321 4029 10333 4032
rect 10367 4029 10379 4063
rect 10428 4060 10456 4100
rect 10505 4097 10517 4131
rect 10551 4097 10563 4131
rect 11333 4131 11391 4137
rect 11333 4128 11345 4131
rect 10505 4091 10563 4097
rect 10796 4100 11345 4128
rect 10686 4060 10692 4072
rect 10428 4032 10692 4060
rect 10321 4023 10379 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 8527 3964 9260 3992
rect 8527 3961 8539 3964
rect 8481 3955 8539 3961
rect 9398 3952 9404 4004
rect 9456 3992 9462 4004
rect 10796 3992 10824 4100
rect 11333 4097 11345 4100
rect 11379 4097 11391 4131
rect 11333 4091 11391 4097
rect 11606 4088 11612 4140
rect 11664 4128 11670 4140
rect 11885 4131 11943 4137
rect 11885 4128 11897 4131
rect 11664 4100 11897 4128
rect 11664 4088 11670 4100
rect 11885 4097 11897 4100
rect 11931 4097 11943 4131
rect 12636 4128 12664 4168
rect 13538 4156 13544 4168
rect 13596 4156 13602 4208
rect 13648 4196 13676 4236
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 14182 4224 14188 4276
rect 14240 4264 14246 4276
rect 14458 4264 14464 4276
rect 14240 4236 14464 4264
rect 14240 4224 14246 4236
rect 14458 4224 14464 4236
rect 14516 4264 14522 4276
rect 15565 4267 15623 4273
rect 15565 4264 15577 4267
rect 14516 4236 15577 4264
rect 14516 4224 14522 4236
rect 15565 4233 15577 4236
rect 15611 4233 15623 4267
rect 15565 4227 15623 4233
rect 14737 4199 14795 4205
rect 13648 4168 14412 4196
rect 14274 4128 14280 4140
rect 12636 4100 13768 4128
rect 14235 4100 14280 4128
rect 11885 4091 11943 4097
rect 13556 4072 13584 4100
rect 9456 3964 10824 3992
rect 10888 4032 11744 4060
rect 9456 3952 9462 3964
rect 8297 3927 8355 3933
rect 8297 3893 8309 3927
rect 8343 3893 8355 3927
rect 8297 3887 8355 3893
rect 8386 3884 8392 3936
rect 8444 3924 8450 3936
rect 8573 3927 8631 3933
rect 8573 3924 8585 3927
rect 8444 3896 8585 3924
rect 8444 3884 8450 3896
rect 8573 3893 8585 3896
rect 8619 3893 8631 3927
rect 8573 3887 8631 3893
rect 8846 3884 8852 3936
rect 8904 3924 8910 3936
rect 9030 3924 9036 3936
rect 8904 3896 9036 3924
rect 8904 3884 8910 3896
rect 9030 3884 9036 3896
rect 9088 3924 9094 3936
rect 9950 3924 9956 3936
rect 9088 3896 9956 3924
rect 9088 3884 9094 3896
rect 9950 3884 9956 3896
rect 10008 3884 10014 3936
rect 10137 3927 10195 3933
rect 10137 3893 10149 3927
rect 10183 3924 10195 3927
rect 10888 3924 10916 4032
rect 11054 3952 11060 4004
rect 11112 3992 11118 4004
rect 11149 3995 11207 4001
rect 11149 3992 11161 3995
rect 11112 3964 11161 3992
rect 11112 3952 11118 3964
rect 11149 3961 11161 3964
rect 11195 3961 11207 3995
rect 11716 3992 11744 4032
rect 11790 4020 11796 4072
rect 11848 4060 11854 4072
rect 11977 4063 12035 4069
rect 11977 4060 11989 4063
rect 11848 4032 11989 4060
rect 11848 4020 11854 4032
rect 11977 4029 11989 4032
rect 12023 4029 12035 4063
rect 11977 4023 12035 4029
rect 12066 4020 12072 4072
rect 12124 4060 12130 4072
rect 12434 4060 12440 4072
rect 12124 4032 12169 4060
rect 12395 4032 12440 4060
rect 12124 4020 12130 4032
rect 12434 4020 12440 4032
rect 12492 4020 12498 4072
rect 12621 4063 12679 4069
rect 12621 4029 12633 4063
rect 12667 4060 12679 4063
rect 12667 4032 13492 4060
rect 12667 4029 12679 4032
rect 12621 4023 12679 4029
rect 11716 3964 12756 3992
rect 11149 3955 11207 3961
rect 10183 3896 10916 3924
rect 10965 3927 11023 3933
rect 10183 3893 10195 3896
rect 10137 3887 10195 3893
rect 10965 3893 10977 3927
rect 11011 3924 11023 3927
rect 12434 3924 12440 3936
rect 11011 3896 12440 3924
rect 11011 3893 11023 3896
rect 10965 3887 11023 3893
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 12728 3924 12756 3964
rect 12802 3952 12808 4004
rect 12860 3992 12866 4004
rect 13173 3995 13231 4001
rect 13173 3992 13185 3995
rect 12860 3964 13185 3992
rect 12860 3952 12866 3964
rect 13173 3961 13185 3964
rect 13219 3961 13231 3995
rect 13173 3955 13231 3961
rect 13262 3924 13268 3936
rect 12728 3896 13268 3924
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 13464 3924 13492 4032
rect 13538 4020 13544 4072
rect 13596 4020 13602 4072
rect 13740 4069 13768 4100
rect 14274 4088 14280 4100
rect 14332 4088 14338 4140
rect 14384 4128 14412 4168
rect 14737 4165 14749 4199
rect 14783 4196 14795 4199
rect 14826 4196 14832 4208
rect 14783 4168 14832 4196
rect 14783 4165 14795 4168
rect 14737 4159 14795 4165
rect 14826 4156 14832 4168
rect 14884 4156 14890 4208
rect 14645 4131 14703 4137
rect 14384 4100 14504 4128
rect 13633 4063 13691 4069
rect 13633 4029 13645 4063
rect 13679 4029 13691 4063
rect 13633 4023 13691 4029
rect 13725 4063 13783 4069
rect 13725 4029 13737 4063
rect 13771 4029 13783 4063
rect 14366 4060 14372 4072
rect 13725 4023 13783 4029
rect 13832 4032 14372 4060
rect 13648 3992 13676 4023
rect 13832 3992 13860 4032
rect 14366 4020 14372 4032
rect 14424 4020 14430 4072
rect 14476 4060 14504 4100
rect 14645 4097 14657 4131
rect 14691 4128 14703 4131
rect 14918 4128 14924 4140
rect 14691 4100 14924 4128
rect 14691 4097 14703 4100
rect 14645 4091 14703 4097
rect 14918 4088 14924 4100
rect 14976 4088 14982 4140
rect 15197 4063 15255 4069
rect 15197 4060 15209 4063
rect 14476 4032 15209 4060
rect 15197 4029 15209 4032
rect 15243 4029 15255 4063
rect 15197 4023 15255 4029
rect 13648 3964 13860 3992
rect 13998 3952 14004 4004
rect 14056 3992 14062 4004
rect 14461 3995 14519 4001
rect 14461 3992 14473 3995
rect 14056 3964 14473 3992
rect 14056 3952 14062 3964
rect 14461 3961 14473 3964
rect 14507 3961 14519 3995
rect 14461 3955 14519 3961
rect 14826 3952 14832 4004
rect 14884 3992 14890 4004
rect 15013 3995 15071 4001
rect 15013 3992 15025 3995
rect 14884 3964 15025 3992
rect 14884 3952 14890 3964
rect 15013 3961 15025 3964
rect 15059 3961 15071 3995
rect 15013 3955 15071 3961
rect 14642 3924 14648 3936
rect 13464 3896 14648 3924
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 14918 3884 14924 3936
rect 14976 3924 14982 3936
rect 15381 3927 15439 3933
rect 15381 3924 15393 3927
rect 14976 3896 15393 3924
rect 14976 3884 14982 3896
rect 15381 3893 15393 3896
rect 15427 3893 15439 3927
rect 15381 3887 15439 3893
rect 1104 3834 16008 3856
rect 1104 3782 2824 3834
rect 2876 3782 2888 3834
rect 2940 3782 2952 3834
rect 3004 3782 3016 3834
rect 3068 3782 3080 3834
rect 3132 3782 6572 3834
rect 6624 3782 6636 3834
rect 6688 3782 6700 3834
rect 6752 3782 6764 3834
rect 6816 3782 6828 3834
rect 6880 3782 10320 3834
rect 10372 3782 10384 3834
rect 10436 3782 10448 3834
rect 10500 3782 10512 3834
rect 10564 3782 10576 3834
rect 10628 3782 14068 3834
rect 14120 3782 14132 3834
rect 14184 3782 14196 3834
rect 14248 3782 14260 3834
rect 14312 3782 14324 3834
rect 14376 3782 16008 3834
rect 1104 3760 16008 3782
rect 1581 3723 1639 3729
rect 1581 3689 1593 3723
rect 1627 3720 1639 3723
rect 3237 3723 3295 3729
rect 1627 3692 3004 3720
rect 1627 3689 1639 3692
rect 1581 3683 1639 3689
rect 2976 3664 3004 3692
rect 3237 3689 3249 3723
rect 3283 3720 3295 3723
rect 3694 3720 3700 3732
rect 3283 3692 3700 3720
rect 3283 3689 3295 3692
rect 3237 3683 3295 3689
rect 3694 3680 3700 3692
rect 3752 3680 3758 3732
rect 3786 3680 3792 3732
rect 3844 3720 3850 3732
rect 5718 3720 5724 3732
rect 3844 3692 5724 3720
rect 3844 3680 3850 3692
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 6454 3680 6460 3732
rect 6512 3720 6518 3732
rect 6825 3723 6883 3729
rect 6825 3720 6837 3723
rect 6512 3692 6837 3720
rect 6512 3680 6518 3692
rect 6825 3689 6837 3692
rect 6871 3689 6883 3723
rect 6825 3683 6883 3689
rect 7006 3680 7012 3732
rect 7064 3680 7070 3732
rect 7653 3723 7711 3729
rect 7653 3689 7665 3723
rect 7699 3720 7711 3723
rect 8662 3720 8668 3732
rect 7699 3692 8668 3720
rect 7699 3689 7711 3692
rect 7653 3683 7711 3689
rect 8662 3680 8668 3692
rect 8720 3680 8726 3732
rect 9214 3720 9220 3732
rect 8772 3692 9220 3720
rect 2958 3612 2964 3664
rect 3016 3612 3022 3664
rect 3050 3612 3056 3664
rect 3108 3652 3114 3664
rect 3326 3652 3332 3664
rect 3108 3624 3332 3652
rect 3108 3612 3114 3624
rect 3326 3612 3332 3624
rect 3384 3612 3390 3664
rect 5169 3655 5227 3661
rect 5169 3621 5181 3655
rect 5215 3621 5227 3655
rect 5169 3615 5227 3621
rect 1854 3584 1860 3596
rect 1815 3556 1860 3584
rect 1854 3544 1860 3556
rect 1912 3544 1918 3596
rect 3789 3587 3847 3593
rect 3789 3584 3801 3587
rect 3252 3556 3801 3584
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 1765 3519 1823 3525
rect 1765 3516 1777 3519
rect 992 3488 1777 3516
rect 992 3476 998 3488
rect 1765 3485 1777 3488
rect 1811 3485 1823 3519
rect 1872 3516 1900 3544
rect 2682 3516 2688 3528
rect 1872 3488 2688 3516
rect 1765 3479 1823 3485
rect 2682 3476 2688 3488
rect 2740 3516 2746 3528
rect 3252 3516 3280 3556
rect 3789 3553 3801 3556
rect 3835 3553 3847 3587
rect 3789 3547 3847 3553
rect 2740 3488 3280 3516
rect 2740 3476 2746 3488
rect 3326 3476 3332 3528
rect 3384 3516 3390 3528
rect 4056 3519 4114 3525
rect 3384 3488 3429 3516
rect 3384 3476 3390 3488
rect 4056 3485 4068 3519
rect 4102 3516 4114 3519
rect 4522 3516 4528 3528
rect 4102 3488 4528 3516
rect 4102 3485 4114 3488
rect 4056 3479 4114 3485
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 5184 3516 5212 3615
rect 5258 3612 5264 3664
rect 5316 3652 5322 3664
rect 5316 3624 5361 3652
rect 5316 3612 5322 3624
rect 6546 3612 6552 3664
rect 6604 3652 6610 3664
rect 7024 3652 7052 3680
rect 8772 3664 8800 3692
rect 9214 3680 9220 3692
rect 9272 3680 9278 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 11238 3720 11244 3732
rect 9640 3692 11244 3720
rect 9640 3680 9646 3692
rect 11238 3680 11244 3692
rect 11296 3720 11302 3732
rect 12526 3720 12532 3732
rect 11296 3692 12532 3720
rect 11296 3680 11302 3692
rect 12526 3680 12532 3692
rect 12584 3680 12590 3732
rect 12802 3720 12808 3732
rect 12636 3692 12808 3720
rect 6604 3624 7052 3652
rect 6604 3612 6610 3624
rect 7098 3612 7104 3664
rect 7156 3652 7162 3664
rect 8386 3652 8392 3664
rect 7156 3624 8392 3652
rect 7156 3612 7162 3624
rect 8386 3612 8392 3624
rect 8444 3612 8450 3664
rect 8481 3655 8539 3661
rect 8481 3621 8493 3655
rect 8527 3621 8539 3655
rect 8754 3652 8760 3664
rect 8715 3624 8760 3652
rect 8481 3615 8539 3621
rect 5442 3584 5448 3596
rect 5403 3556 5448 3584
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 7006 3584 7012 3596
rect 6967 3556 7012 3584
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 7193 3587 7251 3593
rect 7193 3553 7205 3587
rect 7239 3584 7251 3587
rect 7374 3584 7380 3596
rect 7239 3556 7380 3584
rect 7239 3553 7251 3556
rect 7193 3547 7251 3553
rect 7374 3544 7380 3556
rect 7432 3544 7438 3596
rect 7650 3544 7656 3596
rect 7708 3584 7714 3596
rect 7926 3584 7932 3596
rect 7708 3556 7932 3584
rect 7708 3544 7714 3556
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 8021 3587 8079 3593
rect 8021 3553 8033 3587
rect 8067 3584 8079 3587
rect 8110 3584 8116 3596
rect 8067 3556 8116 3584
rect 8067 3553 8079 3556
rect 8021 3547 8079 3553
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 8496 3584 8524 3615
rect 8754 3612 8760 3624
rect 8812 3612 8818 3664
rect 9674 3652 9680 3664
rect 8965 3624 9352 3652
rect 9635 3624 9680 3652
rect 8846 3584 8852 3596
rect 8496 3556 8852 3584
rect 8846 3544 8852 3556
rect 8904 3544 8910 3596
rect 5712 3519 5770 3525
rect 5712 3516 5724 3519
rect 5184 3488 5724 3516
rect 5712 3485 5724 3488
rect 5758 3516 5770 3519
rect 8965 3516 8993 3624
rect 9125 3587 9183 3593
rect 9125 3584 9137 3587
rect 9048 3556 9137 3584
rect 9048 3528 9076 3556
rect 9125 3553 9137 3556
rect 9171 3553 9183 3587
rect 9324 3584 9352 3624
rect 9674 3612 9680 3624
rect 9732 3612 9738 3664
rect 9858 3612 9864 3664
rect 9916 3652 9922 3664
rect 10686 3652 10692 3664
rect 9916 3624 10692 3652
rect 9916 3612 9922 3624
rect 10686 3612 10692 3624
rect 10744 3612 10750 3664
rect 11422 3652 11428 3664
rect 10888 3624 11428 3652
rect 10321 3587 10379 3593
rect 10321 3584 10333 3587
rect 9324 3556 10333 3584
rect 9125 3547 9183 3553
rect 10321 3553 10333 3556
rect 10367 3553 10379 3587
rect 10321 3547 10379 3553
rect 5758 3488 8993 3516
rect 5758 3485 5770 3488
rect 5712 3479 5770 3485
rect 9030 3476 9036 3528
rect 9088 3476 9094 3528
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 10042 3516 10048 3528
rect 9355 3488 10048 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 10137 3519 10195 3525
rect 10137 3485 10149 3519
rect 10183 3516 10195 3519
rect 10888 3516 10916 3624
rect 11422 3612 11428 3624
rect 11480 3612 11486 3664
rect 12250 3612 12256 3664
rect 12308 3652 12314 3664
rect 12636 3652 12664 3692
rect 12802 3680 12808 3692
rect 12860 3680 12866 3732
rect 12894 3680 12900 3732
rect 12952 3720 12958 3732
rect 13081 3723 13139 3729
rect 13081 3720 13093 3723
rect 12952 3692 13093 3720
rect 12952 3680 12958 3692
rect 13081 3689 13093 3692
rect 13127 3689 13139 3723
rect 13081 3683 13139 3689
rect 13446 3680 13452 3732
rect 13504 3720 13510 3732
rect 15286 3720 15292 3732
rect 13504 3692 15292 3720
rect 13504 3680 13510 3692
rect 15286 3680 15292 3692
rect 15344 3680 15350 3732
rect 15378 3680 15384 3732
rect 15436 3720 15442 3732
rect 15565 3723 15623 3729
rect 15565 3720 15577 3723
rect 15436 3692 15577 3720
rect 15436 3680 15442 3692
rect 15565 3689 15577 3692
rect 15611 3689 15623 3723
rect 15565 3683 15623 3689
rect 12308 3624 12664 3652
rect 12308 3612 12314 3624
rect 13538 3612 13544 3664
rect 13596 3652 13602 3664
rect 13596 3624 13676 3652
rect 13596 3612 13602 3624
rect 10962 3544 10968 3596
rect 11020 3584 11026 3596
rect 11149 3587 11207 3593
rect 11149 3584 11161 3587
rect 11020 3556 11161 3584
rect 11020 3544 11026 3556
rect 11149 3553 11161 3556
rect 11195 3553 11207 3587
rect 11149 3547 11207 3553
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 12069 3587 12127 3593
rect 11296 3556 11836 3584
rect 11296 3544 11302 3556
rect 10183 3488 10916 3516
rect 10183 3485 10195 3488
rect 10137 3479 10195 3485
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11514 3516 11520 3528
rect 11112 3488 11520 3516
rect 11112 3476 11118 3488
rect 11514 3476 11520 3488
rect 11572 3476 11578 3528
rect 11808 3525 11836 3556
rect 12069 3553 12081 3587
rect 12115 3584 12127 3587
rect 12342 3584 12348 3596
rect 12115 3556 12348 3584
rect 12115 3553 12127 3556
rect 12069 3547 12127 3553
rect 12342 3544 12348 3556
rect 12400 3544 12406 3596
rect 13648 3593 13676 3624
rect 12897 3587 12955 3593
rect 12897 3553 12909 3587
rect 12943 3553 12955 3587
rect 12897 3547 12955 3553
rect 13633 3587 13691 3593
rect 13633 3553 13645 3587
rect 13679 3553 13691 3587
rect 13633 3547 13691 3553
rect 11793 3519 11851 3525
rect 11793 3485 11805 3519
rect 11839 3485 11851 3519
rect 11793 3479 11851 3485
rect 11974 3476 11980 3528
rect 12032 3516 12038 3528
rect 12621 3519 12679 3525
rect 12621 3516 12633 3519
rect 12032 3488 12633 3516
rect 12032 3476 12038 3488
rect 12621 3485 12633 3488
rect 12667 3485 12679 3519
rect 12621 3479 12679 3485
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 2102 3451 2160 3457
rect 2102 3448 2114 3451
rect 1728 3420 2114 3448
rect 1728 3408 1734 3420
rect 2102 3417 2114 3420
rect 2148 3448 2160 3451
rect 2314 3448 2320 3460
rect 2148 3420 2320 3448
rect 2148 3417 2160 3420
rect 2102 3411 2160 3417
rect 2314 3408 2320 3420
rect 2372 3408 2378 3460
rect 2406 3408 2412 3460
rect 2464 3448 2470 3460
rect 7006 3448 7012 3460
rect 2464 3420 7012 3448
rect 2464 3408 2470 3420
rect 7006 3408 7012 3420
rect 7064 3448 7070 3460
rect 7650 3448 7656 3460
rect 7064 3420 7656 3448
rect 7064 3408 7070 3420
rect 7650 3408 7656 3420
rect 7708 3408 7714 3460
rect 7742 3408 7748 3460
rect 7800 3448 7806 3460
rect 8113 3451 8171 3457
rect 8113 3448 8125 3451
rect 7800 3420 8125 3448
rect 7800 3408 7806 3420
rect 8113 3417 8125 3420
rect 8159 3417 8171 3451
rect 8113 3411 8171 3417
rect 8662 3408 8668 3460
rect 8720 3448 8726 3460
rect 11698 3448 11704 3460
rect 8720 3420 11704 3448
rect 8720 3408 8726 3420
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 11885 3451 11943 3457
rect 11885 3417 11897 3451
rect 11931 3417 11943 3451
rect 12912 3448 12940 3547
rect 13722 3544 13728 3596
rect 13780 3584 13786 3596
rect 15396 3584 15424 3680
rect 13780 3556 15424 3584
rect 13780 3544 13786 3556
rect 13262 3476 13268 3528
rect 13320 3516 13326 3528
rect 13449 3519 13507 3525
rect 13449 3516 13461 3519
rect 13320 3488 13461 3516
rect 13320 3476 13326 3488
rect 13449 3485 13461 3488
rect 13495 3485 13507 3519
rect 13449 3479 13507 3485
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 13596 3488 13641 3516
rect 13596 3476 13602 3488
rect 13906 3476 13912 3528
rect 13964 3516 13970 3528
rect 14936 3525 14964 3556
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 13964 3488 14105 3516
rect 13964 3476 13970 3488
rect 14093 3485 14105 3488
rect 14139 3485 14151 3519
rect 14093 3479 14151 3485
rect 14921 3519 14979 3525
rect 14921 3485 14933 3519
rect 14967 3485 14979 3519
rect 15286 3516 15292 3528
rect 15247 3488 15292 3516
rect 14921 3479 14979 3485
rect 15286 3476 15292 3488
rect 15344 3516 15350 3528
rect 15562 3516 15568 3528
rect 15344 3488 15568 3516
rect 15344 3476 15350 3488
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 14369 3451 14427 3457
rect 12912 3420 13216 3448
rect 11885 3411 11943 3417
rect 2958 3340 2964 3392
rect 3016 3380 3022 3392
rect 3234 3380 3240 3392
rect 3016 3352 3240 3380
rect 3016 3340 3022 3352
rect 3234 3340 3240 3352
rect 3292 3340 3298 3392
rect 3513 3383 3571 3389
rect 3513 3349 3525 3383
rect 3559 3380 3571 3383
rect 4522 3380 4528 3392
rect 3559 3352 4528 3380
rect 3559 3349 3571 3352
rect 3513 3343 3571 3349
rect 4522 3340 4528 3352
rect 4580 3340 4586 3392
rect 5442 3340 5448 3392
rect 5500 3380 5506 3392
rect 5902 3380 5908 3392
rect 5500 3352 5908 3380
rect 5500 3340 5506 3352
rect 5902 3340 5908 3352
rect 5960 3340 5966 3392
rect 6178 3340 6184 3392
rect 6236 3380 6242 3392
rect 6822 3380 6828 3392
rect 6236 3352 6828 3380
rect 6236 3340 6242 3352
rect 6822 3340 6828 3352
rect 6880 3340 6886 3392
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7285 3383 7343 3389
rect 7285 3380 7297 3383
rect 6972 3352 7297 3380
rect 6972 3340 6978 3352
rect 7285 3349 7297 3352
rect 7331 3349 7343 3383
rect 7285 3343 7343 3349
rect 7466 3340 7472 3392
rect 7524 3380 7530 3392
rect 9030 3380 9036 3392
rect 7524 3352 9036 3380
rect 7524 3340 7530 3352
rect 9030 3340 9036 3352
rect 9088 3340 9094 3392
rect 9214 3380 9220 3392
rect 9175 3352 9220 3380
rect 9214 3340 9220 3352
rect 9272 3340 9278 3392
rect 9766 3380 9772 3392
rect 9727 3352 9772 3380
rect 9766 3340 9772 3352
rect 9824 3340 9830 3392
rect 10229 3383 10287 3389
rect 10229 3349 10241 3383
rect 10275 3380 10287 3383
rect 10502 3380 10508 3392
rect 10275 3352 10508 3380
rect 10275 3349 10287 3352
rect 10229 3343 10287 3349
rect 10502 3340 10508 3352
rect 10560 3340 10566 3392
rect 10594 3340 10600 3392
rect 10652 3380 10658 3392
rect 10652 3352 10697 3380
rect 10652 3340 10658 3352
rect 10778 3340 10784 3392
rect 10836 3380 10842 3392
rect 10965 3383 11023 3389
rect 10965 3380 10977 3383
rect 10836 3352 10977 3380
rect 10836 3340 10842 3352
rect 10965 3349 10977 3352
rect 11011 3349 11023 3383
rect 10965 3343 11023 3349
rect 11057 3383 11115 3389
rect 11057 3349 11069 3383
rect 11103 3380 11115 3383
rect 11238 3380 11244 3392
rect 11103 3352 11244 3380
rect 11103 3349 11115 3352
rect 11057 3343 11115 3349
rect 11238 3340 11244 3352
rect 11296 3340 11302 3392
rect 11422 3380 11428 3392
rect 11383 3352 11428 3380
rect 11422 3340 11428 3352
rect 11480 3340 11486 3392
rect 11514 3340 11520 3392
rect 11572 3380 11578 3392
rect 11900 3380 11928 3411
rect 11572 3352 11928 3380
rect 11572 3340 11578 3352
rect 11974 3340 11980 3392
rect 12032 3380 12038 3392
rect 12253 3383 12311 3389
rect 12253 3380 12265 3383
rect 12032 3352 12265 3380
rect 12032 3340 12038 3352
rect 12253 3349 12265 3352
rect 12299 3349 12311 3383
rect 12253 3343 12311 3349
rect 12713 3383 12771 3389
rect 12713 3349 12725 3383
rect 12759 3380 12771 3383
rect 13078 3380 13084 3392
rect 12759 3352 13084 3380
rect 12759 3349 12771 3352
rect 12713 3343 12771 3349
rect 13078 3340 13084 3352
rect 13136 3340 13142 3392
rect 13188 3380 13216 3420
rect 14369 3417 14381 3451
rect 14415 3448 14427 3451
rect 14642 3448 14648 3460
rect 14415 3420 14648 3448
rect 14415 3417 14427 3420
rect 14369 3411 14427 3417
rect 14642 3408 14648 3420
rect 14700 3408 14706 3460
rect 13262 3380 13268 3392
rect 13188 3352 13268 3380
rect 13262 3340 13268 3352
rect 13320 3340 13326 3392
rect 13538 3340 13544 3392
rect 13596 3380 13602 3392
rect 14737 3383 14795 3389
rect 14737 3380 14749 3383
rect 13596 3352 14749 3380
rect 13596 3340 13602 3352
rect 14737 3349 14749 3352
rect 14783 3349 14795 3383
rect 15102 3380 15108 3392
rect 15063 3352 15108 3380
rect 14737 3343 14795 3349
rect 15102 3340 15108 3352
rect 15160 3340 15166 3392
rect 1104 3290 16008 3312
rect 1104 3238 4698 3290
rect 4750 3238 4762 3290
rect 4814 3238 4826 3290
rect 4878 3238 4890 3290
rect 4942 3238 4954 3290
rect 5006 3238 8446 3290
rect 8498 3238 8510 3290
rect 8562 3238 8574 3290
rect 8626 3238 8638 3290
rect 8690 3238 8702 3290
rect 8754 3238 12194 3290
rect 12246 3238 12258 3290
rect 12310 3238 12322 3290
rect 12374 3238 12386 3290
rect 12438 3238 12450 3290
rect 12502 3238 16008 3290
rect 1104 3216 16008 3238
rect 1670 3136 1676 3188
rect 1728 3176 1734 3188
rect 2225 3179 2283 3185
rect 2225 3176 2237 3179
rect 1728 3148 2237 3176
rect 1728 3136 1734 3148
rect 2225 3145 2237 3148
rect 2271 3176 2283 3179
rect 2590 3176 2596 3188
rect 2271 3148 2596 3176
rect 2271 3145 2283 3148
rect 2225 3139 2283 3145
rect 2590 3136 2596 3148
rect 2648 3136 2654 3188
rect 2685 3179 2743 3185
rect 2685 3145 2697 3179
rect 2731 3176 2743 3179
rect 6178 3176 6184 3188
rect 2731 3148 6184 3176
rect 2731 3145 2743 3148
rect 2685 3139 2743 3145
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 6362 3176 6368 3188
rect 6323 3148 6368 3176
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 7466 3176 7472 3188
rect 6748 3148 6914 3176
rect 7427 3148 7472 3176
rect 1581 3111 1639 3117
rect 1581 3077 1593 3111
rect 1627 3108 1639 3111
rect 3142 3108 3148 3120
rect 1627 3080 3148 3108
rect 1627 3077 1639 3080
rect 1581 3071 1639 3077
rect 3142 3068 3148 3080
rect 3200 3068 3206 3120
rect 3786 3068 3792 3120
rect 3844 3108 3850 3120
rect 4154 3108 4160 3120
rect 3844 3080 4160 3108
rect 3844 3068 3850 3080
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 5442 3108 5448 3120
rect 4540 3080 5448 3108
rect 1854 3040 1860 3052
rect 1815 3012 1860 3040
rect 1854 3000 1860 3012
rect 1912 3000 1918 3052
rect 2130 3000 2136 3052
rect 2188 3040 2194 3052
rect 2317 3043 2375 3049
rect 2317 3040 2329 3043
rect 2188 3012 2329 3040
rect 2188 3000 2194 3012
rect 2317 3009 2329 3012
rect 2363 3040 2375 3043
rect 2590 3040 2596 3052
rect 2363 3012 2596 3040
rect 2363 3009 2375 3012
rect 2317 3003 2375 3009
rect 2590 3000 2596 3012
rect 2648 3000 2654 3052
rect 2682 3000 2688 3052
rect 2740 3040 2746 3052
rect 2777 3043 2835 3049
rect 2777 3040 2789 3043
rect 2740 3012 2789 3040
rect 2740 3000 2746 3012
rect 2777 3009 2789 3012
rect 2823 3009 2835 3043
rect 3033 3043 3091 3049
rect 3033 3040 3045 3043
rect 2777 3003 2835 3009
rect 2884 3012 3045 3040
rect 2038 2972 2044 2984
rect 1999 2944 2044 2972
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 2884 2972 2912 3012
rect 3033 3009 3045 3012
rect 3079 3040 3091 3043
rect 3326 3040 3332 3052
rect 3079 3012 3332 3040
rect 3079 3009 3091 3012
rect 3033 3003 3091 3009
rect 3326 3000 3332 3012
rect 3384 3000 3390 3052
rect 4540 3049 4568 3080
rect 5442 3068 5448 3080
rect 5500 3068 5506 3120
rect 5721 3111 5779 3117
rect 5721 3077 5733 3111
rect 5767 3108 5779 3111
rect 5902 3108 5908 3120
rect 5767 3080 5908 3108
rect 5767 3077 5779 3080
rect 5721 3071 5779 3077
rect 5902 3068 5908 3080
rect 5960 3068 5966 3120
rect 6454 3068 6460 3120
rect 6512 3108 6518 3120
rect 6748 3117 6776 3148
rect 6733 3111 6791 3117
rect 6733 3108 6745 3111
rect 6512 3080 6745 3108
rect 6512 3068 6518 3080
rect 6733 3077 6745 3080
rect 6779 3077 6791 3111
rect 6886 3108 6914 3148
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 7558 3136 7564 3188
rect 7616 3176 7622 3188
rect 7929 3179 7987 3185
rect 7616 3148 7661 3176
rect 7616 3136 7622 3148
rect 7929 3145 7941 3179
rect 7975 3176 7987 3179
rect 10597 3179 10655 3185
rect 7975 3148 10456 3176
rect 7975 3145 7987 3148
rect 7929 3139 7987 3145
rect 8297 3111 8355 3117
rect 8297 3108 8309 3111
rect 6886 3080 8309 3108
rect 6733 3071 6791 3077
rect 8297 3077 8309 3080
rect 8343 3077 8355 3111
rect 8938 3108 8944 3120
rect 8899 3080 8944 3108
rect 8297 3071 8355 3077
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 9309 3111 9367 3117
rect 9309 3108 9321 3111
rect 9048 3080 9321 3108
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4893 3043 4951 3049
rect 4893 3040 4905 3043
rect 4672 3012 4905 3040
rect 4672 3000 4678 3012
rect 4893 3009 4905 3012
rect 4939 3009 4951 3043
rect 4893 3003 4951 3009
rect 4982 3000 4988 3052
rect 5040 3040 5046 3052
rect 5810 3040 5816 3052
rect 5040 3012 5085 3040
rect 5771 3012 5816 3040
rect 5040 3000 5046 3012
rect 5810 3000 5816 3012
rect 5868 3000 5874 3052
rect 8386 3040 8392 3052
rect 8347 3012 8392 3040
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 8662 3000 8668 3052
rect 8720 3040 8726 3052
rect 9048 3040 9076 3080
rect 9309 3077 9321 3080
rect 9355 3077 9367 3111
rect 9309 3071 9367 3077
rect 9398 3068 9404 3120
rect 9456 3108 9462 3120
rect 10226 3108 10232 3120
rect 9456 3080 9501 3108
rect 10187 3080 10232 3108
rect 9456 3068 9462 3080
rect 10226 3068 10232 3080
rect 10284 3068 10290 3120
rect 10318 3040 10324 3052
rect 8720 3012 9076 3040
rect 9140 3012 10324 3040
rect 8720 3000 8726 3012
rect 4706 2972 4712 2984
rect 2148 2944 2912 2972
rect 4667 2944 4712 2972
rect 658 2796 664 2848
rect 716 2836 722 2848
rect 2148 2836 2176 2944
rect 4706 2932 4712 2944
rect 4764 2972 4770 2984
rect 5537 2975 5595 2981
rect 5537 2972 5549 2975
rect 4764 2944 5549 2972
rect 4764 2932 4770 2944
rect 5537 2941 5549 2944
rect 5583 2941 5595 2975
rect 5537 2935 5595 2941
rect 6086 2932 6092 2984
rect 6144 2972 6150 2984
rect 6362 2972 6368 2984
rect 6144 2944 6368 2972
rect 6144 2932 6150 2944
rect 6362 2932 6368 2944
rect 6420 2972 6426 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6420 2944 6837 2972
rect 6420 2932 6426 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 6914 2932 6920 2984
rect 6972 2972 6978 2984
rect 6972 2944 7017 2972
rect 6972 2932 6978 2944
rect 7190 2932 7196 2984
rect 7248 2972 7254 2984
rect 7285 2975 7343 2981
rect 7285 2972 7297 2975
rect 7248 2944 7297 2972
rect 7248 2932 7254 2944
rect 7285 2941 7297 2944
rect 7331 2941 7343 2975
rect 7285 2935 7343 2941
rect 8113 2975 8171 2981
rect 8113 2941 8125 2975
rect 8159 2941 8171 2975
rect 8113 2935 8171 2941
rect 4341 2907 4399 2913
rect 4341 2904 4353 2907
rect 3712 2876 4353 2904
rect 716 2808 2176 2836
rect 716 2796 722 2808
rect 2314 2796 2320 2848
rect 2372 2836 2378 2848
rect 3712 2836 3740 2876
rect 4341 2873 4353 2876
rect 4387 2873 4399 2907
rect 4341 2867 4399 2873
rect 5353 2907 5411 2913
rect 5353 2873 5365 2907
rect 5399 2904 5411 2907
rect 5626 2904 5632 2916
rect 5399 2876 5632 2904
rect 5399 2873 5411 2876
rect 5353 2867 5411 2873
rect 5626 2864 5632 2876
rect 5684 2864 5690 2916
rect 6181 2907 6239 2913
rect 6181 2873 6193 2907
rect 6227 2904 6239 2907
rect 6546 2904 6552 2916
rect 6227 2876 6552 2904
rect 6227 2873 6239 2876
rect 6181 2867 6239 2873
rect 6546 2864 6552 2876
rect 6604 2864 6610 2916
rect 6730 2864 6736 2916
rect 6788 2904 6794 2916
rect 8128 2904 8156 2935
rect 8754 2904 8760 2916
rect 6788 2876 8156 2904
rect 8715 2876 8760 2904
rect 6788 2864 6794 2876
rect 8754 2864 8760 2876
rect 8812 2864 8818 2916
rect 2372 2808 3740 2836
rect 4157 2839 4215 2845
rect 2372 2796 2378 2808
rect 4157 2805 4169 2839
rect 4203 2836 4215 2839
rect 9140 2836 9168 3012
rect 10060 2981 10088 3012
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 10428 3040 10456 3148
rect 10597 3145 10609 3179
rect 10643 3145 10655 3179
rect 10597 3139 10655 3145
rect 10612 3108 10640 3139
rect 11054 3136 11060 3188
rect 11112 3176 11118 3188
rect 11241 3179 11299 3185
rect 11241 3176 11253 3179
rect 11112 3148 11253 3176
rect 11112 3136 11118 3148
rect 11241 3145 11253 3148
rect 11287 3145 11299 3179
rect 11241 3139 11299 3145
rect 11517 3179 11575 3185
rect 11517 3145 11529 3179
rect 11563 3176 11575 3179
rect 11790 3176 11796 3188
rect 11563 3148 11796 3176
rect 11563 3145 11575 3148
rect 11517 3139 11575 3145
rect 11790 3136 11796 3148
rect 11848 3136 11854 3188
rect 11974 3136 11980 3188
rect 12032 3136 12038 3188
rect 12713 3179 12771 3185
rect 12713 3176 12725 3179
rect 12176 3148 12725 3176
rect 11992 3108 12020 3136
rect 12176 3120 12204 3148
rect 12713 3145 12725 3148
rect 12759 3145 12771 3179
rect 12713 3139 12771 3145
rect 13170 3136 13176 3188
rect 13228 3136 13234 3188
rect 13262 3136 13268 3188
rect 13320 3176 13326 3188
rect 14458 3176 14464 3188
rect 13320 3148 14464 3176
rect 13320 3136 13326 3148
rect 14458 3136 14464 3148
rect 14516 3136 14522 3188
rect 15194 3176 15200 3188
rect 14568 3148 15200 3176
rect 10612 3080 11100 3108
rect 11072 3052 11100 3080
rect 11716 3080 12020 3108
rect 10778 3040 10784 3052
rect 10428 3012 10784 3040
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 11054 3000 11060 3052
rect 11112 3000 11118 3052
rect 11149 3043 11207 3049
rect 11149 3009 11161 3043
rect 11195 3040 11207 3043
rect 11716 3040 11744 3080
rect 12158 3068 12164 3120
rect 12216 3068 12222 3120
rect 12250 3068 12256 3120
rect 12308 3108 12314 3120
rect 12618 3108 12624 3120
rect 12308 3080 12624 3108
rect 12308 3068 12314 3080
rect 12618 3068 12624 3080
rect 12676 3068 12682 3120
rect 13188 3108 13216 3136
rect 12728 3080 13216 3108
rect 11195 3012 11744 3040
rect 11885 3043 11943 3049
rect 11195 3009 11207 3012
rect 11149 3003 11207 3009
rect 11885 3009 11897 3043
rect 11931 3009 11943 3043
rect 11885 3003 11943 3009
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3040 12035 3043
rect 12728 3040 12756 3080
rect 12023 3012 12756 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2941 9275 2975
rect 9217 2935 9275 2941
rect 10045 2975 10103 2981
rect 10045 2941 10057 2975
rect 10091 2941 10103 2975
rect 10045 2935 10103 2941
rect 10137 2975 10195 2981
rect 10137 2941 10149 2975
rect 10183 2972 10195 2975
rect 10594 2972 10600 2984
rect 10183 2944 10600 2972
rect 10183 2941 10195 2944
rect 10137 2935 10195 2941
rect 9232 2904 9260 2935
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 10686 2932 10692 2984
rect 10744 2972 10750 2984
rect 10965 2975 11023 2981
rect 10965 2972 10977 2975
rect 10744 2944 10977 2972
rect 10744 2932 10750 2944
rect 10965 2941 10977 2944
rect 11011 2941 11023 2975
rect 10965 2935 11023 2941
rect 11698 2932 11704 2984
rect 11756 2972 11762 2984
rect 11900 2972 11928 3003
rect 12802 3000 12808 3052
rect 12860 3040 12866 3052
rect 13173 3043 13231 3049
rect 13173 3040 13185 3043
rect 12860 3012 13185 3040
rect 12860 3000 12866 3012
rect 13173 3009 13185 3012
rect 13219 3009 13231 3043
rect 13173 3003 13231 3009
rect 13446 3000 13452 3052
rect 13504 3040 13510 3052
rect 14568 3049 14596 3148
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 15378 3136 15384 3188
rect 15436 3176 15442 3188
rect 16666 3176 16672 3188
rect 15436 3148 16672 3176
rect 15436 3136 15442 3148
rect 16666 3136 16672 3148
rect 16724 3136 16730 3188
rect 14921 3111 14979 3117
rect 14921 3077 14933 3111
rect 14967 3108 14979 3111
rect 16942 3108 16948 3120
rect 14967 3080 16948 3108
rect 14967 3077 14979 3080
rect 14921 3071 14979 3077
rect 16942 3068 16948 3080
rect 17000 3068 17006 3120
rect 13725 3043 13783 3049
rect 13725 3040 13737 3043
rect 13504 3012 13737 3040
rect 13504 3000 13510 3012
rect 13725 3009 13737 3012
rect 13771 3009 13783 3043
rect 13725 3003 13783 3009
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3009 14703 3043
rect 14645 3003 14703 3009
rect 11756 2944 11928 2972
rect 12161 2975 12219 2981
rect 11756 2932 11762 2944
rect 12161 2941 12173 2975
rect 12207 2972 12219 2975
rect 12250 2972 12256 2984
rect 12207 2944 12256 2972
rect 12207 2941 12219 2944
rect 12161 2935 12219 2941
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 12437 2975 12495 2981
rect 12437 2941 12449 2975
rect 12483 2941 12495 2975
rect 12437 2935 12495 2941
rect 12621 2975 12679 2981
rect 12621 2941 12633 2975
rect 12667 2941 12679 2975
rect 13357 2975 13415 2981
rect 13357 2972 13369 2975
rect 12621 2935 12679 2941
rect 13188 2944 13369 2972
rect 9490 2904 9496 2916
rect 9232 2876 9496 2904
rect 9490 2864 9496 2876
rect 9548 2904 9554 2916
rect 12452 2904 12480 2935
rect 9548 2876 12480 2904
rect 9548 2864 9554 2876
rect 4203 2808 9168 2836
rect 9769 2839 9827 2845
rect 4203 2805 4215 2808
rect 4157 2799 4215 2805
rect 9769 2805 9781 2839
rect 9815 2836 9827 2839
rect 10042 2836 10048 2848
rect 9815 2808 10048 2836
rect 9815 2805 9827 2808
rect 9769 2799 9827 2805
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 10962 2796 10968 2848
rect 11020 2836 11026 2848
rect 12636 2836 12664 2935
rect 13188 2916 13216 2944
rect 13357 2941 13369 2944
rect 13403 2941 13415 2975
rect 13357 2935 13415 2941
rect 13630 2932 13636 2984
rect 13688 2972 13694 2984
rect 13814 2972 13820 2984
rect 13688 2944 13820 2972
rect 13688 2932 13694 2944
rect 13814 2932 13820 2944
rect 13872 2932 13878 2984
rect 14001 2975 14059 2981
rect 14001 2941 14013 2975
rect 14047 2972 14059 2975
rect 14458 2972 14464 2984
rect 14047 2944 14464 2972
rect 14047 2941 14059 2944
rect 14001 2935 14059 2941
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 14660 2972 14688 3003
rect 14826 3000 14832 3052
rect 14884 3040 14890 3052
rect 15197 3043 15255 3049
rect 15197 3040 15209 3043
rect 14884 3012 15209 3040
rect 14884 3000 14890 3012
rect 15197 3009 15209 3012
rect 15243 3040 15255 3043
rect 15838 3040 15844 3052
rect 15243 3012 15844 3040
rect 15243 3009 15255 3012
rect 15197 3003 15255 3009
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 15378 2972 15384 2984
rect 14660 2944 15384 2972
rect 15378 2932 15384 2944
rect 15436 2932 15442 2984
rect 15473 2975 15531 2981
rect 15473 2941 15485 2975
rect 15519 2972 15531 2975
rect 16574 2972 16580 2984
rect 15519 2944 16580 2972
rect 15519 2941 15531 2944
rect 15473 2935 15531 2941
rect 16574 2932 16580 2944
rect 16632 2932 16638 2984
rect 13170 2864 13176 2916
rect 13228 2864 13234 2916
rect 13446 2864 13452 2916
rect 13504 2904 13510 2916
rect 15930 2904 15936 2916
rect 13504 2876 15936 2904
rect 13504 2864 13510 2876
rect 15930 2864 15936 2876
rect 15988 2864 15994 2916
rect 13078 2836 13084 2848
rect 11020 2808 12664 2836
rect 13039 2808 13084 2836
rect 11020 2796 11026 2808
rect 13078 2796 13084 2808
rect 13136 2796 13142 2848
rect 14369 2839 14427 2845
rect 14369 2805 14381 2839
rect 14415 2836 14427 2839
rect 14458 2836 14464 2848
rect 14415 2808 14464 2836
rect 14415 2805 14427 2808
rect 14369 2799 14427 2805
rect 14458 2796 14464 2808
rect 14516 2796 14522 2848
rect 1104 2746 16008 2768
rect 1104 2694 2824 2746
rect 2876 2694 2888 2746
rect 2940 2694 2952 2746
rect 3004 2694 3016 2746
rect 3068 2694 3080 2746
rect 3132 2694 6572 2746
rect 6624 2694 6636 2746
rect 6688 2694 6700 2746
rect 6752 2694 6764 2746
rect 6816 2694 6828 2746
rect 6880 2694 10320 2746
rect 10372 2694 10384 2746
rect 10436 2694 10448 2746
rect 10500 2694 10512 2746
rect 10564 2694 10576 2746
rect 10628 2694 14068 2746
rect 14120 2694 14132 2746
rect 14184 2694 14196 2746
rect 14248 2694 14260 2746
rect 14312 2694 14324 2746
rect 14376 2694 16008 2746
rect 1104 2672 16008 2694
rect 1486 2592 1492 2644
rect 1544 2632 1550 2644
rect 4246 2632 4252 2644
rect 1544 2604 4252 2632
rect 1544 2592 1550 2604
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4522 2632 4528 2644
rect 4483 2604 4528 2632
rect 4522 2592 4528 2604
rect 4580 2592 4586 2644
rect 5353 2635 5411 2641
rect 5353 2601 5365 2635
rect 5399 2601 5411 2635
rect 5353 2595 5411 2601
rect 3142 2564 3148 2576
rect 1688 2536 3148 2564
rect 1688 2505 1716 2536
rect 3142 2524 3148 2536
rect 3200 2524 3206 2576
rect 4338 2564 4344 2576
rect 3988 2536 4344 2564
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2465 1731 2499
rect 1673 2459 1731 2465
rect 1946 2456 1952 2508
rect 2004 2496 2010 2508
rect 2133 2499 2191 2505
rect 2133 2496 2145 2499
rect 2004 2468 2145 2496
rect 2004 2456 2010 2468
rect 2133 2465 2145 2468
rect 2179 2465 2191 2499
rect 2314 2496 2320 2508
rect 2275 2468 2320 2496
rect 2133 2459 2191 2465
rect 2314 2456 2320 2468
rect 2372 2456 2378 2508
rect 2682 2456 2688 2508
rect 2740 2496 2746 2508
rect 3988 2505 4016 2536
rect 4338 2524 4344 2536
rect 4396 2524 4402 2576
rect 2961 2499 3019 2505
rect 2961 2496 2973 2499
rect 2740 2468 2973 2496
rect 2740 2456 2746 2468
rect 2961 2465 2973 2468
rect 3007 2465 3019 2499
rect 2961 2459 3019 2465
rect 3973 2499 4031 2505
rect 3973 2465 3985 2499
rect 4019 2465 4031 2499
rect 3973 2459 4031 2465
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4801 2499 4859 2505
rect 4120 2468 4165 2496
rect 4120 2456 4126 2468
rect 4801 2465 4813 2499
rect 4847 2496 4859 2499
rect 5074 2496 5080 2508
rect 4847 2468 5080 2496
rect 4847 2465 4859 2468
rect 4801 2459 4859 2465
rect 5074 2456 5080 2468
rect 5132 2456 5138 2508
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2428 1915 2431
rect 3142 2428 3148 2440
rect 1903 2400 3148 2428
rect 1903 2397 1915 2400
rect 1857 2391 1915 2397
rect 3142 2388 3148 2400
rect 3200 2388 3206 2440
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 3786 2428 3792 2440
rect 3283 2400 3792 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 4890 2428 4896 2440
rect 4264 2400 4896 2428
rect 2038 2320 2044 2372
rect 2096 2360 2102 2372
rect 2409 2363 2467 2369
rect 2409 2360 2421 2363
rect 2096 2332 2421 2360
rect 2096 2320 2102 2332
rect 2409 2329 2421 2332
rect 2455 2329 2467 2363
rect 2409 2323 2467 2329
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 4157 2363 4215 2369
rect 4157 2360 4169 2363
rect 2648 2332 4169 2360
rect 2648 2320 2654 2332
rect 4157 2329 4169 2332
rect 4203 2329 4215 2363
rect 4157 2323 4215 2329
rect 2777 2295 2835 2301
rect 2777 2261 2789 2295
rect 2823 2292 2835 2295
rect 3050 2292 3056 2304
rect 2823 2264 3056 2292
rect 2823 2261 2835 2264
rect 2777 2255 2835 2261
rect 3050 2252 3056 2264
rect 3108 2252 3114 2304
rect 3145 2295 3203 2301
rect 3145 2261 3157 2295
rect 3191 2292 3203 2295
rect 3510 2292 3516 2304
rect 3191 2264 3516 2292
rect 3191 2261 3203 2264
rect 3145 2255 3203 2261
rect 3510 2252 3516 2264
rect 3568 2252 3574 2304
rect 3605 2295 3663 2301
rect 3605 2261 3617 2295
rect 3651 2292 3663 2295
rect 4264 2292 4292 2400
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 4522 2320 4528 2372
rect 4580 2360 4586 2372
rect 4985 2363 5043 2369
rect 4985 2360 4997 2363
rect 4580 2332 4997 2360
rect 4580 2320 4586 2332
rect 4985 2329 4997 2332
rect 5031 2329 5043 2363
rect 5368 2360 5396 2595
rect 6914 2592 6920 2644
rect 6972 2632 6978 2644
rect 8754 2632 8760 2644
rect 6972 2604 8760 2632
rect 6972 2592 6978 2604
rect 8754 2592 8760 2604
rect 8812 2632 8818 2644
rect 8938 2632 8944 2644
rect 8812 2604 8944 2632
rect 8812 2592 8818 2604
rect 8938 2592 8944 2604
rect 8996 2592 9002 2644
rect 9030 2592 9036 2644
rect 9088 2592 9094 2644
rect 9306 2632 9312 2644
rect 9232 2604 9312 2632
rect 5445 2567 5503 2573
rect 5445 2533 5457 2567
rect 5491 2533 5503 2567
rect 6822 2564 6828 2576
rect 5445 2527 5503 2533
rect 6012 2536 6828 2564
rect 5460 2440 5488 2527
rect 5902 2496 5908 2508
rect 5863 2468 5908 2496
rect 5902 2456 5908 2468
rect 5960 2456 5966 2508
rect 6012 2505 6040 2536
rect 6822 2524 6828 2536
rect 6880 2524 6886 2576
rect 9048 2564 9076 2592
rect 7852 2536 9076 2564
rect 5997 2499 6055 2505
rect 5997 2465 6009 2499
rect 6043 2465 6055 2499
rect 5997 2459 6055 2465
rect 6086 2456 6092 2508
rect 6144 2496 6150 2508
rect 6457 2499 6515 2505
rect 6457 2496 6469 2499
rect 6144 2468 6469 2496
rect 6144 2456 6150 2468
rect 6457 2465 6469 2468
rect 6503 2465 6515 2499
rect 6457 2459 6515 2465
rect 6641 2499 6699 2505
rect 6641 2465 6653 2499
rect 6687 2496 6699 2499
rect 7098 2496 7104 2508
rect 6687 2468 7104 2496
rect 6687 2465 6699 2468
rect 6641 2459 6699 2465
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 7377 2499 7435 2505
rect 7377 2465 7389 2499
rect 7423 2465 7435 2499
rect 7377 2459 7435 2465
rect 7469 2499 7527 2505
rect 7469 2465 7481 2499
rect 7515 2496 7527 2499
rect 7742 2496 7748 2508
rect 7515 2468 7748 2496
rect 7515 2465 7527 2468
rect 7469 2459 7527 2465
rect 5442 2388 5448 2440
rect 5500 2388 5506 2440
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6733 2431 6791 2437
rect 6733 2397 6745 2431
rect 6779 2428 6791 2431
rect 6914 2428 6920 2440
rect 6779 2400 6920 2428
rect 6779 2397 6791 2400
rect 6733 2391 6791 2397
rect 6914 2388 6920 2400
rect 6972 2388 6978 2440
rect 7392 2428 7420 2459
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 7852 2428 7880 2536
rect 8205 2499 8263 2505
rect 8205 2465 8217 2499
rect 8251 2496 8263 2499
rect 8294 2496 8300 2508
rect 8251 2468 8300 2496
rect 8251 2465 8263 2468
rect 8205 2459 8263 2465
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 8478 2456 8484 2508
rect 8536 2496 8542 2508
rect 8754 2496 8760 2508
rect 8536 2468 8760 2496
rect 8536 2456 8542 2468
rect 8754 2456 8760 2468
rect 8812 2456 8818 2508
rect 9232 2505 9260 2604
rect 9306 2592 9312 2604
rect 9364 2592 9370 2644
rect 9398 2592 9404 2644
rect 9456 2632 9462 2644
rect 9677 2635 9735 2641
rect 9677 2632 9689 2635
rect 9456 2604 9689 2632
rect 9456 2592 9462 2604
rect 9677 2601 9689 2604
rect 9723 2601 9735 2635
rect 9677 2595 9735 2601
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 10100 2604 12664 2632
rect 10100 2592 10106 2604
rect 10962 2564 10968 2576
rect 9600 2536 10968 2564
rect 9033 2499 9091 2505
rect 9033 2465 9045 2499
rect 9079 2465 9091 2499
rect 9033 2459 9091 2465
rect 9217 2499 9275 2505
rect 9217 2465 9229 2499
rect 9263 2465 9275 2499
rect 9217 2459 9275 2465
rect 7392 2400 7880 2428
rect 7926 2388 7932 2440
rect 7984 2428 7990 2440
rect 9048 2428 9076 2459
rect 7984 2400 9076 2428
rect 7984 2388 7990 2400
rect 8389 2363 8447 2369
rect 8389 2360 8401 2363
rect 5368 2332 8401 2360
rect 4985 2323 5043 2329
rect 8389 2329 8401 2332
rect 8435 2329 8447 2363
rect 8389 2323 8447 2329
rect 8478 2320 8484 2372
rect 8536 2320 8542 2372
rect 8662 2320 8668 2372
rect 8720 2360 8726 2372
rect 8720 2332 8892 2360
rect 8720 2320 8726 2332
rect 3651 2264 4292 2292
rect 3651 2261 3663 2264
rect 3605 2255 3663 2261
rect 4338 2252 4344 2304
rect 4396 2292 4402 2304
rect 4893 2295 4951 2301
rect 4893 2292 4905 2295
rect 4396 2264 4905 2292
rect 4396 2252 4402 2264
rect 4893 2261 4905 2264
rect 4939 2292 4951 2295
rect 6454 2292 6460 2304
rect 4939 2264 6460 2292
rect 4939 2261 4951 2264
rect 4893 2255 4951 2261
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 7098 2292 7104 2304
rect 7059 2264 7104 2292
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 7558 2292 7564 2304
rect 7519 2264 7564 2292
rect 7558 2252 7564 2264
rect 7616 2252 7622 2304
rect 7926 2292 7932 2304
rect 7887 2264 7932 2292
rect 7926 2252 7932 2264
rect 7984 2252 7990 2304
rect 8294 2292 8300 2304
rect 8255 2264 8300 2292
rect 8294 2252 8300 2264
rect 8352 2252 8358 2304
rect 8496 2292 8524 2320
rect 8757 2295 8815 2301
rect 8757 2292 8769 2295
rect 8496 2264 8769 2292
rect 8757 2261 8769 2264
rect 8803 2261 8815 2295
rect 8864 2292 8892 2332
rect 8938 2320 8944 2372
rect 8996 2360 9002 2372
rect 9600 2360 9628 2536
rect 10962 2524 10968 2536
rect 11020 2524 11026 2576
rect 11790 2524 11796 2576
rect 11848 2564 11854 2576
rect 12345 2567 12403 2573
rect 12345 2564 12357 2567
rect 11848 2536 12357 2564
rect 11848 2524 11854 2536
rect 12345 2533 12357 2536
rect 12391 2533 12403 2567
rect 12636 2564 12664 2604
rect 12710 2592 12716 2644
rect 12768 2632 12774 2644
rect 13906 2632 13912 2644
rect 12768 2604 13584 2632
rect 13867 2604 13912 2632
rect 12768 2592 12774 2604
rect 13556 2564 13584 2604
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 15565 2635 15623 2641
rect 15565 2632 15577 2635
rect 14016 2604 15577 2632
rect 14016 2564 14044 2604
rect 15565 2601 15577 2604
rect 15611 2601 15623 2635
rect 15565 2595 15623 2601
rect 12636 2536 13492 2564
rect 13556 2536 14044 2564
rect 12345 2527 12403 2533
rect 9950 2496 9956 2508
rect 9911 2468 9956 2496
rect 9950 2456 9956 2468
rect 10008 2456 10014 2508
rect 10042 2456 10048 2508
rect 10100 2496 10106 2508
rect 11054 2496 11060 2508
rect 10100 2468 10145 2496
rect 11015 2468 11060 2496
rect 10100 2456 10106 2468
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2465 11207 2499
rect 11149 2459 11207 2465
rect 10226 2388 10232 2440
rect 10284 2428 10290 2440
rect 11164 2428 11192 2459
rect 11330 2456 11336 2508
rect 11388 2496 11394 2508
rect 12069 2499 12127 2505
rect 12069 2496 12081 2499
rect 11388 2468 12081 2496
rect 11388 2456 11394 2468
rect 12069 2465 12081 2468
rect 12115 2465 12127 2499
rect 12894 2496 12900 2508
rect 12855 2468 12900 2496
rect 12069 2459 12127 2465
rect 12894 2456 12900 2468
rect 12952 2456 12958 2508
rect 13262 2496 13268 2508
rect 13223 2468 13268 2496
rect 13262 2456 13268 2468
rect 13320 2456 13326 2508
rect 13464 2505 13492 2536
rect 14090 2524 14096 2576
rect 14148 2564 14154 2576
rect 14185 2567 14243 2573
rect 14185 2564 14197 2567
rect 14148 2536 14197 2564
rect 14148 2524 14154 2536
rect 14185 2533 14197 2536
rect 14231 2533 14243 2567
rect 15654 2564 15660 2576
rect 14185 2527 14243 2533
rect 14384 2536 15660 2564
rect 13449 2499 13507 2505
rect 13449 2465 13461 2499
rect 13495 2465 13507 2499
rect 13449 2459 13507 2465
rect 10284 2400 11192 2428
rect 10284 2388 10290 2400
rect 11238 2388 11244 2440
rect 11296 2428 11302 2440
rect 11514 2428 11520 2440
rect 11296 2400 11520 2428
rect 11296 2388 11302 2400
rect 11514 2388 11520 2400
rect 11572 2388 11578 2440
rect 11882 2428 11888 2440
rect 11843 2400 11888 2428
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 12526 2388 12532 2440
rect 12584 2428 12590 2440
rect 12805 2431 12863 2437
rect 12805 2428 12817 2431
rect 12584 2400 12817 2428
rect 12584 2388 12590 2400
rect 12805 2397 12817 2400
rect 12851 2397 12863 2431
rect 12805 2391 12863 2397
rect 13078 2388 13084 2440
rect 13136 2428 13142 2440
rect 14384 2437 14412 2536
rect 15654 2524 15660 2536
rect 15712 2524 15718 2576
rect 14737 2499 14795 2505
rect 14737 2465 14749 2499
rect 14783 2496 14795 2499
rect 15562 2496 15568 2508
rect 14783 2468 15568 2496
rect 14783 2465 14795 2468
rect 14737 2459 14795 2465
rect 15562 2456 15568 2468
rect 15620 2456 15626 2508
rect 13541 2431 13599 2437
rect 13541 2428 13553 2431
rect 13136 2400 13553 2428
rect 13136 2388 13142 2400
rect 13541 2397 13553 2400
rect 13587 2397 13599 2431
rect 13541 2391 13599 2397
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2428 15071 2431
rect 15746 2428 15752 2440
rect 15059 2400 15752 2428
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 8996 2332 9628 2360
rect 8996 2320 9002 2332
rect 9674 2320 9680 2372
rect 9732 2360 9738 2372
rect 9858 2360 9864 2372
rect 9732 2332 9864 2360
rect 9732 2320 9738 2332
rect 9858 2320 9864 2332
rect 9916 2320 9922 2372
rect 10137 2363 10195 2369
rect 10137 2329 10149 2363
rect 10183 2360 10195 2363
rect 10318 2360 10324 2372
rect 10183 2332 10324 2360
rect 10183 2329 10195 2332
rect 10137 2323 10195 2329
rect 10318 2320 10324 2332
rect 10376 2320 10382 2372
rect 11977 2363 12035 2369
rect 10520 2332 11836 2360
rect 9122 2292 9128 2304
rect 8864 2264 9128 2292
rect 8757 2255 8815 2261
rect 9122 2252 9128 2264
rect 9180 2252 9186 2304
rect 9306 2292 9312 2304
rect 9219 2264 9312 2292
rect 9306 2252 9312 2264
rect 9364 2292 9370 2304
rect 10410 2292 10416 2304
rect 9364 2264 10416 2292
rect 9364 2252 9370 2264
rect 10410 2252 10416 2264
rect 10468 2252 10474 2304
rect 10520 2301 10548 2332
rect 10505 2295 10563 2301
rect 10505 2261 10517 2295
rect 10551 2261 10563 2295
rect 10505 2255 10563 2261
rect 10594 2252 10600 2304
rect 10652 2292 10658 2304
rect 10962 2292 10968 2304
rect 10652 2264 10697 2292
rect 10923 2264 10968 2292
rect 10652 2252 10658 2264
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 11514 2292 11520 2304
rect 11475 2264 11520 2292
rect 11514 2252 11520 2264
rect 11572 2252 11578 2304
rect 11808 2292 11836 2332
rect 11977 2329 11989 2363
rect 12023 2360 12035 2363
rect 12618 2360 12624 2372
rect 12023 2332 12624 2360
rect 12023 2329 12035 2332
rect 11977 2323 12035 2329
rect 12618 2320 12624 2332
rect 12676 2320 12682 2372
rect 12713 2363 12771 2369
rect 12713 2329 12725 2363
rect 12759 2329 12771 2363
rect 12713 2323 12771 2329
rect 12728 2292 12756 2323
rect 14274 2320 14280 2372
rect 14332 2360 14338 2372
rect 14476 2360 14504 2391
rect 14332 2332 14504 2360
rect 14332 2320 14338 2332
rect 14734 2320 14740 2372
rect 14792 2360 14798 2372
rect 15028 2360 15056 2391
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 14792 2332 15056 2360
rect 15289 2363 15347 2369
rect 14792 2320 14798 2332
rect 15289 2329 15301 2363
rect 15335 2360 15347 2363
rect 15930 2360 15936 2372
rect 15335 2332 15936 2360
rect 15335 2329 15347 2332
rect 15289 2323 15347 2329
rect 15930 2320 15936 2332
rect 15988 2320 15994 2372
rect 11808 2264 12756 2292
rect 12802 2252 12808 2304
rect 12860 2292 12866 2304
rect 16482 2292 16488 2304
rect 12860 2264 16488 2292
rect 12860 2252 12866 2264
rect 16482 2252 16488 2264
rect 16540 2252 16546 2304
rect 1104 2202 16008 2224
rect 1104 2150 4698 2202
rect 4750 2150 4762 2202
rect 4814 2150 4826 2202
rect 4878 2150 4890 2202
rect 4942 2150 4954 2202
rect 5006 2150 8446 2202
rect 8498 2150 8510 2202
rect 8562 2150 8574 2202
rect 8626 2150 8638 2202
rect 8690 2150 8702 2202
rect 8754 2150 12194 2202
rect 12246 2150 12258 2202
rect 12310 2150 12322 2202
rect 12374 2150 12386 2202
rect 12438 2150 12450 2202
rect 12502 2150 16008 2202
rect 1104 2128 16008 2150
rect 3050 2048 3056 2100
rect 3108 2088 3114 2100
rect 10962 2088 10968 2100
rect 3108 2060 10968 2088
rect 3108 2048 3114 2060
rect 10962 2048 10968 2060
rect 11020 2048 11026 2100
rect 11146 2048 11152 2100
rect 11204 2088 11210 2100
rect 12066 2088 12072 2100
rect 11204 2060 12072 2088
rect 11204 2048 11210 2060
rect 12066 2048 12072 2060
rect 12124 2048 12130 2100
rect 12618 2048 12624 2100
rect 12676 2088 12682 2100
rect 15010 2088 15016 2100
rect 12676 2060 15016 2088
rect 12676 2048 12682 2060
rect 15010 2048 15016 2060
rect 15068 2048 15074 2100
rect 3142 1980 3148 2032
rect 3200 2020 3206 2032
rect 6822 2020 6828 2032
rect 3200 1992 6828 2020
rect 3200 1980 3206 1992
rect 6822 1980 6828 1992
rect 6880 1980 6886 2032
rect 7033 1992 8248 2020
rect 4430 1912 4436 1964
rect 4488 1952 4494 1964
rect 7033 1952 7061 1992
rect 4488 1924 7061 1952
rect 4488 1912 4494 1924
rect 7098 1912 7104 1964
rect 7156 1952 7162 1964
rect 7156 1924 8156 1952
rect 7156 1912 7162 1924
rect 4062 1776 4068 1828
rect 4120 1816 4126 1828
rect 6914 1816 6920 1828
rect 4120 1788 6920 1816
rect 4120 1776 4126 1788
rect 6914 1776 6920 1788
rect 6972 1776 6978 1828
rect 8128 1816 8156 1924
rect 8220 1884 8248 1992
rect 8846 1980 8852 2032
rect 8904 2020 8910 2032
rect 11606 2020 11612 2032
rect 8904 1992 11612 2020
rect 8904 1980 8910 1992
rect 11606 1980 11612 1992
rect 11664 1980 11670 2032
rect 8294 1912 8300 1964
rect 8352 1952 8358 1964
rect 11422 1952 11428 1964
rect 8352 1924 11428 1952
rect 8352 1912 8358 1924
rect 11422 1912 11428 1924
rect 11480 1912 11486 1964
rect 11514 1912 11520 1964
rect 11572 1952 11578 1964
rect 13262 1952 13268 1964
rect 11572 1924 13268 1952
rect 11572 1912 11578 1924
rect 13262 1912 13268 1924
rect 13320 1912 13326 1964
rect 9674 1884 9680 1896
rect 8220 1856 9680 1884
rect 9674 1844 9680 1856
rect 9732 1844 9738 1896
rect 9766 1844 9772 1896
rect 9824 1884 9830 1896
rect 10042 1884 10048 1896
rect 9824 1856 10048 1884
rect 9824 1844 9830 1856
rect 10042 1844 10048 1856
rect 10100 1884 10106 1896
rect 14918 1884 14924 1896
rect 10100 1856 14924 1884
rect 10100 1844 10106 1856
rect 14918 1844 14924 1856
rect 14976 1844 14982 1896
rect 11698 1816 11704 1828
rect 8128 1788 11704 1816
rect 11698 1776 11704 1788
rect 11756 1776 11762 1828
rect 6362 1708 6368 1760
rect 6420 1748 6426 1760
rect 7650 1748 7656 1760
rect 6420 1720 7656 1748
rect 6420 1708 6426 1720
rect 7650 1708 7656 1720
rect 7708 1708 7714 1760
rect 7742 1708 7748 1760
rect 7800 1748 7806 1760
rect 11054 1748 11060 1760
rect 7800 1720 11060 1748
rect 7800 1708 7806 1720
rect 11054 1708 11060 1720
rect 11112 1708 11118 1760
rect 2222 1640 2228 1692
rect 2280 1680 2286 1692
rect 2280 1652 2774 1680
rect 2280 1640 2286 1652
rect 2746 1612 2774 1652
rect 7558 1640 7564 1692
rect 7616 1680 7622 1692
rect 11422 1680 11428 1692
rect 7616 1652 11428 1680
rect 7616 1640 7622 1652
rect 11422 1640 11428 1652
rect 11480 1640 11486 1692
rect 10502 1612 10508 1624
rect 2746 1584 10508 1612
rect 10502 1572 10508 1584
rect 10560 1572 10566 1624
rect 10686 1572 10692 1624
rect 10744 1612 10750 1624
rect 13722 1612 13728 1624
rect 10744 1584 13728 1612
rect 10744 1572 10750 1584
rect 13722 1572 13728 1584
rect 13780 1572 13786 1624
rect 4522 1504 4528 1556
rect 4580 1544 4586 1556
rect 8938 1544 8944 1556
rect 4580 1516 8944 1544
rect 4580 1504 4586 1516
rect 8938 1504 8944 1516
rect 8996 1504 9002 1556
rect 9030 1504 9036 1556
rect 9088 1544 9094 1556
rect 9674 1544 9680 1556
rect 9088 1516 9680 1544
rect 9088 1504 9094 1516
rect 9674 1504 9680 1516
rect 9732 1504 9738 1556
rect 10134 1504 10140 1556
rect 10192 1544 10198 1556
rect 16298 1544 16304 1556
rect 10192 1516 16304 1544
rect 10192 1504 10198 1516
rect 16298 1504 16304 1516
rect 16356 1504 16362 1556
rect 5350 1436 5356 1488
rect 5408 1476 5414 1488
rect 10594 1476 10600 1488
rect 5408 1448 10600 1476
rect 5408 1436 5414 1448
rect 10594 1436 10600 1448
rect 10652 1436 10658 1488
rect 10778 1436 10784 1488
rect 10836 1476 10842 1488
rect 13446 1476 13452 1488
rect 10836 1448 13452 1476
rect 10836 1436 10842 1448
rect 13446 1436 13452 1448
rect 13504 1436 13510 1488
rect 2774 1368 2780 1420
rect 2832 1408 2838 1420
rect 3418 1408 3424 1420
rect 2832 1380 3424 1408
rect 2832 1368 2838 1380
rect 3418 1368 3424 1380
rect 3476 1368 3482 1420
rect 3602 1368 3608 1420
rect 3660 1408 3666 1420
rect 8018 1408 8024 1420
rect 3660 1380 8024 1408
rect 3660 1368 3666 1380
rect 8018 1368 8024 1380
rect 8076 1368 8082 1420
rect 8110 1368 8116 1420
rect 8168 1408 8174 1420
rect 8662 1408 8668 1420
rect 8168 1380 8668 1408
rect 8168 1368 8174 1380
rect 8662 1368 8668 1380
rect 8720 1368 8726 1420
rect 6822 1300 6828 1352
rect 6880 1340 6886 1352
rect 11790 1340 11796 1352
rect 6880 1312 11796 1340
rect 6880 1300 6886 1312
rect 11790 1300 11796 1312
rect 11848 1300 11854 1352
rect 3510 1232 3516 1284
rect 3568 1272 3574 1284
rect 14642 1272 14648 1284
rect 3568 1244 14648 1272
rect 3568 1232 3574 1244
rect 14642 1232 14648 1244
rect 14700 1232 14706 1284
rect 6178 1164 6184 1216
rect 6236 1204 6242 1216
rect 11238 1204 11244 1216
rect 6236 1176 11244 1204
rect 6236 1164 6242 1176
rect 11238 1164 11244 1176
rect 11296 1164 11302 1216
rect 14458 1204 14464 1216
rect 11348 1176 14464 1204
rect 3970 1096 3976 1148
rect 4028 1136 4034 1148
rect 11348 1136 11376 1176
rect 14458 1164 14464 1176
rect 14516 1164 14522 1216
rect 4028 1108 11376 1136
rect 4028 1096 4034 1108
rect 11514 1096 11520 1148
rect 11572 1136 11578 1148
rect 13078 1136 13084 1148
rect 11572 1108 13084 1136
rect 11572 1096 11578 1108
rect 13078 1096 13084 1108
rect 13136 1096 13142 1148
rect 5902 1028 5908 1080
rect 5960 1068 5966 1080
rect 6822 1068 6828 1080
rect 5960 1040 6828 1068
rect 5960 1028 5966 1040
rect 6822 1028 6828 1040
rect 6880 1028 6886 1080
rect 7374 1028 7380 1080
rect 7432 1068 7438 1080
rect 10686 1068 10692 1080
rect 7432 1040 10692 1068
rect 7432 1028 7438 1040
rect 10686 1028 10692 1040
rect 10744 1028 10750 1080
rect 106 960 112 1012
rect 164 1000 170 1012
rect 15102 1000 15108 1012
rect 164 972 15108 1000
rect 164 960 170 972
rect 15102 960 15108 972
rect 15160 960 15166 1012
rect 6086 892 6092 944
rect 6144 932 6150 944
rect 10226 932 10232 944
rect 6144 904 10232 932
rect 6144 892 6150 904
rect 10226 892 10232 904
rect 10284 892 10290 944
rect 3602 824 3608 876
rect 3660 864 3666 876
rect 12986 864 12992 876
rect 3660 836 12992 864
rect 3660 824 3666 836
rect 12986 824 12992 836
rect 13044 824 13050 876
rect 5626 756 5632 808
rect 5684 796 5690 808
rect 10870 796 10876 808
rect 5684 768 10876 796
rect 5684 756 5690 768
rect 10870 756 10876 768
rect 10928 756 10934 808
rect 3694 688 3700 740
rect 3752 728 3758 740
rect 11514 728 11520 740
rect 3752 700 11520 728
rect 3752 688 3758 700
rect 11514 688 11520 700
rect 11572 688 11578 740
rect 6822 212 6828 264
rect 6880 252 6886 264
rect 9766 252 9772 264
rect 6880 224 9772 252
rect 6880 212 6886 224
rect 9766 212 9772 224
rect 9824 212 9830 264
rect 4430 144 4436 196
rect 4488 184 4494 196
rect 15378 184 15384 196
rect 4488 156 15384 184
rect 4488 144 4494 156
rect 15378 144 15384 156
rect 15436 144 15442 196
rect 1854 76 1860 128
rect 1912 116 1918 128
rect 14366 116 14372 128
rect 1912 88 14372 116
rect 1912 76 1918 88
rect 14366 76 14372 88
rect 14424 76 14430 128
rect 842 8 848 60
rect 900 48 906 60
rect 13630 48 13636 60
rect 900 20 13636 48
rect 900 8 906 20
rect 13630 8 13636 20
rect 13688 8 13694 60
<< via1 >>
rect 4068 17960 4120 18012
rect 6368 17960 6420 18012
rect 13912 17824 13964 17876
rect 15476 17824 15528 17876
rect 4698 17382 4750 17434
rect 4762 17382 4814 17434
rect 4826 17382 4878 17434
rect 4890 17382 4942 17434
rect 4954 17382 5006 17434
rect 8446 17382 8498 17434
rect 8510 17382 8562 17434
rect 8574 17382 8626 17434
rect 8638 17382 8690 17434
rect 8702 17382 8754 17434
rect 12194 17382 12246 17434
rect 12258 17382 12310 17434
rect 12322 17382 12374 17434
rect 12386 17382 12438 17434
rect 12450 17382 12502 17434
rect 940 17212 992 17264
rect 3148 17144 3200 17196
rect 1952 16940 2004 16992
rect 13084 17008 13136 17060
rect 14004 17008 14056 17060
rect 2824 16838 2876 16890
rect 2888 16838 2940 16890
rect 2952 16838 3004 16890
rect 3016 16838 3068 16890
rect 3080 16838 3132 16890
rect 6572 16838 6624 16890
rect 6636 16838 6688 16890
rect 6700 16838 6752 16890
rect 6764 16838 6816 16890
rect 6828 16838 6880 16890
rect 10320 16838 10372 16890
rect 10384 16838 10436 16890
rect 10448 16838 10500 16890
rect 10512 16838 10564 16890
rect 10576 16838 10628 16890
rect 14068 16838 14120 16890
rect 14132 16838 14184 16890
rect 14196 16838 14248 16890
rect 14260 16838 14312 16890
rect 14324 16838 14376 16890
rect 1584 16736 1636 16788
rect 9772 16736 9824 16788
rect 1768 16668 1820 16720
rect 6184 16532 6236 16584
rect 8208 16532 8260 16584
rect 10048 16532 10100 16584
rect 2320 16396 2372 16448
rect 7748 16396 7800 16448
rect 4698 16294 4750 16346
rect 4762 16294 4814 16346
rect 4826 16294 4878 16346
rect 4890 16294 4942 16346
rect 4954 16294 5006 16346
rect 8446 16294 8498 16346
rect 8510 16294 8562 16346
rect 8574 16294 8626 16346
rect 8638 16294 8690 16346
rect 8702 16294 8754 16346
rect 12194 16294 12246 16346
rect 12258 16294 12310 16346
rect 12322 16294 12374 16346
rect 12386 16294 12438 16346
rect 12450 16294 12502 16346
rect 5356 16235 5408 16244
rect 5356 16201 5365 16235
rect 5365 16201 5399 16235
rect 5399 16201 5408 16235
rect 5356 16192 5408 16201
rect 2044 16124 2096 16176
rect 7840 16056 7892 16108
rect 12900 16056 12952 16108
rect 2504 15988 2556 16040
rect 5540 15988 5592 16040
rect 5816 15988 5868 16040
rect 9404 15988 9456 16040
rect 5632 15920 5684 15972
rect 10232 15920 10284 15972
rect 13820 15920 13872 15972
rect 1032 15852 1084 15904
rect 1676 15852 1728 15904
rect 3700 15895 3752 15904
rect 3700 15861 3709 15895
rect 3709 15861 3743 15895
rect 3743 15861 3752 15895
rect 3700 15852 3752 15861
rect 9404 15852 9456 15904
rect 15108 15852 15160 15904
rect 15752 15852 15804 15904
rect 2824 15750 2876 15802
rect 2888 15750 2940 15802
rect 2952 15750 3004 15802
rect 3016 15750 3068 15802
rect 3080 15750 3132 15802
rect 6572 15750 6624 15802
rect 6636 15750 6688 15802
rect 6700 15750 6752 15802
rect 6764 15750 6816 15802
rect 6828 15750 6880 15802
rect 10320 15750 10372 15802
rect 10384 15750 10436 15802
rect 10448 15750 10500 15802
rect 10512 15750 10564 15802
rect 10576 15750 10628 15802
rect 14068 15750 14120 15802
rect 14132 15750 14184 15802
rect 14196 15750 14248 15802
rect 14260 15750 14312 15802
rect 14324 15750 14376 15802
rect 3240 15648 3292 15700
rect 3516 15648 3568 15700
rect 5356 15648 5408 15700
rect 7012 15691 7064 15700
rect 7012 15657 7021 15691
rect 7021 15657 7055 15691
rect 7055 15657 7064 15691
rect 7012 15648 7064 15657
rect 7748 15648 7800 15700
rect 2412 15580 2464 15632
rect 3608 15580 3660 15632
rect 3056 15512 3108 15564
rect 9956 15648 10008 15700
rect 10876 15648 10928 15700
rect 9220 15580 9272 15632
rect 11796 15580 11848 15632
rect 14556 15580 14608 15632
rect 3976 15555 4028 15564
rect 3976 15521 3985 15555
rect 3985 15521 4019 15555
rect 4019 15521 4028 15555
rect 3976 15512 4028 15521
rect 5356 15512 5408 15564
rect 5540 15512 5592 15564
rect 4344 15444 4396 15496
rect 6000 15444 6052 15496
rect 6276 15444 6328 15496
rect 8024 15444 8076 15496
rect 9036 15444 9088 15496
rect 9680 15512 9732 15564
rect 15568 15512 15620 15564
rect 10692 15444 10744 15496
rect 3700 15376 3752 15428
rect 4436 15376 4488 15428
rect 4528 15376 4580 15428
rect 10140 15376 10192 15428
rect 3240 15308 3292 15360
rect 4344 15308 4396 15360
rect 5540 15351 5592 15360
rect 5540 15317 5549 15351
rect 5549 15317 5583 15351
rect 5583 15317 5592 15351
rect 5540 15308 5592 15317
rect 6184 15308 6236 15360
rect 7748 15351 7800 15360
rect 7748 15317 7757 15351
rect 7757 15317 7791 15351
rect 7791 15317 7800 15351
rect 7748 15308 7800 15317
rect 8116 15308 8168 15360
rect 9772 15308 9824 15360
rect 15200 15308 15252 15360
rect 4698 15206 4750 15258
rect 4762 15206 4814 15258
rect 4826 15206 4878 15258
rect 4890 15206 4942 15258
rect 4954 15206 5006 15258
rect 8446 15206 8498 15258
rect 8510 15206 8562 15258
rect 8574 15206 8626 15258
rect 8638 15206 8690 15258
rect 8702 15206 8754 15258
rect 12194 15206 12246 15258
rect 12258 15206 12310 15258
rect 12322 15206 12374 15258
rect 12386 15206 12438 15258
rect 12450 15206 12502 15258
rect 3056 15147 3108 15156
rect 3056 15113 3065 15147
rect 3065 15113 3099 15147
rect 3099 15113 3108 15147
rect 3056 15104 3108 15113
rect 3240 15147 3292 15156
rect 3240 15113 3249 15147
rect 3249 15113 3283 15147
rect 3283 15113 3292 15147
rect 3240 15104 3292 15113
rect 3608 15147 3660 15156
rect 3608 15113 3617 15147
rect 3617 15113 3651 15147
rect 3651 15113 3660 15147
rect 3608 15104 3660 15113
rect 756 15036 808 15088
rect 3332 15036 3384 15088
rect 3700 14968 3752 15020
rect 3792 15011 3844 15020
rect 3792 14977 3801 15011
rect 3801 14977 3835 15011
rect 3835 14977 3844 15011
rect 4344 15036 4396 15088
rect 4528 15104 4580 15156
rect 5356 15104 5408 15156
rect 5724 15104 5776 15156
rect 6368 15147 6420 15156
rect 6368 15113 6377 15147
rect 6377 15113 6411 15147
rect 6411 15113 6420 15147
rect 6368 15104 6420 15113
rect 7288 15104 7340 15156
rect 6092 15036 6144 15088
rect 3792 14968 3844 14977
rect 5172 15011 5224 15020
rect 5172 14977 5181 15011
rect 5181 14977 5215 15011
rect 5215 14977 5224 15011
rect 5172 14968 5224 14977
rect 5448 15011 5500 15020
rect 5448 14977 5457 15011
rect 5457 14977 5491 15011
rect 5491 14977 5500 15011
rect 5448 14968 5500 14977
rect 6184 15011 6236 15020
rect 6184 14977 6193 15011
rect 6193 14977 6227 15011
rect 6227 14977 6236 15011
rect 6184 14968 6236 14977
rect 7564 14968 7616 15020
rect 7748 14968 7800 15020
rect 4436 14900 4488 14952
rect 3056 14832 3108 14884
rect 3240 14832 3292 14884
rect 3976 14832 4028 14884
rect 5356 14900 5408 14952
rect 5540 14900 5592 14952
rect 7012 14943 7064 14952
rect 7012 14909 7021 14943
rect 7021 14909 7055 14943
rect 7055 14909 7064 14943
rect 7012 14900 7064 14909
rect 7104 14943 7156 14952
rect 7104 14909 7113 14943
rect 7113 14909 7147 14943
rect 7147 14909 7156 14943
rect 7104 14900 7156 14909
rect 6092 14832 6144 14884
rect 7196 14832 7248 14884
rect 8484 14900 8536 14952
rect 12808 14900 12860 14952
rect 1124 14764 1176 14816
rect 2688 14764 2740 14816
rect 5356 14764 5408 14816
rect 7380 14764 7432 14816
rect 8484 14807 8536 14816
rect 8484 14773 8493 14807
rect 8493 14773 8527 14807
rect 8527 14773 8536 14807
rect 8484 14764 8536 14773
rect 8668 14807 8720 14816
rect 8668 14773 8677 14807
rect 8677 14773 8711 14807
rect 8711 14773 8720 14807
rect 8668 14764 8720 14773
rect 8852 14807 8904 14816
rect 8852 14773 8861 14807
rect 8861 14773 8895 14807
rect 8895 14773 8904 14807
rect 8852 14764 8904 14773
rect 9680 14764 9732 14816
rect 12072 14764 12124 14816
rect 2824 14662 2876 14714
rect 2888 14662 2940 14714
rect 2952 14662 3004 14714
rect 3016 14662 3068 14714
rect 3080 14662 3132 14714
rect 6572 14662 6624 14714
rect 6636 14662 6688 14714
rect 6700 14662 6752 14714
rect 6764 14662 6816 14714
rect 6828 14662 6880 14714
rect 10320 14662 10372 14714
rect 10384 14662 10436 14714
rect 10448 14662 10500 14714
rect 10512 14662 10564 14714
rect 10576 14662 10628 14714
rect 14068 14662 14120 14714
rect 14132 14662 14184 14714
rect 14196 14662 14248 14714
rect 14260 14662 14312 14714
rect 14324 14662 14376 14714
rect 1216 14560 1268 14612
rect 4528 14560 4580 14612
rect 4620 14560 4672 14612
rect 848 14492 900 14544
rect 2504 14492 2556 14544
rect 3332 14535 3384 14544
rect 3332 14501 3341 14535
rect 3341 14501 3375 14535
rect 3375 14501 3384 14535
rect 3332 14492 3384 14501
rect 3608 14535 3660 14544
rect 3608 14501 3617 14535
rect 3617 14501 3651 14535
rect 3651 14501 3660 14535
rect 3608 14492 3660 14501
rect 4160 14492 4212 14544
rect 1952 14467 2004 14476
rect 1952 14433 1961 14467
rect 1961 14433 1995 14467
rect 1995 14433 2004 14467
rect 1952 14424 2004 14433
rect 2228 14467 2280 14476
rect 2228 14433 2237 14467
rect 2237 14433 2271 14467
rect 2271 14433 2280 14467
rect 2228 14424 2280 14433
rect 3608 14356 3660 14408
rect 3792 14399 3844 14408
rect 3792 14365 3801 14399
rect 3801 14365 3835 14399
rect 3835 14365 3844 14399
rect 3792 14356 3844 14365
rect 4068 14424 4120 14476
rect 7656 14560 7708 14612
rect 8208 14560 8260 14612
rect 8852 14560 8904 14612
rect 14648 14560 14700 14612
rect 5448 14492 5500 14544
rect 5724 14492 5776 14544
rect 7840 14492 7892 14544
rect 9220 14492 9272 14544
rect 9404 14535 9456 14544
rect 9404 14501 9413 14535
rect 9413 14501 9447 14535
rect 9447 14501 9456 14535
rect 9404 14492 9456 14501
rect 12624 14492 12676 14544
rect 6092 14467 6144 14476
rect 6092 14433 6101 14467
rect 6101 14433 6135 14467
rect 6135 14433 6144 14467
rect 6092 14424 6144 14433
rect 4344 14356 4396 14408
rect 2044 14288 2096 14340
rect 2688 14288 2740 14340
rect 3332 14288 3384 14340
rect 3516 14288 3568 14340
rect 3700 14288 3752 14340
rect 4252 14288 4304 14340
rect 4620 14356 4672 14408
rect 5172 14356 5224 14408
rect 5540 14356 5592 14408
rect 5908 14399 5960 14408
rect 5908 14365 5917 14399
rect 5917 14365 5951 14399
rect 5951 14365 5960 14399
rect 5908 14356 5960 14365
rect 940 14220 992 14272
rect 4160 14220 4212 14272
rect 5632 14288 5684 14340
rect 7472 14424 7524 14476
rect 8208 14424 8260 14476
rect 6828 14399 6880 14408
rect 6828 14365 6837 14399
rect 6837 14365 6871 14399
rect 6871 14365 6880 14399
rect 6828 14356 6880 14365
rect 7380 14356 7432 14408
rect 7932 14356 7984 14408
rect 8484 14356 8536 14408
rect 7288 14288 7340 14340
rect 7564 14331 7616 14340
rect 7564 14297 7573 14331
rect 7573 14297 7607 14331
rect 7607 14297 7616 14331
rect 7564 14288 7616 14297
rect 11704 14424 11756 14476
rect 9588 14399 9640 14408
rect 9588 14365 9597 14399
rect 9597 14365 9631 14399
rect 9631 14365 9640 14399
rect 9588 14356 9640 14365
rect 11796 14356 11848 14408
rect 12992 14356 13044 14408
rect 5172 14220 5224 14272
rect 5540 14263 5592 14272
rect 5540 14229 5549 14263
rect 5549 14229 5583 14263
rect 5583 14229 5592 14263
rect 5540 14220 5592 14229
rect 6000 14263 6052 14272
rect 6000 14229 6009 14263
rect 6009 14229 6043 14263
rect 6043 14229 6052 14263
rect 6000 14220 6052 14229
rect 6184 14220 6236 14272
rect 9312 14220 9364 14272
rect 9404 14220 9456 14272
rect 13636 14288 13688 14340
rect 4698 14118 4750 14170
rect 4762 14118 4814 14170
rect 4826 14118 4878 14170
rect 4890 14118 4942 14170
rect 4954 14118 5006 14170
rect 8446 14118 8498 14170
rect 8510 14118 8562 14170
rect 8574 14118 8626 14170
rect 8638 14118 8690 14170
rect 8702 14118 8754 14170
rect 12194 14118 12246 14170
rect 12258 14118 12310 14170
rect 12322 14118 12374 14170
rect 12386 14118 12438 14170
rect 12450 14118 12502 14170
rect 1492 14059 1544 14068
rect 1492 14025 1501 14059
rect 1501 14025 1535 14059
rect 1535 14025 1544 14059
rect 1492 14016 1544 14025
rect 1952 14016 2004 14068
rect 3884 14016 3936 14068
rect 2136 13948 2188 14000
rect 3424 13948 3476 14000
rect 3516 13948 3568 14000
rect 4160 13991 4212 14000
rect 4160 13957 4169 13991
rect 4169 13957 4203 13991
rect 4203 13957 4212 13991
rect 4160 13948 4212 13957
rect 5540 13948 5592 14000
rect 2044 13880 2096 13932
rect 2412 13923 2464 13932
rect 1400 13812 1452 13864
rect 1860 13744 1912 13796
rect 2412 13889 2421 13923
rect 2421 13889 2455 13923
rect 2455 13889 2464 13923
rect 2412 13880 2464 13889
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 3240 13923 3292 13932
rect 3240 13889 3249 13923
rect 3249 13889 3283 13923
rect 3283 13889 3292 13923
rect 3240 13880 3292 13889
rect 3332 13812 3384 13864
rect 3516 13812 3568 13864
rect 4344 13855 4396 13864
rect 4344 13821 4353 13855
rect 4353 13821 4387 13855
rect 4387 13821 4396 13855
rect 4344 13812 4396 13821
rect 5172 13880 5224 13932
rect 5448 13880 5500 13932
rect 6368 13948 6420 14000
rect 6736 13948 6788 14000
rect 8208 13948 8260 14000
rect 5540 13812 5592 13864
rect 5908 13880 5960 13932
rect 7104 13880 7156 13932
rect 7564 13880 7616 13932
rect 8668 13880 8720 13932
rect 6092 13855 6144 13864
rect 6092 13821 6101 13855
rect 6101 13821 6135 13855
rect 6135 13821 6144 13855
rect 6092 13812 6144 13821
rect 7012 13812 7064 13864
rect 9128 14016 9180 14068
rect 8944 13948 8996 14000
rect 9404 14016 9456 14068
rect 10232 13948 10284 14000
rect 9588 13923 9640 13932
rect 9588 13889 9597 13923
rect 9597 13889 9631 13923
rect 9631 13889 9640 13923
rect 9588 13880 9640 13889
rect 2688 13744 2740 13796
rect 4436 13744 4488 13796
rect 5172 13744 5224 13796
rect 6644 13744 6696 13796
rect 7196 13744 7248 13796
rect 9128 13744 9180 13796
rect 9772 13812 9824 13864
rect 10048 13812 10100 13864
rect 15476 13812 15528 13864
rect 9588 13744 9640 13796
rect 10140 13744 10192 13796
rect 11152 13744 11204 13796
rect 4528 13676 4580 13728
rect 4896 13676 4948 13728
rect 6368 13676 6420 13728
rect 8944 13676 8996 13728
rect 13268 13676 13320 13728
rect 2824 13574 2876 13626
rect 2888 13574 2940 13626
rect 2952 13574 3004 13626
rect 3016 13574 3068 13626
rect 3080 13574 3132 13626
rect 6572 13574 6624 13626
rect 6636 13574 6688 13626
rect 6700 13574 6752 13626
rect 6764 13574 6816 13626
rect 6828 13574 6880 13626
rect 10320 13574 10372 13626
rect 10384 13574 10436 13626
rect 10448 13574 10500 13626
rect 10512 13574 10564 13626
rect 10576 13574 10628 13626
rect 14068 13574 14120 13626
rect 14132 13574 14184 13626
rect 14196 13574 14248 13626
rect 14260 13574 14312 13626
rect 14324 13574 14376 13626
rect 2688 13515 2740 13524
rect 2688 13481 2697 13515
rect 2697 13481 2731 13515
rect 2731 13481 2740 13515
rect 2688 13472 2740 13481
rect 3608 13472 3660 13524
rect 4436 13472 4488 13524
rect 6000 13472 6052 13524
rect 7104 13472 7156 13524
rect 8300 13472 8352 13524
rect 9036 13515 9088 13524
rect 9036 13481 9045 13515
rect 9045 13481 9079 13515
rect 9079 13481 9088 13515
rect 9496 13515 9548 13524
rect 9036 13472 9088 13481
rect 9496 13481 9505 13515
rect 9505 13481 9539 13515
rect 9539 13481 9548 13515
rect 9496 13472 9548 13481
rect 9588 13472 9640 13524
rect 10048 13472 10100 13524
rect 10140 13472 10192 13524
rect 10692 13515 10744 13524
rect 10692 13481 10701 13515
rect 10701 13481 10735 13515
rect 10735 13481 10744 13515
rect 10692 13472 10744 13481
rect 11520 13472 11572 13524
rect 1676 13379 1728 13388
rect 1676 13345 1685 13379
rect 1685 13345 1719 13379
rect 1719 13345 1728 13379
rect 1676 13336 1728 13345
rect 3424 13336 3476 13388
rect 3792 13336 3844 13388
rect 4436 13379 4488 13388
rect 4436 13345 4445 13379
rect 4445 13345 4479 13379
rect 4479 13345 4488 13379
rect 4436 13336 4488 13345
rect 4896 13336 4948 13388
rect 5264 13336 5316 13388
rect 3240 13268 3292 13320
rect 9220 13404 9272 13456
rect 9956 13404 10008 13456
rect 6552 13336 6604 13388
rect 7380 13336 7432 13388
rect 7564 13379 7616 13388
rect 7564 13345 7573 13379
rect 7573 13345 7607 13379
rect 7607 13345 7616 13379
rect 7564 13336 7616 13345
rect 5816 13268 5868 13320
rect 6920 13311 6972 13320
rect 6920 13277 6929 13311
rect 6929 13277 6963 13311
rect 6963 13277 6972 13311
rect 6920 13268 6972 13277
rect 7840 13336 7892 13388
rect 7932 13336 7984 13388
rect 8300 13336 8352 13388
rect 2228 13243 2280 13252
rect 2228 13209 2237 13243
rect 2237 13209 2271 13243
rect 2271 13209 2280 13243
rect 2228 13200 2280 13209
rect 2688 13132 2740 13184
rect 3332 13132 3384 13184
rect 4620 13132 4672 13184
rect 6736 13200 6788 13252
rect 7840 13200 7892 13252
rect 7932 13200 7984 13252
rect 5448 13132 5500 13184
rect 7104 13132 7156 13184
rect 7196 13132 7248 13184
rect 7748 13132 7800 13184
rect 11336 13336 11388 13388
rect 9404 13268 9456 13320
rect 10784 13268 10836 13320
rect 10876 13311 10928 13320
rect 10876 13277 10885 13311
rect 10885 13277 10919 13311
rect 10919 13277 10928 13311
rect 10876 13268 10928 13277
rect 11244 13200 11296 13252
rect 11612 13200 11664 13252
rect 14832 13200 14884 13252
rect 9588 13132 9640 13184
rect 10600 13132 10652 13184
rect 10692 13132 10744 13184
rect 13176 13132 13228 13184
rect 4698 13030 4750 13082
rect 4762 13030 4814 13082
rect 4826 13030 4878 13082
rect 4890 13030 4942 13082
rect 4954 13030 5006 13082
rect 8446 13030 8498 13082
rect 8510 13030 8562 13082
rect 8574 13030 8626 13082
rect 8638 13030 8690 13082
rect 8702 13030 8754 13082
rect 12194 13030 12246 13082
rect 12258 13030 12310 13082
rect 12322 13030 12374 13082
rect 12386 13030 12438 13082
rect 12450 13030 12502 13082
rect 1768 12928 1820 12980
rect 2136 12971 2188 12980
rect 2136 12937 2145 12971
rect 2145 12937 2179 12971
rect 2179 12937 2188 12971
rect 2136 12928 2188 12937
rect 2320 12971 2372 12980
rect 2320 12937 2329 12971
rect 2329 12937 2363 12971
rect 2363 12937 2372 12971
rect 2320 12928 2372 12937
rect 2964 12928 3016 12980
rect 3792 12928 3844 12980
rect 4620 12971 4672 12980
rect 4620 12937 4629 12971
rect 4629 12937 4663 12971
rect 4663 12937 4672 12971
rect 4620 12928 4672 12937
rect 6000 12928 6052 12980
rect 6460 12928 6512 12980
rect 6736 12928 6788 12980
rect 9220 12928 9272 12980
rect 9588 12928 9640 12980
rect 1768 12835 1820 12844
rect 1768 12801 1777 12835
rect 1777 12801 1811 12835
rect 1811 12801 1820 12835
rect 1768 12792 1820 12801
rect 7012 12860 7064 12912
rect 11612 12928 11664 12980
rect 11796 12928 11848 12980
rect 15844 12928 15896 12980
rect 4988 12835 5040 12844
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 5448 12792 5500 12844
rect 5264 12767 5316 12776
rect 5264 12733 5273 12767
rect 5273 12733 5307 12767
rect 5307 12733 5316 12767
rect 5264 12724 5316 12733
rect 5724 12724 5776 12776
rect 4252 12656 4304 12708
rect 5172 12656 5224 12708
rect 2504 12631 2556 12640
rect 2504 12597 2513 12631
rect 2513 12597 2547 12631
rect 2547 12597 2556 12631
rect 2504 12588 2556 12597
rect 5908 12792 5960 12844
rect 6368 12792 6420 12844
rect 8024 12835 8076 12844
rect 7472 12767 7524 12776
rect 7472 12733 7481 12767
rect 7481 12733 7515 12767
rect 7515 12733 7524 12767
rect 7472 12724 7524 12733
rect 7748 12767 7800 12776
rect 7748 12733 7757 12767
rect 7757 12733 7791 12767
rect 7791 12733 7800 12767
rect 7748 12724 7800 12733
rect 5908 12656 5960 12708
rect 7196 12656 7248 12708
rect 6276 12588 6328 12640
rect 8024 12801 8033 12835
rect 8033 12801 8067 12835
rect 8067 12801 8076 12835
rect 8024 12792 8076 12801
rect 8300 12792 8352 12844
rect 8208 12724 8260 12776
rect 8300 12656 8352 12708
rect 9496 12792 9548 12844
rect 9864 12860 9916 12912
rect 10232 12860 10284 12912
rect 10600 12903 10652 12912
rect 10600 12869 10609 12903
rect 10609 12869 10643 12903
rect 10643 12869 10652 12903
rect 10600 12860 10652 12869
rect 16212 12860 16264 12912
rect 11152 12792 11204 12844
rect 8760 12724 8812 12776
rect 9036 12767 9088 12776
rect 9036 12733 9045 12767
rect 9045 12733 9079 12767
rect 9079 12733 9088 12767
rect 9864 12767 9916 12776
rect 9036 12724 9088 12733
rect 9864 12733 9873 12767
rect 9873 12733 9907 12767
rect 9907 12733 9916 12767
rect 9864 12724 9916 12733
rect 9220 12656 9272 12708
rect 10692 12724 10744 12776
rect 10968 12724 11020 12776
rect 11520 12656 11572 12708
rect 11704 12656 11756 12708
rect 11796 12699 11848 12708
rect 11796 12665 11805 12699
rect 11805 12665 11839 12699
rect 11839 12665 11848 12699
rect 11796 12656 11848 12665
rect 12532 12656 12584 12708
rect 9588 12588 9640 12640
rect 9772 12588 9824 12640
rect 10692 12588 10744 12640
rect 12348 12588 12400 12640
rect 2824 12486 2876 12538
rect 2888 12486 2940 12538
rect 2952 12486 3004 12538
rect 3016 12486 3068 12538
rect 3080 12486 3132 12538
rect 6572 12486 6624 12538
rect 6636 12486 6688 12538
rect 6700 12486 6752 12538
rect 6764 12486 6816 12538
rect 6828 12486 6880 12538
rect 10320 12486 10372 12538
rect 10384 12486 10436 12538
rect 10448 12486 10500 12538
rect 10512 12486 10564 12538
rect 10576 12486 10628 12538
rect 14068 12486 14120 12538
rect 14132 12486 14184 12538
rect 14196 12486 14248 12538
rect 14260 12486 14312 12538
rect 14324 12486 14376 12538
rect 3240 12384 3292 12436
rect 5080 12384 5132 12436
rect 2780 12316 2832 12368
rect 5632 12316 5684 12368
rect 1584 12248 1636 12300
rect 2228 12291 2280 12300
rect 2228 12257 2237 12291
rect 2237 12257 2271 12291
rect 2271 12257 2280 12291
rect 2228 12248 2280 12257
rect 2688 12248 2740 12300
rect 3056 12248 3108 12300
rect 3424 12291 3476 12300
rect 3424 12257 3433 12291
rect 3433 12257 3467 12291
rect 3467 12257 3476 12291
rect 3424 12248 3476 12257
rect 3976 12248 4028 12300
rect 7196 12384 7248 12436
rect 8024 12384 8076 12436
rect 9404 12384 9456 12436
rect 9496 12384 9548 12436
rect 11796 12384 11848 12436
rect 11980 12427 12032 12436
rect 11980 12393 11989 12427
rect 11989 12393 12023 12427
rect 12023 12393 12032 12427
rect 11980 12384 12032 12393
rect 8944 12316 8996 12368
rect 10692 12316 10744 12368
rect 10876 12316 10928 12368
rect 3792 12223 3844 12232
rect 3792 12189 3801 12223
rect 3801 12189 3835 12223
rect 3835 12189 3844 12223
rect 3792 12180 3844 12189
rect 4528 12180 4580 12232
rect 5080 12180 5132 12232
rect 664 12044 716 12096
rect 1124 12044 1176 12096
rect 3148 12044 3200 12096
rect 3608 12044 3660 12096
rect 6276 12180 6328 12232
rect 5632 12112 5684 12164
rect 6552 12112 6604 12164
rect 6828 12180 6880 12232
rect 7564 12180 7616 12232
rect 9680 12248 9732 12300
rect 9864 12248 9916 12300
rect 8116 12180 8168 12232
rect 6736 12112 6788 12164
rect 9220 12180 9272 12232
rect 9404 12223 9456 12232
rect 9404 12189 9413 12223
rect 9413 12189 9447 12223
rect 9447 12189 9456 12223
rect 9404 12180 9456 12189
rect 10048 12180 10100 12232
rect 11152 12248 11204 12300
rect 11612 12316 11664 12368
rect 12440 12384 12492 12436
rect 12348 12316 12400 12368
rect 13544 12384 13596 12436
rect 13820 12384 13872 12436
rect 13452 12316 13504 12368
rect 16948 12316 17000 12368
rect 11980 12248 12032 12300
rect 12532 12291 12584 12300
rect 12532 12257 12541 12291
rect 12541 12257 12575 12291
rect 12575 12257 12584 12291
rect 12532 12248 12584 12257
rect 14096 12248 14148 12300
rect 14464 12291 14516 12300
rect 14464 12257 14473 12291
rect 14473 12257 14507 12291
rect 14507 12257 14516 12291
rect 14464 12248 14516 12257
rect 5724 12044 5776 12096
rect 6000 12044 6052 12096
rect 6920 12044 6972 12096
rect 8208 12044 8260 12096
rect 9864 12112 9916 12164
rect 10876 12112 10928 12164
rect 9220 12044 9272 12096
rect 9588 12044 9640 12096
rect 13268 12180 13320 12232
rect 11520 12112 11572 12164
rect 13360 12112 13412 12164
rect 11796 12044 11848 12096
rect 12624 12087 12676 12096
rect 12624 12053 12633 12087
rect 12633 12053 12667 12087
rect 12667 12053 12676 12087
rect 12624 12044 12676 12053
rect 13452 12087 13504 12096
rect 13452 12053 13461 12087
rect 13461 12053 13495 12087
rect 13495 12053 13504 12087
rect 13452 12044 13504 12053
rect 14004 12044 14056 12096
rect 14556 12112 14608 12164
rect 16488 12112 16540 12164
rect 14188 12044 14240 12096
rect 16672 12044 16724 12096
rect 4698 11942 4750 11994
rect 4762 11942 4814 11994
rect 4826 11942 4878 11994
rect 4890 11942 4942 11994
rect 4954 11942 5006 11994
rect 8446 11942 8498 11994
rect 8510 11942 8562 11994
rect 8574 11942 8626 11994
rect 8638 11942 8690 11994
rect 8702 11942 8754 11994
rect 12194 11942 12246 11994
rect 12258 11942 12310 11994
rect 12322 11942 12374 11994
rect 12386 11942 12438 11994
rect 12450 11942 12502 11994
rect 1124 11840 1176 11892
rect 1308 11840 1360 11892
rect 1584 11840 1636 11892
rect 2412 11840 2464 11892
rect 2688 11883 2740 11892
rect 2688 11849 2697 11883
rect 2697 11849 2731 11883
rect 2731 11849 2740 11883
rect 2688 11840 2740 11849
rect 3056 11883 3108 11892
rect 3056 11849 3065 11883
rect 3065 11849 3099 11883
rect 3099 11849 3108 11883
rect 3056 11840 3108 11849
rect 3884 11883 3936 11892
rect 3884 11849 3893 11883
rect 3893 11849 3927 11883
rect 3927 11849 3936 11883
rect 3884 11840 3936 11849
rect 4344 11840 4396 11892
rect 5724 11840 5776 11892
rect 6276 11840 6328 11892
rect 2596 11772 2648 11824
rect 4068 11772 4120 11824
rect 1860 11747 1912 11756
rect 1860 11713 1869 11747
rect 1869 11713 1903 11747
rect 1903 11713 1912 11747
rect 1860 11704 1912 11713
rect 3976 11704 4028 11756
rect 4620 11704 4672 11756
rect 1584 11679 1636 11688
rect 1584 11645 1593 11679
rect 1593 11645 1627 11679
rect 1627 11645 1636 11679
rect 1584 11636 1636 11645
rect 2596 11679 2648 11688
rect 2596 11645 2605 11679
rect 2605 11645 2639 11679
rect 2639 11645 2648 11679
rect 2596 11636 2648 11645
rect 3608 11636 3660 11688
rect 4068 11636 4120 11688
rect 4528 11568 4580 11620
rect 6736 11772 6788 11824
rect 6368 11679 6420 11688
rect 4160 11500 4212 11552
rect 4712 11500 4764 11552
rect 6368 11645 6377 11679
rect 6377 11645 6411 11679
rect 6411 11645 6420 11679
rect 6368 11636 6420 11645
rect 8116 11772 8168 11824
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 10048 11840 10100 11892
rect 10416 11840 10468 11892
rect 11520 11883 11572 11892
rect 11520 11849 11529 11883
rect 11529 11849 11563 11883
rect 11563 11849 11572 11883
rect 11520 11840 11572 11849
rect 12900 11840 12952 11892
rect 13912 11840 13964 11892
rect 14556 11883 14608 11892
rect 14556 11849 14565 11883
rect 14565 11849 14599 11883
rect 14599 11849 14608 11883
rect 14556 11840 14608 11849
rect 14740 11840 14792 11892
rect 8668 11704 8720 11756
rect 8852 11704 8904 11756
rect 8300 11636 8352 11688
rect 6092 11568 6144 11620
rect 6276 11568 6328 11620
rect 5172 11500 5224 11552
rect 5448 11500 5500 11552
rect 7472 11500 7524 11552
rect 8208 11500 8260 11552
rect 9588 11704 9640 11756
rect 11796 11772 11848 11824
rect 11980 11772 12032 11824
rect 8944 11568 8996 11620
rect 9680 11636 9732 11688
rect 10600 11704 10652 11756
rect 11152 11747 11204 11756
rect 11152 11713 11161 11747
rect 11161 11713 11195 11747
rect 11195 11713 11204 11747
rect 11152 11704 11204 11713
rect 11244 11704 11296 11756
rect 9772 11568 9824 11620
rect 9864 11568 9916 11620
rect 10232 11636 10284 11688
rect 10416 11636 10468 11688
rect 12440 11772 12492 11824
rect 13084 11772 13136 11824
rect 16212 11772 16264 11824
rect 13360 11704 13412 11756
rect 16304 11704 16356 11756
rect 11520 11636 11572 11688
rect 11980 11636 12032 11688
rect 12348 11636 12400 11688
rect 12532 11636 12584 11688
rect 13912 11636 13964 11688
rect 15108 11636 15160 11688
rect 15384 11636 15436 11688
rect 15936 11636 15988 11688
rect 9404 11543 9456 11552
rect 9404 11509 9413 11543
rect 9413 11509 9447 11543
rect 9447 11509 9456 11543
rect 9404 11500 9456 11509
rect 10876 11500 10928 11552
rect 11244 11500 11296 11552
rect 14096 11568 14148 11620
rect 14280 11568 14332 11620
rect 16028 11568 16080 11620
rect 12256 11500 12308 11552
rect 13084 11543 13136 11552
rect 13084 11509 13093 11543
rect 13093 11509 13127 11543
rect 13127 11509 13136 11543
rect 13084 11500 13136 11509
rect 13360 11543 13412 11552
rect 13360 11509 13369 11543
rect 13369 11509 13403 11543
rect 13403 11509 13412 11543
rect 13360 11500 13412 11509
rect 15016 11500 15068 11552
rect 15384 11500 15436 11552
rect 15568 11543 15620 11552
rect 15568 11509 15577 11543
rect 15577 11509 15611 11543
rect 15611 11509 15620 11543
rect 15568 11500 15620 11509
rect 2824 11398 2876 11450
rect 2888 11398 2940 11450
rect 2952 11398 3004 11450
rect 3016 11398 3068 11450
rect 3080 11398 3132 11450
rect 6572 11398 6624 11450
rect 6636 11398 6688 11450
rect 6700 11398 6752 11450
rect 6764 11398 6816 11450
rect 6828 11398 6880 11450
rect 10320 11398 10372 11450
rect 10384 11398 10436 11450
rect 10448 11398 10500 11450
rect 10512 11398 10564 11450
rect 10576 11398 10628 11450
rect 14068 11398 14120 11450
rect 14132 11398 14184 11450
rect 14196 11398 14248 11450
rect 14260 11398 14312 11450
rect 14324 11398 14376 11450
rect 3516 11296 3568 11348
rect 4160 11296 4212 11348
rect 4344 11296 4396 11348
rect 4620 11339 4672 11348
rect 4620 11305 4629 11339
rect 4629 11305 4663 11339
rect 4663 11305 4672 11339
rect 4620 11296 4672 11305
rect 5448 11296 5500 11348
rect 1676 11203 1728 11212
rect 1676 11169 1685 11203
rect 1685 11169 1719 11203
rect 1719 11169 1728 11203
rect 1676 11160 1728 11169
rect 2228 11203 2280 11212
rect 2228 11169 2237 11203
rect 2237 11169 2271 11203
rect 2271 11169 2280 11203
rect 2228 11160 2280 11169
rect 1952 11135 2004 11144
rect 1952 11101 1961 11135
rect 1961 11101 1995 11135
rect 1995 11101 2004 11135
rect 1952 11092 2004 11101
rect 6092 11228 6144 11280
rect 7196 11296 7248 11348
rect 7288 11296 7340 11348
rect 9036 11296 9088 11348
rect 9312 11296 9364 11348
rect 10140 11296 10192 11348
rect 3332 11203 3384 11212
rect 3332 11169 3341 11203
rect 3341 11169 3375 11203
rect 3375 11169 3384 11203
rect 3332 11160 3384 11169
rect 3792 11160 3844 11212
rect 4068 11203 4120 11212
rect 4068 11169 4077 11203
rect 4077 11169 4111 11203
rect 4111 11169 4120 11203
rect 4068 11160 4120 11169
rect 5080 11160 5132 11212
rect 7932 11160 7984 11212
rect 8852 11160 8904 11212
rect 11980 11296 12032 11348
rect 12440 11339 12492 11348
rect 12440 11305 12449 11339
rect 12449 11305 12483 11339
rect 12483 11305 12492 11339
rect 12440 11296 12492 11305
rect 12716 11339 12768 11348
rect 12716 11305 12725 11339
rect 12725 11305 12759 11339
rect 12759 11305 12768 11339
rect 12716 11296 12768 11305
rect 12900 11339 12952 11348
rect 12900 11305 12909 11339
rect 12909 11305 12943 11339
rect 12943 11305 12952 11339
rect 12900 11296 12952 11305
rect 12992 11296 13044 11348
rect 13544 11296 13596 11348
rect 14556 11339 14608 11348
rect 14556 11305 14565 11339
rect 14565 11305 14599 11339
rect 14599 11305 14608 11339
rect 14556 11296 14608 11305
rect 2320 11067 2372 11076
rect 2320 11033 2329 11067
rect 2329 11033 2363 11067
rect 2363 11033 2372 11067
rect 2320 11024 2372 11033
rect 1584 10956 1636 11008
rect 6000 11092 6052 11144
rect 6368 11092 6420 11144
rect 7748 11092 7800 11144
rect 7840 11092 7892 11144
rect 8024 11092 8076 11144
rect 8392 11092 8444 11144
rect 9220 11092 9272 11144
rect 10324 11203 10376 11212
rect 10324 11169 10333 11203
rect 10333 11169 10367 11203
rect 10367 11169 10376 11203
rect 10324 11160 10376 11169
rect 4528 11024 4580 11076
rect 2596 10956 2648 11008
rect 4252 10999 4304 11008
rect 4252 10965 4261 10999
rect 4261 10965 4295 10999
rect 4295 10965 4304 10999
rect 4896 11024 4948 11076
rect 5448 11024 5500 11076
rect 5816 11067 5868 11076
rect 5816 11033 5834 11067
rect 5834 11033 5868 11067
rect 5816 11024 5868 11033
rect 7656 11024 7708 11076
rect 9036 11024 9088 11076
rect 9864 11092 9916 11144
rect 11520 11228 11572 11280
rect 10600 11092 10652 11144
rect 11612 11160 11664 11212
rect 12164 11228 12216 11280
rect 14372 11228 14424 11280
rect 15384 11296 15436 11348
rect 15568 11296 15620 11348
rect 15844 11296 15896 11348
rect 9956 11024 10008 11076
rect 10508 11024 10560 11076
rect 10968 11067 11020 11076
rect 10968 11033 10977 11067
rect 10977 11033 11011 11067
rect 11011 11033 11020 11067
rect 10968 11024 11020 11033
rect 11152 11024 11204 11076
rect 4252 10956 4304 10965
rect 6828 10956 6880 11008
rect 7472 10956 7524 11008
rect 7748 10956 7800 11008
rect 10140 10956 10192 11008
rect 10324 10956 10376 11008
rect 12348 11092 12400 11144
rect 11612 11024 11664 11076
rect 12256 11067 12308 11076
rect 12256 11033 12265 11067
rect 12265 11033 12299 11067
rect 12299 11033 12308 11067
rect 12256 11024 12308 11033
rect 12808 11092 12860 11144
rect 13452 11160 13504 11212
rect 14004 11160 14056 11212
rect 16580 11228 16632 11280
rect 13176 11092 13228 11144
rect 11428 10999 11480 11008
rect 11428 10965 11437 10999
rect 11437 10965 11471 10999
rect 11471 10965 11480 10999
rect 11428 10956 11480 10965
rect 11704 10956 11756 11008
rect 12900 10956 12952 11008
rect 13360 10956 13412 11008
rect 13636 10956 13688 11008
rect 13912 11092 13964 11144
rect 14648 11092 14700 11144
rect 14924 11092 14976 11144
rect 15384 11092 15436 11144
rect 14096 11024 14148 11076
rect 15568 11067 15620 11076
rect 15568 11033 15577 11067
rect 15577 11033 15611 11067
rect 15611 11033 15620 11067
rect 15568 11024 15620 11033
rect 15752 11024 15804 11076
rect 14188 10956 14240 11008
rect 14740 10999 14792 11008
rect 14740 10965 14749 10999
rect 14749 10965 14783 10999
rect 14783 10965 14792 10999
rect 14740 10956 14792 10965
rect 15108 10956 15160 11008
rect 4698 10854 4750 10906
rect 4762 10854 4814 10906
rect 4826 10854 4878 10906
rect 4890 10854 4942 10906
rect 4954 10854 5006 10906
rect 8446 10854 8498 10906
rect 8510 10854 8562 10906
rect 8574 10854 8626 10906
rect 8638 10854 8690 10906
rect 8702 10854 8754 10906
rect 12194 10854 12246 10906
rect 12258 10854 12310 10906
rect 12322 10854 12374 10906
rect 12386 10854 12438 10906
rect 12450 10854 12502 10906
rect 1584 10795 1636 10804
rect 1584 10761 1593 10795
rect 1593 10761 1627 10795
rect 1627 10761 1636 10795
rect 1584 10752 1636 10761
rect 2136 10752 2188 10804
rect 3332 10752 3384 10804
rect 2780 10727 2832 10736
rect 2780 10693 2789 10727
rect 2789 10693 2823 10727
rect 2823 10693 2832 10727
rect 2780 10684 2832 10693
rect 3056 10684 3108 10736
rect 5632 10752 5684 10804
rect 2504 10616 2556 10668
rect 2688 10591 2740 10600
rect 2688 10557 2697 10591
rect 2697 10557 2731 10591
rect 2731 10557 2740 10591
rect 2688 10548 2740 10557
rect 3056 10480 3108 10532
rect 5172 10684 5224 10736
rect 5264 10684 5316 10736
rect 6920 10752 6972 10804
rect 7012 10752 7064 10804
rect 9128 10752 9180 10804
rect 10048 10752 10100 10804
rect 10968 10795 11020 10804
rect 10968 10761 10977 10795
rect 10977 10761 11011 10795
rect 11011 10761 11020 10795
rect 11520 10795 11572 10804
rect 10968 10752 11020 10761
rect 11520 10761 11529 10795
rect 11529 10761 11563 10795
rect 11563 10761 11572 10795
rect 11520 10752 11572 10761
rect 11888 10752 11940 10804
rect 12992 10752 13044 10804
rect 13176 10752 13228 10804
rect 14004 10795 14056 10804
rect 3884 10616 3936 10668
rect 4804 10616 4856 10668
rect 6644 10659 6696 10668
rect 6644 10625 6678 10659
rect 6678 10625 6696 10659
rect 6644 10616 6696 10625
rect 8944 10684 8996 10736
rect 8116 10616 8168 10668
rect 10876 10616 10928 10668
rect 11152 10616 11204 10668
rect 13360 10684 13412 10736
rect 14004 10761 14013 10795
rect 14013 10761 14047 10795
rect 14047 10761 14056 10795
rect 14004 10752 14056 10761
rect 14096 10795 14148 10804
rect 14096 10761 14105 10795
rect 14105 10761 14139 10795
rect 14139 10761 14148 10795
rect 14096 10752 14148 10761
rect 14280 10795 14332 10804
rect 14280 10761 14289 10795
rect 14289 10761 14323 10795
rect 14323 10761 14332 10795
rect 14280 10752 14332 10761
rect 15108 10752 15160 10804
rect 16212 10752 16264 10804
rect 14372 10684 14424 10736
rect 12440 10616 12492 10668
rect 6368 10591 6420 10600
rect 6368 10557 6377 10591
rect 6377 10557 6411 10591
rect 6411 10557 6420 10591
rect 6368 10548 6420 10557
rect 3332 10480 3384 10532
rect 4344 10412 4396 10464
rect 4620 10412 4672 10464
rect 4804 10455 4856 10464
rect 4804 10421 4813 10455
rect 4813 10421 4847 10455
rect 4847 10421 4856 10455
rect 7840 10548 7892 10600
rect 7932 10548 7984 10600
rect 9312 10548 9364 10600
rect 10140 10591 10192 10600
rect 7656 10480 7708 10532
rect 10140 10557 10149 10591
rect 10149 10557 10183 10591
rect 10183 10557 10192 10591
rect 10140 10548 10192 10557
rect 4804 10412 4856 10421
rect 8392 10412 8444 10464
rect 9956 10480 10008 10532
rect 10324 10548 10376 10600
rect 11704 10548 11756 10600
rect 12348 10548 12400 10600
rect 13452 10616 13504 10668
rect 11888 10480 11940 10532
rect 14096 10548 14148 10600
rect 14556 10548 14608 10600
rect 13452 10480 13504 10532
rect 14188 10480 14240 10532
rect 16580 10480 16632 10532
rect 10140 10412 10192 10464
rect 10692 10412 10744 10464
rect 11520 10412 11572 10464
rect 11980 10412 12032 10464
rect 12716 10412 12768 10464
rect 13636 10412 13688 10464
rect 14740 10455 14792 10464
rect 14740 10421 14749 10455
rect 14749 10421 14783 10455
rect 14783 10421 14792 10455
rect 14740 10412 14792 10421
rect 2824 10310 2876 10362
rect 2888 10310 2940 10362
rect 2952 10310 3004 10362
rect 3016 10310 3068 10362
rect 3080 10310 3132 10362
rect 6572 10310 6624 10362
rect 6636 10310 6688 10362
rect 6700 10310 6752 10362
rect 6764 10310 6816 10362
rect 6828 10310 6880 10362
rect 10320 10310 10372 10362
rect 10384 10310 10436 10362
rect 10448 10310 10500 10362
rect 10512 10310 10564 10362
rect 10576 10310 10628 10362
rect 14068 10310 14120 10362
rect 14132 10310 14184 10362
rect 14196 10310 14248 10362
rect 14260 10310 14312 10362
rect 14324 10310 14376 10362
rect 6920 10208 6972 10260
rect 8116 10208 8168 10260
rect 2136 10183 2188 10192
rect 2136 10149 2145 10183
rect 2145 10149 2179 10183
rect 2179 10149 2188 10183
rect 2136 10140 2188 10149
rect 4160 10140 4212 10192
rect 5448 10140 5500 10192
rect 1584 9936 1636 9988
rect 1952 10072 2004 10124
rect 5172 10115 5224 10124
rect 5172 10081 5181 10115
rect 5181 10081 5215 10115
rect 5215 10081 5224 10115
rect 5172 10072 5224 10081
rect 7748 10072 7800 10124
rect 2228 10047 2280 10056
rect 2228 10013 2237 10047
rect 2237 10013 2271 10047
rect 2271 10013 2280 10047
rect 2228 10004 2280 10013
rect 3240 10004 3292 10056
rect 2596 9936 2648 9988
rect 2780 9936 2832 9988
rect 4344 10004 4396 10056
rect 4620 10004 4672 10056
rect 6736 10004 6788 10056
rect 7380 10004 7432 10056
rect 8852 10072 8904 10124
rect 10140 10208 10192 10260
rect 11244 10251 11296 10260
rect 11244 10217 11253 10251
rect 11253 10217 11287 10251
rect 11287 10217 11296 10251
rect 11244 10208 11296 10217
rect 10048 10140 10100 10192
rect 12716 10208 12768 10260
rect 11980 10140 12032 10192
rect 13820 10208 13872 10260
rect 15660 10251 15712 10260
rect 15660 10217 15669 10251
rect 15669 10217 15703 10251
rect 15703 10217 15712 10251
rect 15660 10208 15712 10217
rect 8944 10047 8996 10056
rect 3424 9936 3476 9988
rect 4528 9936 4580 9988
rect 5816 9936 5868 9988
rect 5908 9936 5960 9988
rect 1768 9911 1820 9920
rect 1768 9877 1777 9911
rect 1777 9877 1811 9911
rect 1811 9877 1820 9911
rect 1768 9868 1820 9877
rect 2044 9868 2096 9920
rect 3240 9868 3292 9920
rect 3884 9868 3936 9920
rect 4068 9868 4120 9920
rect 4620 9868 4672 9920
rect 6368 9868 6420 9920
rect 8392 9936 8444 9988
rect 8944 10013 8953 10047
rect 8953 10013 8987 10047
rect 8987 10013 8996 10047
rect 8944 10004 8996 10013
rect 10784 10072 10836 10124
rect 10600 10004 10652 10056
rect 11704 10072 11756 10124
rect 11888 10115 11940 10124
rect 11888 10081 11897 10115
rect 11897 10081 11931 10115
rect 11931 10081 11940 10115
rect 12624 10115 12676 10124
rect 11888 10072 11940 10081
rect 12624 10081 12633 10115
rect 12633 10081 12667 10115
rect 12667 10081 12676 10115
rect 12624 10072 12676 10081
rect 13084 10072 13136 10124
rect 14188 10140 14240 10192
rect 13176 10004 13228 10056
rect 13636 10072 13688 10124
rect 13820 10004 13872 10056
rect 10600 9868 10652 9920
rect 11152 9868 11204 9920
rect 11704 9911 11756 9920
rect 11704 9877 11713 9911
rect 11713 9877 11747 9911
rect 11747 9877 11756 9911
rect 11704 9868 11756 9877
rect 12072 9911 12124 9920
rect 12072 9877 12081 9911
rect 12081 9877 12115 9911
rect 12115 9877 12124 9911
rect 12072 9868 12124 9877
rect 12808 9868 12860 9920
rect 13360 9979 13412 9988
rect 13360 9945 13369 9979
rect 13369 9945 13403 9979
rect 13403 9945 13412 9979
rect 13360 9936 13412 9945
rect 14556 9936 14608 9988
rect 13636 9868 13688 9920
rect 14096 9911 14148 9920
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 14188 9868 14240 9920
rect 4698 9766 4750 9818
rect 4762 9766 4814 9818
rect 4826 9766 4878 9818
rect 4890 9766 4942 9818
rect 4954 9766 5006 9818
rect 8446 9766 8498 9818
rect 8510 9766 8562 9818
rect 8574 9766 8626 9818
rect 8638 9766 8690 9818
rect 8702 9766 8754 9818
rect 12194 9766 12246 9818
rect 12258 9766 12310 9818
rect 12322 9766 12374 9818
rect 12386 9766 12438 9818
rect 12450 9766 12502 9818
rect 2504 9664 2556 9716
rect 4344 9664 4396 9716
rect 2688 9528 2740 9580
rect 2964 9571 3016 9580
rect 2964 9537 2982 9571
rect 2982 9537 3016 9571
rect 2964 9528 3016 9537
rect 3424 9528 3476 9580
rect 4160 9528 4212 9580
rect 4436 9528 4488 9580
rect 5172 9596 5224 9648
rect 6460 9596 6512 9648
rect 6368 9571 6420 9580
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 6920 9664 6972 9716
rect 7932 9664 7984 9716
rect 9036 9664 9088 9716
rect 9864 9664 9916 9716
rect 11428 9664 11480 9716
rect 6736 9596 6788 9648
rect 7380 9596 7432 9648
rect 7748 9596 7800 9648
rect 8208 9528 8260 9580
rect 8668 9528 8720 9580
rect 9128 9528 9180 9580
rect 9956 9528 10008 9580
rect 1676 9392 1728 9444
rect 1860 9435 1912 9444
rect 1860 9401 1869 9435
rect 1869 9401 1903 9435
rect 1903 9401 1912 9435
rect 1860 9392 1912 9401
rect 10600 9460 10652 9512
rect 11428 9528 11480 9580
rect 12532 9664 12584 9716
rect 13360 9664 13412 9716
rect 14188 9664 14240 9716
rect 14740 9664 14792 9716
rect 14832 9707 14884 9716
rect 14832 9673 14841 9707
rect 14841 9673 14875 9707
rect 14875 9673 14884 9707
rect 14832 9664 14884 9673
rect 15108 9664 15160 9716
rect 12440 9596 12492 9648
rect 12532 9528 12584 9580
rect 12992 9528 13044 9580
rect 13452 9528 13504 9580
rect 7656 9392 7708 9444
rect 4252 9324 4304 9376
rect 4436 9324 4488 9376
rect 5448 9324 5500 9376
rect 5816 9324 5868 9376
rect 7104 9324 7156 9376
rect 8944 9324 8996 9376
rect 9680 9324 9732 9376
rect 9956 9324 10008 9376
rect 10784 9392 10836 9444
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 10692 9324 10744 9333
rect 11888 9460 11940 9512
rect 12072 9503 12124 9512
rect 12072 9469 12081 9503
rect 12081 9469 12115 9503
rect 12115 9469 12124 9503
rect 12900 9503 12952 9512
rect 12072 9460 12124 9469
rect 12900 9469 12909 9503
rect 12909 9469 12943 9503
rect 12943 9469 12952 9503
rect 12900 9460 12952 9469
rect 13084 9460 13136 9512
rect 11796 9392 11848 9444
rect 14648 9528 14700 9580
rect 14832 9528 14884 9580
rect 14556 9503 14608 9512
rect 13176 9367 13228 9376
rect 13176 9333 13185 9367
rect 13185 9333 13219 9367
rect 13219 9333 13228 9367
rect 13176 9324 13228 9333
rect 13728 9324 13780 9376
rect 14556 9469 14565 9503
rect 14565 9469 14599 9503
rect 14599 9469 14608 9503
rect 14556 9460 14608 9469
rect 14464 9392 14516 9444
rect 14832 9392 14884 9444
rect 15292 9324 15344 9376
rect 2824 9222 2876 9274
rect 2888 9222 2940 9274
rect 2952 9222 3004 9274
rect 3016 9222 3068 9274
rect 3080 9222 3132 9274
rect 6572 9222 6624 9274
rect 6636 9222 6688 9274
rect 6700 9222 6752 9274
rect 6764 9222 6816 9274
rect 6828 9222 6880 9274
rect 10320 9222 10372 9274
rect 10384 9222 10436 9274
rect 10448 9222 10500 9274
rect 10512 9222 10564 9274
rect 10576 9222 10628 9274
rect 14068 9222 14120 9274
rect 14132 9222 14184 9274
rect 14196 9222 14248 9274
rect 14260 9222 14312 9274
rect 14324 9222 14376 9274
rect 3516 9120 3568 9172
rect 3792 9120 3844 9172
rect 4252 9120 4304 9172
rect 4620 9120 4672 9172
rect 6920 9120 6972 9172
rect 9036 9120 9088 9172
rect 9404 9120 9456 9172
rect 11244 9163 11296 9172
rect 11244 9129 11253 9163
rect 11253 9129 11287 9163
rect 11287 9129 11296 9163
rect 11244 9120 11296 9129
rect 11704 9120 11756 9172
rect 2136 9095 2188 9104
rect 2136 9061 2145 9095
rect 2145 9061 2179 9095
rect 2179 9061 2188 9095
rect 2136 9052 2188 9061
rect 3884 9052 3936 9104
rect 5908 9095 5960 9104
rect 5908 9061 5917 9095
rect 5917 9061 5951 9095
rect 5951 9061 5960 9095
rect 5908 9052 5960 9061
rect 6184 9052 6236 9104
rect 10692 9052 10744 9104
rect 14556 9120 14608 9172
rect 15476 9120 15528 9172
rect 12900 9095 12952 9104
rect 12900 9061 12909 9095
rect 12909 9061 12943 9095
rect 12943 9061 12952 9095
rect 12900 9052 12952 9061
rect 13636 9052 13688 9104
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 2228 9027 2280 9036
rect 1676 8984 1728 8993
rect 2228 8993 2237 9027
rect 2237 8993 2271 9027
rect 2271 8993 2280 9027
rect 2228 8984 2280 8993
rect 3976 9027 4028 9036
rect 3976 8993 3985 9027
rect 3985 8993 4019 9027
rect 4019 8993 4028 9027
rect 3976 8984 4028 8993
rect 1124 8916 1176 8968
rect 5540 8959 5592 8968
rect 3148 8848 3200 8900
rect 4252 8780 4304 8832
rect 5080 8780 5132 8832
rect 5540 8925 5558 8959
rect 5558 8925 5592 8959
rect 5540 8916 5592 8925
rect 8392 8984 8444 9036
rect 6184 8916 6236 8968
rect 9128 8916 9180 8968
rect 9496 8916 9548 8968
rect 11888 9027 11940 9036
rect 11888 8993 11897 9027
rect 11897 8993 11931 9027
rect 11931 8993 11940 9027
rect 11888 8984 11940 8993
rect 12716 9027 12768 9036
rect 12716 8993 12725 9027
rect 12725 8993 12759 9027
rect 12759 8993 12768 9027
rect 12716 8984 12768 8993
rect 13268 8984 13320 9036
rect 14464 9052 14516 9104
rect 14556 9027 14608 9036
rect 10508 8916 10560 8968
rect 10784 8916 10836 8968
rect 11060 8916 11112 8968
rect 11796 8916 11848 8968
rect 12072 8916 12124 8968
rect 12164 8916 12216 8968
rect 12808 8916 12860 8968
rect 14556 8993 14565 9027
rect 14565 8993 14599 9027
rect 14599 8993 14608 9027
rect 14556 8984 14608 8993
rect 14832 9052 14884 9104
rect 15292 9052 15344 9104
rect 16120 9052 16172 9104
rect 16580 9052 16632 9104
rect 7012 8891 7064 8900
rect 7012 8857 7030 8891
rect 7030 8857 7064 8891
rect 7012 8848 7064 8857
rect 7196 8848 7248 8900
rect 5724 8780 5776 8832
rect 8852 8780 8904 8832
rect 9680 8848 9732 8900
rect 10232 8848 10284 8900
rect 13084 8848 13136 8900
rect 13544 8848 13596 8900
rect 10784 8823 10836 8832
rect 10784 8789 10793 8823
rect 10793 8789 10827 8823
rect 10827 8789 10836 8823
rect 10784 8780 10836 8789
rect 11244 8780 11296 8832
rect 15660 8848 15712 8900
rect 13820 8780 13872 8832
rect 16212 8780 16264 8832
rect 16396 8780 16448 8832
rect 4698 8678 4750 8730
rect 4762 8678 4814 8730
rect 4826 8678 4878 8730
rect 4890 8678 4942 8730
rect 4954 8678 5006 8730
rect 8446 8678 8498 8730
rect 8510 8678 8562 8730
rect 8574 8678 8626 8730
rect 8638 8678 8690 8730
rect 8702 8678 8754 8730
rect 12194 8678 12246 8730
rect 12258 8678 12310 8730
rect 12322 8678 12374 8730
rect 12386 8678 12438 8730
rect 12450 8678 12502 8730
rect 2412 8576 2464 8628
rect 3332 8576 3384 8628
rect 1952 8440 2004 8492
rect 1400 8304 1452 8356
rect 4160 8440 4212 8492
rect 4436 8483 4488 8492
rect 4436 8449 4454 8483
rect 4454 8449 4488 8483
rect 4436 8440 4488 8449
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 2596 8236 2648 8288
rect 3424 8236 3476 8288
rect 6000 8576 6052 8628
rect 7748 8619 7800 8628
rect 7748 8585 7757 8619
rect 7757 8585 7791 8619
rect 7791 8585 7800 8619
rect 7748 8576 7800 8585
rect 9128 8619 9180 8628
rect 9128 8585 9137 8619
rect 9137 8585 9171 8619
rect 9171 8585 9180 8619
rect 9128 8576 9180 8585
rect 5816 8508 5868 8560
rect 7012 8508 7064 8560
rect 11244 8576 11296 8628
rect 11520 8619 11572 8628
rect 11520 8585 11529 8619
rect 11529 8585 11563 8619
rect 11563 8585 11572 8619
rect 11520 8576 11572 8585
rect 11796 8576 11848 8628
rect 13176 8619 13228 8628
rect 13176 8585 13185 8619
rect 13185 8585 13219 8619
rect 13219 8585 13228 8619
rect 13176 8576 13228 8585
rect 13912 8576 13964 8628
rect 14464 8576 14516 8628
rect 14740 8576 14792 8628
rect 15200 8619 15252 8628
rect 15200 8585 15209 8619
rect 15209 8585 15243 8619
rect 15243 8585 15252 8619
rect 15200 8576 15252 8585
rect 15568 8576 15620 8628
rect 5448 8440 5500 8492
rect 7104 8440 7156 8492
rect 7840 8483 7892 8492
rect 7840 8449 7849 8483
rect 7849 8449 7883 8483
rect 7883 8449 7892 8483
rect 7840 8440 7892 8449
rect 10232 8508 10284 8560
rect 10416 8508 10468 8560
rect 11704 8508 11756 8560
rect 12164 8508 12216 8560
rect 12992 8508 13044 8560
rect 13360 8508 13412 8560
rect 6184 8415 6236 8424
rect 6184 8381 6193 8415
rect 6193 8381 6227 8415
rect 6227 8381 6236 8415
rect 6184 8372 6236 8381
rect 7380 8372 7432 8424
rect 11612 8440 11664 8492
rect 12256 8440 12308 8492
rect 12348 8440 12400 8492
rect 12716 8483 12768 8492
rect 12716 8449 12725 8483
rect 12725 8449 12759 8483
rect 12759 8449 12768 8483
rect 12716 8440 12768 8449
rect 13176 8440 13228 8492
rect 14556 8440 14608 8492
rect 14832 8440 14884 8492
rect 10692 8372 10744 8424
rect 11796 8372 11848 8424
rect 12624 8372 12676 8424
rect 12992 8372 13044 8424
rect 13544 8372 13596 8424
rect 13636 8372 13688 8424
rect 14004 8372 14056 8424
rect 5448 8236 5500 8288
rect 14556 8304 14608 8356
rect 15660 8372 15712 8424
rect 11060 8279 11112 8288
rect 11060 8245 11069 8279
rect 11069 8245 11103 8279
rect 11103 8245 11112 8279
rect 11060 8236 11112 8245
rect 11704 8236 11756 8288
rect 12532 8236 12584 8288
rect 12900 8236 12952 8288
rect 16764 8236 16816 8288
rect 2824 8134 2876 8186
rect 2888 8134 2940 8186
rect 2952 8134 3004 8186
rect 3016 8134 3068 8186
rect 3080 8134 3132 8186
rect 6572 8134 6624 8186
rect 6636 8134 6688 8186
rect 6700 8134 6752 8186
rect 6764 8134 6816 8186
rect 6828 8134 6880 8186
rect 10320 8134 10372 8186
rect 10384 8134 10436 8186
rect 10448 8134 10500 8186
rect 10512 8134 10564 8186
rect 10576 8134 10628 8186
rect 14068 8134 14120 8186
rect 14132 8134 14184 8186
rect 14196 8134 14248 8186
rect 14260 8134 14312 8186
rect 14324 8134 14376 8186
rect 1860 8075 1912 8084
rect 1860 8041 1869 8075
rect 1869 8041 1903 8075
rect 1903 8041 1912 8075
rect 1860 8032 1912 8041
rect 2228 8032 2280 8084
rect 4712 8032 4764 8084
rect 5172 8032 5224 8084
rect 5724 8032 5776 8084
rect 10692 8032 10744 8084
rect 10784 8032 10836 8084
rect 12256 8032 12308 8084
rect 13360 8032 13412 8084
rect 16120 8032 16172 8084
rect 2136 7896 2188 7948
rect 5172 7896 5224 7948
rect 5632 7896 5684 7948
rect 3608 7871 3660 7880
rect 3608 7837 3617 7871
rect 3617 7837 3651 7871
rect 3651 7837 3660 7871
rect 3608 7828 3660 7837
rect 3700 7828 3752 7880
rect 4068 7828 4120 7880
rect 5356 7828 5408 7880
rect 6460 7828 6512 7880
rect 7840 7828 7892 7880
rect 9312 7828 9364 7880
rect 9772 7828 9824 7880
rect 10232 7828 10284 7880
rect 12164 7896 12216 7948
rect 12348 7939 12400 7948
rect 12348 7905 12357 7939
rect 12357 7905 12391 7939
rect 12391 7905 12400 7939
rect 12348 7896 12400 7905
rect 14004 7964 14056 8016
rect 15384 7964 15436 8016
rect 3424 7735 3476 7744
rect 3424 7701 3433 7735
rect 3433 7701 3467 7735
rect 3467 7701 3476 7735
rect 3424 7692 3476 7701
rect 5632 7692 5684 7744
rect 9036 7760 9088 7812
rect 9404 7760 9456 7812
rect 11796 7828 11848 7880
rect 13544 7896 13596 7948
rect 15108 7896 15160 7948
rect 15476 7939 15528 7948
rect 15476 7905 15485 7939
rect 15485 7905 15519 7939
rect 15519 7905 15528 7939
rect 15476 7896 15528 7905
rect 14004 7828 14056 7880
rect 15660 7828 15712 7880
rect 10692 7803 10744 7812
rect 10692 7769 10726 7803
rect 10726 7769 10744 7803
rect 10692 7760 10744 7769
rect 7840 7692 7892 7744
rect 7932 7692 7984 7744
rect 12624 7760 12676 7812
rect 13728 7760 13780 7812
rect 13820 7760 13872 7812
rect 14096 7760 14148 7812
rect 14648 7760 14700 7812
rect 15108 7760 15160 7812
rect 15200 7760 15252 7812
rect 16120 7760 16172 7812
rect 11244 7692 11296 7744
rect 11796 7735 11848 7744
rect 11796 7701 11805 7735
rect 11805 7701 11839 7735
rect 11839 7701 11848 7735
rect 11796 7692 11848 7701
rect 11888 7735 11940 7744
rect 11888 7701 11897 7735
rect 11897 7701 11931 7735
rect 11931 7701 11940 7735
rect 12992 7735 13044 7744
rect 11888 7692 11940 7701
rect 12992 7701 13001 7735
rect 13001 7701 13035 7735
rect 13035 7701 13044 7735
rect 12992 7692 13044 7701
rect 13268 7692 13320 7744
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 13912 7692 13964 7744
rect 14464 7735 14516 7744
rect 14464 7701 14473 7735
rect 14473 7701 14507 7735
rect 14507 7701 14516 7735
rect 14464 7692 14516 7701
rect 14740 7692 14792 7744
rect 15292 7735 15344 7744
rect 15292 7701 15301 7735
rect 15301 7701 15335 7735
rect 15335 7701 15344 7735
rect 15292 7692 15344 7701
rect 15660 7692 15712 7744
rect 4698 7590 4750 7642
rect 4762 7590 4814 7642
rect 4826 7590 4878 7642
rect 4890 7590 4942 7642
rect 4954 7590 5006 7642
rect 8446 7590 8498 7642
rect 8510 7590 8562 7642
rect 8574 7590 8626 7642
rect 8638 7590 8690 7642
rect 8702 7590 8754 7642
rect 12194 7590 12246 7642
rect 12258 7590 12310 7642
rect 12322 7590 12374 7642
rect 12386 7590 12438 7642
rect 12450 7590 12502 7642
rect 2136 7488 2188 7540
rect 4528 7488 4580 7540
rect 5080 7488 5132 7540
rect 4160 7420 4212 7472
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 1860 7395 1912 7404
rect 1860 7361 1869 7395
rect 1869 7361 1903 7395
rect 1903 7361 1912 7395
rect 1860 7352 1912 7361
rect 2504 7352 2556 7404
rect 4620 7352 4672 7404
rect 5172 7420 5224 7472
rect 8024 7488 8076 7540
rect 5448 7352 5500 7404
rect 10048 7488 10100 7540
rect 10968 7488 11020 7540
rect 11152 7531 11204 7540
rect 11152 7497 11161 7531
rect 11161 7497 11195 7531
rect 11195 7497 11204 7531
rect 11152 7488 11204 7497
rect 11244 7420 11296 7472
rect 6920 7352 6972 7404
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 8024 7352 8076 7404
rect 9036 7352 9088 7404
rect 9496 7352 9548 7404
rect 6184 7327 6236 7336
rect 6184 7293 6193 7327
rect 6193 7293 6227 7327
rect 6227 7293 6236 7327
rect 6184 7284 6236 7293
rect 9312 7284 9364 7336
rect 9772 7352 9824 7404
rect 9956 7395 10008 7404
rect 9956 7361 9990 7395
rect 9990 7361 10008 7395
rect 9956 7352 10008 7361
rect 11152 7352 11204 7404
rect 13268 7488 13320 7540
rect 13728 7488 13780 7540
rect 14924 7488 14976 7540
rect 12256 7420 12308 7472
rect 11980 7395 12032 7404
rect 11980 7361 11989 7395
rect 11989 7361 12023 7395
rect 12023 7361 12032 7395
rect 11980 7352 12032 7361
rect 12440 7352 12492 7404
rect 12716 7395 12768 7404
rect 12716 7361 12725 7395
rect 12725 7361 12759 7395
rect 12759 7361 12768 7395
rect 12716 7352 12768 7361
rect 12992 7420 13044 7472
rect 15200 7463 15252 7472
rect 15200 7429 15209 7463
rect 15209 7429 15243 7463
rect 15243 7429 15252 7463
rect 15200 7420 15252 7429
rect 10692 7284 10744 7336
rect 10968 7284 11020 7336
rect 11244 7284 11296 7336
rect 3056 7216 3108 7268
rect 2228 7148 2280 7200
rect 3332 7148 3384 7200
rect 6460 7148 6512 7200
rect 8208 7216 8260 7268
rect 9404 7216 9456 7268
rect 11520 7259 11572 7268
rect 11520 7225 11529 7259
rect 11529 7225 11563 7259
rect 11563 7225 11572 7259
rect 11520 7216 11572 7225
rect 13544 7352 13596 7404
rect 14372 7352 14424 7404
rect 14556 7352 14608 7404
rect 15016 7352 15068 7404
rect 7840 7148 7892 7200
rect 10692 7148 10744 7200
rect 11060 7191 11112 7200
rect 11060 7157 11069 7191
rect 11069 7157 11103 7191
rect 11103 7157 11112 7191
rect 11060 7148 11112 7157
rect 11152 7148 11204 7200
rect 12348 7216 12400 7268
rect 12624 7216 12676 7268
rect 12716 7216 12768 7268
rect 13728 7284 13780 7336
rect 12532 7148 12584 7200
rect 12808 7148 12860 7200
rect 15292 7327 15344 7336
rect 15292 7293 15301 7327
rect 15301 7293 15335 7327
rect 15335 7293 15344 7327
rect 15292 7284 15344 7293
rect 14004 7259 14056 7268
rect 14004 7225 14013 7259
rect 14013 7225 14047 7259
rect 14047 7225 14056 7259
rect 14004 7216 14056 7225
rect 15200 7216 15252 7268
rect 15016 7148 15068 7200
rect 2824 7046 2876 7098
rect 2888 7046 2940 7098
rect 2952 7046 3004 7098
rect 3016 7046 3068 7098
rect 3080 7046 3132 7098
rect 6572 7046 6624 7098
rect 6636 7046 6688 7098
rect 6700 7046 6752 7098
rect 6764 7046 6816 7098
rect 6828 7046 6880 7098
rect 10320 7046 10372 7098
rect 10384 7046 10436 7098
rect 10448 7046 10500 7098
rect 10512 7046 10564 7098
rect 10576 7046 10628 7098
rect 14068 7046 14120 7098
rect 14132 7046 14184 7098
rect 14196 7046 14248 7098
rect 14260 7046 14312 7098
rect 14324 7046 14376 7098
rect 3884 6944 3936 6996
rect 7104 6944 7156 6996
rect 7656 6944 7708 6996
rect 9680 6944 9732 6996
rect 9956 6944 10008 6996
rect 10784 6944 10836 6996
rect 11152 6944 11204 6996
rect 11888 6944 11940 6996
rect 6276 6876 6328 6928
rect 10968 6876 11020 6928
rect 11336 6876 11388 6928
rect 12164 6944 12216 6996
rect 12256 6876 12308 6928
rect 13268 6876 13320 6928
rect 2596 6808 2648 6860
rect 3976 6851 4028 6860
rect 3976 6817 3985 6851
rect 3985 6817 4019 6851
rect 4019 6817 4028 6851
rect 3976 6808 4028 6817
rect 6184 6808 6236 6860
rect 9312 6808 9364 6860
rect 848 6740 900 6792
rect 1492 6740 1544 6792
rect 3516 6740 3568 6792
rect 4160 6740 4212 6792
rect 5172 6740 5224 6792
rect 1676 6647 1728 6656
rect 1676 6613 1685 6647
rect 1685 6613 1719 6647
rect 1719 6613 1728 6647
rect 1676 6604 1728 6613
rect 2412 6604 2464 6656
rect 4436 6647 4488 6656
rect 4436 6613 4445 6647
rect 4445 6613 4479 6647
rect 4479 6613 4488 6647
rect 4436 6604 4488 6613
rect 5264 6604 5316 6656
rect 5448 6604 5500 6656
rect 7012 6715 7064 6724
rect 7012 6681 7030 6715
rect 7030 6681 7064 6715
rect 7012 6672 7064 6681
rect 7748 6740 7800 6792
rect 8116 6740 8168 6792
rect 9864 6672 9916 6724
rect 7840 6604 7892 6656
rect 7932 6604 7984 6656
rect 9128 6604 9180 6656
rect 9404 6604 9456 6656
rect 9496 6604 9548 6656
rect 9772 6604 9824 6656
rect 10232 6740 10284 6792
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10692 6808 10744 6860
rect 11520 6808 11572 6860
rect 11796 6808 11848 6860
rect 11888 6851 11940 6860
rect 11888 6817 11897 6851
rect 11897 6817 11931 6851
rect 11931 6817 11940 6851
rect 11888 6808 11940 6817
rect 12716 6808 12768 6860
rect 12900 6808 12952 6860
rect 13360 6851 13412 6860
rect 13360 6817 13369 6851
rect 13369 6817 13403 6851
rect 13403 6817 13412 6851
rect 13360 6808 13412 6817
rect 13636 6944 13688 6996
rect 13728 6944 13780 6996
rect 15568 6944 15620 6996
rect 14280 6876 14332 6928
rect 14648 6851 14700 6860
rect 14648 6817 14657 6851
rect 14657 6817 14691 6851
rect 14691 6817 14700 6851
rect 14648 6808 14700 6817
rect 15200 6808 15252 6860
rect 10324 6740 10376 6749
rect 10416 6672 10468 6724
rect 10968 6672 11020 6724
rect 11612 6783 11664 6792
rect 11612 6749 11621 6783
rect 11621 6749 11655 6783
rect 11655 6749 11664 6783
rect 11612 6740 11664 6749
rect 12440 6783 12492 6792
rect 12440 6749 12449 6783
rect 12449 6749 12483 6783
rect 12483 6749 12492 6783
rect 12440 6740 12492 6749
rect 10600 6604 10652 6656
rect 10876 6604 10928 6656
rect 11796 6604 11848 6656
rect 13084 6672 13136 6724
rect 13728 6740 13780 6792
rect 14556 6740 14608 6792
rect 14832 6672 14884 6724
rect 13544 6604 13596 6656
rect 13912 6604 13964 6656
rect 14096 6647 14148 6656
rect 14096 6613 14105 6647
rect 14105 6613 14139 6647
rect 14139 6613 14148 6647
rect 14096 6604 14148 6613
rect 14188 6604 14240 6656
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14924 6647 14976 6656
rect 14556 6604 14608 6613
rect 14924 6613 14933 6647
rect 14933 6613 14967 6647
rect 14967 6613 14976 6647
rect 14924 6604 14976 6613
rect 15108 6604 15160 6656
rect 4698 6502 4750 6554
rect 4762 6502 4814 6554
rect 4826 6502 4878 6554
rect 4890 6502 4942 6554
rect 4954 6502 5006 6554
rect 8446 6502 8498 6554
rect 8510 6502 8562 6554
rect 8574 6502 8626 6554
rect 8638 6502 8690 6554
rect 8702 6502 8754 6554
rect 12194 6502 12246 6554
rect 12258 6502 12310 6554
rect 12322 6502 12374 6554
rect 12386 6502 12438 6554
rect 12450 6502 12502 6554
rect 3608 6400 3660 6452
rect 4620 6400 4672 6452
rect 6092 6400 6144 6452
rect 8116 6400 8168 6452
rect 8300 6400 8352 6452
rect 10784 6400 10836 6452
rect 2228 6332 2280 6384
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 1860 6307 1912 6316
rect 1860 6273 1869 6307
rect 1869 6273 1903 6307
rect 1903 6273 1912 6307
rect 2136 6307 2188 6316
rect 1860 6264 1912 6273
rect 2136 6273 2170 6307
rect 2170 6273 2188 6307
rect 2136 6264 2188 6273
rect 4160 6332 4212 6384
rect 4528 6264 4580 6316
rect 4804 6307 4856 6316
rect 4804 6273 4813 6307
rect 4813 6273 4847 6307
rect 4847 6273 4856 6307
rect 4804 6264 4856 6273
rect 5356 6264 5408 6316
rect 7196 6332 7248 6384
rect 6460 6264 6512 6316
rect 7012 6264 7064 6316
rect 7748 6264 7800 6316
rect 8484 6264 8536 6316
rect 9404 6332 9456 6384
rect 9680 6332 9732 6384
rect 10140 6332 10192 6384
rect 11520 6332 11572 6384
rect 12164 6332 12216 6384
rect 9864 6264 9916 6316
rect 11612 6264 11664 6316
rect 11704 6264 11756 6316
rect 12900 6332 12952 6384
rect 13544 6443 13596 6452
rect 13268 6332 13320 6384
rect 13544 6409 13553 6443
rect 13553 6409 13587 6443
rect 13587 6409 13596 6443
rect 13544 6400 13596 6409
rect 14004 6443 14056 6452
rect 14004 6409 14013 6443
rect 14013 6409 14047 6443
rect 14047 6409 14056 6443
rect 14004 6400 14056 6409
rect 14096 6400 14148 6452
rect 14648 6400 14700 6452
rect 14924 6332 14976 6384
rect 9312 6239 9364 6248
rect 9312 6205 9321 6239
rect 9321 6205 9355 6239
rect 9355 6205 9364 6239
rect 9312 6196 9364 6205
rect 10784 6196 10836 6248
rect 11152 6196 11204 6248
rect 12072 6239 12124 6248
rect 12072 6205 12081 6239
rect 12081 6205 12115 6239
rect 12115 6205 12124 6239
rect 12072 6196 12124 6205
rect 13912 6264 13964 6316
rect 12256 6196 12308 6248
rect 12808 6196 12860 6248
rect 12900 6196 12952 6248
rect 13084 6196 13136 6248
rect 13820 6239 13872 6248
rect 13820 6205 13829 6239
rect 13829 6205 13863 6239
rect 13863 6205 13872 6239
rect 13820 6196 13872 6205
rect 14464 6239 14516 6248
rect 14464 6205 14473 6239
rect 14473 6205 14507 6239
rect 14507 6205 14516 6239
rect 14464 6196 14516 6205
rect 16028 6264 16080 6316
rect 14832 6239 14884 6248
rect 14832 6205 14841 6239
rect 14841 6205 14875 6239
rect 14875 6205 14884 6239
rect 14832 6196 14884 6205
rect 9036 6128 9088 6180
rect 4528 6060 4580 6112
rect 5908 6060 5960 6112
rect 6184 6103 6236 6112
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 7104 6060 7156 6112
rect 7564 6060 7616 6112
rect 9128 6060 9180 6112
rect 9312 6060 9364 6112
rect 11612 6128 11664 6180
rect 14188 6128 14240 6180
rect 14280 6128 14332 6180
rect 14648 6128 14700 6180
rect 15660 6128 15712 6180
rect 16028 6128 16080 6180
rect 10784 6060 10836 6112
rect 10968 6060 11020 6112
rect 11428 6060 11480 6112
rect 12900 6060 12952 6112
rect 13176 6103 13228 6112
rect 13176 6069 13185 6103
rect 13185 6069 13219 6103
rect 13219 6069 13228 6103
rect 13176 6060 13228 6069
rect 13820 6060 13872 6112
rect 14924 6060 14976 6112
rect 15936 6060 15988 6112
rect 2824 5958 2876 6010
rect 2888 5958 2940 6010
rect 2952 5958 3004 6010
rect 3016 5958 3068 6010
rect 3080 5958 3132 6010
rect 6572 5958 6624 6010
rect 6636 5958 6688 6010
rect 6700 5958 6752 6010
rect 6764 5958 6816 6010
rect 6828 5958 6880 6010
rect 10320 5958 10372 6010
rect 10384 5958 10436 6010
rect 10448 5958 10500 6010
rect 10512 5958 10564 6010
rect 10576 5958 10628 6010
rect 14068 5958 14120 6010
rect 14132 5958 14184 6010
rect 14196 5958 14248 6010
rect 14260 5958 14312 6010
rect 14324 5958 14376 6010
rect 1952 5856 2004 5908
rect 2136 5856 2188 5908
rect 4160 5856 4212 5908
rect 7380 5856 7432 5908
rect 7472 5856 7524 5908
rect 7840 5856 7892 5908
rect 3792 5788 3844 5840
rect 8484 5831 8536 5840
rect 8484 5797 8493 5831
rect 8493 5797 8527 5831
rect 8527 5797 8536 5831
rect 8484 5788 8536 5797
rect 4804 5652 4856 5704
rect 1860 5559 1912 5568
rect 1860 5525 1869 5559
rect 1869 5525 1903 5559
rect 1903 5525 1912 5559
rect 1860 5516 1912 5525
rect 5080 5584 5132 5636
rect 5264 5516 5316 5568
rect 5632 5652 5684 5704
rect 7748 5652 7800 5704
rect 8944 5720 8996 5772
rect 9220 5763 9272 5772
rect 9220 5729 9229 5763
rect 9229 5729 9263 5763
rect 9263 5729 9272 5763
rect 9220 5720 9272 5729
rect 9956 5788 10008 5840
rect 10140 5788 10192 5840
rect 11060 5720 11112 5772
rect 11796 5856 11848 5908
rect 12440 5856 12492 5908
rect 12900 5856 12952 5908
rect 11704 5788 11756 5840
rect 12164 5788 12216 5840
rect 12624 5788 12676 5840
rect 12808 5788 12860 5840
rect 6460 5584 6512 5636
rect 8668 5652 8720 5704
rect 10968 5652 11020 5704
rect 11612 5652 11664 5704
rect 12532 5652 12584 5704
rect 12716 5720 12768 5772
rect 12900 5763 12952 5772
rect 12900 5729 12909 5763
rect 12909 5729 12943 5763
rect 12943 5729 12952 5763
rect 13268 5788 13320 5840
rect 14004 5788 14056 5840
rect 12900 5720 12952 5729
rect 13544 5695 13596 5704
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 8576 5584 8628 5636
rect 12072 5584 12124 5636
rect 14096 5584 14148 5636
rect 14924 5856 14976 5908
rect 16580 5856 16632 5908
rect 14832 5831 14884 5840
rect 14832 5797 14841 5831
rect 14841 5797 14875 5831
rect 14875 5797 14884 5831
rect 14832 5788 14884 5797
rect 16304 5788 16356 5840
rect 15752 5720 15804 5772
rect 15844 5652 15896 5704
rect 14832 5584 14884 5636
rect 15752 5584 15804 5636
rect 16028 5584 16080 5636
rect 6552 5559 6604 5568
rect 6552 5525 6561 5559
rect 6561 5525 6595 5559
rect 6595 5525 6604 5559
rect 6552 5516 6604 5525
rect 8208 5516 8260 5568
rect 9128 5516 9180 5568
rect 9680 5559 9732 5568
rect 9680 5525 9689 5559
rect 9689 5525 9723 5559
rect 9723 5525 9732 5559
rect 9680 5516 9732 5525
rect 9772 5516 9824 5568
rect 10508 5516 10560 5568
rect 10784 5516 10836 5568
rect 11244 5516 11296 5568
rect 11428 5516 11480 5568
rect 11520 5516 11572 5568
rect 11796 5516 11848 5568
rect 11980 5516 12032 5568
rect 12532 5516 12584 5568
rect 12624 5516 12676 5568
rect 12992 5516 13044 5568
rect 16764 5516 16816 5568
rect 4698 5414 4750 5466
rect 4762 5414 4814 5466
rect 4826 5414 4878 5466
rect 4890 5414 4942 5466
rect 4954 5414 5006 5466
rect 8446 5414 8498 5466
rect 8510 5414 8562 5466
rect 8574 5414 8626 5466
rect 8638 5414 8690 5466
rect 8702 5414 8754 5466
rect 12194 5414 12246 5466
rect 12258 5414 12310 5466
rect 12322 5414 12374 5466
rect 12386 5414 12438 5466
rect 12450 5414 12502 5466
rect 1676 5312 1728 5364
rect 2136 5355 2188 5364
rect 2136 5321 2145 5355
rect 2145 5321 2179 5355
rect 2179 5321 2188 5355
rect 2136 5312 2188 5321
rect 4344 5355 4396 5364
rect 3792 5244 3844 5296
rect 4344 5321 4353 5355
rect 4353 5321 4387 5355
rect 4387 5321 4396 5355
rect 4344 5312 4396 5321
rect 5080 5312 5132 5364
rect 8024 5312 8076 5364
rect 8944 5312 8996 5364
rect 10600 5355 10652 5364
rect 10600 5321 10609 5355
rect 10609 5321 10643 5355
rect 10643 5321 10652 5355
rect 10600 5312 10652 5321
rect 5448 5244 5500 5296
rect 6092 5244 6144 5296
rect 6276 5244 6328 5296
rect 7196 5244 7248 5296
rect 7656 5244 7708 5296
rect 2228 5219 2280 5228
rect 2228 5185 2237 5219
rect 2237 5185 2271 5219
rect 2271 5185 2280 5219
rect 2228 5176 2280 5185
rect 2320 5176 2372 5228
rect 3240 5176 3292 5228
rect 5172 5176 5224 5228
rect 7748 5219 7800 5228
rect 7748 5185 7757 5219
rect 7757 5185 7791 5219
rect 7791 5185 7800 5219
rect 7748 5176 7800 5185
rect 1308 5040 1360 5092
rect 4436 5108 4488 5160
rect 4252 5040 4304 5092
rect 5080 5040 5132 5092
rect 4620 4972 4672 5024
rect 4804 4972 4856 5024
rect 5448 4972 5500 5024
rect 6552 5108 6604 5160
rect 8852 5244 8904 5296
rect 10324 5244 10376 5296
rect 10416 5244 10468 5296
rect 8116 5219 8168 5228
rect 8116 5185 8150 5219
rect 8150 5185 8168 5219
rect 8116 5176 8168 5185
rect 10508 5176 10560 5228
rect 11060 5176 11112 5228
rect 11980 5355 12032 5364
rect 11980 5321 11989 5355
rect 11989 5321 12023 5355
rect 12023 5321 12032 5355
rect 11980 5312 12032 5321
rect 11796 5244 11848 5296
rect 12532 5244 12584 5296
rect 12900 5312 12952 5364
rect 11612 5176 11664 5228
rect 6368 5083 6420 5092
rect 6368 5049 6377 5083
rect 6377 5049 6411 5083
rect 6411 5049 6420 5083
rect 6368 5040 6420 5049
rect 6276 4972 6328 5024
rect 9220 5108 9272 5160
rect 7840 4972 7892 5024
rect 9864 5151 9916 5160
rect 9864 5117 9873 5151
rect 9873 5117 9907 5151
rect 9907 5117 9916 5151
rect 9864 5108 9916 5117
rect 10232 5108 10284 5160
rect 12256 5176 12308 5228
rect 12164 5151 12216 5160
rect 12164 5117 12173 5151
rect 12173 5117 12207 5151
rect 12207 5117 12216 5151
rect 12164 5108 12216 5117
rect 12808 5176 12860 5228
rect 13084 5244 13136 5296
rect 13728 5312 13780 5364
rect 15292 5312 15344 5364
rect 15476 5312 15528 5364
rect 14004 5287 14056 5296
rect 14004 5253 14013 5287
rect 14013 5253 14047 5287
rect 14047 5253 14056 5287
rect 14004 5244 14056 5253
rect 13636 5176 13688 5228
rect 13728 5176 13780 5228
rect 14648 5244 14700 5296
rect 15568 5244 15620 5296
rect 14280 5219 14332 5228
rect 14280 5185 14289 5219
rect 14289 5185 14323 5219
rect 14323 5185 14332 5219
rect 14280 5176 14332 5185
rect 14832 5176 14884 5228
rect 9220 5015 9272 5024
rect 9220 4981 9229 5015
rect 9229 4981 9263 5015
rect 9263 4981 9272 5015
rect 9220 4972 9272 4981
rect 9588 4972 9640 5024
rect 11980 5040 12032 5092
rect 12348 5040 12400 5092
rect 12256 4972 12308 5024
rect 14188 5108 14240 5160
rect 16120 5176 16172 5228
rect 15476 5108 15528 5160
rect 12532 4972 12584 5024
rect 14280 5040 14332 5092
rect 15292 5040 15344 5092
rect 13360 4972 13412 5024
rect 13820 4972 13872 5024
rect 14648 4972 14700 5024
rect 15568 5015 15620 5024
rect 15568 4981 15577 5015
rect 15577 4981 15611 5015
rect 15611 4981 15620 5015
rect 15568 4972 15620 4981
rect 16396 4972 16448 5024
rect 2824 4870 2876 4922
rect 2888 4870 2940 4922
rect 2952 4870 3004 4922
rect 3016 4870 3068 4922
rect 3080 4870 3132 4922
rect 6572 4870 6624 4922
rect 6636 4870 6688 4922
rect 6700 4870 6752 4922
rect 6764 4870 6816 4922
rect 6828 4870 6880 4922
rect 10320 4870 10372 4922
rect 10384 4870 10436 4922
rect 10448 4870 10500 4922
rect 10512 4870 10564 4922
rect 10576 4870 10628 4922
rect 14068 4870 14120 4922
rect 14132 4870 14184 4922
rect 14196 4870 14248 4922
rect 14260 4870 14312 4922
rect 14324 4870 14376 4922
rect 1584 4675 1636 4684
rect 1584 4641 1593 4675
rect 1593 4641 1627 4675
rect 1627 4641 1636 4675
rect 1584 4632 1636 4641
rect 2228 4768 2280 4820
rect 4436 4768 4488 4820
rect 8116 4768 8168 4820
rect 8208 4768 8260 4820
rect 8668 4768 8720 4820
rect 9128 4768 9180 4820
rect 9864 4768 9916 4820
rect 7012 4700 7064 4752
rect 8484 4700 8536 4752
rect 10784 4768 10836 4820
rect 11152 4768 11204 4820
rect 11612 4768 11664 4820
rect 12440 4768 12492 4820
rect 14648 4768 14700 4820
rect 14832 4811 14884 4820
rect 14832 4777 14841 4811
rect 14841 4777 14875 4811
rect 14875 4777 14884 4811
rect 14832 4768 14884 4777
rect 14924 4811 14976 4820
rect 14924 4777 14933 4811
rect 14933 4777 14967 4811
rect 14967 4777 14976 4811
rect 14924 4768 14976 4777
rect 15108 4768 15160 4820
rect 15292 4768 15344 4820
rect 5172 4632 5224 4684
rect 7288 4632 7340 4684
rect 8852 4632 8904 4684
rect 1768 4564 1820 4616
rect 2412 4564 2464 4616
rect 3516 4564 3568 4616
rect 4804 4564 4856 4616
rect 756 4428 808 4480
rect 1768 4471 1820 4480
rect 1768 4437 1777 4471
rect 1777 4437 1811 4471
rect 1811 4437 1820 4471
rect 1768 4428 1820 4437
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 3792 4428 3844 4480
rect 5264 4539 5316 4548
rect 5264 4505 5273 4539
rect 5273 4505 5307 4539
rect 5307 4505 5316 4539
rect 5264 4496 5316 4505
rect 6092 4564 6144 4616
rect 6736 4564 6788 4616
rect 6920 4564 6972 4616
rect 7748 4564 7800 4616
rect 8668 4564 8720 4616
rect 9404 4564 9456 4616
rect 9680 4564 9732 4616
rect 6368 4496 6420 4548
rect 8116 4496 8168 4548
rect 8208 4539 8260 4548
rect 8208 4505 8226 4539
rect 8226 4505 8260 4539
rect 10324 4632 10376 4684
rect 8208 4496 8260 4505
rect 6092 4428 6144 4480
rect 7012 4428 7064 4480
rect 9220 4471 9272 4480
rect 9220 4437 9229 4471
rect 9229 4437 9263 4471
rect 9263 4437 9272 4471
rect 9220 4428 9272 4437
rect 9312 4428 9364 4480
rect 9588 4428 9640 4480
rect 10508 4564 10560 4616
rect 10416 4496 10468 4548
rect 10784 4675 10836 4684
rect 10784 4641 10793 4675
rect 10793 4641 10827 4675
rect 10827 4641 10836 4675
rect 10784 4632 10836 4641
rect 11244 4632 11296 4684
rect 10968 4607 11020 4616
rect 10968 4573 10977 4607
rect 10977 4573 11011 4607
rect 11011 4573 11020 4607
rect 10968 4564 11020 4573
rect 11428 4700 11480 4752
rect 13636 4700 13688 4752
rect 15476 4700 15528 4752
rect 11612 4564 11664 4616
rect 11888 4632 11940 4684
rect 11244 4428 11296 4480
rect 11704 4428 11756 4480
rect 11888 4428 11940 4480
rect 12992 4632 13044 4684
rect 12072 4564 12124 4616
rect 14924 4632 14976 4684
rect 15660 4632 15712 4684
rect 13268 4564 13320 4616
rect 14188 4564 14240 4616
rect 15108 4564 15160 4616
rect 15384 4564 15436 4616
rect 15292 4539 15344 4548
rect 15292 4505 15301 4539
rect 15301 4505 15335 4539
rect 15335 4505 15344 4539
rect 15292 4496 15344 4505
rect 12072 4428 12124 4480
rect 12532 4471 12584 4480
rect 12532 4437 12541 4471
rect 12541 4437 12575 4471
rect 12575 4437 12584 4471
rect 12532 4428 12584 4437
rect 13084 4428 13136 4480
rect 13268 4428 13320 4480
rect 15752 4428 15804 4480
rect 16488 4428 16540 4480
rect 4698 4326 4750 4378
rect 4762 4326 4814 4378
rect 4826 4326 4878 4378
rect 4890 4326 4942 4378
rect 4954 4326 5006 4378
rect 8446 4326 8498 4378
rect 8510 4326 8562 4378
rect 8574 4326 8626 4378
rect 8638 4326 8690 4378
rect 8702 4326 8754 4378
rect 12194 4326 12246 4378
rect 12258 4326 12310 4378
rect 12322 4326 12374 4378
rect 12386 4326 12438 4378
rect 12450 4326 12502 4378
rect 1124 4224 1176 4276
rect 1676 4267 1728 4276
rect 1676 4233 1685 4267
rect 1685 4233 1719 4267
rect 1719 4233 1728 4267
rect 1676 4224 1728 4233
rect 2044 4224 2096 4276
rect 2320 4224 2372 4276
rect 2688 4224 2740 4276
rect 3240 4224 3292 4276
rect 3884 4224 3936 4276
rect 4436 4224 4488 4276
rect 2412 4156 2464 4208
rect 1860 4088 1912 4140
rect 2964 4131 3016 4140
rect 2964 4097 2982 4131
rect 2982 4097 3016 4131
rect 8852 4224 8904 4276
rect 2964 4088 3016 4097
rect 5080 4131 5132 4140
rect 5080 4097 5114 4131
rect 5114 4097 5132 4131
rect 5080 4088 5132 4097
rect 6276 4088 6328 4140
rect 6828 4131 6880 4140
rect 6828 4097 6837 4131
rect 6837 4097 6871 4131
rect 6871 4097 6880 4131
rect 6828 4088 6880 4097
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 7748 4156 7800 4208
rect 8024 4156 8076 4208
rect 10508 4224 10560 4276
rect 12624 4224 12676 4276
rect 13084 4267 13136 4276
rect 7656 4088 7708 4140
rect 6552 4063 6604 4072
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 8392 4088 8444 4140
rect 8300 4020 8352 4072
rect 8760 4088 8812 4140
rect 1768 3884 1820 3936
rect 3516 3884 3568 3936
rect 6276 3884 6328 3936
rect 8208 3884 8260 3936
rect 9404 4156 9456 4208
rect 10324 4156 10376 4208
rect 10140 4088 10192 4140
rect 11060 4156 11112 4208
rect 11152 4156 11204 4208
rect 11244 4156 11296 4208
rect 13084 4233 13093 4267
rect 13093 4233 13127 4267
rect 13127 4233 13136 4267
rect 13084 4224 13136 4233
rect 14096 4267 14148 4276
rect 13544 4199 13596 4208
rect 9588 4063 9640 4072
rect 9588 4029 9597 4063
rect 9597 4029 9631 4063
rect 9631 4029 9640 4063
rect 9588 4020 9640 4029
rect 9956 4020 10008 4072
rect 10692 4020 10744 4072
rect 9404 3952 9456 4004
rect 11612 4088 11664 4140
rect 13544 4165 13553 4199
rect 13553 4165 13587 4199
rect 13587 4165 13596 4199
rect 13544 4156 13596 4165
rect 14096 4233 14105 4267
rect 14105 4233 14139 4267
rect 14139 4233 14148 4267
rect 14096 4224 14148 4233
rect 14188 4224 14240 4276
rect 14464 4224 14516 4276
rect 14280 4131 14332 4140
rect 8392 3884 8444 3936
rect 8852 3884 8904 3936
rect 9036 3884 9088 3936
rect 9956 3884 10008 3936
rect 11060 3952 11112 4004
rect 11796 4020 11848 4072
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12440 4063 12492 4072
rect 12072 4020 12124 4029
rect 12440 4029 12449 4063
rect 12449 4029 12483 4063
rect 12483 4029 12492 4063
rect 12440 4020 12492 4029
rect 12440 3884 12492 3936
rect 12808 3952 12860 4004
rect 13268 3884 13320 3936
rect 13544 4020 13596 4072
rect 14280 4097 14289 4131
rect 14289 4097 14323 4131
rect 14323 4097 14332 4131
rect 14280 4088 14332 4097
rect 14832 4156 14884 4208
rect 14372 4020 14424 4072
rect 14924 4088 14976 4140
rect 14004 3952 14056 4004
rect 14832 3952 14884 4004
rect 14648 3884 14700 3936
rect 14924 3884 14976 3936
rect 2824 3782 2876 3834
rect 2888 3782 2940 3834
rect 2952 3782 3004 3834
rect 3016 3782 3068 3834
rect 3080 3782 3132 3834
rect 6572 3782 6624 3834
rect 6636 3782 6688 3834
rect 6700 3782 6752 3834
rect 6764 3782 6816 3834
rect 6828 3782 6880 3834
rect 10320 3782 10372 3834
rect 10384 3782 10436 3834
rect 10448 3782 10500 3834
rect 10512 3782 10564 3834
rect 10576 3782 10628 3834
rect 14068 3782 14120 3834
rect 14132 3782 14184 3834
rect 14196 3782 14248 3834
rect 14260 3782 14312 3834
rect 14324 3782 14376 3834
rect 3700 3680 3752 3732
rect 3792 3680 3844 3732
rect 5724 3680 5776 3732
rect 6460 3680 6512 3732
rect 7012 3680 7064 3732
rect 8668 3680 8720 3732
rect 2964 3612 3016 3664
rect 3056 3612 3108 3664
rect 3332 3612 3384 3664
rect 1860 3587 1912 3596
rect 1860 3553 1869 3587
rect 1869 3553 1903 3587
rect 1903 3553 1912 3587
rect 1860 3544 1912 3553
rect 940 3476 992 3528
rect 2688 3476 2740 3528
rect 3332 3519 3384 3528
rect 3332 3485 3341 3519
rect 3341 3485 3375 3519
rect 3375 3485 3384 3519
rect 3332 3476 3384 3485
rect 4528 3476 4580 3528
rect 5264 3655 5316 3664
rect 5264 3621 5273 3655
rect 5273 3621 5307 3655
rect 5307 3621 5316 3655
rect 5264 3612 5316 3621
rect 6552 3612 6604 3664
rect 9220 3680 9272 3732
rect 9588 3680 9640 3732
rect 11244 3680 11296 3732
rect 12532 3680 12584 3732
rect 7104 3612 7156 3664
rect 8392 3612 8444 3664
rect 8760 3655 8812 3664
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 7012 3587 7064 3596
rect 7012 3553 7021 3587
rect 7021 3553 7055 3587
rect 7055 3553 7064 3587
rect 7012 3544 7064 3553
rect 7380 3544 7432 3596
rect 7656 3544 7708 3596
rect 7932 3587 7984 3596
rect 7932 3553 7941 3587
rect 7941 3553 7975 3587
rect 7975 3553 7984 3587
rect 7932 3544 7984 3553
rect 8116 3544 8168 3596
rect 8760 3621 8769 3655
rect 8769 3621 8803 3655
rect 8803 3621 8812 3655
rect 8760 3612 8812 3621
rect 9680 3655 9732 3664
rect 8852 3544 8904 3596
rect 9680 3621 9689 3655
rect 9689 3621 9723 3655
rect 9723 3621 9732 3655
rect 9680 3612 9732 3621
rect 9864 3612 9916 3664
rect 10692 3612 10744 3664
rect 9036 3476 9088 3528
rect 10048 3476 10100 3528
rect 11428 3612 11480 3664
rect 12256 3612 12308 3664
rect 12808 3680 12860 3732
rect 12900 3680 12952 3732
rect 13452 3680 13504 3732
rect 15292 3680 15344 3732
rect 15384 3723 15436 3732
rect 15384 3689 15393 3723
rect 15393 3689 15427 3723
rect 15427 3689 15436 3723
rect 15384 3680 15436 3689
rect 13544 3612 13596 3664
rect 10968 3544 11020 3596
rect 11244 3544 11296 3596
rect 11060 3476 11112 3528
rect 11520 3476 11572 3528
rect 12348 3544 12400 3596
rect 11980 3476 12032 3528
rect 1676 3408 1728 3460
rect 2320 3408 2372 3460
rect 2412 3408 2464 3460
rect 7012 3408 7064 3460
rect 7656 3408 7708 3460
rect 7748 3408 7800 3460
rect 8668 3408 8720 3460
rect 11704 3408 11756 3460
rect 13728 3544 13780 3596
rect 13268 3476 13320 3528
rect 13544 3519 13596 3528
rect 13544 3485 13553 3519
rect 13553 3485 13587 3519
rect 13587 3485 13596 3519
rect 13544 3476 13596 3485
rect 13912 3476 13964 3528
rect 15292 3519 15344 3528
rect 15292 3485 15301 3519
rect 15301 3485 15335 3519
rect 15335 3485 15344 3519
rect 15292 3476 15344 3485
rect 15568 3476 15620 3528
rect 2964 3340 3016 3392
rect 3240 3340 3292 3392
rect 4528 3340 4580 3392
rect 5448 3340 5500 3392
rect 5908 3340 5960 3392
rect 6184 3340 6236 3392
rect 6828 3340 6880 3392
rect 6920 3340 6972 3392
rect 7472 3340 7524 3392
rect 9036 3340 9088 3392
rect 9220 3383 9272 3392
rect 9220 3349 9229 3383
rect 9229 3349 9263 3383
rect 9263 3349 9272 3383
rect 9220 3340 9272 3349
rect 9772 3383 9824 3392
rect 9772 3349 9781 3383
rect 9781 3349 9815 3383
rect 9815 3349 9824 3383
rect 9772 3340 9824 3349
rect 10508 3340 10560 3392
rect 10600 3383 10652 3392
rect 10600 3349 10609 3383
rect 10609 3349 10643 3383
rect 10643 3349 10652 3383
rect 10600 3340 10652 3349
rect 10784 3340 10836 3392
rect 11244 3340 11296 3392
rect 11428 3383 11480 3392
rect 11428 3349 11437 3383
rect 11437 3349 11471 3383
rect 11471 3349 11480 3383
rect 11428 3340 11480 3349
rect 11520 3340 11572 3392
rect 11980 3340 12032 3392
rect 13084 3340 13136 3392
rect 14648 3408 14700 3460
rect 13268 3340 13320 3392
rect 13544 3340 13596 3392
rect 15108 3383 15160 3392
rect 15108 3349 15117 3383
rect 15117 3349 15151 3383
rect 15151 3349 15160 3383
rect 15108 3340 15160 3349
rect 4698 3238 4750 3290
rect 4762 3238 4814 3290
rect 4826 3238 4878 3290
rect 4890 3238 4942 3290
rect 4954 3238 5006 3290
rect 8446 3238 8498 3290
rect 8510 3238 8562 3290
rect 8574 3238 8626 3290
rect 8638 3238 8690 3290
rect 8702 3238 8754 3290
rect 12194 3238 12246 3290
rect 12258 3238 12310 3290
rect 12322 3238 12374 3290
rect 12386 3238 12438 3290
rect 12450 3238 12502 3290
rect 1676 3136 1728 3188
rect 2596 3136 2648 3188
rect 6184 3136 6236 3188
rect 6368 3179 6420 3188
rect 6368 3145 6377 3179
rect 6377 3145 6411 3179
rect 6411 3145 6420 3179
rect 6368 3136 6420 3145
rect 7472 3179 7524 3188
rect 3148 3068 3200 3120
rect 3792 3068 3844 3120
rect 4160 3068 4212 3120
rect 1860 3043 1912 3052
rect 1860 3009 1869 3043
rect 1869 3009 1903 3043
rect 1903 3009 1912 3043
rect 1860 3000 1912 3009
rect 2136 3000 2188 3052
rect 2596 3000 2648 3052
rect 2688 3000 2740 3052
rect 2044 2975 2096 2984
rect 2044 2941 2053 2975
rect 2053 2941 2087 2975
rect 2087 2941 2096 2975
rect 2044 2932 2096 2941
rect 3332 3000 3384 3052
rect 5448 3068 5500 3120
rect 5908 3068 5960 3120
rect 6460 3068 6512 3120
rect 7472 3145 7481 3179
rect 7481 3145 7515 3179
rect 7515 3145 7524 3179
rect 7472 3136 7524 3145
rect 7564 3179 7616 3188
rect 7564 3145 7573 3179
rect 7573 3145 7607 3179
rect 7607 3145 7616 3179
rect 7564 3136 7616 3145
rect 8944 3111 8996 3120
rect 8944 3077 8953 3111
rect 8953 3077 8987 3111
rect 8987 3077 8996 3111
rect 8944 3068 8996 3077
rect 4620 3000 4672 3052
rect 4988 3043 5040 3052
rect 4988 3009 4997 3043
rect 4997 3009 5031 3043
rect 5031 3009 5040 3043
rect 5816 3043 5868 3052
rect 4988 3000 5040 3009
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 8668 3000 8720 3052
rect 9404 3111 9456 3120
rect 9404 3077 9413 3111
rect 9413 3077 9447 3111
rect 9447 3077 9456 3111
rect 10232 3111 10284 3120
rect 9404 3068 9456 3077
rect 10232 3077 10241 3111
rect 10241 3077 10275 3111
rect 10275 3077 10284 3111
rect 10232 3068 10284 3077
rect 4712 2975 4764 2984
rect 664 2796 716 2848
rect 4712 2941 4721 2975
rect 4721 2941 4755 2975
rect 4755 2941 4764 2975
rect 4712 2932 4764 2941
rect 6092 2932 6144 2984
rect 6368 2932 6420 2984
rect 6920 2975 6972 2984
rect 6920 2941 6929 2975
rect 6929 2941 6963 2975
rect 6963 2941 6972 2975
rect 6920 2932 6972 2941
rect 7196 2932 7248 2984
rect 2320 2796 2372 2848
rect 5632 2864 5684 2916
rect 6552 2864 6604 2916
rect 6736 2864 6788 2916
rect 8760 2907 8812 2916
rect 8760 2873 8769 2907
rect 8769 2873 8803 2907
rect 8803 2873 8812 2907
rect 8760 2864 8812 2873
rect 10324 3000 10376 3052
rect 11060 3136 11112 3188
rect 11796 3136 11848 3188
rect 11980 3136 12032 3188
rect 13176 3136 13228 3188
rect 13268 3136 13320 3188
rect 14464 3136 14516 3188
rect 10784 3000 10836 3052
rect 11060 3000 11112 3052
rect 12164 3068 12216 3120
rect 12256 3068 12308 3120
rect 12624 3068 12676 3120
rect 10600 2932 10652 2984
rect 10692 2932 10744 2984
rect 11704 2932 11756 2984
rect 12808 3000 12860 3052
rect 13452 3000 13504 3052
rect 15200 3136 15252 3188
rect 15384 3136 15436 3188
rect 16672 3136 16724 3188
rect 16948 3068 17000 3120
rect 12256 2932 12308 2984
rect 9496 2864 9548 2916
rect 10048 2796 10100 2848
rect 10968 2796 11020 2848
rect 13636 2932 13688 2984
rect 13820 2932 13872 2984
rect 14464 2932 14516 2984
rect 14832 3000 14884 3052
rect 15844 3000 15896 3052
rect 15384 2932 15436 2984
rect 16580 2932 16632 2984
rect 13176 2864 13228 2916
rect 13452 2864 13504 2916
rect 15936 2864 15988 2916
rect 13084 2839 13136 2848
rect 13084 2805 13093 2839
rect 13093 2805 13127 2839
rect 13127 2805 13136 2839
rect 13084 2796 13136 2805
rect 14464 2796 14516 2848
rect 2824 2694 2876 2746
rect 2888 2694 2940 2746
rect 2952 2694 3004 2746
rect 3016 2694 3068 2746
rect 3080 2694 3132 2746
rect 6572 2694 6624 2746
rect 6636 2694 6688 2746
rect 6700 2694 6752 2746
rect 6764 2694 6816 2746
rect 6828 2694 6880 2746
rect 10320 2694 10372 2746
rect 10384 2694 10436 2746
rect 10448 2694 10500 2746
rect 10512 2694 10564 2746
rect 10576 2694 10628 2746
rect 14068 2694 14120 2746
rect 14132 2694 14184 2746
rect 14196 2694 14248 2746
rect 14260 2694 14312 2746
rect 14324 2694 14376 2746
rect 1492 2592 1544 2644
rect 4252 2592 4304 2644
rect 4528 2635 4580 2644
rect 4528 2601 4537 2635
rect 4537 2601 4571 2635
rect 4571 2601 4580 2635
rect 4528 2592 4580 2601
rect 3148 2524 3200 2576
rect 1952 2456 2004 2508
rect 2320 2499 2372 2508
rect 2320 2465 2329 2499
rect 2329 2465 2363 2499
rect 2363 2465 2372 2499
rect 2320 2456 2372 2465
rect 2688 2456 2740 2508
rect 4344 2524 4396 2576
rect 4068 2499 4120 2508
rect 4068 2465 4077 2499
rect 4077 2465 4111 2499
rect 4111 2465 4120 2499
rect 4068 2456 4120 2465
rect 5080 2456 5132 2508
rect 3148 2388 3200 2440
rect 3792 2388 3844 2440
rect 2044 2320 2096 2372
rect 2596 2320 2648 2372
rect 3056 2252 3108 2304
rect 3516 2252 3568 2304
rect 4896 2388 4948 2440
rect 4528 2320 4580 2372
rect 6920 2592 6972 2644
rect 8760 2592 8812 2644
rect 8944 2592 8996 2644
rect 9036 2592 9088 2644
rect 5908 2499 5960 2508
rect 5908 2465 5917 2499
rect 5917 2465 5951 2499
rect 5951 2465 5960 2499
rect 5908 2456 5960 2465
rect 6828 2524 6880 2576
rect 6092 2456 6144 2508
rect 7104 2456 7156 2508
rect 5448 2388 5500 2440
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 6920 2388 6972 2440
rect 7748 2456 7800 2508
rect 8300 2456 8352 2508
rect 8484 2456 8536 2508
rect 8760 2456 8812 2508
rect 9312 2592 9364 2644
rect 9404 2592 9456 2644
rect 10048 2592 10100 2644
rect 7932 2388 7984 2440
rect 8484 2320 8536 2372
rect 8668 2320 8720 2372
rect 4344 2252 4396 2304
rect 6460 2252 6512 2304
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 7104 2252 7156 2261
rect 7564 2295 7616 2304
rect 7564 2261 7573 2295
rect 7573 2261 7607 2295
rect 7607 2261 7616 2295
rect 7564 2252 7616 2261
rect 7932 2295 7984 2304
rect 7932 2261 7941 2295
rect 7941 2261 7975 2295
rect 7975 2261 7984 2295
rect 7932 2252 7984 2261
rect 8300 2295 8352 2304
rect 8300 2261 8309 2295
rect 8309 2261 8343 2295
rect 8343 2261 8352 2295
rect 8300 2252 8352 2261
rect 8944 2320 8996 2372
rect 10968 2524 11020 2576
rect 11796 2524 11848 2576
rect 12716 2592 12768 2644
rect 13912 2635 13964 2644
rect 13912 2601 13921 2635
rect 13921 2601 13955 2635
rect 13955 2601 13964 2635
rect 13912 2592 13964 2601
rect 9956 2499 10008 2508
rect 9956 2465 9965 2499
rect 9965 2465 9999 2499
rect 9999 2465 10008 2499
rect 9956 2456 10008 2465
rect 10048 2499 10100 2508
rect 10048 2465 10057 2499
rect 10057 2465 10091 2499
rect 10091 2465 10100 2499
rect 11060 2499 11112 2508
rect 10048 2456 10100 2465
rect 11060 2465 11069 2499
rect 11069 2465 11103 2499
rect 11103 2465 11112 2499
rect 11060 2456 11112 2465
rect 10232 2388 10284 2440
rect 11336 2456 11388 2508
rect 12900 2499 12952 2508
rect 12900 2465 12909 2499
rect 12909 2465 12943 2499
rect 12943 2465 12952 2499
rect 12900 2456 12952 2465
rect 13268 2499 13320 2508
rect 13268 2465 13277 2499
rect 13277 2465 13311 2499
rect 13311 2465 13320 2499
rect 13268 2456 13320 2465
rect 14096 2524 14148 2576
rect 11244 2388 11296 2440
rect 11520 2388 11572 2440
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 11888 2388 11940 2397
rect 12532 2388 12584 2440
rect 13084 2388 13136 2440
rect 15660 2524 15712 2576
rect 15568 2456 15620 2508
rect 9680 2320 9732 2372
rect 9864 2320 9916 2372
rect 10324 2320 10376 2372
rect 9128 2252 9180 2304
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 10416 2252 10468 2304
rect 10600 2295 10652 2304
rect 10600 2261 10609 2295
rect 10609 2261 10643 2295
rect 10643 2261 10652 2295
rect 10968 2295 11020 2304
rect 10600 2252 10652 2261
rect 10968 2261 10977 2295
rect 10977 2261 11011 2295
rect 11011 2261 11020 2295
rect 10968 2252 11020 2261
rect 11520 2295 11572 2304
rect 11520 2261 11529 2295
rect 11529 2261 11563 2295
rect 11563 2261 11572 2295
rect 11520 2252 11572 2261
rect 12624 2320 12676 2372
rect 14280 2320 14332 2372
rect 14740 2320 14792 2372
rect 15752 2388 15804 2440
rect 15936 2320 15988 2372
rect 12808 2252 12860 2304
rect 16488 2252 16540 2304
rect 4698 2150 4750 2202
rect 4762 2150 4814 2202
rect 4826 2150 4878 2202
rect 4890 2150 4942 2202
rect 4954 2150 5006 2202
rect 8446 2150 8498 2202
rect 8510 2150 8562 2202
rect 8574 2150 8626 2202
rect 8638 2150 8690 2202
rect 8702 2150 8754 2202
rect 12194 2150 12246 2202
rect 12258 2150 12310 2202
rect 12322 2150 12374 2202
rect 12386 2150 12438 2202
rect 12450 2150 12502 2202
rect 3056 2048 3108 2100
rect 10968 2048 11020 2100
rect 11152 2048 11204 2100
rect 12072 2048 12124 2100
rect 12624 2048 12676 2100
rect 15016 2048 15068 2100
rect 3148 1980 3200 2032
rect 6828 1980 6880 2032
rect 4436 1912 4488 1964
rect 7104 1912 7156 1964
rect 4068 1776 4120 1828
rect 6920 1776 6972 1828
rect 8852 1980 8904 2032
rect 11612 1980 11664 2032
rect 8300 1912 8352 1964
rect 11428 1912 11480 1964
rect 11520 1912 11572 1964
rect 13268 1912 13320 1964
rect 9680 1844 9732 1896
rect 9772 1844 9824 1896
rect 10048 1844 10100 1896
rect 14924 1844 14976 1896
rect 11704 1776 11756 1828
rect 6368 1708 6420 1760
rect 7656 1708 7708 1760
rect 7748 1708 7800 1760
rect 11060 1708 11112 1760
rect 2228 1640 2280 1692
rect 7564 1640 7616 1692
rect 11428 1640 11480 1692
rect 10508 1572 10560 1624
rect 10692 1572 10744 1624
rect 13728 1572 13780 1624
rect 4528 1504 4580 1556
rect 8944 1504 8996 1556
rect 9036 1504 9088 1556
rect 9680 1504 9732 1556
rect 10140 1504 10192 1556
rect 16304 1504 16356 1556
rect 5356 1436 5408 1488
rect 10600 1436 10652 1488
rect 10784 1436 10836 1488
rect 13452 1436 13504 1488
rect 2780 1368 2832 1420
rect 3424 1368 3476 1420
rect 3608 1368 3660 1420
rect 8024 1368 8076 1420
rect 8116 1368 8168 1420
rect 8668 1368 8720 1420
rect 6828 1300 6880 1352
rect 11796 1300 11848 1352
rect 3516 1232 3568 1284
rect 14648 1232 14700 1284
rect 6184 1164 6236 1216
rect 11244 1164 11296 1216
rect 3976 1096 4028 1148
rect 14464 1164 14516 1216
rect 11520 1096 11572 1148
rect 13084 1096 13136 1148
rect 5908 1028 5960 1080
rect 6828 1028 6880 1080
rect 7380 1028 7432 1080
rect 10692 1028 10744 1080
rect 112 960 164 1012
rect 15108 960 15160 1012
rect 6092 892 6144 944
rect 10232 892 10284 944
rect 3608 824 3660 876
rect 12992 824 13044 876
rect 5632 756 5684 808
rect 10876 756 10928 808
rect 3700 688 3752 740
rect 11520 688 11572 740
rect 6828 212 6880 264
rect 9772 212 9824 264
rect 4436 144 4488 196
rect 15384 144 15436 196
rect 1860 76 1912 128
rect 14372 76 14424 128
rect 848 8 900 60
rect 13636 8 13688 60
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 938 19200 994 20000
rect 1306 19200 1362 20000
rect 1674 19200 1730 20000
rect 2042 19200 2098 20000
rect 2410 19200 2466 20000
rect 2778 19200 2834 20000
rect 2884 19230 3096 19258
rect 216 15745 244 19200
rect 584 15881 612 19200
rect 952 17270 980 19200
rect 1320 17898 1348 19200
rect 1398 17912 1454 17921
rect 1320 17870 1398 17898
rect 1398 17847 1454 17856
rect 940 17264 992 17270
rect 940 17206 992 17212
rect 1584 16788 1636 16794
rect 1584 16730 1636 16736
rect 1032 15904 1084 15910
rect 570 15872 626 15881
rect 1032 15846 1084 15852
rect 570 15807 626 15816
rect 202 15736 258 15745
rect 202 15671 258 15680
rect 756 15088 808 15094
rect 756 15030 808 15036
rect 664 12096 716 12102
rect 664 12038 716 12044
rect 676 2854 704 12038
rect 768 4486 796 15030
rect 848 14544 900 14550
rect 848 14486 900 14492
rect 860 6798 888 14486
rect 940 14272 992 14278
rect 940 14214 992 14220
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 756 4480 808 4486
rect 756 4422 808 4428
rect 952 3534 980 14214
rect 1044 7993 1072 15846
rect 1490 15600 1546 15609
rect 1490 15535 1546 15544
rect 1124 14816 1176 14822
rect 1124 14758 1176 14764
rect 1136 12102 1164 14758
rect 1216 14612 1268 14618
rect 1216 14554 1268 14560
rect 1124 12096 1176 12102
rect 1124 12038 1176 12044
rect 1124 11892 1176 11898
rect 1124 11834 1176 11840
rect 1136 8974 1164 11834
rect 1124 8968 1176 8974
rect 1124 8910 1176 8916
rect 1030 7984 1086 7993
rect 1030 7919 1086 7928
rect 1136 4282 1164 8910
rect 1124 4276 1176 4282
rect 1124 4218 1176 4224
rect 940 3528 992 3534
rect 940 3470 992 3476
rect 664 2848 716 2854
rect 664 2790 716 2796
rect 1228 2145 1256 14554
rect 1504 14074 1532 15535
rect 1596 14657 1624 16730
rect 1688 15910 1716 19200
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1768 16720 1820 16726
rect 1768 16662 1820 16668
rect 1676 15904 1728 15910
rect 1676 15846 1728 15852
rect 1582 14648 1638 14657
rect 1582 14583 1638 14592
rect 1674 14376 1730 14385
rect 1674 14311 1730 14320
rect 1492 14068 1544 14074
rect 1492 14010 1544 14016
rect 1306 13968 1362 13977
rect 1306 13903 1362 13912
rect 1320 11898 1348 13903
rect 1400 13864 1452 13870
rect 1400 13806 1452 13812
rect 1308 11892 1360 11898
rect 1308 11834 1360 11840
rect 1306 11792 1362 11801
rect 1306 11727 1362 11736
rect 1320 5098 1348 11727
rect 1412 9489 1440 13806
rect 1398 9480 1454 9489
rect 1398 9415 1454 9424
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1308 5092 1360 5098
rect 1308 5034 1360 5040
rect 1214 2136 1270 2145
rect 1214 2071 1270 2080
rect 386 1048 442 1057
rect 112 1012 164 1018
rect 386 983 442 992
rect 112 954 164 960
rect 124 800 152 954
rect 400 800 428 983
rect 768 870 888 898
rect 768 800 796 870
rect 110 0 166 800
rect 386 0 442 800
rect 754 0 810 800
rect 860 66 888 870
rect 1136 870 1256 898
rect 1136 800 1164 870
rect 848 60 900 66
rect 848 2 900 8
rect 1122 0 1178 800
rect 1228 105 1256 870
rect 1412 800 1440 8298
rect 1504 7410 1532 14010
rect 1582 13424 1638 13433
rect 1688 13394 1716 14311
rect 1582 13359 1638 13368
rect 1676 13388 1728 13394
rect 1596 12306 1624 13359
rect 1676 13330 1728 13336
rect 1780 12986 1808 16662
rect 1964 14521 1992 16934
rect 2056 16182 2084 19200
rect 2134 16552 2190 16561
rect 2134 16487 2190 16496
rect 2044 16176 2096 16182
rect 2044 16118 2096 16124
rect 1950 14512 2006 14521
rect 1950 14447 1952 14456
rect 2004 14447 2006 14456
rect 1952 14418 2004 14424
rect 1964 14387 1992 14418
rect 2044 14340 2096 14346
rect 2044 14282 2096 14288
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 1860 13796 1912 13802
rect 1860 13738 1912 13744
rect 1768 12980 1820 12986
rect 1768 12922 1820 12928
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1780 12617 1808 12786
rect 1766 12608 1822 12617
rect 1766 12543 1822 12552
rect 1872 12434 1900 13738
rect 1780 12406 1900 12434
rect 1584 12300 1636 12306
rect 1584 12242 1636 12248
rect 1582 11928 1638 11937
rect 1582 11863 1584 11872
rect 1636 11863 1638 11872
rect 1584 11834 1636 11840
rect 1584 11688 1636 11694
rect 1584 11630 1636 11636
rect 1596 11098 1624 11630
rect 1674 11384 1730 11393
rect 1674 11319 1730 11328
rect 1688 11218 1716 11319
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1596 11070 1716 11098
rect 1584 11008 1636 11014
rect 1584 10950 1636 10956
rect 1596 10810 1624 10950
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1584 9988 1636 9994
rect 1584 9930 1636 9936
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1492 6792 1544 6798
rect 1492 6734 1544 6740
rect 1504 2650 1532 6734
rect 1596 4808 1624 9930
rect 1688 9450 1716 11070
rect 1780 10962 1808 12406
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1872 11121 1900 11698
rect 1964 11150 1992 14010
rect 2056 13938 2084 14282
rect 2148 14006 2176 16487
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2226 15464 2282 15473
rect 2226 15399 2282 15408
rect 2240 14482 2268 15399
rect 2228 14476 2280 14482
rect 2228 14418 2280 14424
rect 2136 14000 2188 14006
rect 2136 13942 2188 13948
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 1952 11144 2004 11150
rect 1858 11112 1914 11121
rect 1952 11086 2004 11092
rect 1858 11047 1914 11056
rect 2056 10962 2084 13874
rect 2228 13252 2280 13258
rect 2228 13194 2280 13200
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2148 12889 2176 12922
rect 2134 12880 2190 12889
rect 2134 12815 2190 12824
rect 2134 12744 2190 12753
rect 2134 12679 2190 12688
rect 1780 10934 1900 10962
rect 1768 9920 1820 9926
rect 1768 9862 1820 9868
rect 1676 9444 1728 9450
rect 1676 9386 1728 9392
rect 1674 9072 1730 9081
rect 1674 9007 1676 9016
rect 1728 9007 1730 9016
rect 1676 8978 1728 8984
rect 1780 8242 1808 9862
rect 1872 9674 1900 10934
rect 1964 10934 2084 10962
rect 1964 10130 1992 10934
rect 2148 10810 2176 12679
rect 2240 12481 2268 13194
rect 2332 12986 2360 16390
rect 2424 15638 2452 19200
rect 2792 19122 2820 19200
rect 2884 19122 2912 19230
rect 2792 19094 2912 19122
rect 2594 17776 2650 17785
rect 2594 17711 2650 17720
rect 2504 16040 2556 16046
rect 2504 15982 2556 15988
rect 2412 15632 2464 15638
rect 2412 15574 2464 15580
rect 2516 14550 2544 15982
rect 2504 14544 2556 14550
rect 2504 14486 2556 14492
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2226 12472 2282 12481
rect 2226 12407 2282 12416
rect 2228 12300 2280 12306
rect 2228 12242 2280 12248
rect 2240 12209 2268 12242
rect 2226 12200 2282 12209
rect 2226 12135 2282 12144
rect 2240 11370 2268 12135
rect 2424 11898 2452 13874
rect 2504 12640 2556 12646
rect 2504 12582 2556 12588
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2240 11342 2452 11370
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2240 11121 2268 11154
rect 2226 11112 2282 11121
rect 2226 11047 2282 11056
rect 2320 11076 2372 11082
rect 2320 11018 2372 11024
rect 2136 10804 2188 10810
rect 2056 10764 2136 10792
rect 1952 10124 2004 10130
rect 1952 10066 2004 10072
rect 2056 9926 2084 10764
rect 2136 10746 2188 10752
rect 2134 10568 2190 10577
rect 2134 10503 2190 10512
rect 2148 10198 2176 10503
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 2228 10056 2280 10062
rect 2332 10033 2360 11018
rect 2228 9998 2280 10004
rect 2318 10024 2374 10033
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 1872 9646 1992 9674
rect 1860 9444 1912 9450
rect 1860 9386 1912 9392
rect 1872 8945 1900 9386
rect 1858 8936 1914 8945
rect 1858 8871 1914 8880
rect 1964 8498 1992 9646
rect 2134 9480 2190 9489
rect 2134 9415 2190 9424
rect 2148 9110 2176 9415
rect 2136 9104 2188 9110
rect 2136 9046 2188 9052
rect 2240 9042 2268 9998
rect 2318 9959 2374 9968
rect 2228 9036 2280 9042
rect 2228 8978 2280 8984
rect 1952 8492 2004 8498
rect 2004 8452 2176 8480
rect 1952 8434 2004 8440
rect 1780 8214 2084 8242
rect 1860 8084 1912 8090
rect 1860 8026 1912 8032
rect 1872 7410 1900 8026
rect 1860 7404 1912 7410
rect 1860 7346 1912 7352
rect 1766 6896 1822 6905
rect 1766 6831 1822 6840
rect 1676 6656 1728 6662
rect 1676 6598 1728 6604
rect 1688 5370 1716 6598
rect 1780 6322 1808 6831
rect 1872 6322 1900 7346
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1676 5364 1728 5370
rect 1728 5324 1808 5352
rect 1676 5306 1728 5312
rect 1596 4780 1716 4808
rect 1582 4720 1638 4729
rect 1582 4655 1584 4664
rect 1636 4655 1638 4664
rect 1584 4626 1636 4632
rect 1688 4282 1716 4780
rect 1780 4622 1808 5324
rect 1768 4616 1820 4622
rect 1768 4558 1820 4564
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1676 4276 1728 4282
rect 1596 4236 1676 4264
rect 1596 3176 1624 4236
rect 1676 4218 1728 4224
rect 1674 4040 1730 4049
rect 1674 3975 1730 3984
rect 1688 3466 1716 3975
rect 1780 3942 1808 4422
rect 1872 4146 1900 5510
rect 1860 4140 1912 4146
rect 1860 4082 1912 4088
rect 1768 3936 1820 3942
rect 1768 3878 1820 3884
rect 1872 3602 1900 4082
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 1676 3188 1728 3194
rect 1596 3148 1676 3176
rect 1676 3130 1728 3136
rect 1860 3052 1912 3058
rect 1860 2994 1912 3000
rect 1492 2644 1544 2650
rect 1492 2586 1544 2592
rect 1872 2281 1900 2994
rect 1964 2514 1992 5850
rect 2056 5250 2084 8214
rect 2148 7954 2176 8452
rect 2240 8090 2268 8978
rect 2424 8634 2452 11342
rect 2516 10674 2544 12582
rect 2608 11830 2636 17711
rect 3068 17354 3096 19230
rect 3146 19200 3202 20000
rect 3514 19200 3570 20000
rect 3882 19200 3938 20000
rect 4066 19408 4122 19417
rect 4066 19343 4122 19352
rect 3160 17490 3188 19200
rect 3160 17462 3372 17490
rect 3068 17326 3280 17354
rect 3148 17196 3200 17202
rect 3148 17138 3200 17144
rect 2824 16892 3132 16912
rect 2824 16890 2830 16892
rect 2886 16890 2910 16892
rect 2966 16890 2990 16892
rect 3046 16890 3070 16892
rect 3126 16890 3132 16892
rect 2886 16838 2888 16890
rect 3068 16838 3070 16890
rect 2824 16836 2830 16838
rect 2886 16836 2910 16838
rect 2966 16836 2990 16838
rect 3046 16836 3070 16838
rect 3126 16836 3132 16838
rect 2824 16816 3132 16836
rect 2824 15804 3132 15824
rect 2824 15802 2830 15804
rect 2886 15802 2910 15804
rect 2966 15802 2990 15804
rect 3046 15802 3070 15804
rect 3126 15802 3132 15804
rect 2886 15750 2888 15802
rect 3068 15750 3070 15802
rect 2824 15748 2830 15750
rect 2886 15748 2910 15750
rect 2966 15748 2990 15750
rect 3046 15748 3070 15750
rect 3126 15748 3132 15750
rect 2824 15728 3132 15748
rect 3056 15564 3108 15570
rect 3056 15506 3108 15512
rect 3068 15162 3096 15506
rect 3056 15156 3108 15162
rect 3056 15098 3108 15104
rect 3068 14890 3096 15098
rect 3056 14884 3108 14890
rect 3056 14826 3108 14832
rect 2688 14816 2740 14822
rect 2688 14758 2740 14764
rect 2700 14346 2728 14758
rect 2824 14716 3132 14736
rect 2824 14714 2830 14716
rect 2886 14714 2910 14716
rect 2966 14714 2990 14716
rect 3046 14714 3070 14716
rect 3126 14714 3132 14716
rect 2886 14662 2888 14714
rect 3068 14662 3070 14714
rect 2824 14660 2830 14662
rect 2886 14660 2910 14662
rect 2966 14660 2990 14662
rect 3046 14660 3070 14662
rect 3126 14660 3132 14662
rect 2824 14640 3132 14660
rect 3054 14376 3110 14385
rect 2688 14340 2740 14346
rect 3054 14311 3110 14320
rect 2688 14282 2740 14288
rect 3068 13938 3096 14311
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 2688 13796 2740 13802
rect 2688 13738 2740 13744
rect 2700 13530 2728 13738
rect 2824 13628 3132 13648
rect 2824 13626 2830 13628
rect 2886 13626 2910 13628
rect 2966 13626 2990 13628
rect 3046 13626 3070 13628
rect 3126 13626 3132 13628
rect 2886 13574 2888 13626
rect 3068 13574 3070 13626
rect 2824 13572 2830 13574
rect 2886 13572 2910 13574
rect 2966 13572 2990 13574
rect 3046 13572 3070 13574
rect 3126 13572 3132 13574
rect 2824 13552 3132 13572
rect 2688 13524 2740 13530
rect 3160 13512 3188 17138
rect 3252 15706 3280 17326
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3240 15360 3292 15366
rect 3240 15302 3292 15308
rect 3252 15162 3280 15302
rect 3240 15156 3292 15162
rect 3240 15098 3292 15104
rect 3344 15094 3372 17462
rect 3422 16416 3478 16425
rect 3422 16351 3478 16360
rect 3332 15088 3384 15094
rect 3332 15030 3384 15036
rect 3240 14884 3292 14890
rect 3240 14826 3292 14832
rect 3252 13938 3280 14826
rect 3330 14648 3386 14657
rect 3330 14583 3386 14592
rect 3344 14550 3372 14583
rect 3332 14544 3384 14550
rect 3332 14486 3384 14492
rect 3332 14340 3384 14346
rect 3332 14282 3384 14288
rect 3344 14113 3372 14282
rect 3330 14104 3386 14113
rect 3330 14039 3386 14048
rect 3240 13932 3292 13938
rect 3240 13874 3292 13880
rect 2740 13484 2820 13512
rect 2688 13466 2740 13472
rect 2688 13184 2740 13190
rect 2688 13126 2740 13132
rect 2700 12306 2728 13126
rect 2792 12753 2820 13484
rect 2976 13484 3188 13512
rect 2976 12986 3004 13484
rect 3252 13410 3280 13874
rect 3344 13870 3372 14039
rect 3436 14006 3464 16351
rect 3528 15706 3556 19200
rect 3790 16144 3846 16153
rect 3790 16079 3846 16088
rect 3700 15904 3752 15910
rect 3700 15846 3752 15852
rect 3516 15700 3568 15706
rect 3516 15642 3568 15648
rect 3608 15632 3660 15638
rect 3608 15574 3660 15580
rect 3514 15192 3570 15201
rect 3620 15162 3648 15574
rect 3712 15434 3740 15846
rect 3700 15428 3752 15434
rect 3700 15370 3752 15376
rect 3514 15127 3570 15136
rect 3608 15156 3660 15162
rect 3528 14346 3556 15127
rect 3608 15098 3660 15104
rect 3698 15056 3754 15065
rect 3804 15026 3832 16079
rect 3698 14991 3700 15000
rect 3752 14991 3754 15000
rect 3792 15020 3844 15026
rect 3700 14962 3752 14968
rect 3896 15008 3924 19200
rect 3974 18456 4030 18465
rect 3974 18391 4030 18400
rect 3988 15570 4016 18391
rect 4080 18018 4108 19343
rect 4250 19200 4306 20000
rect 4618 19200 4674 20000
rect 4986 19200 5042 20000
rect 5354 19200 5410 20000
rect 5722 19200 5778 20000
rect 6182 19200 6238 20000
rect 6550 19200 6606 20000
rect 6918 19200 6974 20000
rect 7024 19230 7236 19258
rect 4068 18012 4120 18018
rect 4068 17954 4120 17960
rect 3976 15564 4028 15570
rect 3976 15506 4028 15512
rect 3896 14980 4200 15008
rect 3792 14962 3844 14968
rect 3882 14920 3938 14929
rect 3882 14855 3938 14864
rect 3976 14884 4028 14890
rect 3606 14784 3662 14793
rect 3606 14719 3662 14728
rect 3620 14550 3648 14719
rect 3608 14544 3660 14550
rect 3608 14486 3660 14492
rect 3608 14408 3660 14414
rect 3608 14350 3660 14356
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 3516 14340 3568 14346
rect 3516 14282 3568 14288
rect 3514 14240 3570 14249
rect 3514 14175 3570 14184
rect 3528 14006 3556 14175
rect 3424 14000 3476 14006
rect 3516 14000 3568 14006
rect 3424 13942 3476 13948
rect 3514 13968 3516 13977
rect 3568 13968 3570 13977
rect 3514 13903 3570 13912
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3516 13864 3568 13870
rect 3516 13806 3568 13812
rect 3068 13382 3280 13410
rect 3330 13424 3386 13433
rect 2964 12980 3016 12986
rect 2964 12922 3016 12928
rect 2778 12744 2834 12753
rect 2778 12679 2834 12688
rect 3068 12628 3096 13382
rect 3330 13359 3386 13368
rect 3424 13388 3476 13394
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 3068 12600 3188 12628
rect 2824 12540 3132 12560
rect 2824 12538 2830 12540
rect 2886 12538 2910 12540
rect 2966 12538 2990 12540
rect 3046 12538 3070 12540
rect 3126 12538 3132 12540
rect 2886 12486 2888 12538
rect 3068 12486 3070 12538
rect 2824 12484 2830 12486
rect 2886 12484 2910 12486
rect 2966 12484 2990 12486
rect 3046 12484 3070 12486
rect 3126 12484 3132 12486
rect 2824 12464 3132 12484
rect 2780 12368 2832 12374
rect 2780 12310 2832 12316
rect 2688 12300 2740 12306
rect 2688 12242 2740 12248
rect 2792 12209 2820 12310
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 2778 12200 2834 12209
rect 2778 12135 2834 12144
rect 2686 11928 2742 11937
rect 3068 11898 3096 12242
rect 3160 12186 3188 12600
rect 3252 12442 3280 13262
rect 3344 13190 3372 13359
rect 3424 13330 3476 13336
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3436 12696 3464 13330
rect 3344 12668 3464 12696
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3160 12158 3280 12186
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 2686 11863 2688 11872
rect 2740 11863 2742 11872
rect 3056 11892 3108 11898
rect 2688 11834 2740 11840
rect 3056 11834 3108 11840
rect 2596 11824 2648 11830
rect 2596 11766 2648 11772
rect 2596 11688 2648 11694
rect 2596 11630 2648 11636
rect 2608 11014 2636 11630
rect 2824 11452 3132 11472
rect 2824 11450 2830 11452
rect 2886 11450 2910 11452
rect 2966 11450 2990 11452
rect 3046 11450 3070 11452
rect 3126 11450 3132 11452
rect 2886 11398 2888 11450
rect 3068 11398 3070 11450
rect 2824 11396 2830 11398
rect 2886 11396 2910 11398
rect 2966 11396 2990 11398
rect 3046 11396 3070 11398
rect 3126 11396 3132 11398
rect 2824 11376 3132 11396
rect 2596 11008 2648 11014
rect 2596 10950 2648 10956
rect 2594 10840 2650 10849
rect 2594 10775 2650 10784
rect 2778 10840 2834 10849
rect 2778 10775 2834 10784
rect 2504 10668 2556 10674
rect 2504 10610 2556 10616
rect 2516 9722 2544 10610
rect 2608 10112 2636 10775
rect 2792 10742 2820 10775
rect 2780 10736 2832 10742
rect 2780 10678 2832 10684
rect 3056 10736 3108 10742
rect 3056 10678 3108 10684
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2700 10248 2728 10542
rect 3068 10538 3096 10678
rect 3056 10532 3108 10538
rect 3056 10474 3108 10480
rect 2824 10364 3132 10384
rect 2824 10362 2830 10364
rect 2886 10362 2910 10364
rect 2966 10362 2990 10364
rect 3046 10362 3070 10364
rect 3126 10362 3132 10364
rect 2886 10310 2888 10362
rect 3068 10310 3070 10362
rect 2824 10308 2830 10310
rect 2886 10308 2910 10310
rect 2966 10308 2990 10310
rect 3046 10308 3070 10310
rect 3126 10308 3132 10310
rect 2824 10288 3132 10308
rect 2700 10220 2820 10248
rect 2608 10084 2728 10112
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 2608 9897 2636 9930
rect 2594 9888 2650 9897
rect 2594 9823 2650 9832
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2700 9586 2728 10084
rect 2792 9994 2820 10220
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2962 9616 3018 9625
rect 2688 9580 2740 9586
rect 2962 9551 2964 9560
rect 2688 9522 2740 9528
rect 3016 9551 3018 9560
rect 2964 9522 3016 9528
rect 2412 8628 2464 8634
rect 2412 8570 2464 8576
rect 2318 8528 2374 8537
rect 2318 8463 2374 8472
rect 2228 8084 2280 8090
rect 2228 8026 2280 8032
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2148 6322 2176 7482
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2240 6633 2268 7142
rect 2226 6624 2282 6633
rect 2226 6559 2282 6568
rect 2228 6384 2280 6390
rect 2228 6326 2280 6332
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2148 5914 2176 6258
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2134 5536 2190 5545
rect 2134 5471 2190 5480
rect 2148 5370 2176 5471
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2056 5222 2176 5250
rect 2240 5234 2268 6326
rect 2332 5681 2360 8463
rect 2596 8288 2648 8294
rect 2596 8230 2648 8236
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2410 6760 2466 6769
rect 2410 6695 2466 6704
rect 2424 6662 2452 6695
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2318 5672 2374 5681
rect 2318 5607 2374 5616
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 2056 2990 2084 4218
rect 2148 3058 2176 5222
rect 2228 5228 2280 5234
rect 2228 5170 2280 5176
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2240 4826 2268 5170
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2226 4448 2282 4457
rect 2226 4383 2282 4392
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 2134 2816 2190 2825
rect 2134 2751 2190 2760
rect 2042 2544 2098 2553
rect 1952 2508 2004 2514
rect 2042 2479 2098 2488
rect 1952 2450 2004 2456
rect 1858 2272 1914 2281
rect 1858 2207 1914 2216
rect 1964 1737 1992 2450
rect 2056 2378 2084 2479
rect 2044 2372 2096 2378
rect 2044 2314 2096 2320
rect 1950 1728 2006 1737
rect 1950 1663 2006 1672
rect 1780 870 1900 898
rect 1780 800 1808 870
rect 1214 96 1270 105
rect 1214 31 1270 40
rect 1398 0 1454 800
rect 1766 0 1822 800
rect 1872 134 1900 870
rect 2148 800 2176 2751
rect 2240 1698 2268 4383
rect 2332 4282 2360 5170
rect 2424 4622 2452 6598
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2516 4457 2544 7346
rect 2608 6866 2636 8230
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2594 6624 2650 6633
rect 2594 6559 2650 6568
rect 2502 4448 2558 4457
rect 2502 4383 2558 4392
rect 2320 4276 2372 4282
rect 2320 4218 2372 4224
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 2424 3466 2452 4150
rect 2608 3618 2636 6559
rect 2700 4282 2728 9522
rect 2824 9276 3132 9296
rect 2824 9274 2830 9276
rect 2886 9274 2910 9276
rect 2966 9274 2990 9276
rect 3046 9274 3070 9276
rect 3126 9274 3132 9276
rect 2886 9222 2888 9274
rect 3068 9222 3070 9274
rect 2824 9220 2830 9222
rect 2886 9220 2910 9222
rect 2966 9220 2990 9222
rect 3046 9220 3070 9222
rect 3126 9220 3132 9222
rect 2824 9200 3132 9220
rect 3160 8906 3188 12038
rect 3252 10062 3280 12158
rect 3344 11393 3372 12668
rect 3424 12300 3476 12306
rect 3424 12242 3476 12248
rect 3330 11384 3386 11393
rect 3330 11319 3386 11328
rect 3332 11212 3384 11218
rect 3332 11154 3384 11160
rect 3344 10810 3372 11154
rect 3332 10804 3384 10810
rect 3332 10746 3384 10752
rect 3330 10704 3386 10713
rect 3330 10639 3386 10648
rect 3344 10538 3372 10639
rect 3332 10532 3384 10538
rect 3332 10474 3384 10480
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 3436 9994 3464 12242
rect 3528 11354 3556 13806
rect 3620 13530 3648 14350
rect 3700 14340 3752 14346
rect 3700 14282 3752 14288
rect 3608 13524 3660 13530
rect 3608 13466 3660 13472
rect 3606 13288 3662 13297
rect 3606 13223 3662 13232
rect 3620 12102 3648 13223
rect 3712 12481 3740 14282
rect 3804 13841 3832 14350
rect 3896 14249 3924 14855
rect 3976 14826 4028 14832
rect 3882 14240 3938 14249
rect 3882 14175 3938 14184
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 3790 13832 3846 13841
rect 3790 13767 3846 13776
rect 3790 13696 3846 13705
rect 3790 13631 3846 13640
rect 3804 13394 3832 13631
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 3792 12980 3844 12986
rect 3792 12922 3844 12928
rect 3698 12472 3754 12481
rect 3698 12407 3754 12416
rect 3698 12336 3754 12345
rect 3698 12271 3754 12280
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3514 11248 3570 11257
rect 3514 11183 3570 11192
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3148 8900 3200 8906
rect 3148 8842 3200 8848
rect 2824 8188 3132 8208
rect 2824 8186 2830 8188
rect 2886 8186 2910 8188
rect 2966 8186 2990 8188
rect 3046 8186 3070 8188
rect 3126 8186 3132 8188
rect 2886 8134 2888 8186
rect 3068 8134 3070 8186
rect 2824 8132 2830 8134
rect 2886 8132 2910 8134
rect 2966 8132 2990 8134
rect 3046 8132 3070 8134
rect 3126 8132 3132 8134
rect 2824 8112 3132 8132
rect 3146 7440 3202 7449
rect 3146 7375 3202 7384
rect 3054 7304 3110 7313
rect 3054 7239 3056 7248
rect 3108 7239 3110 7248
rect 3056 7210 3108 7216
rect 2824 7100 3132 7120
rect 2824 7098 2830 7100
rect 2886 7098 2910 7100
rect 2966 7098 2990 7100
rect 3046 7098 3070 7100
rect 3126 7098 3132 7100
rect 2886 7046 2888 7098
rect 3068 7046 3070 7098
rect 2824 7044 2830 7046
rect 2886 7044 2910 7046
rect 2966 7044 2990 7046
rect 3046 7044 3070 7046
rect 3126 7044 3132 7046
rect 2824 7024 3132 7044
rect 2824 6012 3132 6032
rect 2824 6010 2830 6012
rect 2886 6010 2910 6012
rect 2966 6010 2990 6012
rect 3046 6010 3070 6012
rect 3126 6010 3132 6012
rect 2886 5958 2888 6010
rect 3068 5958 3070 6010
rect 2824 5956 2830 5958
rect 2886 5956 2910 5958
rect 2966 5956 2990 5958
rect 3046 5956 3070 5958
rect 3126 5956 3132 5958
rect 2824 5936 3132 5956
rect 2824 4924 3132 4944
rect 2824 4922 2830 4924
rect 2886 4922 2910 4924
rect 2966 4922 2990 4924
rect 3046 4922 3070 4924
rect 3126 4922 3132 4924
rect 2886 4870 2888 4922
rect 3068 4870 3070 4922
rect 2824 4868 2830 4870
rect 2886 4868 2910 4870
rect 2966 4868 2990 4870
rect 3046 4868 3070 4870
rect 3126 4868 3132 4870
rect 2824 4848 3132 4868
rect 2962 4720 3018 4729
rect 2962 4655 3018 4664
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2976 4146 3004 4655
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 2824 3836 3132 3856
rect 2824 3834 2830 3836
rect 2886 3834 2910 3836
rect 2966 3834 2990 3836
rect 3046 3834 3070 3836
rect 3126 3834 3132 3836
rect 2886 3782 2888 3834
rect 3068 3782 3070 3834
rect 2824 3780 2830 3782
rect 2886 3780 2910 3782
rect 2966 3780 2990 3782
rect 3046 3780 3070 3782
rect 3126 3780 3132 3782
rect 2824 3760 3132 3780
rect 2516 3590 2636 3618
rect 2964 3664 3016 3670
rect 2964 3606 3016 3612
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 2320 3460 2372 3466
rect 2320 3402 2372 3408
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 2332 2961 2360 3402
rect 2318 2952 2374 2961
rect 2318 2887 2374 2896
rect 2320 2848 2372 2854
rect 2318 2816 2320 2825
rect 2372 2816 2374 2825
rect 2318 2751 2374 2760
rect 2318 2544 2374 2553
rect 2318 2479 2320 2488
rect 2372 2479 2374 2488
rect 2320 2450 2372 2456
rect 2228 1692 2280 1698
rect 2228 1634 2280 1640
rect 2516 800 2544 3590
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2594 3360 2650 3369
rect 2594 3295 2650 3304
rect 2608 3194 2636 3295
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2700 3058 2728 3470
rect 2976 3398 3004 3606
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2778 3224 2834 3233
rect 2778 3159 2834 3168
rect 2596 3052 2648 3058
rect 2596 2994 2648 3000
rect 2688 3052 2740 3058
rect 2688 2994 2740 3000
rect 2608 2378 2636 2994
rect 2792 2836 2820 3159
rect 3068 2972 3096 3606
rect 3160 3126 3188 7375
rect 3252 5234 3280 9862
rect 3528 9674 3556 11183
rect 3344 9646 3556 9674
rect 3344 8634 3372 9646
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 3344 7206 3372 8570
rect 3436 8294 3464 9522
rect 3516 9172 3568 9178
rect 3620 9160 3648 11630
rect 3568 9132 3648 9160
rect 3516 9114 3568 9120
rect 3712 9058 3740 12271
rect 3804 12238 3832 12922
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3896 11898 3924 14010
rect 3988 12306 4016 14826
rect 4172 14550 4200 14980
rect 4160 14544 4212 14550
rect 4160 14486 4212 14492
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 4080 11830 4108 14418
rect 4264 14346 4292 19200
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4356 15366 4384 15438
rect 4436 15428 4488 15434
rect 4436 15370 4488 15376
rect 4528 15428 4580 15434
rect 4528 15370 4580 15376
rect 4344 15360 4396 15366
rect 4344 15302 4396 15308
rect 4344 15088 4396 15094
rect 4344 15030 4396 15036
rect 4356 14414 4384 15030
rect 4448 14958 4476 15370
rect 4540 15162 4568 15370
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4436 14952 4488 14958
rect 4436 14894 4488 14900
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 4252 14340 4304 14346
rect 4252 14282 4304 14288
rect 4160 14272 4212 14278
rect 4158 14240 4160 14249
rect 4212 14240 4214 14249
rect 4158 14175 4214 14184
rect 4160 14000 4212 14006
rect 4158 13968 4160 13977
rect 4212 13968 4214 13977
rect 4158 13903 4214 13912
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 4158 13560 4214 13569
rect 4158 13495 4214 13504
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 3804 9178 3832 11154
rect 3882 11112 3938 11121
rect 3882 11047 3938 11056
rect 3896 10674 3924 11047
rect 3988 10713 4016 11698
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4080 11529 4108 11630
rect 4172 11558 4200 13495
rect 4252 12708 4304 12714
rect 4252 12650 4304 12656
rect 4160 11552 4212 11558
rect 4066 11520 4122 11529
rect 4160 11494 4212 11500
rect 4066 11455 4122 11464
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 3974 10704 4030 10713
rect 3884 10668 3936 10674
rect 3974 10639 4030 10648
rect 3884 10610 3936 10616
rect 3974 10160 4030 10169
rect 3974 10095 4030 10104
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 9217 3924 9862
rect 3882 9208 3938 9217
rect 3792 9172 3844 9178
rect 3882 9143 3938 9152
rect 3792 9114 3844 9120
rect 3528 9030 3740 9058
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3424 7744 3476 7750
rect 3424 7686 3476 7692
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3330 6488 3386 6497
rect 3330 6423 3386 6432
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3240 4480 3292 4486
rect 3238 4448 3240 4457
rect 3292 4448 3294 4457
rect 3238 4383 3294 4392
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3252 3641 3280 4218
rect 3344 3670 3372 6423
rect 3332 3664 3384 3670
rect 3238 3632 3294 3641
rect 3332 3606 3384 3612
rect 3238 3567 3294 3576
rect 3252 3516 3280 3567
rect 3332 3528 3384 3534
rect 3252 3488 3332 3516
rect 3332 3470 3384 3476
rect 3240 3392 3292 3398
rect 3240 3334 3292 3340
rect 3148 3120 3200 3126
rect 3148 3062 3200 3068
rect 3068 2944 3188 2972
rect 2700 2808 2820 2836
rect 2700 2514 2728 2808
rect 2824 2748 3132 2768
rect 2824 2746 2830 2748
rect 2886 2746 2910 2748
rect 2966 2746 2990 2748
rect 3046 2746 3070 2748
rect 3126 2746 3132 2748
rect 2886 2694 2888 2746
rect 3068 2694 3070 2746
rect 2824 2692 2830 2694
rect 2886 2692 2910 2694
rect 2966 2692 2990 2694
rect 3046 2692 3070 2694
rect 3126 2692 3132 2694
rect 2824 2672 3132 2692
rect 3160 2582 3188 2944
rect 3148 2576 3200 2582
rect 3148 2518 3200 2524
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 3068 2106 3096 2246
rect 3056 2100 3108 2106
rect 3056 2042 3108 2048
rect 3160 2038 3188 2382
rect 3148 2032 3200 2038
rect 3148 1974 3200 1980
rect 3252 1442 3280 3334
rect 3332 3052 3384 3058
rect 3332 2994 3384 3000
rect 2780 1420 2832 1426
rect 2780 1362 2832 1368
rect 3160 1414 3280 1442
rect 2792 800 2820 1362
rect 3160 800 3188 1414
rect 1860 128 1912 134
rect 1860 70 1912 76
rect 2134 0 2190 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3344 490 3372 2994
rect 3436 1426 3464 7686
rect 3528 6798 3556 9030
rect 3606 8256 3662 8265
rect 3606 8191 3662 8200
rect 3620 7886 3648 8191
rect 3608 7880 3660 7886
rect 3608 7822 3660 7828
rect 3700 7880 3752 7886
rect 3700 7822 3752 7828
rect 3606 7712 3662 7721
rect 3606 7647 3662 7656
rect 3516 6792 3568 6798
rect 3516 6734 3568 6740
rect 3620 6644 3648 7647
rect 3528 6616 3648 6644
rect 3528 4622 3556 6616
rect 3608 6452 3660 6458
rect 3608 6394 3660 6400
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 3528 2310 3556 3878
rect 3620 3584 3648 6394
rect 3712 5409 3740 7822
rect 3790 7032 3846 7041
rect 3896 7002 3924 9046
rect 3988 9042 4016 10095
rect 4080 9926 4108 11154
rect 4172 10198 4200 11290
rect 4264 11234 4292 12650
rect 4356 11898 4384 13806
rect 4448 13802 4476 14894
rect 4632 14618 4660 19200
rect 5000 17626 5028 19200
rect 5170 18048 5226 18057
rect 5170 17983 5226 17992
rect 5000 17598 5120 17626
rect 4698 17436 5006 17456
rect 4698 17434 4704 17436
rect 4760 17434 4784 17436
rect 4840 17434 4864 17436
rect 4920 17434 4944 17436
rect 5000 17434 5006 17436
rect 4760 17382 4762 17434
rect 4942 17382 4944 17434
rect 4698 17380 4704 17382
rect 4760 17380 4784 17382
rect 4840 17380 4864 17382
rect 4920 17380 4944 17382
rect 5000 17380 5006 17382
rect 4698 17360 5006 17380
rect 4698 16348 5006 16368
rect 4698 16346 4704 16348
rect 4760 16346 4784 16348
rect 4840 16346 4864 16348
rect 4920 16346 4944 16348
rect 5000 16346 5006 16348
rect 4760 16294 4762 16346
rect 4942 16294 4944 16346
rect 4698 16292 4704 16294
rect 4760 16292 4784 16294
rect 4840 16292 4864 16294
rect 4920 16292 4944 16294
rect 5000 16292 5006 16294
rect 4698 16272 5006 16292
rect 4698 15260 5006 15280
rect 4698 15258 4704 15260
rect 4760 15258 4784 15260
rect 4840 15258 4864 15260
rect 4920 15258 4944 15260
rect 5000 15258 5006 15260
rect 4760 15206 4762 15258
rect 4942 15206 4944 15258
rect 4698 15204 4704 15206
rect 4760 15204 4784 15206
rect 4840 15204 4864 15206
rect 4920 15204 4944 15206
rect 5000 15204 5006 15206
rect 4698 15184 5006 15204
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4620 14612 4672 14618
rect 4620 14554 4672 14560
rect 4540 14396 4568 14554
rect 4620 14408 4672 14414
rect 4540 14368 4620 14396
rect 4620 14350 4672 14356
rect 4698 14172 5006 14192
rect 4698 14170 4704 14172
rect 4760 14170 4784 14172
rect 4840 14170 4864 14172
rect 4920 14170 4944 14172
rect 5000 14170 5006 14172
rect 4760 14118 4762 14170
rect 4942 14118 4944 14170
rect 4698 14116 4704 14118
rect 4760 14116 4784 14118
rect 4840 14116 4864 14118
rect 4920 14116 4944 14118
rect 5000 14116 5006 14118
rect 4698 14096 5006 14116
rect 4436 13796 4488 13802
rect 4436 13738 4488 13744
rect 4448 13530 4476 13738
rect 4528 13728 4580 13734
rect 4528 13670 4580 13676
rect 4896 13728 4948 13734
rect 4896 13670 4948 13676
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4436 13388 4488 13394
rect 4436 13330 4488 13336
rect 4344 11892 4396 11898
rect 4344 11834 4396 11840
rect 4356 11354 4384 11834
rect 4344 11348 4396 11354
rect 4344 11290 4396 11296
rect 4264 11206 4384 11234
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4160 10192 4212 10198
rect 4160 10134 4212 10140
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 4172 8498 4200 9522
rect 4264 9382 4292 10950
rect 4356 10470 4384 11206
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4342 10296 4398 10305
rect 4342 10231 4398 10240
rect 4356 10062 4384 10231
rect 4344 10056 4396 10062
rect 4344 9998 4396 10004
rect 4344 9716 4396 9722
rect 4344 9658 4396 9664
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4252 9172 4304 9178
rect 4252 9114 4304 9120
rect 4264 8838 4292 9114
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3974 8392 4030 8401
rect 3974 8327 4030 8336
rect 3790 6967 3846 6976
rect 3884 6996 3936 7002
rect 3804 5846 3832 6967
rect 3884 6938 3936 6944
rect 3988 6866 4016 8327
rect 4068 7880 4120 7886
rect 4068 7822 4120 7828
rect 3976 6860 4028 6866
rect 3976 6802 4028 6808
rect 4080 6202 4108 7822
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 4172 6798 4200 7414
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4172 6390 4200 6734
rect 4160 6384 4212 6390
rect 4160 6326 4212 6332
rect 3896 6174 4108 6202
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3698 5400 3754 5409
rect 3698 5335 3754 5344
rect 3792 5296 3844 5302
rect 3790 5264 3792 5273
rect 3844 5264 3846 5273
rect 3790 5199 3846 5208
rect 3698 5128 3754 5137
rect 3698 5063 3754 5072
rect 3712 3738 3740 5063
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3804 3738 3832 4422
rect 3896 4282 3924 6174
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4172 5794 4200 5850
rect 4080 5766 4200 5794
rect 3884 4276 3936 4282
rect 3884 4218 3936 4224
rect 3700 3732 3752 3738
rect 3700 3674 3752 3680
rect 3792 3732 3844 3738
rect 3792 3674 3844 3680
rect 3620 3556 3924 3584
rect 3606 3496 3662 3505
rect 3606 3431 3662 3440
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3528 1884 3556 2246
rect 3620 1986 3648 3431
rect 3792 3120 3844 3126
rect 3792 3062 3844 3068
rect 3804 2446 3832 3062
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3620 1958 3740 1986
rect 3528 1856 3648 1884
rect 3514 1456 3570 1465
rect 3424 1420 3476 1426
rect 3620 1426 3648 1856
rect 3514 1391 3570 1400
rect 3608 1420 3660 1426
rect 3424 1362 3476 1368
rect 3528 1290 3556 1391
rect 3608 1362 3660 1368
rect 3516 1284 3568 1290
rect 3516 1226 3568 1232
rect 3528 882 3648 898
rect 3528 876 3660 882
rect 3528 870 3608 876
rect 3528 800 3556 870
rect 3608 818 3660 824
rect 3422 504 3478 513
rect 3344 462 3422 490
rect 3422 439 3478 448
rect 3514 0 3570 800
rect 3712 746 3740 1958
rect 3896 800 3924 3556
rect 3974 3360 4030 3369
rect 3974 3295 4030 3304
rect 3988 2496 4016 3295
rect 4080 2774 4108 5766
rect 4356 5370 4384 9658
rect 4448 9586 4476 13330
rect 4540 12238 4568 13670
rect 4908 13394 4936 13670
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4620 13184 4672 13190
rect 4620 13126 4672 13132
rect 4632 12986 4660 13126
rect 4698 13084 5006 13104
rect 4698 13082 4704 13084
rect 4760 13082 4784 13084
rect 4840 13082 4864 13084
rect 4920 13082 4944 13084
rect 5000 13082 5006 13084
rect 4760 13030 4762 13082
rect 4942 13030 4944 13082
rect 4698 13028 4704 13030
rect 4760 13028 4784 13030
rect 4840 13028 4864 13030
rect 4920 13028 4944 13030
rect 5000 13028 5006 13030
rect 4698 13008 5006 13028
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4528 12232 4580 12238
rect 5000 12209 5028 12786
rect 5092 12442 5120 17598
rect 5184 15026 5212 17983
rect 5368 17513 5396 19200
rect 5354 17504 5410 17513
rect 5354 17439 5410 17448
rect 5262 17368 5318 17377
rect 5262 17303 5318 17312
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 5184 14414 5212 14962
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5172 14272 5224 14278
rect 5172 14214 5224 14220
rect 5184 14113 5212 14214
rect 5170 14104 5226 14113
rect 5170 14039 5226 14048
rect 5172 13932 5224 13938
rect 5276 13920 5304 17303
rect 5354 17096 5410 17105
rect 5354 17031 5410 17040
rect 5368 16250 5396 17031
rect 5356 16244 5408 16250
rect 5356 16186 5408 16192
rect 5368 15706 5396 16186
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5356 15700 5408 15706
rect 5356 15642 5408 15648
rect 5368 15570 5396 15642
rect 5552 15570 5580 15982
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5356 15564 5408 15570
rect 5356 15506 5408 15512
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5354 15464 5410 15473
rect 5552 15450 5580 15506
rect 5644 15473 5672 15914
rect 5354 15399 5410 15408
rect 5460 15422 5580 15450
rect 5630 15464 5686 15473
rect 5368 15162 5396 15399
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 5460 15026 5488 15422
rect 5630 15399 5686 15408
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 5552 14958 5580 15302
rect 5630 15192 5686 15201
rect 5736 15162 5764 19200
rect 6196 16590 6224 19200
rect 6368 18012 6420 18018
rect 6368 17954 6420 17960
rect 6184 16584 6236 16590
rect 6184 16526 6236 16532
rect 5816 16040 5868 16046
rect 5816 15982 5868 15988
rect 5630 15127 5686 15136
rect 5724 15156 5776 15162
rect 5356 14952 5408 14958
rect 5356 14894 5408 14900
rect 5540 14952 5592 14958
rect 5540 14894 5592 14900
rect 5368 14822 5396 14894
rect 5356 14816 5408 14822
rect 5356 14758 5408 14764
rect 5448 14544 5500 14550
rect 5224 13892 5304 13920
rect 5368 14504 5448 14532
rect 5172 13874 5224 13880
rect 5368 13841 5396 14504
rect 5448 14486 5500 14492
rect 5552 14414 5580 14894
rect 5644 14793 5672 15127
rect 5724 15098 5776 15104
rect 5630 14784 5686 14793
rect 5630 14719 5686 14728
rect 5828 14657 5856 15982
rect 6090 15736 6146 15745
rect 6090 15671 6146 15680
rect 6000 15496 6052 15502
rect 5906 15464 5962 15473
rect 6000 15438 6052 15444
rect 5906 15399 5962 15408
rect 5814 14648 5870 14657
rect 5814 14583 5870 14592
rect 5724 14544 5776 14550
rect 5724 14486 5776 14492
rect 5540 14408 5592 14414
rect 5538 14376 5540 14385
rect 5592 14376 5594 14385
rect 5538 14311 5594 14320
rect 5632 14340 5684 14346
rect 5632 14282 5684 14288
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 14006 5580 14214
rect 5540 14000 5592 14006
rect 5446 13968 5502 13977
rect 5540 13942 5592 13948
rect 5446 13903 5448 13912
rect 5500 13903 5502 13912
rect 5448 13874 5500 13880
rect 5540 13864 5592 13870
rect 5354 13832 5410 13841
rect 5172 13796 5224 13802
rect 5540 13806 5592 13812
rect 5354 13767 5410 13776
rect 5172 13738 5224 13744
rect 5184 12714 5212 13738
rect 5264 13388 5316 13394
rect 5264 13330 5316 13336
rect 5276 12782 5304 13330
rect 5446 13288 5502 13297
rect 5446 13223 5502 13232
rect 5460 13190 5488 13223
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5448 12844 5500 12850
rect 5448 12786 5500 12792
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5172 12708 5224 12714
rect 5172 12650 5224 12656
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 5080 12232 5132 12238
rect 4528 12174 4580 12180
rect 4986 12200 5042 12209
rect 5080 12174 5132 12180
rect 4986 12135 5042 12144
rect 5092 12073 5120 12174
rect 5078 12064 5134 12073
rect 4698 11996 5006 12016
rect 5276 12050 5304 12718
rect 5078 11999 5134 12008
rect 5184 12022 5304 12050
rect 5354 12064 5410 12073
rect 4698 11994 4704 11996
rect 4760 11994 4784 11996
rect 4840 11994 4864 11996
rect 4920 11994 4944 11996
rect 5000 11994 5006 11996
rect 4760 11942 4762 11994
rect 4942 11942 4944 11994
rect 4698 11940 4704 11942
rect 4760 11940 4784 11942
rect 4840 11940 4864 11942
rect 4920 11940 4944 11942
rect 5000 11940 5006 11942
rect 4698 11920 5006 11940
rect 4620 11756 4672 11762
rect 4672 11716 4844 11744
rect 4620 11698 4672 11704
rect 4528 11620 4580 11626
rect 4528 11562 4580 11568
rect 4540 11082 4568 11562
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4618 11384 4674 11393
rect 4618 11319 4620 11328
rect 4672 11319 4674 11328
rect 4620 11290 4672 11296
rect 4724 11234 4752 11494
rect 4816 11257 4844 11716
rect 5184 11642 5212 12022
rect 5354 11999 5410 12008
rect 5262 11928 5318 11937
rect 5262 11863 5318 11872
rect 5276 11665 5304 11863
rect 4908 11614 5212 11642
rect 5262 11656 5318 11665
rect 4632 11206 4752 11234
rect 4802 11248 4858 11257
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 4632 10962 4660 11206
rect 4802 11183 4858 11192
rect 4908 11082 4936 11614
rect 5262 11591 5318 11600
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5080 11212 5132 11218
rect 5080 11154 5132 11160
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4540 10934 4660 10962
rect 4540 9994 4568 10934
rect 4698 10908 5006 10928
rect 4698 10906 4704 10908
rect 4760 10906 4784 10908
rect 4840 10906 4864 10908
rect 4920 10906 4944 10908
rect 5000 10906 5006 10908
rect 4760 10854 4762 10906
rect 4942 10854 4944 10906
rect 4698 10852 4704 10854
rect 4760 10852 4784 10854
rect 4840 10852 4864 10854
rect 4920 10852 4944 10854
rect 5000 10852 5006 10854
rect 4698 10832 5006 10852
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4816 10470 4844 10610
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4632 10062 4660 10406
rect 4816 10305 4844 10406
rect 4802 10296 4858 10305
rect 4802 10231 4858 10240
rect 4620 10056 4672 10062
rect 4620 9998 4672 10004
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4448 8498 4476 9318
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4540 7546 4568 9930
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4632 9178 4660 9862
rect 4698 9820 5006 9840
rect 4698 9818 4704 9820
rect 4760 9818 4784 9820
rect 4840 9818 4864 9820
rect 4920 9818 4944 9820
rect 5000 9818 5006 9820
rect 4760 9766 4762 9818
rect 4942 9766 4944 9818
rect 4698 9764 4704 9766
rect 4760 9764 4784 9766
rect 4840 9764 4864 9766
rect 4920 9764 4944 9766
rect 5000 9764 5006 9766
rect 4698 9744 5006 9764
rect 5092 9761 5120 11154
rect 5184 10742 5212 11494
rect 5172 10736 5224 10742
rect 5172 10678 5224 10684
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5184 10130 5212 10678
rect 5172 10124 5224 10130
rect 5172 10066 5224 10072
rect 5078 9752 5134 9761
rect 5078 9687 5134 9696
rect 5184 9654 5212 10066
rect 5172 9648 5224 9654
rect 5172 9590 5224 9596
rect 4620 9172 4672 9178
rect 4620 9114 4672 9120
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4698 8732 5006 8752
rect 4698 8730 4704 8732
rect 4760 8730 4784 8732
rect 4840 8730 4864 8732
rect 4920 8730 4944 8732
rect 5000 8730 5006 8732
rect 4760 8678 4762 8730
rect 4942 8678 4944 8730
rect 4698 8676 4704 8678
rect 4760 8676 4784 8678
rect 4840 8676 4864 8678
rect 4920 8676 4944 8678
rect 5000 8676 5006 8678
rect 4698 8656 5006 8676
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4724 8090 4752 8434
rect 4712 8084 4764 8090
rect 4712 8026 4764 8032
rect 4698 7644 5006 7664
rect 4698 7642 4704 7644
rect 4760 7642 4784 7644
rect 4840 7642 4864 7644
rect 4920 7642 4944 7644
rect 5000 7642 5006 7644
rect 4760 7590 4762 7642
rect 4942 7590 4944 7642
rect 4698 7588 4704 7590
rect 4760 7588 4784 7590
rect 4840 7588 4864 7590
rect 4920 7588 4944 7590
rect 5000 7588 5006 7590
rect 4698 7568 5006 7588
rect 5092 7546 5120 8774
rect 5184 8090 5212 9590
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5184 7478 5212 7890
rect 5172 7472 5224 7478
rect 5172 7414 5224 7420
rect 4620 7404 4672 7410
rect 4620 7346 4672 7352
rect 4526 7032 4582 7041
rect 4526 6967 4582 6976
rect 4434 6896 4490 6905
rect 4434 6831 4490 6840
rect 4448 6662 4476 6831
rect 4436 6656 4488 6662
rect 4436 6598 4488 6604
rect 4540 6322 4568 6967
rect 4632 6458 4660 7346
rect 5172 6792 5224 6798
rect 5172 6734 5224 6740
rect 4698 6556 5006 6576
rect 4698 6554 4704 6556
rect 4760 6554 4784 6556
rect 4840 6554 4864 6556
rect 4920 6554 4944 6556
rect 5000 6554 5006 6556
rect 4760 6502 4762 6554
rect 4942 6502 4944 6554
rect 4698 6500 4704 6502
rect 4760 6500 4784 6502
rect 4840 6500 4864 6502
rect 4920 6500 4944 6502
rect 5000 6500 5006 6502
rect 4698 6480 5006 6500
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4528 6316 4580 6322
rect 4448 6276 4528 6304
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4448 5166 4476 6276
rect 4528 6258 4580 6264
rect 4528 6112 4580 6118
rect 4528 6054 4580 6060
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 4158 4176 4214 4185
rect 4158 4111 4214 4120
rect 4172 3126 4200 4111
rect 4264 3233 4292 5034
rect 4436 4820 4488 4826
rect 4356 4780 4436 4808
rect 4250 3224 4306 3233
rect 4250 3159 4306 3168
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4080 2746 4200 2774
rect 4068 2508 4120 2514
rect 3988 2468 4068 2496
rect 4068 2450 4120 2456
rect 3974 2408 4030 2417
rect 3974 2343 4030 2352
rect 3988 1154 4016 2343
rect 4080 1834 4108 2450
rect 4068 1828 4120 1834
rect 4068 1770 4120 1776
rect 3976 1148 4028 1154
rect 3976 1090 4028 1096
rect 4172 800 4200 2746
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4264 2292 4292 2586
rect 4356 2582 4384 4780
rect 4436 4762 4488 4768
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4344 2576 4396 2582
rect 4344 2518 4396 2524
rect 4344 2304 4396 2310
rect 4264 2264 4344 2292
rect 4344 2246 4396 2252
rect 4448 1970 4476 4218
rect 4540 3534 4568 6054
rect 4632 5953 4660 6394
rect 4894 6352 4950 6361
rect 4804 6316 4856 6322
rect 4894 6287 4950 6296
rect 4804 6258 4856 6264
rect 4618 5944 4674 5953
rect 4618 5879 4674 5888
rect 4816 5710 4844 6258
rect 4908 5817 4936 6287
rect 4894 5808 4950 5817
rect 4894 5743 4950 5752
rect 5078 5808 5134 5817
rect 5078 5743 5134 5752
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 5092 5642 5120 5743
rect 5184 5658 5212 6734
rect 5276 6662 5304 10678
rect 5368 7886 5396 11999
rect 5460 11665 5488 12786
rect 5552 12617 5580 13806
rect 5644 13569 5672 14282
rect 5630 13560 5686 13569
rect 5630 13495 5686 13504
rect 5736 13433 5764 14486
rect 5920 14414 5948 15399
rect 6012 14634 6040 15438
rect 6104 15094 6132 15671
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6184 15360 6236 15366
rect 6184 15302 6236 15308
rect 6092 15088 6144 15094
rect 6092 15030 6144 15036
rect 6196 15026 6224 15302
rect 6184 15020 6236 15026
rect 6184 14962 6236 14968
rect 6092 14884 6144 14890
rect 6092 14826 6144 14832
rect 6104 14793 6132 14826
rect 6090 14784 6146 14793
rect 6090 14719 6146 14728
rect 6012 14606 6224 14634
rect 6092 14476 6144 14482
rect 6092 14418 6144 14424
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5920 13705 5948 13874
rect 6012 13841 6040 14214
rect 6104 13954 6132 14418
rect 6196 14278 6224 14606
rect 6184 14272 6236 14278
rect 6184 14214 6236 14220
rect 6104 13926 6224 13954
rect 6092 13864 6144 13870
rect 5998 13832 6054 13841
rect 6196 13841 6224 13926
rect 6288 13852 6316 15438
rect 6380 15162 6408 17954
rect 6564 17082 6592 19200
rect 6932 19122 6960 19200
rect 7024 19122 7052 19230
rect 6932 19094 7052 19122
rect 6472 17054 6592 17082
rect 6368 15156 6420 15162
rect 6368 15098 6420 15104
rect 6380 14006 6408 15098
rect 6368 14000 6420 14006
rect 6368 13942 6420 13948
rect 6092 13806 6144 13812
rect 6182 13832 6238 13841
rect 5998 13767 6054 13776
rect 5906 13696 5962 13705
rect 5906 13631 5962 13640
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 5722 13424 5778 13433
rect 5722 13359 5778 13368
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5538 12608 5594 12617
rect 5538 12543 5594 12552
rect 5632 12368 5684 12374
rect 5538 12336 5594 12345
rect 5632 12310 5684 12316
rect 5538 12271 5594 12280
rect 5446 11656 5502 11665
rect 5446 11591 5502 11600
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 11354 5488 11494
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5460 10198 5488 11018
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5460 9382 5488 10134
rect 5552 9489 5580 12271
rect 5644 12170 5672 12310
rect 5736 12186 5764 12718
rect 5828 12481 5856 13262
rect 5906 13016 5962 13025
rect 6012 12986 6040 13466
rect 5906 12951 5962 12960
rect 6000 12980 6052 12986
rect 5920 12850 5948 12951
rect 6000 12922 6052 12928
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 5908 12708 5960 12714
rect 5908 12650 5960 12656
rect 5814 12472 5870 12481
rect 5814 12407 5870 12416
rect 5632 12164 5684 12170
rect 5736 12158 5856 12186
rect 5632 12106 5684 12112
rect 5644 11121 5672 12106
rect 5724 12096 5776 12102
rect 5722 12064 5724 12073
rect 5776 12064 5778 12073
rect 5722 11999 5778 12008
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5630 11112 5686 11121
rect 5630 11047 5686 11056
rect 5630 10840 5686 10849
rect 5630 10775 5632 10784
rect 5684 10775 5686 10784
rect 5632 10746 5684 10752
rect 5538 9480 5594 9489
rect 5538 9415 5594 9424
rect 5448 9376 5500 9382
rect 5448 9318 5500 9324
rect 5446 9208 5502 9217
rect 5446 9143 5502 9152
rect 5460 8498 5488 9143
rect 5540 8968 5592 8974
rect 5644 8956 5672 10746
rect 5592 8928 5672 8956
rect 5540 8910 5592 8916
rect 5736 8838 5764 11834
rect 5828 11393 5856 12158
rect 5814 11384 5870 11393
rect 5814 11319 5870 11328
rect 5816 11076 5868 11082
rect 5920 11064 5948 12650
rect 6012 12345 6040 12922
rect 5998 12336 6054 12345
rect 5998 12271 6054 12280
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11150 6040 12038
rect 6104 11626 6132 13806
rect 6288 13824 6408 13852
rect 6182 13767 6238 13776
rect 6380 13734 6408 13824
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6380 12850 6408 13670
rect 6472 12986 6500 17054
rect 6572 16892 6880 16912
rect 6572 16890 6578 16892
rect 6634 16890 6658 16892
rect 6714 16890 6738 16892
rect 6794 16890 6818 16892
rect 6874 16890 6880 16892
rect 6634 16838 6636 16890
rect 6816 16838 6818 16890
rect 6572 16836 6578 16838
rect 6634 16836 6658 16838
rect 6714 16836 6738 16838
rect 6794 16836 6818 16838
rect 6874 16836 6880 16838
rect 6572 16816 6880 16836
rect 7010 16008 7066 16017
rect 7010 15943 7066 15952
rect 6572 15804 6880 15824
rect 6572 15802 6578 15804
rect 6634 15802 6658 15804
rect 6714 15802 6738 15804
rect 6794 15802 6818 15804
rect 6874 15802 6880 15804
rect 6634 15750 6636 15802
rect 6816 15750 6818 15802
rect 6572 15748 6578 15750
rect 6634 15748 6658 15750
rect 6714 15748 6738 15750
rect 6794 15748 6818 15750
rect 6874 15748 6880 15750
rect 6572 15728 6880 15748
rect 7024 15706 7052 15943
rect 7012 15700 7064 15706
rect 7012 15642 7064 15648
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 6572 14716 6880 14736
rect 6572 14714 6578 14716
rect 6634 14714 6658 14716
rect 6714 14714 6738 14716
rect 6794 14714 6818 14716
rect 6874 14714 6880 14716
rect 6634 14662 6636 14714
rect 6816 14662 6818 14714
rect 6572 14660 6578 14662
rect 6634 14660 6658 14662
rect 6714 14660 6738 14662
rect 6794 14660 6818 14662
rect 6874 14660 6880 14662
rect 6572 14640 6880 14660
rect 6828 14408 6880 14414
rect 6734 14376 6790 14385
rect 6828 14350 6880 14356
rect 6918 14376 6974 14385
rect 6734 14311 6790 14320
rect 6642 14240 6698 14249
rect 6642 14175 6698 14184
rect 6656 13802 6684 14175
rect 6748 14006 6776 14311
rect 6840 14249 6868 14350
rect 6918 14311 6974 14320
rect 6826 14240 6882 14249
rect 6826 14175 6882 14184
rect 6736 14000 6788 14006
rect 6736 13942 6788 13948
rect 6644 13796 6696 13802
rect 6644 13738 6696 13744
rect 6572 13628 6880 13648
rect 6572 13626 6578 13628
rect 6634 13626 6658 13628
rect 6714 13626 6738 13628
rect 6794 13626 6818 13628
rect 6874 13626 6880 13628
rect 6634 13574 6636 13626
rect 6816 13574 6818 13626
rect 6572 13572 6578 13574
rect 6634 13572 6658 13574
rect 6714 13572 6738 13574
rect 6794 13572 6818 13574
rect 6874 13572 6880 13574
rect 6572 13552 6880 13572
rect 6932 13512 6960 14311
rect 7024 13977 7052 14894
rect 7010 13968 7066 13977
rect 7116 13938 7144 14894
rect 7208 14890 7236 19230
rect 7286 19200 7342 20000
rect 7654 19200 7710 20000
rect 8022 19200 8078 20000
rect 8390 19200 8446 20000
rect 8758 19200 8814 20000
rect 9126 19200 9182 20000
rect 9494 19200 9550 20000
rect 9862 19200 9918 20000
rect 10230 19200 10286 20000
rect 10598 19200 10654 20000
rect 10966 19200 11022 20000
rect 11072 19230 11284 19258
rect 7300 15162 7328 19200
rect 7562 17776 7618 17785
rect 7562 17711 7618 17720
rect 7576 17241 7604 17711
rect 7562 17232 7618 17241
rect 7562 17167 7618 17176
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7378 15056 7434 15065
rect 7378 14991 7434 15000
rect 7564 15020 7616 15026
rect 7196 14884 7248 14890
rect 7196 14826 7248 14832
rect 7392 14822 7420 14991
rect 7564 14962 7616 14968
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7392 14414 7420 14758
rect 7472 14476 7524 14482
rect 7472 14418 7524 14424
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7288 14340 7340 14346
rect 7288 14282 7340 14288
rect 7010 13903 7066 13912
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7012 13864 7064 13870
rect 7012 13806 7064 13812
rect 6840 13484 6960 13512
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6564 12866 6592 13330
rect 6736 13252 6788 13258
rect 6736 13194 6788 13200
rect 6748 12986 6776 13194
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6472 12838 6592 12866
rect 6380 12753 6408 12786
rect 6366 12744 6422 12753
rect 6366 12679 6422 12688
rect 6276 12640 6328 12646
rect 6276 12582 6328 12588
rect 6288 12322 6316 12582
rect 6196 12294 6316 12322
rect 6092 11620 6144 11626
rect 6092 11562 6144 11568
rect 6090 11520 6146 11529
rect 6090 11455 6146 11464
rect 6104 11286 6132 11455
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 6000 11144 6052 11150
rect 6000 11086 6052 11092
rect 6090 11112 6146 11121
rect 5868 11036 5948 11064
rect 6090 11047 6146 11056
rect 5816 11018 5868 11024
rect 5920 9994 5948 11036
rect 5998 10976 6054 10985
rect 5998 10911 6054 10920
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5828 9382 5856 9930
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5920 9110 5948 9930
rect 5908 9104 5960 9110
rect 5908 9046 5960 9052
rect 5814 8936 5870 8945
rect 5814 8871 5870 8880
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5828 8566 5856 8871
rect 6012 8634 6040 10911
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 5448 8492 5500 8498
rect 5448 8434 5500 8440
rect 5538 8392 5594 8401
rect 5538 8327 5594 8336
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5460 7410 5488 8230
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5264 6656 5316 6662
rect 5264 6598 5316 6604
rect 5448 6656 5500 6662
rect 5448 6598 5500 6604
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5368 6089 5396 6258
rect 5354 6080 5410 6089
rect 5354 6015 5410 6024
rect 5080 5636 5132 5642
rect 5184 5630 5396 5658
rect 5080 5578 5132 5584
rect 4698 5468 5006 5488
rect 4698 5466 4704 5468
rect 4760 5466 4784 5468
rect 4840 5466 4864 5468
rect 4920 5466 4944 5468
rect 5000 5466 5006 5468
rect 4760 5414 4762 5466
rect 4942 5414 4944 5466
rect 4698 5412 4704 5414
rect 4760 5412 4784 5414
rect 4840 5412 4864 5414
rect 4920 5412 4944 5414
rect 5000 5412 5006 5414
rect 4698 5392 5006 5412
rect 5092 5370 5120 5578
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 4620 5024 4672 5030
rect 4620 4966 4672 4972
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4528 3392 4580 3398
rect 4528 3334 4580 3340
rect 4540 2774 4568 3334
rect 4632 3058 4660 4966
rect 4816 4622 4844 4966
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4698 4380 5006 4400
rect 4698 4378 4704 4380
rect 4760 4378 4784 4380
rect 4840 4378 4864 4380
rect 4920 4378 4944 4380
rect 5000 4378 5006 4380
rect 4760 4326 4762 4378
rect 4942 4326 4944 4378
rect 4698 4324 4704 4326
rect 4760 4324 4784 4326
rect 4840 4324 4864 4326
rect 4920 4324 4944 4326
rect 5000 4324 5006 4326
rect 4698 4304 5006 4324
rect 5092 4146 5120 5034
rect 5184 4690 5212 5170
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5170 4584 5226 4593
rect 5276 4554 5304 5510
rect 5170 4519 5226 4528
rect 5264 4548 5316 4554
rect 5080 4140 5132 4146
rect 5080 4082 5132 4088
rect 4698 3292 5006 3312
rect 4698 3290 4704 3292
rect 4760 3290 4784 3292
rect 4840 3290 4864 3292
rect 4920 3290 4944 3292
rect 5000 3290 5006 3292
rect 4760 3238 4762 3290
rect 4942 3238 4944 3290
rect 4698 3236 4704 3238
rect 4760 3236 4784 3238
rect 4840 3236 4864 3238
rect 4920 3236 4944 3238
rect 5000 3236 5006 3238
rect 4698 3216 5006 3236
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4724 2825 4752 2926
rect 4710 2816 4766 2825
rect 4540 2746 4660 2774
rect 4710 2751 4766 2760
rect 4526 2680 4582 2689
rect 4526 2615 4528 2624
rect 4580 2615 4582 2624
rect 4528 2586 4580 2592
rect 4528 2372 4580 2378
rect 4528 2314 4580 2320
rect 4540 2145 4568 2314
rect 4526 2136 4582 2145
rect 4526 2071 4582 2080
rect 4436 1964 4488 1970
rect 4436 1906 4488 1912
rect 4540 1562 4568 2071
rect 4528 1556 4580 1562
rect 4528 1498 4580 1504
rect 4448 870 4568 898
rect 3700 740 3752 746
rect 3700 682 3752 688
rect 3882 0 3938 800
rect 4158 0 4214 800
rect 4448 202 4476 870
rect 4540 800 4568 870
rect 4436 196 4488 202
rect 4436 138 4488 144
rect 4526 0 4582 800
rect 4632 762 4660 2746
rect 4896 2440 4948 2446
rect 5000 2428 5028 2994
rect 5092 2514 5120 4082
rect 5080 2508 5132 2514
rect 5080 2450 5132 2456
rect 4948 2400 5028 2428
rect 4896 2382 4948 2388
rect 4698 2204 5006 2224
rect 4698 2202 4704 2204
rect 4760 2202 4784 2204
rect 4840 2202 4864 2204
rect 4920 2202 4944 2204
rect 5000 2202 5006 2204
rect 4760 2150 4762 2202
rect 4942 2150 4944 2202
rect 4698 2148 4704 2150
rect 4760 2148 4784 2150
rect 4840 2148 4864 2150
rect 4920 2148 4944 2150
rect 5000 2148 5006 2150
rect 4698 2128 5006 2148
rect 5184 1394 5212 4519
rect 5264 4490 5316 4496
rect 5262 4448 5318 4457
rect 5262 4383 5318 4392
rect 5276 3670 5304 4383
rect 5264 3664 5316 3670
rect 5264 3606 5316 3612
rect 5368 1494 5396 5630
rect 5460 5302 5488 6598
rect 5552 5681 5580 8327
rect 5814 8120 5870 8129
rect 5724 8084 5776 8090
rect 5814 8055 5870 8064
rect 5724 8026 5776 8032
rect 5630 7984 5686 7993
rect 5630 7919 5632 7928
rect 5684 7919 5686 7928
rect 5632 7890 5684 7896
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5644 5710 5672 7686
rect 5632 5704 5684 5710
rect 5538 5672 5594 5681
rect 5632 5646 5684 5652
rect 5538 5607 5594 5616
rect 5736 5556 5764 8026
rect 5552 5528 5764 5556
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5460 3602 5488 4966
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5460 3126 5488 3334
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5552 2825 5580 5528
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5630 3496 5686 3505
rect 5630 3431 5686 3440
rect 5644 2922 5672 3431
rect 5632 2916 5684 2922
rect 5632 2858 5684 2864
rect 5538 2816 5594 2825
rect 5538 2751 5594 2760
rect 5446 2544 5502 2553
rect 5446 2479 5502 2488
rect 5460 2446 5488 2479
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 5356 1488 5408 1494
rect 5356 1430 5408 1436
rect 5184 1366 5304 1394
rect 4816 870 4936 898
rect 4816 762 4844 870
rect 4908 800 4936 870
rect 5276 800 5304 1366
rect 5736 1170 5764 3674
rect 5828 3369 5856 8055
rect 5906 7848 5962 7857
rect 5906 7783 5962 7792
rect 5920 6118 5948 7783
rect 5998 7712 6054 7721
rect 5998 7647 6054 7656
rect 5908 6112 5960 6118
rect 5908 6054 5960 6060
rect 6012 5692 6040 7647
rect 6104 6905 6132 11047
rect 6196 9110 6224 12294
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6288 11898 6316 12174
rect 6366 12064 6422 12073
rect 6366 11999 6422 12008
rect 6472 12050 6500 12838
rect 6840 12628 6868 13484
rect 6918 13424 6974 13433
rect 6918 13359 6974 13368
rect 6932 13326 6960 13359
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 7024 12918 7052 13806
rect 7196 13796 7248 13802
rect 7196 13738 7248 13744
rect 7102 13560 7158 13569
rect 7102 13495 7104 13504
rect 7156 13495 7158 13504
rect 7104 13466 7156 13472
rect 7208 13410 7236 13738
rect 7116 13382 7236 13410
rect 7116 13190 7144 13382
rect 7104 13184 7156 13190
rect 7104 13126 7156 13132
rect 7196 13184 7248 13190
rect 7196 13126 7248 13132
rect 7012 12912 7064 12918
rect 7208 12889 7236 13126
rect 7012 12854 7064 12860
rect 7194 12880 7250 12889
rect 6840 12600 6960 12628
rect 6572 12540 6880 12560
rect 6572 12538 6578 12540
rect 6634 12538 6658 12540
rect 6714 12538 6738 12540
rect 6794 12538 6818 12540
rect 6874 12538 6880 12540
rect 6634 12486 6636 12538
rect 6816 12486 6818 12538
rect 6572 12484 6578 12486
rect 6634 12484 6658 12486
rect 6714 12484 6738 12486
rect 6794 12484 6818 12486
rect 6874 12484 6880 12486
rect 6572 12464 6880 12484
rect 6932 12322 6960 12600
rect 6564 12294 6960 12322
rect 6564 12170 6592 12294
rect 6828 12232 6880 12238
rect 6828 12174 6880 12180
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6748 12050 6776 12106
rect 6840 12073 6868 12174
rect 6920 12096 6972 12102
rect 6472 12022 6776 12050
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6380 11694 6408 11999
rect 6368 11688 6420 11694
rect 6368 11630 6420 11636
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 6288 9897 6316 11562
rect 6380 11150 6408 11630
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6380 10606 6408 11086
rect 6368 10600 6420 10606
rect 6368 10542 6420 10548
rect 6380 9926 6408 10542
rect 6368 9920 6420 9926
rect 6274 9888 6330 9897
rect 6368 9862 6420 9868
rect 6274 9823 6330 9832
rect 6380 9586 6408 9862
rect 6472 9654 6500 12022
rect 6748 11830 6776 12022
rect 6826 12064 6882 12073
rect 6920 12038 6972 12044
rect 6826 11999 6882 12008
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6572 11452 6880 11472
rect 6572 11450 6578 11452
rect 6634 11450 6658 11452
rect 6714 11450 6738 11452
rect 6794 11450 6818 11452
rect 6874 11450 6880 11452
rect 6634 11398 6636 11450
rect 6816 11398 6818 11450
rect 6572 11396 6578 11398
rect 6634 11396 6658 11398
rect 6714 11396 6738 11398
rect 6794 11396 6818 11398
rect 6874 11396 6880 11398
rect 6572 11376 6880 11396
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6840 10849 6868 10950
rect 6826 10840 6882 10849
rect 6932 10810 6960 12038
rect 7024 10810 7052 12854
rect 7194 12815 7250 12824
rect 7194 12744 7250 12753
rect 7194 12679 7196 12688
rect 7248 12679 7250 12688
rect 7196 12650 7248 12656
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7102 12200 7158 12209
rect 7102 12135 7158 12144
rect 6826 10775 6882 10784
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6644 10668 6696 10674
rect 6696 10628 6868 10656
rect 6644 10610 6696 10616
rect 6840 10588 6868 10628
rect 6840 10560 6960 10588
rect 6572 10364 6880 10384
rect 6572 10362 6578 10364
rect 6634 10362 6658 10364
rect 6714 10362 6738 10364
rect 6794 10362 6818 10364
rect 6874 10362 6880 10364
rect 6634 10310 6636 10362
rect 6816 10310 6818 10362
rect 6572 10308 6578 10310
rect 6634 10308 6658 10310
rect 6714 10308 6738 10310
rect 6794 10308 6818 10310
rect 6874 10308 6880 10310
rect 6572 10288 6880 10308
rect 6932 10266 6960 10560
rect 7116 10441 7144 12135
rect 7208 11801 7236 12378
rect 7194 11792 7250 11801
rect 7194 11727 7250 11736
rect 7300 11354 7328 14282
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7288 11348 7340 11354
rect 7288 11290 7340 11296
rect 7208 11234 7236 11290
rect 7392 11234 7420 13330
rect 7484 12782 7512 14418
rect 7576 14346 7604 14962
rect 7668 14618 7696 19200
rect 7748 16448 7800 16454
rect 7748 16390 7800 16396
rect 7760 15745 7788 16390
rect 7840 16108 7892 16114
rect 7840 16050 7892 16056
rect 7746 15736 7802 15745
rect 7746 15671 7748 15680
rect 7800 15671 7802 15680
rect 7748 15642 7800 15648
rect 7748 15360 7800 15366
rect 7852 15337 7880 16050
rect 8036 15502 8064 19200
rect 8404 17626 8432 19200
rect 8312 17598 8432 17626
rect 8772 17626 8800 19200
rect 8772 17598 8984 17626
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 8116 15360 8168 15366
rect 7748 15302 7800 15308
rect 7838 15328 7894 15337
rect 7760 15026 7788 15302
rect 8116 15302 8168 15308
rect 7838 15263 7894 15272
rect 7838 15192 7894 15201
rect 7838 15127 7894 15136
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7760 14793 7788 14962
rect 7746 14784 7802 14793
rect 7746 14719 7802 14728
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7760 14498 7788 14719
rect 7852 14657 7880 15127
rect 7838 14648 7894 14657
rect 7838 14583 7894 14592
rect 8022 14648 8078 14657
rect 8022 14583 8078 14592
rect 7668 14470 7788 14498
rect 7840 14544 7892 14550
rect 7840 14486 7892 14492
rect 7564 14340 7616 14346
rect 7564 14282 7616 14288
rect 7576 13938 7604 14282
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7564 13388 7616 13394
rect 7564 13330 7616 13336
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 7576 12238 7604 13330
rect 7564 12232 7616 12238
rect 7564 12174 7616 12180
rect 7472 11552 7524 11558
rect 7576 11540 7604 12174
rect 7524 11512 7604 11540
rect 7472 11494 7524 11500
rect 7208 11206 7420 11234
rect 7102 10432 7158 10441
rect 7102 10367 7158 10376
rect 7010 10296 7066 10305
rect 6920 10260 6972 10266
rect 7010 10231 7066 10240
rect 6920 10202 6972 10208
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6748 9654 6776 9998
rect 6932 9722 6960 10202
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6460 9648 6512 9654
rect 6460 9590 6512 9596
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6918 9480 6974 9489
rect 6918 9415 6974 9424
rect 6572 9276 6880 9296
rect 6572 9274 6578 9276
rect 6634 9274 6658 9276
rect 6714 9274 6738 9276
rect 6794 9274 6818 9276
rect 6874 9274 6880 9276
rect 6634 9222 6636 9274
rect 6816 9222 6818 9274
rect 6572 9220 6578 9222
rect 6634 9220 6658 9222
rect 6714 9220 6738 9222
rect 6794 9220 6818 9222
rect 6874 9220 6880 9222
rect 6572 9200 6880 9220
rect 6932 9178 6960 9415
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6184 8968 6236 8974
rect 6184 8910 6236 8916
rect 6196 8430 6224 8910
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6196 7342 6224 8366
rect 6572 8188 6880 8208
rect 6572 8186 6578 8188
rect 6634 8186 6658 8188
rect 6714 8186 6738 8188
rect 6794 8186 6818 8188
rect 6874 8186 6880 8188
rect 6634 8134 6636 8186
rect 6816 8134 6818 8186
rect 6572 8132 6578 8134
rect 6634 8132 6658 8134
rect 6714 8132 6738 8134
rect 6794 8132 6818 8134
rect 6874 8132 6880 8134
rect 6572 8112 6880 8132
rect 6460 7880 6512 7886
rect 6288 7840 6460 7868
rect 6184 7336 6236 7342
rect 6184 7278 6236 7284
rect 6090 6896 6146 6905
rect 6196 6866 6224 7278
rect 6288 6934 6316 7840
rect 6460 7822 6512 7828
rect 6932 7410 6960 9114
rect 7024 8945 7052 10231
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7010 8936 7066 8945
rect 7010 8871 7012 8880
rect 7064 8871 7066 8880
rect 7012 8842 7064 8848
rect 7012 8560 7064 8566
rect 7012 8502 7064 8508
rect 6920 7404 6972 7410
rect 6920 7346 6972 7352
rect 6458 7304 6514 7313
rect 6458 7239 6514 7248
rect 6918 7304 6974 7313
rect 6918 7239 6974 7248
rect 6472 7206 6500 7239
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6572 7100 6880 7120
rect 6572 7098 6578 7100
rect 6634 7098 6658 7100
rect 6714 7098 6738 7100
rect 6794 7098 6818 7100
rect 6874 7098 6880 7100
rect 6634 7046 6636 7098
rect 6816 7046 6818 7098
rect 6572 7044 6578 7046
rect 6634 7044 6658 7046
rect 6714 7044 6738 7046
rect 6794 7044 6818 7046
rect 6874 7044 6880 7046
rect 6572 7024 6880 7044
rect 6276 6928 6328 6934
rect 6276 6870 6328 6876
rect 6090 6831 6146 6840
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 5920 5664 6040 5692
rect 5920 3398 5948 5664
rect 6104 5302 6132 6394
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 6104 4622 6132 5238
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6092 4480 6144 4486
rect 6092 4422 6144 4428
rect 5908 3392 5960 3398
rect 5814 3360 5870 3369
rect 5908 3334 5960 3340
rect 5814 3295 5870 3304
rect 5828 3058 5856 3295
rect 5906 3224 5962 3233
rect 5906 3159 5962 3168
rect 5920 3126 5948 3159
rect 5908 3120 5960 3126
rect 5908 3062 5960 3068
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 6104 2990 6132 4422
rect 6196 3398 6224 6054
rect 6288 5302 6316 6870
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6472 5896 6500 6258
rect 6572 6012 6880 6032
rect 6572 6010 6578 6012
rect 6634 6010 6658 6012
rect 6714 6010 6738 6012
rect 6794 6010 6818 6012
rect 6874 6010 6880 6012
rect 6634 5958 6636 6010
rect 6816 5958 6818 6010
rect 6572 5956 6578 5958
rect 6634 5956 6658 5958
rect 6714 5956 6738 5958
rect 6794 5956 6818 5958
rect 6874 5956 6880 5958
rect 6572 5936 6880 5956
rect 6472 5868 6592 5896
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6368 5092 6420 5098
rect 6368 5034 6420 5040
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6288 4146 6316 4966
rect 6380 4554 6408 5034
rect 6368 4548 6420 4554
rect 6368 4490 6420 4496
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6276 3936 6328 3942
rect 6276 3878 6328 3884
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6092 2984 6144 2990
rect 6092 2926 6144 2932
rect 6090 2816 6146 2825
rect 6090 2751 6146 2760
rect 5906 2680 5962 2689
rect 5906 2615 5962 2624
rect 5814 2544 5870 2553
rect 5920 2514 5948 2615
rect 6104 2514 6132 2751
rect 5814 2479 5870 2488
rect 5908 2508 5960 2514
rect 5828 2446 5856 2479
rect 5908 2450 5960 2456
rect 6092 2508 6144 2514
rect 6092 2450 6144 2456
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6090 2272 6146 2281
rect 6090 2207 6146 2216
rect 5736 1142 6040 1170
rect 5908 1080 5960 1086
rect 5908 1022 5960 1028
rect 5552 870 5672 898
rect 5552 800 5580 870
rect 5644 814 5672 870
rect 5632 808 5684 814
rect 4632 734 4844 762
rect 4894 0 4950 800
rect 5262 0 5318 800
rect 5538 0 5594 800
rect 5920 800 5948 1022
rect 5632 750 5684 756
rect 5906 0 5962 800
rect 6012 762 6040 1142
rect 6104 950 6132 2207
rect 6196 1222 6224 3130
rect 6288 2961 6316 3878
rect 6472 3738 6500 5578
rect 6564 5574 6592 5868
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6564 5166 6592 5510
rect 6932 5273 6960 7239
rect 7024 6730 7052 8502
rect 7116 8498 7144 9318
rect 7208 8906 7236 11206
rect 7484 11014 7512 11494
rect 7668 11370 7696 14470
rect 7746 14104 7802 14113
rect 7746 14039 7802 14048
rect 7760 13705 7788 14039
rect 7746 13696 7802 13705
rect 7746 13631 7802 13640
rect 7760 13190 7788 13631
rect 7852 13394 7880 14486
rect 7932 14408 7984 14414
rect 7932 14350 7984 14356
rect 7944 13394 7972 14350
rect 7840 13388 7892 13394
rect 7840 13330 7892 13336
rect 7932 13388 7984 13394
rect 7932 13330 7984 13336
rect 7840 13252 7892 13258
rect 7840 13194 7892 13200
rect 7932 13252 7984 13258
rect 7932 13194 7984 13200
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7760 11393 7788 12718
rect 7576 11342 7696 11370
rect 7746 11384 7802 11393
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7380 10056 7432 10062
rect 7380 9998 7432 10004
rect 7392 9654 7420 9998
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7286 9344 7342 9353
rect 7286 9279 7342 9288
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7300 7721 7328 9279
rect 7470 8936 7526 8945
rect 7470 8871 7526 8880
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7286 7712 7342 7721
rect 7286 7647 7342 7656
rect 7286 7168 7342 7177
rect 7286 7103 7342 7112
rect 7102 7032 7158 7041
rect 7102 6967 7104 6976
rect 7156 6967 7158 6976
rect 7104 6938 7156 6944
rect 7012 6724 7064 6730
rect 7012 6666 7064 6672
rect 7024 6440 7052 6666
rect 7024 6412 7144 6440
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6918 5264 6974 5273
rect 6918 5199 6974 5208
rect 6552 5160 6604 5166
rect 6552 5102 6604 5108
rect 6572 4924 6880 4944
rect 6572 4922 6578 4924
rect 6634 4922 6658 4924
rect 6714 4922 6738 4924
rect 6794 4922 6818 4924
rect 6874 4922 6880 4924
rect 6634 4870 6636 4922
rect 6816 4870 6818 4922
rect 6572 4868 6578 4870
rect 6634 4868 6658 4870
rect 6714 4868 6738 4870
rect 6794 4868 6818 4870
rect 6874 4868 6880 4870
rect 6572 4848 6880 4868
rect 7024 4758 7052 6258
rect 7116 6118 7144 6412
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7208 5930 7236 6326
rect 7116 5902 7236 5930
rect 7116 5137 7144 5902
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 7102 5128 7158 5137
rect 7102 5063 7158 5072
rect 7102 4856 7158 4865
rect 7102 4791 7158 4800
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 6736 4616 6788 4622
rect 6736 4558 6788 4564
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6552 4072 6604 4078
rect 6550 4040 6552 4049
rect 6604 4040 6606 4049
rect 6550 3975 6606 3984
rect 6748 3924 6776 4558
rect 6932 4146 6960 4558
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 7024 4185 7052 4422
rect 7010 4176 7066 4185
rect 6828 4140 6880 4146
rect 6828 4082 6880 4088
rect 6920 4140 6972 4146
rect 7010 4111 7066 4120
rect 6920 4082 6972 4088
rect 6840 4049 6868 4082
rect 6826 4040 6882 4049
rect 6826 3975 6882 3984
rect 6748 3896 6960 3924
rect 6572 3836 6880 3856
rect 6572 3834 6578 3836
rect 6634 3834 6658 3836
rect 6714 3834 6738 3836
rect 6794 3834 6818 3836
rect 6874 3834 6880 3836
rect 6634 3782 6636 3834
rect 6816 3782 6818 3834
rect 6572 3780 6578 3782
rect 6634 3780 6658 3782
rect 6714 3780 6738 3782
rect 6794 3780 6818 3782
rect 6874 3780 6880 3782
rect 6572 3760 6880 3780
rect 6460 3732 6512 3738
rect 6460 3674 6512 3680
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6380 3097 6408 3130
rect 6460 3120 6512 3126
rect 6366 3088 6422 3097
rect 6460 3062 6512 3068
rect 6366 3023 6422 3032
rect 6368 2984 6420 2990
rect 6274 2952 6330 2961
rect 6368 2926 6420 2932
rect 6274 2887 6330 2896
rect 6380 1766 6408 2926
rect 6472 2310 6500 3062
rect 6564 2922 6592 3606
rect 6932 3482 6960 3896
rect 7116 3754 7144 4791
rect 7024 3738 7144 3754
rect 7012 3732 7144 3738
rect 7064 3726 7144 3732
rect 7012 3674 7064 3680
rect 7104 3664 7156 3670
rect 7104 3606 7156 3612
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6748 3454 6960 3482
rect 7024 3466 7052 3538
rect 7012 3460 7064 3466
rect 6748 2922 6776 3454
rect 7012 3402 7064 3408
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6840 2972 6868 3334
rect 6932 3074 6960 3334
rect 6932 3046 7052 3074
rect 6920 2984 6972 2990
rect 6840 2944 6920 2972
rect 6920 2926 6972 2932
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6572 2748 6880 2768
rect 6572 2746 6578 2748
rect 6634 2746 6658 2748
rect 6714 2746 6738 2748
rect 6794 2746 6818 2748
rect 6874 2746 6880 2748
rect 6634 2694 6636 2746
rect 6816 2694 6818 2746
rect 6572 2692 6578 2694
rect 6634 2692 6658 2694
rect 6714 2692 6738 2694
rect 6794 2692 6818 2694
rect 6874 2692 6880 2694
rect 6572 2672 6880 2692
rect 6920 2644 6972 2650
rect 6920 2586 6972 2592
rect 6828 2576 6880 2582
rect 6826 2544 6828 2553
rect 6880 2544 6882 2553
rect 6826 2479 6882 2488
rect 6932 2446 6960 2586
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6828 2032 6880 2038
rect 6828 1974 6880 1980
rect 6368 1760 6420 1766
rect 6368 1702 6420 1708
rect 6840 1358 6868 1974
rect 7024 1873 7052 3046
rect 7116 2514 7144 3606
rect 7208 2990 7236 5238
rect 7300 5001 7328 7103
rect 7392 5953 7420 8366
rect 7484 6361 7512 8871
rect 7470 6352 7526 6361
rect 7470 6287 7526 6296
rect 7576 6118 7604 11342
rect 7746 11319 7802 11328
rect 7852 11234 7880 13194
rect 7944 11370 7972 13194
rect 8036 13025 8064 14583
rect 8022 13016 8078 13025
rect 8022 12951 8078 12960
rect 8036 12850 8064 12951
rect 8024 12844 8076 12850
rect 8024 12786 8076 12792
rect 8024 12436 8076 12442
rect 8024 12378 8076 12384
rect 8036 12345 8064 12378
rect 8022 12336 8078 12345
rect 8022 12271 8078 12280
rect 8128 12238 8156 15302
rect 8220 14618 8248 16526
rect 8208 14612 8260 14618
rect 8208 14554 8260 14560
rect 8208 14476 8260 14482
rect 8208 14418 8260 14424
rect 8220 14006 8248 14418
rect 8208 14000 8260 14006
rect 8208 13942 8260 13948
rect 8220 12782 8248 13942
rect 8312 13530 8340 17598
rect 8446 17436 8754 17456
rect 8446 17434 8452 17436
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8748 17434 8754 17436
rect 8508 17382 8510 17434
rect 8690 17382 8692 17434
rect 8446 17380 8452 17382
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8748 17380 8754 17382
rect 8446 17360 8754 17380
rect 8446 16348 8754 16368
rect 8446 16346 8452 16348
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8748 16346 8754 16348
rect 8508 16294 8510 16346
rect 8690 16294 8692 16346
rect 8446 16292 8452 16294
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8748 16292 8754 16294
rect 8446 16272 8754 16292
rect 8446 15260 8754 15280
rect 8446 15258 8452 15260
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8748 15258 8754 15260
rect 8508 15206 8510 15258
rect 8690 15206 8692 15258
rect 8446 15204 8452 15206
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8748 15204 8754 15206
rect 8446 15184 8754 15204
rect 8484 14952 8536 14958
rect 8484 14894 8536 14900
rect 8496 14822 8524 14894
rect 8484 14816 8536 14822
rect 8484 14758 8536 14764
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8496 14414 8524 14758
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8680 14260 8708 14758
rect 8864 14618 8892 14758
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8680 14232 8892 14260
rect 8446 14172 8754 14192
rect 8446 14170 8452 14172
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8748 14170 8754 14172
rect 8508 14118 8510 14170
rect 8690 14118 8692 14170
rect 8446 14116 8452 14118
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8748 14116 8754 14118
rect 8446 14096 8754 14116
rect 8668 13932 8720 13938
rect 8864 13920 8892 14232
rect 8956 14006 8984 17598
rect 9036 15496 9088 15502
rect 9036 15438 9088 15444
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8720 13892 8892 13920
rect 8668 13874 8720 13880
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8312 12850 8340 13330
rect 8446 13084 8754 13104
rect 8446 13082 8452 13084
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8748 13082 8754 13084
rect 8508 13030 8510 13082
rect 8690 13030 8692 13082
rect 8446 13028 8452 13030
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8748 13028 8754 13030
rect 8446 13008 8754 13028
rect 8300 12844 8352 12850
rect 8300 12786 8352 12792
rect 8208 12776 8260 12782
rect 8208 12718 8260 12724
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8300 12708 8352 12714
rect 8300 12650 8352 12656
rect 8206 12472 8262 12481
rect 8206 12407 8262 12416
rect 8116 12232 8168 12238
rect 8116 12174 8168 12180
rect 8220 12102 8248 12407
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8116 11824 8168 11830
rect 8114 11792 8116 11801
rect 8168 11792 8170 11801
rect 8312 11778 8340 12650
rect 8772 12345 8800 12718
rect 8758 12336 8814 12345
rect 8758 12271 8814 12280
rect 8446 11996 8754 12016
rect 8446 11994 8452 11996
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8748 11994 8754 11996
rect 8508 11942 8510 11994
rect 8690 11942 8692 11994
rect 8446 11940 8452 11942
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8748 11940 8754 11942
rect 8446 11920 8754 11940
rect 8574 11792 8630 11801
rect 8312 11750 8432 11778
rect 8114 11727 8170 11736
rect 8300 11688 8352 11694
rect 8300 11630 8352 11636
rect 8208 11552 8260 11558
rect 8208 11494 8260 11500
rect 8114 11384 8170 11393
rect 7944 11342 8064 11370
rect 7760 11206 7880 11234
rect 7932 11212 7984 11218
rect 7760 11150 7788 11206
rect 7932 11154 7984 11160
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7656 11076 7708 11082
rect 7656 11018 7708 11024
rect 7668 10538 7696 11018
rect 7748 11008 7800 11014
rect 7748 10950 7800 10956
rect 7656 10532 7708 10538
rect 7656 10474 7708 10480
rect 7668 9450 7696 10474
rect 7760 10130 7788 10950
rect 7852 10606 7880 11086
rect 7944 10962 7972 11154
rect 8036 11150 8064 11342
rect 8114 11319 8170 11328
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 8128 10985 8156 11319
rect 8114 10976 8170 10985
rect 7944 10934 8064 10962
rect 7840 10600 7892 10606
rect 7932 10600 7984 10606
rect 7840 10542 7892 10548
rect 7930 10568 7932 10577
rect 7984 10568 7986 10577
rect 7930 10503 7986 10512
rect 7748 10124 7800 10130
rect 7748 10066 7800 10072
rect 7930 9888 7986 9897
rect 7930 9823 7986 9832
rect 7944 9722 7972 9823
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 7748 9648 7800 9654
rect 7748 9590 7800 9596
rect 7656 9444 7708 9450
rect 7656 9386 7708 9392
rect 7760 8634 7788 9590
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7852 7886 7880 8434
rect 7840 7880 7892 7886
rect 7840 7822 7892 7828
rect 7852 7750 7880 7822
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7852 7410 7880 7686
rect 7840 7404 7892 7410
rect 7840 7346 7892 7352
rect 7944 7313 7972 7686
rect 8036 7546 8064 10934
rect 8114 10911 8170 10920
rect 8114 10840 8170 10849
rect 8114 10775 8170 10784
rect 8128 10674 8156 10775
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 8116 10260 8168 10266
rect 8220 10248 8248 11494
rect 8168 10220 8248 10248
rect 8116 10202 8168 10208
rect 8114 9752 8170 9761
rect 8114 9687 8170 9696
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 7930 7304 7986 7313
rect 7930 7239 7986 7248
rect 7840 7200 7892 7206
rect 7840 7142 7892 7148
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7378 5944 7434 5953
rect 7378 5879 7380 5888
rect 7432 5879 7434 5888
rect 7472 5908 7524 5914
rect 7380 5850 7432 5856
rect 7472 5850 7524 5856
rect 7484 5148 7512 5850
rect 7392 5120 7512 5148
rect 7286 4992 7342 5001
rect 7286 4927 7342 4936
rect 7288 4684 7340 4690
rect 7288 4626 7340 4632
rect 7196 2984 7248 2990
rect 7196 2926 7248 2932
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7116 1970 7144 2246
rect 7104 1964 7156 1970
rect 7104 1906 7156 1912
rect 7010 1864 7066 1873
rect 6920 1828 6972 1834
rect 7010 1799 7066 1808
rect 6920 1770 6972 1776
rect 6828 1352 6880 1358
rect 6828 1294 6880 1300
rect 6184 1216 6236 1222
rect 6184 1158 6236 1164
rect 6828 1080 6880 1086
rect 6828 1022 6880 1028
rect 6092 944 6144 950
rect 6092 886 6144 892
rect 6196 870 6316 898
rect 6196 762 6224 870
rect 6288 800 6316 870
rect 6656 870 6776 898
rect 6656 800 6684 870
rect 6012 734 6224 762
rect 6274 0 6330 800
rect 6642 0 6698 800
rect 6748 241 6776 870
rect 6840 270 6868 1022
rect 6932 800 6960 1770
rect 7300 800 7328 4626
rect 7392 3890 7420 5120
rect 7470 4992 7526 5001
rect 7470 4927 7526 4936
rect 7484 4049 7512 4927
rect 7470 4040 7526 4049
rect 7470 3975 7526 3984
rect 7392 3862 7512 3890
rect 7378 3768 7434 3777
rect 7378 3703 7434 3712
rect 7392 3602 7420 3703
rect 7380 3596 7432 3602
rect 7380 3538 7432 3544
rect 7484 3398 7512 3862
rect 7472 3392 7524 3398
rect 7378 3360 7434 3369
rect 7472 3334 7524 3340
rect 7378 3295 7434 3304
rect 7392 1086 7420 3295
rect 7470 3224 7526 3233
rect 7576 3194 7604 6054
rect 7668 5302 7696 6938
rect 7748 6792 7800 6798
rect 7748 6734 7800 6740
rect 7760 6322 7788 6734
rect 7852 6662 7880 7142
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7760 5710 7788 6258
rect 7852 5914 7880 6598
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7656 5296 7708 5302
rect 7656 5238 7708 5244
rect 7668 4146 7696 5238
rect 7760 5234 7788 5646
rect 7748 5228 7800 5234
rect 7748 5170 7800 5176
rect 7760 4622 7788 5170
rect 7840 5024 7892 5030
rect 7840 4966 7892 4972
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7748 4208 7800 4214
rect 7746 4176 7748 4185
rect 7800 4176 7802 4185
rect 7656 4140 7708 4146
rect 7746 4111 7802 4120
rect 7656 4082 7708 4088
rect 7746 4040 7802 4049
rect 7746 3975 7802 3984
rect 7656 3596 7708 3602
rect 7656 3538 7708 3544
rect 7668 3466 7696 3538
rect 7760 3466 7788 3975
rect 7656 3460 7708 3466
rect 7656 3402 7708 3408
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7470 3159 7472 3168
rect 7524 3159 7526 3168
rect 7564 3188 7616 3194
rect 7472 3130 7524 3136
rect 7564 3130 7616 3136
rect 7576 3040 7604 3130
rect 7576 3012 7696 3040
rect 7470 2952 7526 2961
rect 7470 2887 7526 2896
rect 7484 2689 7512 2887
rect 7470 2680 7526 2689
rect 7470 2615 7526 2624
rect 7564 2304 7616 2310
rect 7564 2246 7616 2252
rect 7576 1698 7604 2246
rect 7668 1850 7696 3012
rect 7852 2774 7880 4966
rect 7944 3602 7972 6598
rect 8036 5370 8064 7346
rect 8128 6798 8156 9687
rect 8220 9586 8248 10220
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8312 9024 8340 11630
rect 8404 11150 8432 11750
rect 8864 11762 8892 13892
rect 8944 13728 8996 13734
rect 8944 13670 8996 13676
rect 8956 12374 8984 13670
rect 9048 13530 9076 15438
rect 9140 14074 9168 19200
rect 9404 16040 9456 16046
rect 9404 15982 9456 15988
rect 9416 15910 9444 15982
rect 9404 15904 9456 15910
rect 9404 15846 9456 15852
rect 9220 15632 9272 15638
rect 9220 15574 9272 15580
rect 9232 14550 9260 15574
rect 9402 14920 9458 14929
rect 9402 14855 9458 14864
rect 9416 14550 9444 14855
rect 9220 14544 9272 14550
rect 9220 14486 9272 14492
rect 9404 14544 9456 14550
rect 9404 14486 9456 14492
rect 9402 14376 9458 14385
rect 9402 14311 9458 14320
rect 9416 14278 9444 14311
rect 9312 14272 9364 14278
rect 9312 14214 9364 14220
rect 9404 14272 9456 14278
rect 9404 14214 9456 14220
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9128 13796 9180 13802
rect 9128 13738 9180 13744
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9036 12776 9088 12782
rect 9036 12718 9088 12724
rect 8944 12368 8996 12374
rect 9048 12345 9076 12718
rect 8944 12310 8996 12316
rect 9034 12336 9090 12345
rect 8956 11880 8984 12310
rect 9034 12271 9090 12280
rect 9140 11937 9168 13738
rect 9220 13456 9272 13462
rect 9220 13398 9272 13404
rect 9232 12986 9260 13398
rect 9220 12980 9272 12986
rect 9220 12922 9272 12928
rect 9324 12730 9352 14214
rect 9402 14104 9458 14113
rect 9402 14039 9404 14048
rect 9456 14039 9458 14048
rect 9404 14010 9456 14016
rect 9508 13530 9536 19200
rect 9876 18034 9904 19200
rect 9876 18006 9996 18034
rect 9678 17912 9734 17921
rect 9678 17847 9734 17856
rect 9862 17912 9918 17921
rect 9862 17847 9918 17856
rect 9692 15570 9720 17847
rect 9772 16788 9824 16794
rect 9772 16730 9824 16736
rect 9680 15564 9732 15570
rect 9680 15506 9732 15512
rect 9784 15366 9812 16730
rect 9876 16697 9904 17847
rect 9862 16688 9918 16697
rect 9862 16623 9918 16632
rect 9968 15706 9996 18006
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 9772 15360 9824 15366
rect 9772 15302 9824 15308
rect 9586 15056 9642 15065
rect 9586 14991 9642 15000
rect 9600 14414 9628 14991
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9692 14657 9720 14758
rect 9678 14648 9734 14657
rect 9678 14583 9734 14592
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 9588 13932 9640 13938
rect 9692 13920 9720 14583
rect 9640 13892 9720 13920
rect 9588 13874 9640 13880
rect 10060 13870 10088 16526
rect 10244 15978 10272 19200
rect 10612 17048 10640 19200
rect 10980 17954 11008 19200
rect 10888 17926 11008 17954
rect 10612 17020 10732 17048
rect 10320 16892 10628 16912
rect 10320 16890 10326 16892
rect 10382 16890 10406 16892
rect 10462 16890 10486 16892
rect 10542 16890 10566 16892
rect 10622 16890 10628 16892
rect 10382 16838 10384 16890
rect 10564 16838 10566 16890
rect 10320 16836 10326 16838
rect 10382 16836 10406 16838
rect 10462 16836 10486 16838
rect 10542 16836 10566 16838
rect 10622 16836 10628 16838
rect 10320 16816 10628 16836
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10320 15804 10628 15824
rect 10320 15802 10326 15804
rect 10382 15802 10406 15804
rect 10462 15802 10486 15804
rect 10542 15802 10566 15804
rect 10622 15802 10628 15804
rect 10382 15750 10384 15802
rect 10564 15750 10566 15802
rect 10320 15748 10326 15750
rect 10382 15748 10406 15750
rect 10462 15748 10486 15750
rect 10542 15748 10566 15750
rect 10622 15748 10628 15750
rect 10320 15728 10628 15748
rect 10704 15502 10732 17020
rect 10888 16574 10916 17926
rect 10796 16546 10916 16574
rect 10966 16552 11022 16561
rect 10692 15496 10744 15502
rect 10692 15438 10744 15444
rect 10140 15428 10192 15434
rect 10140 15370 10192 15376
rect 9772 13864 9824 13870
rect 9770 13832 9772 13841
rect 10048 13864 10100 13870
rect 9824 13832 9826 13841
rect 9588 13796 9640 13802
rect 9640 13756 9720 13784
rect 10048 13806 10100 13812
rect 10152 13802 10180 15370
rect 10320 14716 10628 14736
rect 10320 14714 10326 14716
rect 10382 14714 10406 14716
rect 10462 14714 10486 14716
rect 10542 14714 10566 14716
rect 10622 14714 10628 14716
rect 10382 14662 10384 14714
rect 10564 14662 10566 14714
rect 10320 14660 10326 14662
rect 10382 14660 10406 14662
rect 10462 14660 10486 14662
rect 10542 14660 10566 14662
rect 10622 14660 10628 14662
rect 10320 14640 10628 14660
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 9770 13767 9826 13776
rect 10140 13796 10192 13802
rect 9588 13738 9640 13744
rect 9496 13524 9548 13530
rect 9496 13466 9548 13472
rect 9588 13524 9640 13530
rect 9588 13466 9640 13472
rect 9404 13320 9456 13326
rect 9402 13288 9404 13297
rect 9456 13288 9458 13297
rect 9600 13274 9628 13466
rect 9402 13223 9458 13232
rect 9508 13246 9628 13274
rect 9508 12850 9536 13246
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9600 12986 9628 13126
rect 9588 12980 9640 12986
rect 9588 12922 9640 12928
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9600 12730 9628 12922
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9324 12702 9628 12730
rect 9232 12238 9260 12650
rect 9220 12232 9272 12238
rect 9324 12220 9352 12702
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9404 12436 9456 12442
rect 9496 12436 9548 12442
rect 9456 12396 9496 12424
rect 9404 12378 9456 12384
rect 9496 12378 9548 12384
rect 9404 12232 9456 12238
rect 9324 12192 9404 12220
rect 9220 12174 9272 12180
rect 9404 12174 9456 12180
rect 9600 12186 9628 12582
rect 9692 12306 9720 13756
rect 10140 13738 10192 13744
rect 10152 13682 10180 13738
rect 10060 13654 10180 13682
rect 10060 13530 10088 13654
rect 10138 13560 10194 13569
rect 10048 13524 10100 13530
rect 10138 13495 10140 13504
rect 10048 13466 10100 13472
rect 10192 13495 10194 13504
rect 10140 13466 10192 13472
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9968 13297 9996 13398
rect 10244 13297 10272 13942
rect 10320 13628 10628 13648
rect 10320 13626 10326 13628
rect 10382 13626 10406 13628
rect 10462 13626 10486 13628
rect 10542 13626 10566 13628
rect 10622 13626 10628 13628
rect 10382 13574 10384 13626
rect 10564 13574 10566 13626
rect 10320 13572 10326 13574
rect 10382 13572 10406 13574
rect 10462 13572 10486 13574
rect 10542 13572 10566 13574
rect 10622 13572 10628 13574
rect 10320 13552 10628 13572
rect 10704 13530 10732 15438
rect 10692 13524 10744 13530
rect 10692 13466 10744 13472
rect 10796 13410 10824 16546
rect 11072 16538 11100 19230
rect 11256 19122 11284 19230
rect 11334 19200 11390 20000
rect 11794 19200 11850 20000
rect 12162 19200 12218 20000
rect 12530 19200 12586 20000
rect 12898 19200 12954 20000
rect 13266 19200 13322 20000
rect 13634 19200 13690 20000
rect 14002 19200 14058 20000
rect 14370 19200 14426 20000
rect 14738 19200 14794 20000
rect 15106 19200 15162 20000
rect 15474 19200 15530 20000
rect 15842 19200 15898 20000
rect 16210 19200 16266 20000
rect 16578 19200 16634 20000
rect 16946 19200 17002 20000
rect 11348 19122 11376 19200
rect 11256 19094 11376 19122
rect 11022 16510 11100 16538
rect 10966 16487 11022 16496
rect 11058 16008 11114 16017
rect 11058 15943 11114 15952
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10704 13382 10824 13410
rect 9954 13288 10010 13297
rect 9954 13223 10010 13232
rect 10230 13288 10286 13297
rect 10230 13223 10286 13232
rect 10244 13002 10272 13223
rect 10704 13190 10732 13382
rect 10888 13326 10916 15642
rect 11072 15065 11100 15943
rect 11808 15638 11836 19200
rect 12176 17626 12204 19200
rect 12084 17598 12204 17626
rect 11796 15632 11848 15638
rect 11796 15574 11848 15580
rect 11058 15056 11114 15065
rect 11058 14991 11114 15000
rect 12084 14822 12112 17598
rect 12194 17436 12502 17456
rect 12194 17434 12200 17436
rect 12256 17434 12280 17436
rect 12336 17434 12360 17436
rect 12416 17434 12440 17436
rect 12496 17434 12502 17436
rect 12256 17382 12258 17434
rect 12438 17382 12440 17434
rect 12194 17380 12200 17382
rect 12256 17380 12280 17382
rect 12336 17380 12360 17382
rect 12416 17380 12440 17382
rect 12496 17380 12502 17382
rect 12194 17360 12502 17380
rect 12194 16348 12502 16368
rect 12194 16346 12200 16348
rect 12256 16346 12280 16348
rect 12336 16346 12360 16348
rect 12416 16346 12440 16348
rect 12496 16346 12502 16348
rect 12256 16294 12258 16346
rect 12438 16294 12440 16346
rect 12194 16292 12200 16294
rect 12256 16292 12280 16294
rect 12336 16292 12360 16294
rect 12416 16292 12440 16294
rect 12496 16292 12502 16294
rect 12194 16272 12502 16292
rect 12544 15609 12572 19200
rect 12912 16114 12940 19200
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 12530 15600 12586 15609
rect 12530 15535 12586 15544
rect 12194 15260 12502 15280
rect 12194 15258 12200 15260
rect 12256 15258 12280 15260
rect 12336 15258 12360 15260
rect 12416 15258 12440 15260
rect 12496 15258 12502 15260
rect 12256 15206 12258 15258
rect 12438 15206 12440 15258
rect 12194 15204 12200 15206
rect 12256 15204 12280 15206
rect 12336 15204 12360 15206
rect 12416 15204 12440 15206
rect 12496 15204 12502 15206
rect 12194 15184 12502 15204
rect 12072 14816 12124 14822
rect 12072 14758 12124 14764
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 10784 13320 10836 13326
rect 10784 13262 10836 13268
rect 10876 13320 10928 13326
rect 10876 13262 10928 13268
rect 10600 13184 10652 13190
rect 10600 13126 10652 13132
rect 10692 13184 10744 13190
rect 10692 13126 10744 13132
rect 9968 12974 10272 13002
rect 9864 12912 9916 12918
rect 9864 12854 9916 12860
rect 9876 12782 9904 12854
rect 9864 12776 9916 12782
rect 9864 12718 9916 12724
rect 9772 12640 9824 12646
rect 9772 12582 9824 12588
rect 9680 12300 9732 12306
rect 9680 12242 9732 12248
rect 9678 12200 9734 12209
rect 9600 12158 9678 12186
rect 9678 12135 9734 12144
rect 9220 12096 9272 12102
rect 9588 12096 9640 12102
rect 9272 12056 9588 12084
rect 9220 12038 9272 12044
rect 9588 12038 9640 12044
rect 9126 11928 9182 11937
rect 9036 11892 9088 11898
rect 8956 11852 9036 11880
rect 9126 11863 9182 11872
rect 9036 11834 9088 11840
rect 9232 11801 9260 12038
rect 8942 11792 8998 11801
rect 8574 11727 8630 11736
rect 8668 11756 8720 11762
rect 8392 11144 8444 11150
rect 8588 11121 8616 11727
rect 8852 11756 8904 11762
rect 8720 11716 8800 11744
rect 8668 11698 8720 11704
rect 8772 11121 8800 11716
rect 8942 11727 8998 11736
rect 9218 11792 9274 11801
rect 9218 11727 9274 11736
rect 9588 11756 9640 11762
rect 8852 11698 8904 11704
rect 8956 11626 8984 11727
rect 9588 11698 9640 11704
rect 9310 11656 9366 11665
rect 8944 11620 8996 11626
rect 9310 11591 9366 11600
rect 8944 11562 8996 11568
rect 9034 11520 9090 11529
rect 9034 11455 9090 11464
rect 9048 11354 9076 11455
rect 9324 11354 9352 11591
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9416 11257 9444 11494
rect 9600 11336 9628 11698
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 9508 11308 9628 11336
rect 9402 11248 9458 11257
rect 8852 11212 8904 11218
rect 9402 11183 9458 11192
rect 8852 11154 8904 11160
rect 8392 11086 8444 11092
rect 8574 11112 8630 11121
rect 8574 11047 8630 11056
rect 8758 11112 8814 11121
rect 8758 11047 8814 11056
rect 8446 10908 8754 10928
rect 8446 10906 8452 10908
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8748 10906 8754 10908
rect 8508 10854 8510 10906
rect 8690 10854 8692 10906
rect 8446 10852 8452 10854
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8748 10852 8754 10854
rect 8446 10832 8754 10852
rect 8390 10568 8446 10577
rect 8390 10503 8446 10512
rect 8404 10470 8432 10503
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 9994 8432 10406
rect 8864 10130 8892 11154
rect 9220 11144 9272 11150
rect 9220 11086 9272 11092
rect 9036 11076 9088 11082
rect 9036 11018 9088 11024
rect 8942 10976 8998 10985
rect 8942 10911 8998 10920
rect 8956 10742 8984 10911
rect 9048 10826 9076 11018
rect 9048 10810 9168 10826
rect 9048 10804 9180 10810
rect 9048 10798 9128 10804
rect 9128 10746 9180 10752
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8956 9874 8984 9998
rect 8956 9846 9168 9874
rect 8446 9820 8754 9840
rect 8446 9818 8452 9820
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8748 9818 8754 9820
rect 8508 9766 8510 9818
rect 8690 9766 8692 9818
rect 8446 9764 8452 9766
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8748 9764 8754 9766
rect 8446 9744 8754 9764
rect 8850 9752 8906 9761
rect 8850 9687 8906 9696
rect 9034 9752 9090 9761
rect 9034 9687 9036 9696
rect 8668 9580 8720 9586
rect 8864 9568 8892 9687
rect 9088 9687 9090 9696
rect 9036 9658 9088 9664
rect 8720 9540 8892 9568
rect 9034 9616 9090 9625
rect 9140 9586 9168 9846
rect 9034 9551 9090 9560
rect 9128 9580 9180 9586
rect 8668 9522 8720 9528
rect 8944 9376 8996 9382
rect 8944 9318 8996 9324
rect 8392 9036 8444 9042
rect 8312 8996 8392 9024
rect 8392 8978 8444 8984
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8446 8732 8754 8752
rect 8446 8730 8452 8732
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8748 8730 8754 8732
rect 8508 8678 8510 8730
rect 8690 8678 8692 8730
rect 8446 8676 8452 8678
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8748 8676 8754 8678
rect 8446 8656 8754 8676
rect 8446 7644 8754 7664
rect 8446 7642 8452 7644
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8748 7642 8754 7644
rect 8508 7590 8510 7642
rect 8690 7590 8692 7642
rect 8446 7588 8452 7590
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8748 7588 8754 7590
rect 8446 7568 8754 7588
rect 8298 7304 8354 7313
rect 8208 7268 8260 7274
rect 8298 7239 8354 7248
rect 8208 7210 8260 7216
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8128 6089 8156 6394
rect 8114 6080 8170 6089
rect 8114 6015 8170 6024
rect 8220 5658 8248 7210
rect 8312 6905 8340 7239
rect 8864 6905 8892 8774
rect 8298 6896 8354 6905
rect 8298 6831 8354 6840
rect 8850 6896 8906 6905
rect 8850 6831 8906 6840
rect 8446 6556 8754 6576
rect 8446 6554 8452 6556
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8748 6554 8754 6556
rect 8508 6502 8510 6554
rect 8690 6502 8692 6554
rect 8446 6500 8452 6502
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8748 6500 8754 6502
rect 8446 6480 8754 6500
rect 8300 6452 8352 6458
rect 8956 6440 8984 9318
rect 9048 9178 9076 9551
rect 9128 9522 9180 9528
rect 9036 9172 9088 9178
rect 9036 9114 9088 9120
rect 9140 8974 9168 9522
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 9034 8800 9090 8809
rect 9034 8735 9090 8744
rect 9048 7818 9076 8735
rect 9140 8634 9168 8910
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9036 7812 9088 7818
rect 9036 7754 9088 7760
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8300 6394 8352 6400
rect 8680 6412 8984 6440
rect 8312 6225 8340 6394
rect 8484 6316 8536 6322
rect 8484 6258 8536 6264
rect 8298 6216 8354 6225
rect 8298 6151 8354 6160
rect 8496 5846 8524 6258
rect 8484 5840 8536 5846
rect 8536 5800 8616 5828
rect 8484 5782 8536 5788
rect 8220 5630 8340 5658
rect 8588 5642 8616 5800
rect 8680 5710 8708 6412
rect 9048 6338 9076 7346
rect 9126 7032 9182 7041
rect 9126 6967 9182 6976
rect 9140 6662 9168 6967
rect 9128 6656 9180 6662
rect 9128 6598 9180 6604
rect 8956 6310 9076 6338
rect 8850 6216 8906 6225
rect 8850 6151 8906 6160
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8022 4992 8078 5001
rect 8022 4927 8078 4936
rect 8036 4457 8064 4927
rect 8128 4826 8156 5170
rect 8220 4826 8248 5510
rect 8116 4820 8168 4826
rect 8116 4762 8168 4768
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 8022 4448 8078 4457
rect 8022 4383 8078 4392
rect 8036 4214 8064 4383
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7760 2746 7880 2774
rect 7760 2514 7788 2746
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7944 2446 7972 3538
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7932 2304 7984 2310
rect 7930 2272 7932 2281
rect 7984 2272 7986 2281
rect 7930 2207 7986 2216
rect 7668 1822 7788 1850
rect 7760 1766 7788 1822
rect 7656 1760 7708 1766
rect 7656 1702 7708 1708
rect 7748 1760 7800 1766
rect 7748 1702 7800 1708
rect 7564 1692 7616 1698
rect 7564 1634 7616 1640
rect 7668 1465 7696 1702
rect 8036 1544 8064 4150
rect 8128 4049 8156 4490
rect 8220 4321 8248 4490
rect 8206 4312 8262 4321
rect 8206 4247 8262 4256
rect 8114 4040 8170 4049
rect 8114 3975 8170 3984
rect 8220 3942 8248 4247
rect 8312 4154 8340 5630
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8446 5468 8754 5488
rect 8446 5466 8452 5468
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8748 5466 8754 5468
rect 8508 5414 8510 5466
rect 8690 5414 8692 5466
rect 8446 5412 8452 5414
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8748 5412 8754 5414
rect 8446 5392 8754 5412
rect 8864 5302 8892 6151
rect 8956 5778 8984 6310
rect 9232 6304 9260 11086
rect 9312 10600 9364 10606
rect 9508 10554 9536 11308
rect 9586 11248 9642 11257
rect 9586 11183 9642 11192
rect 9364 10548 9536 10554
rect 9312 10542 9536 10548
rect 9324 10526 9536 10542
rect 9310 10160 9366 10169
rect 9310 10095 9366 10104
rect 9324 7886 9352 10095
rect 9402 10024 9458 10033
rect 9402 9959 9458 9968
rect 9416 9178 9444 9959
rect 9600 9761 9628 11183
rect 9586 9752 9642 9761
rect 9586 9687 9642 9696
rect 9692 9382 9720 11630
rect 9784 11626 9812 12582
rect 9862 12472 9918 12481
rect 9862 12407 9918 12416
rect 9876 12306 9904 12407
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9864 12164 9916 12170
rect 9864 12106 9916 12112
rect 9876 11626 9904 12106
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9312 7880 9364 7886
rect 9312 7822 9364 7828
rect 9404 7812 9456 7818
rect 9404 7754 9456 7760
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 9324 6866 9352 7278
rect 9416 7274 9444 7754
rect 9508 7410 9536 8910
rect 9680 8900 9732 8906
rect 9680 8842 9732 8848
rect 9692 8809 9720 8842
rect 9678 8800 9734 8809
rect 9678 8735 9734 8744
rect 9784 8072 9812 11562
rect 9968 11506 9996 12974
rect 10612 12918 10640 13126
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10244 12434 10272 12854
rect 10612 12628 10640 12854
rect 10704 12782 10732 13126
rect 10692 12776 10744 12782
rect 10692 12718 10744 12724
rect 10692 12640 10744 12646
rect 10612 12600 10692 12628
rect 10692 12582 10744 12588
rect 10320 12540 10628 12560
rect 10320 12538 10326 12540
rect 10382 12538 10406 12540
rect 10462 12538 10486 12540
rect 10542 12538 10566 12540
rect 10622 12538 10628 12540
rect 10382 12486 10384 12538
rect 10564 12486 10566 12538
rect 10320 12484 10326 12486
rect 10382 12484 10406 12486
rect 10462 12484 10486 12486
rect 10542 12484 10566 12486
rect 10622 12484 10628 12486
rect 10320 12464 10628 12484
rect 10244 12406 10364 12434
rect 10046 12336 10102 12345
rect 10046 12271 10102 12280
rect 10060 12238 10088 12271
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 10048 11892 10100 11898
rect 10048 11834 10100 11840
rect 9876 11478 9996 11506
rect 9876 11150 9904 11478
rect 9954 11384 10010 11393
rect 9954 11319 10010 11328
rect 9864 11144 9916 11150
rect 9864 11086 9916 11092
rect 9876 9722 9904 11086
rect 9968 11082 9996 11319
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 10060 10810 10088 11834
rect 10230 11792 10286 11801
rect 10230 11727 10286 11736
rect 10244 11694 10272 11727
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10336 11540 10364 12406
rect 10692 12368 10744 12374
rect 10692 12310 10744 12316
rect 10598 12064 10654 12073
rect 10598 11999 10654 12008
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10428 11694 10456 11834
rect 10612 11762 10640 11999
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10138 11520 10194 11529
rect 10138 11455 10194 11464
rect 10244 11512 10364 11540
rect 10152 11354 10180 11455
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10152 10606 10180 10950
rect 10140 10600 10192 10606
rect 10138 10568 10140 10577
rect 10192 10568 10194 10577
rect 9956 10532 10008 10538
rect 10138 10503 10194 10512
rect 9956 10474 10008 10480
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9862 9616 9918 9625
rect 9968 9586 9996 10474
rect 10140 10464 10192 10470
rect 10138 10432 10140 10441
rect 10192 10432 10194 10441
rect 10138 10367 10194 10376
rect 10138 10296 10194 10305
rect 10138 10231 10140 10240
rect 10192 10231 10194 10240
rect 10140 10202 10192 10208
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 9862 9551 9918 9560
rect 9956 9580 10008 9586
rect 9876 8401 9904 9551
rect 9956 9522 10008 9528
rect 9956 9376 10008 9382
rect 9956 9318 10008 9324
rect 9862 8392 9918 8401
rect 9862 8327 9918 8336
rect 9968 8129 9996 9318
rect 10060 9081 10088 10134
rect 10244 9489 10272 11512
rect 10320 11452 10628 11472
rect 10320 11450 10326 11452
rect 10382 11450 10406 11452
rect 10462 11450 10486 11452
rect 10542 11450 10566 11452
rect 10622 11450 10628 11452
rect 10382 11398 10384 11450
rect 10564 11398 10566 11450
rect 10320 11396 10326 11398
rect 10382 11396 10406 11398
rect 10462 11396 10486 11398
rect 10542 11396 10566 11398
rect 10622 11396 10628 11398
rect 10320 11376 10628 11396
rect 10322 11248 10378 11257
rect 10322 11183 10324 11192
rect 10376 11183 10378 11192
rect 10598 11248 10654 11257
rect 10598 11183 10654 11192
rect 10324 11154 10376 11160
rect 10336 11014 10364 11154
rect 10612 11150 10640 11183
rect 10600 11144 10652 11150
rect 10600 11086 10652 11092
rect 10508 11076 10560 11082
rect 10508 11018 10560 11024
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10336 10606 10364 10950
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10520 10452 10548 11018
rect 10704 10554 10732 12310
rect 10796 10656 10824 13262
rect 10888 12374 10916 13262
rect 11058 12880 11114 12889
rect 11164 12850 11192 13738
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 11256 12889 11284 13194
rect 11242 12880 11298 12889
rect 11058 12815 11114 12824
rect 11152 12844 11204 12850
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10876 12368 10928 12374
rect 10980 12345 11008 12718
rect 10876 12310 10928 12316
rect 10966 12336 11022 12345
rect 10888 12170 10916 12310
rect 10966 12271 11022 12280
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 10888 11676 10916 12106
rect 10888 11648 11008 11676
rect 10876 11552 10928 11558
rect 10876 11494 10928 11500
rect 10888 10792 10916 11494
rect 10980 11082 11008 11648
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10968 10804 11020 10810
rect 10888 10764 10968 10792
rect 10968 10746 11020 10752
rect 10876 10668 10928 10674
rect 10796 10628 10876 10656
rect 10876 10610 10928 10616
rect 10704 10526 10824 10554
rect 10692 10464 10744 10470
rect 10520 10424 10692 10452
rect 10692 10406 10744 10412
rect 10320 10364 10628 10384
rect 10320 10362 10326 10364
rect 10382 10362 10406 10364
rect 10462 10362 10486 10364
rect 10542 10362 10566 10364
rect 10622 10362 10628 10364
rect 10382 10310 10384 10362
rect 10564 10310 10566 10362
rect 10320 10308 10326 10310
rect 10382 10308 10406 10310
rect 10462 10308 10486 10310
rect 10542 10308 10566 10310
rect 10622 10308 10628 10310
rect 10320 10288 10628 10308
rect 10796 10305 10824 10526
rect 10782 10296 10838 10305
rect 10782 10231 10838 10240
rect 10796 10130 10824 10231
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10600 10056 10652 10062
rect 10600 9998 10652 10004
rect 10690 10024 10746 10033
rect 10612 9926 10640 9998
rect 10690 9959 10746 9968
rect 10600 9920 10652 9926
rect 10600 9862 10652 9868
rect 10598 9616 10654 9625
rect 10598 9551 10654 9560
rect 10704 9568 10732 9959
rect 10612 9518 10640 9551
rect 10704 9540 10824 9568
rect 10600 9512 10652 9518
rect 10230 9480 10286 9489
rect 10600 9454 10652 9460
rect 10690 9480 10746 9489
rect 10230 9415 10286 9424
rect 10796 9450 10824 9540
rect 10690 9415 10746 9424
rect 10784 9444 10836 9450
rect 10704 9382 10732 9415
rect 10784 9386 10836 9392
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10320 9276 10628 9296
rect 10320 9274 10326 9276
rect 10382 9274 10406 9276
rect 10462 9274 10486 9276
rect 10542 9274 10566 9276
rect 10622 9274 10628 9276
rect 10382 9222 10384 9274
rect 10564 9222 10566 9274
rect 10320 9220 10326 9222
rect 10382 9220 10406 9222
rect 10462 9220 10486 9222
rect 10542 9220 10566 9222
rect 10622 9220 10628 9222
rect 10320 9200 10628 9220
rect 10704 9110 10732 9318
rect 10692 9104 10744 9110
rect 10046 9072 10102 9081
rect 10692 9046 10744 9052
rect 10046 9007 10102 9016
rect 10796 8974 10824 9386
rect 10508 8968 10560 8974
rect 10508 8910 10560 8916
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10232 8900 10284 8906
rect 10284 8860 10456 8888
rect 10232 8842 10284 8848
rect 10046 8664 10102 8673
rect 10046 8599 10102 8608
rect 10060 8265 10088 8599
rect 10428 8566 10456 8860
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10416 8560 10468 8566
rect 10416 8502 10468 8508
rect 10138 8392 10194 8401
rect 10138 8327 10194 8336
rect 10046 8256 10102 8265
rect 10046 8191 10102 8200
rect 9600 8044 9812 8072
rect 9954 8120 10010 8129
rect 9954 8055 10010 8064
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9404 7268 9456 7274
rect 9404 7210 9456 7216
rect 9494 7032 9550 7041
rect 9494 6967 9550 6976
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9140 6276 9260 6304
rect 9140 6202 9168 6276
rect 9324 6254 9352 6802
rect 9508 6662 9536 6967
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9496 6656 9548 6662
rect 9496 6598 9548 6604
rect 9416 6390 9444 6598
rect 9404 6384 9456 6390
rect 9456 6344 9536 6372
rect 9404 6326 9456 6332
rect 9312 6248 9364 6254
rect 9036 6180 9088 6186
rect 9140 6174 9229 6202
rect 9312 6190 9364 6196
rect 9402 6216 9458 6225
rect 9201 6168 9229 6174
rect 9201 6140 9260 6168
rect 9402 6151 9458 6160
rect 9036 6122 9088 6128
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8482 4856 8538 4865
rect 8482 4791 8538 4800
rect 8668 4820 8720 4826
rect 8496 4758 8524 4791
rect 8668 4762 8720 4768
rect 8484 4752 8536 4758
rect 8484 4694 8536 4700
rect 8680 4622 8708 4762
rect 8864 4690 8892 5238
rect 8852 4684 8904 4690
rect 8852 4626 8904 4632
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8956 4457 8984 5306
rect 8942 4448 8998 4457
rect 8446 4380 8754 4400
rect 8942 4383 8998 4392
rect 8446 4378 8452 4380
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8748 4378 8754 4380
rect 8508 4326 8510 4378
rect 8690 4326 8692 4378
rect 8446 4324 8452 4326
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8748 4324 8754 4326
rect 8446 4304 8754 4324
rect 8852 4276 8904 4282
rect 8852 4218 8904 4224
rect 8312 4146 8432 4154
rect 8312 4140 8444 4146
rect 8312 4126 8392 4140
rect 8392 4082 8444 4088
rect 8760 4140 8812 4146
rect 8760 4082 8812 4088
rect 8300 4072 8352 4078
rect 8300 4014 8352 4020
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8128 3097 8156 3538
rect 8114 3088 8170 3097
rect 8114 3023 8170 3032
rect 8312 2774 8340 4014
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8404 3670 8432 3878
rect 8772 3754 8800 4082
rect 8864 3942 8892 4218
rect 8852 3936 8904 3942
rect 8852 3878 8904 3884
rect 8956 3754 8984 4383
rect 9048 3942 9076 6122
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9140 5574 9168 6054
rect 9232 5778 9260 6140
rect 9312 6112 9364 6118
rect 9312 6054 9364 6060
rect 9220 5772 9272 5778
rect 9220 5714 9272 5720
rect 9218 5672 9274 5681
rect 9218 5607 9274 5616
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 9140 4826 9168 5510
rect 9232 5166 9260 5607
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9220 5024 9272 5030
rect 9220 4966 9272 4972
rect 9128 4820 9180 4826
rect 9128 4762 9180 4768
rect 9232 4729 9260 4966
rect 9218 4720 9274 4729
rect 9218 4655 9274 4664
rect 9324 4604 9352 6054
rect 9416 4622 9444 6151
rect 9140 4576 9352 4604
rect 9404 4616 9456 4622
rect 9036 3936 9088 3942
rect 9036 3878 9088 3884
rect 8668 3732 8720 3738
rect 8772 3726 8984 3754
rect 8668 3674 8720 3680
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8680 3466 8708 3674
rect 8760 3664 8812 3670
rect 8758 3632 8760 3641
rect 8812 3632 8814 3641
rect 8758 3567 8814 3576
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8446 3292 8754 3312
rect 8446 3290 8452 3292
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8748 3290 8754 3292
rect 8508 3238 8510 3290
rect 8690 3238 8692 3290
rect 8446 3236 8452 3238
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8748 3236 8754 3238
rect 8446 3216 8754 3236
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 8668 3052 8720 3058
rect 8668 2994 8720 3000
rect 8220 2746 8340 2774
rect 8036 1516 8156 1544
rect 7654 1456 7710 1465
rect 8128 1426 8156 1516
rect 7654 1391 7710 1400
rect 8024 1420 8076 1426
rect 7380 1080 7432 1086
rect 7380 1022 7432 1028
rect 7668 800 7696 1391
rect 8024 1362 8076 1368
rect 8116 1420 8168 1426
rect 8116 1362 8168 1368
rect 8220 1394 8248 2746
rect 8298 2680 8354 2689
rect 8298 2615 8354 2624
rect 8312 2514 8340 2615
rect 8404 2553 8432 2994
rect 8390 2544 8446 2553
rect 8300 2508 8352 2514
rect 8390 2479 8446 2488
rect 8484 2508 8536 2514
rect 8300 2450 8352 2456
rect 8484 2450 8536 2456
rect 8496 2378 8524 2450
rect 8680 2378 8708 2994
rect 8758 2952 8814 2961
rect 8758 2887 8760 2896
rect 8812 2887 8814 2896
rect 8760 2858 8812 2864
rect 8758 2680 8814 2689
rect 8758 2615 8760 2624
rect 8812 2615 8814 2624
rect 8760 2586 8812 2592
rect 8760 2508 8812 2514
rect 8760 2450 8812 2456
rect 8484 2372 8536 2378
rect 8484 2314 8536 2320
rect 8668 2372 8720 2378
rect 8668 2314 8720 2320
rect 8300 2304 8352 2310
rect 8772 2292 8800 2450
rect 8864 2394 8892 3538
rect 8956 3126 8984 3726
rect 9140 3618 9168 4576
rect 9404 4558 9456 4564
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9232 3738 9260 4422
rect 9220 3732 9272 3738
rect 9220 3674 9272 3680
rect 9140 3590 9260 3618
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 9048 3398 9076 3470
rect 9232 3398 9260 3590
rect 9036 3392 9088 3398
rect 9036 3334 9088 3340
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 9048 2650 9076 3334
rect 9218 3088 9274 3097
rect 9218 3023 9274 3032
rect 8944 2644 8996 2650
rect 8944 2586 8996 2592
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 8956 2496 8984 2586
rect 8956 2468 9076 2496
rect 8864 2378 8984 2394
rect 8864 2372 8996 2378
rect 8864 2366 8944 2372
rect 8944 2314 8996 2320
rect 8772 2264 8892 2292
rect 8300 2246 8352 2252
rect 8312 1970 8340 2246
rect 8446 2204 8754 2224
rect 8446 2202 8452 2204
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8748 2202 8754 2204
rect 8508 2150 8510 2202
rect 8690 2150 8692 2202
rect 8446 2148 8452 2150
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8748 2148 8754 2150
rect 8446 2128 8754 2148
rect 8864 2038 8892 2264
rect 8852 2032 8904 2038
rect 8852 1974 8904 1980
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 9048 1562 9076 2468
rect 9126 2408 9182 2417
rect 9126 2343 9182 2352
rect 9140 2310 9168 2343
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 8944 1556 8996 1562
rect 8944 1498 8996 1504
rect 9036 1556 9088 1562
rect 9036 1498 9088 1504
rect 8668 1420 8720 1426
rect 8220 1366 8340 1394
rect 8036 800 8064 1362
rect 8312 800 8340 1366
rect 8668 1362 8720 1368
rect 8680 800 8708 1362
rect 8956 1306 8984 1498
rect 9232 1329 9260 3023
rect 9324 2650 9352 4422
rect 9402 4312 9458 4321
rect 9402 4247 9458 4256
rect 9416 4214 9444 4247
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 9404 4004 9456 4010
rect 9404 3946 9456 3952
rect 9416 3777 9444 3946
rect 9402 3768 9458 3777
rect 9402 3703 9458 3712
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9416 2650 9444 3062
rect 9508 2922 9536 6344
rect 9600 5352 9628 8044
rect 9678 7984 9734 7993
rect 9678 7919 9734 7928
rect 9692 7002 9720 7919
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 9784 7410 9812 7822
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 9772 7404 9824 7410
rect 9956 7404 10008 7410
rect 9772 7346 9824 7352
rect 9876 7364 9956 7392
rect 9680 6996 9732 7002
rect 9680 6938 9732 6944
rect 9876 6848 9904 7364
rect 9956 7346 10008 7352
rect 10060 7041 10088 7482
rect 10152 7177 10180 8327
rect 10244 8276 10272 8502
rect 10520 8276 10548 8910
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10692 8424 10744 8430
rect 10796 8401 10824 8774
rect 10692 8366 10744 8372
rect 10782 8392 10838 8401
rect 10244 8248 10548 8276
rect 10244 7886 10272 8248
rect 10320 8188 10628 8208
rect 10320 8186 10326 8188
rect 10382 8186 10406 8188
rect 10462 8186 10486 8188
rect 10542 8186 10566 8188
rect 10622 8186 10628 8188
rect 10382 8134 10384 8186
rect 10564 8134 10566 8186
rect 10320 8132 10326 8134
rect 10382 8132 10406 8134
rect 10462 8132 10486 8134
rect 10542 8132 10566 8134
rect 10622 8132 10628 8134
rect 10320 8112 10628 8132
rect 10704 8090 10732 8366
rect 10782 8327 10838 8336
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10232 7880 10284 7886
rect 10232 7822 10284 7828
rect 10138 7168 10194 7177
rect 10138 7103 10194 7112
rect 10046 7032 10102 7041
rect 9956 6996 10008 7002
rect 10046 6967 10102 6976
rect 10244 6984 10272 7822
rect 10704 7818 10732 8026
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10690 7712 10746 7721
rect 10690 7647 10746 7656
rect 10704 7342 10732 7647
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10704 7206 10732 7237
rect 10692 7200 10744 7206
rect 10796 7154 10824 8026
rect 10744 7148 10824 7154
rect 10692 7142 10824 7148
rect 10704 7126 10824 7142
rect 10320 7100 10628 7120
rect 10320 7098 10326 7100
rect 10382 7098 10406 7100
rect 10462 7098 10486 7100
rect 10542 7098 10566 7100
rect 10622 7098 10628 7100
rect 10382 7046 10384 7098
rect 10564 7046 10566 7098
rect 10320 7044 10326 7046
rect 10382 7044 10406 7046
rect 10462 7044 10486 7046
rect 10542 7044 10566 7046
rect 10622 7044 10628 7046
rect 10320 7024 10628 7044
rect 10244 6956 10364 6984
rect 9956 6938 10008 6944
rect 9692 6820 9904 6848
rect 9692 6390 9720 6820
rect 9864 6724 9916 6730
rect 9864 6666 9916 6672
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9784 5794 9812 6598
rect 9876 6322 9904 6666
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 9692 5766 9812 5794
rect 9692 5574 9720 5766
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9600 5324 9720 5352
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9600 4486 9628 4966
rect 9692 4622 9720 5324
rect 9784 4865 9812 5510
rect 9876 5166 9904 6258
rect 9968 6089 9996 6938
rect 10336 6798 10364 6956
rect 10704 6866 10732 7126
rect 10782 7032 10838 7041
rect 10782 6967 10784 6976
rect 10836 6967 10838 6976
rect 10784 6938 10836 6944
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10232 6792 10284 6798
rect 10060 6752 10232 6780
rect 9954 6080 10010 6089
rect 9954 6015 10010 6024
rect 9968 5846 9996 6015
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 9954 5536 10010 5545
rect 9954 5471 10010 5480
rect 9864 5160 9916 5166
rect 9864 5102 9916 5108
rect 9862 4992 9918 5001
rect 9862 4927 9918 4936
rect 9770 4856 9826 4865
rect 9876 4826 9904 4927
rect 9770 4791 9826 4800
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9588 4480 9640 4486
rect 9692 4468 9720 4558
rect 9692 4440 9812 4468
rect 9588 4422 9640 4428
rect 9588 4072 9640 4078
rect 9586 4040 9588 4049
rect 9640 4040 9642 4049
rect 9586 3975 9642 3984
rect 9678 3768 9734 3777
rect 9588 3732 9640 3738
rect 9678 3703 9734 3712
rect 9588 3674 9640 3680
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9312 2644 9364 2650
rect 9312 2586 9364 2592
rect 9404 2644 9456 2650
rect 9404 2586 9456 2592
rect 9310 2544 9366 2553
rect 9310 2479 9366 2488
rect 9324 2310 9352 2479
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9600 1465 9628 3674
rect 9692 3670 9720 3703
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9784 3516 9812 4440
rect 9968 4321 9996 5471
rect 9954 4312 10010 4321
rect 9954 4247 10010 4256
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 9968 3942 9996 4014
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 9864 3664 9916 3670
rect 9862 3632 9864 3641
rect 9916 3632 9918 3641
rect 9862 3567 9918 3576
rect 9692 3488 9812 3516
rect 9692 2496 9720 3488
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9784 2564 9812 3334
rect 9784 2536 9904 2564
rect 9692 2468 9812 2496
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 9692 1902 9720 2314
rect 9784 1902 9812 2468
rect 9876 2378 9904 2536
rect 9968 2514 9996 3878
rect 10060 3534 10088 6752
rect 10232 6734 10284 6740
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10888 6746 10916 10610
rect 10966 10432 11022 10441
rect 10966 10367 11022 10376
rect 10980 9897 11008 10367
rect 10966 9888 11022 9897
rect 10966 9823 11022 9832
rect 10966 9208 11022 9217
rect 10966 9143 11022 9152
rect 10980 7546 11008 9143
rect 11072 8974 11100 12815
rect 11242 12815 11298 12824
rect 11152 12786 11204 12792
rect 11152 12300 11204 12306
rect 11204 12260 11284 12288
rect 11152 12242 11204 12248
rect 11150 12200 11206 12209
rect 11150 12135 11206 12144
rect 11164 11762 11192 12135
rect 11256 11762 11284 12260
rect 11152 11756 11204 11762
rect 11152 11698 11204 11704
rect 11244 11756 11296 11762
rect 11244 11698 11296 11704
rect 11256 11642 11284 11698
rect 11164 11614 11284 11642
rect 11164 11082 11192 11614
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11256 10962 11284 11494
rect 11164 10934 11284 10962
rect 11164 10674 11192 10934
rect 11242 10704 11298 10713
rect 11152 10668 11204 10674
rect 11242 10639 11298 10648
rect 11152 10610 11204 10616
rect 11256 10266 11284 10639
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11152 9920 11204 9926
rect 11150 9888 11152 9897
rect 11204 9888 11206 9897
rect 11150 9823 11206 9832
rect 11150 9616 11206 9625
rect 11150 9551 11206 9560
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 11060 8288 11112 8294
rect 11060 8230 11112 8236
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 10968 7336 11020 7342
rect 11072 7313 11100 8230
rect 11164 7546 11192 9551
rect 11242 9480 11298 9489
rect 11242 9415 11298 9424
rect 11256 9178 11284 9415
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11256 8634 11284 8774
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11242 7848 11298 7857
rect 11242 7783 11298 7792
rect 11256 7750 11284 7783
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11244 7472 11296 7478
rect 11150 7440 11206 7449
rect 11244 7414 11296 7420
rect 11150 7375 11152 7384
rect 11204 7375 11206 7384
rect 11152 7346 11204 7352
rect 11256 7342 11284 7414
rect 11244 7336 11296 7342
rect 10968 7278 11020 7284
rect 11058 7304 11114 7313
rect 10980 6934 11008 7278
rect 11114 7262 11192 7290
rect 11244 7278 11296 7284
rect 11058 7239 11114 7248
rect 11164 7206 11192 7262
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 11152 7200 11204 7206
rect 11348 7177 11376 13330
rect 11426 13152 11482 13161
rect 11426 13087 11482 13096
rect 11440 11014 11468 13087
rect 11532 12832 11560 13466
rect 11612 13252 11664 13258
rect 11612 13194 11664 13200
rect 11624 12986 11652 13194
rect 11612 12980 11664 12986
rect 11612 12922 11664 12928
rect 11532 12804 11652 12832
rect 11520 12708 11572 12714
rect 11520 12650 11572 12656
rect 11532 12170 11560 12650
rect 11624 12374 11652 12804
rect 11716 12714 11744 14418
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 11808 12986 11836 14350
rect 12084 13569 12112 14758
rect 12194 14172 12502 14192
rect 12194 14170 12200 14172
rect 12256 14170 12280 14172
rect 12336 14170 12360 14172
rect 12416 14170 12440 14172
rect 12496 14170 12502 14172
rect 12256 14118 12258 14170
rect 12438 14118 12440 14170
rect 12194 14116 12200 14118
rect 12256 14116 12280 14118
rect 12336 14116 12360 14118
rect 12416 14116 12440 14118
rect 12496 14116 12502 14118
rect 12194 14096 12502 14116
rect 12070 13560 12126 13569
rect 12070 13495 12126 13504
rect 12070 13424 12126 13433
rect 12070 13359 12126 13368
rect 11796 12980 11848 12986
rect 11796 12922 11848 12928
rect 11808 12714 11836 12922
rect 11886 12744 11942 12753
rect 11704 12708 11756 12714
rect 11704 12650 11756 12656
rect 11796 12708 11848 12714
rect 11886 12679 11942 12688
rect 11796 12650 11848 12656
rect 11612 12368 11664 12374
rect 11612 12310 11664 12316
rect 11520 12164 11572 12170
rect 11572 12124 11652 12152
rect 11520 12106 11572 12112
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11532 11801 11560 11834
rect 11518 11792 11574 11801
rect 11518 11727 11574 11736
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11532 11286 11560 11630
rect 11520 11280 11572 11286
rect 11520 11222 11572 11228
rect 11624 11218 11652 12124
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11518 11112 11574 11121
rect 11518 11047 11574 11056
rect 11612 11076 11664 11082
rect 11428 11008 11480 11014
rect 11428 10950 11480 10956
rect 11532 10810 11560 11047
rect 11612 11018 11664 11024
rect 11520 10804 11572 10810
rect 11520 10746 11572 10752
rect 11624 10690 11652 11018
rect 11716 11014 11744 12650
rect 11808 12442 11836 12650
rect 11796 12436 11848 12442
rect 11796 12378 11848 12384
rect 11796 12096 11848 12102
rect 11794 12064 11796 12073
rect 11848 12064 11850 12073
rect 11794 11999 11850 12008
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11716 10849 11744 10950
rect 11702 10840 11758 10849
rect 11702 10775 11758 10784
rect 11532 10662 11652 10690
rect 11532 10470 11560 10662
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11440 9586 11468 9658
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11152 7142 11204 7148
rect 11334 7168 11390 7177
rect 10968 6928 11020 6934
rect 10968 6870 11020 6876
rect 10888 6730 11008 6746
rect 10416 6724 10468 6730
rect 10888 6724 11020 6730
rect 10888 6718 10968 6724
rect 10416 6666 10468 6672
rect 10968 6666 11020 6672
rect 10140 6384 10192 6390
rect 10140 6326 10192 6332
rect 10152 5953 10180 6326
rect 10428 6100 10456 6666
rect 10600 6656 10652 6662
rect 10876 6656 10928 6662
rect 10652 6616 10732 6644
rect 10600 6598 10652 6604
rect 10244 6072 10456 6100
rect 10138 5944 10194 5953
rect 10138 5879 10194 5888
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10152 4146 10180 5782
rect 10244 5166 10272 6072
rect 10320 6012 10628 6032
rect 10320 6010 10326 6012
rect 10382 6010 10406 6012
rect 10462 6010 10486 6012
rect 10542 6010 10566 6012
rect 10622 6010 10628 6012
rect 10382 5958 10384 6010
rect 10564 5958 10566 6010
rect 10320 5956 10326 5958
rect 10382 5956 10406 5958
rect 10462 5956 10486 5958
rect 10542 5956 10566 5958
rect 10622 5956 10628 5958
rect 10320 5936 10628 5956
rect 10704 5930 10732 6616
rect 10876 6598 10928 6604
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10796 6254 10824 6394
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10784 6112 10836 6118
rect 10782 6080 10784 6089
rect 10836 6080 10838 6089
rect 10782 6015 10838 6024
rect 10782 5944 10838 5953
rect 10704 5902 10782 5930
rect 10782 5879 10838 5888
rect 10690 5672 10746 5681
rect 10690 5607 10746 5616
rect 10508 5568 10560 5574
rect 10508 5510 10560 5516
rect 10598 5536 10654 5545
rect 10324 5296 10376 5302
rect 10322 5264 10324 5273
rect 10416 5296 10468 5302
rect 10376 5264 10378 5273
rect 10416 5238 10468 5244
rect 10322 5199 10378 5208
rect 10232 5160 10284 5166
rect 10428 5137 10456 5238
rect 10520 5234 10548 5510
rect 10598 5471 10654 5480
rect 10612 5370 10640 5471
rect 10600 5364 10652 5370
rect 10600 5306 10652 5312
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10232 5102 10284 5108
rect 10414 5128 10470 5137
rect 10244 4321 10272 5102
rect 10414 5063 10470 5072
rect 10320 4924 10628 4944
rect 10320 4922 10326 4924
rect 10382 4922 10406 4924
rect 10462 4922 10486 4924
rect 10542 4922 10566 4924
rect 10622 4922 10628 4924
rect 10382 4870 10384 4922
rect 10564 4870 10566 4922
rect 10320 4868 10326 4870
rect 10382 4868 10406 4870
rect 10462 4868 10486 4870
rect 10542 4868 10566 4870
rect 10622 4868 10628 4870
rect 10320 4848 10628 4868
rect 10324 4684 10376 4690
rect 10704 4672 10732 5607
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10796 4826 10824 5510
rect 10888 5352 10916 6598
rect 10980 6236 11008 6666
rect 11072 6372 11100 7142
rect 11334 7103 11390 7112
rect 11152 6996 11204 7002
rect 11152 6938 11204 6944
rect 11164 6497 11192 6938
rect 11336 6928 11388 6934
rect 11336 6870 11388 6876
rect 11242 6760 11298 6769
rect 11242 6695 11298 6704
rect 11150 6488 11206 6497
rect 11150 6423 11206 6432
rect 11072 6344 11192 6372
rect 11164 6254 11192 6344
rect 11152 6248 11204 6254
rect 10980 6208 11100 6236
rect 10968 6112 11020 6118
rect 11072 6089 11100 6208
rect 11152 6190 11204 6196
rect 10968 6054 11020 6060
rect 11058 6080 11114 6089
rect 10980 5710 11008 6054
rect 11058 6015 11114 6024
rect 11058 5944 11114 5953
rect 11058 5879 11114 5888
rect 11072 5778 11100 5879
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 10968 5704 11020 5710
rect 11256 5681 11284 6695
rect 10968 5646 11020 5652
rect 11242 5672 11298 5681
rect 11242 5607 11298 5616
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11256 5409 11284 5510
rect 11242 5400 11298 5409
rect 10888 5324 11192 5352
rect 11242 5335 11298 5344
rect 11060 5228 11112 5234
rect 11164 5216 11192 5324
rect 11164 5188 11284 5216
rect 11060 5170 11112 5176
rect 10966 4992 11022 5001
rect 10966 4927 11022 4936
rect 10874 4856 10930 4865
rect 10784 4820 10836 4826
rect 10874 4791 10930 4800
rect 10784 4762 10836 4768
rect 10784 4684 10836 4690
rect 10704 4644 10784 4672
rect 10324 4626 10376 4632
rect 10784 4626 10836 4632
rect 10230 4312 10286 4321
rect 10230 4247 10286 4256
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10244 3720 10272 4247
rect 10336 4214 10364 4626
rect 10508 4616 10560 4622
rect 10888 4570 10916 4791
rect 10980 4622 11008 4927
rect 10560 4564 10916 4570
rect 10508 4558 10916 4564
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10416 4548 10468 4554
rect 10520 4542 10916 4558
rect 10416 4490 10468 4496
rect 10428 4264 10456 4490
rect 10508 4276 10560 4282
rect 10428 4236 10508 4264
rect 10508 4218 10560 4224
rect 11072 4214 11100 5170
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11164 4298 11192 4762
rect 11256 4690 11284 5188
rect 11244 4684 11296 4690
rect 11244 4626 11296 4632
rect 11242 4584 11298 4593
rect 11242 4519 11298 4528
rect 11256 4486 11284 4519
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11164 4270 11284 4298
rect 11256 4214 11284 4270
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 10336 4049 10364 4150
rect 10692 4072 10744 4078
rect 10322 4040 10378 4049
rect 10874 4040 10930 4049
rect 10744 4020 10874 4026
rect 10692 4014 10874 4020
rect 10704 3998 10874 4014
rect 10322 3975 10378 3984
rect 10874 3975 10930 3984
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10320 3836 10628 3856
rect 10320 3834 10326 3836
rect 10382 3834 10406 3836
rect 10462 3834 10486 3836
rect 10542 3834 10566 3836
rect 10622 3834 10628 3836
rect 10382 3782 10384 3834
rect 10564 3782 10566 3834
rect 10320 3780 10326 3782
rect 10382 3780 10406 3782
rect 10462 3780 10486 3782
rect 10542 3780 10566 3782
rect 10622 3780 10628 3782
rect 10320 3760 10628 3780
rect 11072 3720 11100 3946
rect 10244 3692 10364 3720
rect 10230 3632 10286 3641
rect 10230 3567 10286 3576
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10244 3126 10272 3567
rect 10232 3120 10284 3126
rect 10232 3062 10284 3068
rect 10336 3058 10364 3692
rect 10888 3692 11100 3720
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10428 3556 10640 3584
rect 10428 3097 10456 3556
rect 10506 3496 10562 3505
rect 10506 3431 10562 3440
rect 10520 3398 10548 3431
rect 10612 3398 10640 3556
rect 10508 3392 10560 3398
rect 10508 3334 10560 3340
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10704 3097 10732 3606
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10414 3088 10470 3097
rect 10324 3052 10376 3058
rect 10414 3023 10470 3032
rect 10690 3088 10746 3097
rect 10796 3058 10824 3334
rect 10690 3023 10746 3032
rect 10784 3052 10836 3058
rect 10324 2994 10376 3000
rect 10784 2994 10836 3000
rect 10600 2984 10652 2990
rect 10138 2952 10194 2961
rect 10138 2887 10194 2896
rect 10598 2952 10600 2961
rect 10692 2984 10744 2990
rect 10652 2952 10654 2961
rect 10692 2926 10744 2932
rect 10598 2887 10654 2896
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10060 2650 10088 2790
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10046 2544 10102 2553
rect 9956 2508 10008 2514
rect 10046 2479 10048 2488
rect 9956 2450 10008 2456
rect 10100 2479 10102 2488
rect 10048 2450 10100 2456
rect 9864 2372 9916 2378
rect 9864 2314 9916 2320
rect 9680 1896 9732 1902
rect 9680 1838 9732 1844
rect 9772 1896 9824 1902
rect 9772 1838 9824 1844
rect 10048 1896 10100 1902
rect 10048 1838 10100 1844
rect 9680 1556 9732 1562
rect 9680 1498 9732 1504
rect 9586 1456 9642 1465
rect 9586 1391 9642 1400
rect 9218 1320 9274 1329
rect 8956 1278 9076 1306
rect 9048 800 9076 1278
rect 9218 1255 9274 1264
rect 9232 836 9352 864
rect 6828 264 6880 270
rect 6734 232 6790 241
rect 6828 206 6880 212
rect 6734 167 6790 176
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7654 0 7710 800
rect 8022 0 8078 800
rect 8298 0 8354 800
rect 8666 0 8722 800
rect 9034 0 9090 800
rect 9126 776 9182 785
rect 9232 762 9260 836
rect 9324 800 9352 836
rect 9692 800 9720 1498
rect 10060 800 10088 1838
rect 10152 1562 10180 2887
rect 10695 2836 10723 2926
rect 10695 2808 10732 2836
rect 10320 2748 10628 2768
rect 10320 2746 10326 2748
rect 10382 2746 10406 2748
rect 10462 2746 10486 2748
rect 10542 2746 10566 2748
rect 10622 2746 10628 2748
rect 10382 2694 10384 2746
rect 10564 2694 10566 2746
rect 10320 2692 10326 2694
rect 10382 2692 10406 2694
rect 10462 2692 10486 2694
rect 10542 2692 10566 2694
rect 10622 2692 10628 2694
rect 10320 2672 10628 2692
rect 10322 2544 10378 2553
rect 10322 2479 10378 2488
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10140 1556 10192 1562
rect 10140 1498 10192 1504
rect 10244 950 10272 2382
rect 10336 2378 10364 2479
rect 10704 2394 10732 2808
rect 10782 2816 10838 2825
rect 10782 2751 10838 2760
rect 10324 2372 10376 2378
rect 10324 2314 10376 2320
rect 10520 2366 10732 2394
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 10232 944 10284 950
rect 10232 886 10284 892
rect 10428 800 10456 2246
rect 10520 1630 10548 2366
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10508 1624 10560 1630
rect 10508 1566 10560 1572
rect 10612 1494 10640 2246
rect 10692 1624 10744 1630
rect 10692 1566 10744 1572
rect 10600 1488 10652 1494
rect 10600 1430 10652 1436
rect 10704 1086 10732 1566
rect 10796 1494 10824 2751
rect 10784 1488 10836 1494
rect 10784 1430 10836 1436
rect 10692 1080 10744 1086
rect 10692 1022 10744 1028
rect 10704 800 10732 1022
rect 10888 814 10916 3692
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10980 3233 11008 3538
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 10966 3224 11022 3233
rect 11072 3194 11100 3470
rect 10966 3159 11022 3168
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 10980 2582 11008 2790
rect 11072 2689 11100 2994
rect 11058 2680 11114 2689
rect 11058 2615 11114 2624
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 11060 2508 11112 2514
rect 11164 2496 11192 4150
rect 11244 3732 11296 3738
rect 11244 3674 11296 3680
rect 11256 3602 11284 3674
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11244 3392 11296 3398
rect 11244 3334 11296 3340
rect 11256 3233 11284 3334
rect 11242 3224 11298 3233
rect 11242 3159 11298 3168
rect 11348 2632 11376 6870
rect 11440 6118 11468 9522
rect 11532 9353 11560 10406
rect 11716 10130 11744 10542
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11704 9920 11756 9926
rect 11610 9888 11666 9897
rect 11704 9862 11756 9868
rect 11610 9823 11666 9832
rect 11518 9344 11574 9353
rect 11518 9279 11574 9288
rect 11520 8628 11572 8634
rect 11520 8570 11572 8576
rect 11532 8537 11560 8570
rect 11518 8528 11574 8537
rect 11624 8498 11652 9823
rect 11716 9178 11744 9862
rect 11808 9450 11836 11766
rect 11900 10810 11928 12679
rect 11978 12472 12034 12481
rect 11978 12407 11980 12416
rect 12032 12407 12034 12416
rect 11980 12378 12032 12384
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11992 11830 12020 12242
rect 11980 11824 12032 11830
rect 11980 11766 12032 11772
rect 11980 11688 12032 11694
rect 11978 11656 11980 11665
rect 12032 11656 12034 11665
rect 11978 11591 12034 11600
rect 11978 11384 12034 11393
rect 11978 11319 11980 11328
rect 12032 11319 12034 11328
rect 11980 11290 12032 11296
rect 11978 11248 12034 11257
rect 11978 11183 12034 11192
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11900 10130 11928 10474
rect 11992 10470 12020 11183
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11980 10192 12032 10198
rect 11980 10134 12032 10140
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11886 10024 11942 10033
rect 11886 9959 11942 9968
rect 11900 9518 11928 9959
rect 11992 9897 12020 10134
rect 12084 9926 12112 13359
rect 12194 13084 12502 13104
rect 12194 13082 12200 13084
rect 12256 13082 12280 13084
rect 12336 13082 12360 13084
rect 12416 13082 12440 13084
rect 12496 13082 12502 13084
rect 12256 13030 12258 13082
rect 12438 13030 12440 13082
rect 12194 13028 12200 13030
rect 12256 13028 12280 13030
rect 12336 13028 12360 13030
rect 12416 13028 12440 13030
rect 12496 13028 12502 13030
rect 12194 13008 12502 13028
rect 12544 12889 12572 15535
rect 12808 14952 12860 14958
rect 12808 14894 12860 14900
rect 12624 14544 12676 14550
rect 12624 14486 12676 14492
rect 12530 12880 12586 12889
rect 12530 12815 12586 12824
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12348 12640 12400 12646
rect 12348 12582 12400 12588
rect 12360 12374 12388 12582
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 12452 12084 12480 12378
rect 12544 12306 12572 12650
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12636 12102 12664 14486
rect 12714 13288 12770 13297
rect 12714 13223 12770 13232
rect 12624 12096 12676 12102
rect 12452 12056 12572 12084
rect 12194 11996 12502 12016
rect 12194 11994 12200 11996
rect 12256 11994 12280 11996
rect 12336 11994 12360 11996
rect 12416 11994 12440 11996
rect 12496 11994 12502 11996
rect 12256 11942 12258 11994
rect 12438 11942 12440 11994
rect 12194 11940 12200 11942
rect 12256 11940 12280 11942
rect 12336 11940 12360 11942
rect 12416 11940 12440 11942
rect 12496 11940 12502 11942
rect 12194 11920 12502 11940
rect 12440 11824 12492 11830
rect 12440 11766 12492 11772
rect 12348 11688 12400 11694
rect 12162 11656 12218 11665
rect 12348 11630 12400 11636
rect 12162 11591 12218 11600
rect 12176 11286 12204 11591
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12164 11280 12216 11286
rect 12164 11222 12216 11228
rect 12268 11082 12296 11494
rect 12360 11150 12388 11630
rect 12452 11354 12480 11766
rect 12544 11694 12572 12056
rect 12622 12064 12624 12073
rect 12676 12064 12678 12073
rect 12622 11999 12678 12008
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12622 11384 12678 11393
rect 12440 11348 12492 11354
rect 12728 11354 12756 13223
rect 12820 11393 12848 14894
rect 12912 12481 12940 16050
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 12898 12472 12954 12481
rect 12898 12407 12954 12416
rect 12898 12200 12954 12209
rect 12898 12135 12954 12144
rect 12912 11898 12940 12135
rect 12900 11892 12952 11898
rect 12900 11834 12952 11840
rect 12806 11384 12862 11393
rect 12622 11319 12678 11328
rect 12716 11348 12768 11354
rect 12440 11290 12492 11296
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12256 11076 12308 11082
rect 12256 11018 12308 11024
rect 12360 10996 12388 11086
rect 12360 10968 12572 10996
rect 12194 10908 12502 10928
rect 12194 10906 12200 10908
rect 12256 10906 12280 10908
rect 12336 10906 12360 10908
rect 12416 10906 12440 10908
rect 12496 10906 12502 10908
rect 12256 10854 12258 10906
rect 12438 10854 12440 10906
rect 12194 10852 12200 10854
rect 12256 10852 12280 10854
rect 12336 10852 12360 10854
rect 12416 10852 12440 10854
rect 12496 10852 12502 10854
rect 12194 10832 12502 10852
rect 12544 10792 12572 10968
rect 12360 10764 12572 10792
rect 12360 10606 12388 10764
rect 12438 10704 12494 10713
rect 12438 10639 12440 10648
rect 12492 10639 12494 10648
rect 12440 10610 12492 10616
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12636 10248 12664 11319
rect 12912 11354 12940 11834
rect 13004 11354 13032 14350
rect 13096 11830 13124 17002
rect 13280 13734 13308 19200
rect 13648 17954 13676 19200
rect 13556 17926 13676 17954
rect 13556 16574 13584 17926
rect 13912 17876 13964 17882
rect 13912 17818 13964 17824
rect 13372 16546 13584 16574
rect 13268 13728 13320 13734
rect 13268 13670 13320 13676
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 13084 11824 13136 11830
rect 13084 11766 13136 11772
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 12806 11319 12862 11328
rect 12900 11348 12952 11354
rect 12716 11290 12768 11296
rect 12900 11290 12952 11296
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12728 10470 12756 11290
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12898 11112 12954 11121
rect 12716 10464 12768 10470
rect 12716 10406 12768 10412
rect 12544 10220 12664 10248
rect 12716 10260 12768 10266
rect 12072 9920 12124 9926
rect 11978 9888 12034 9897
rect 12072 9862 12124 9868
rect 11978 9823 12034 9832
rect 12194 9820 12502 9840
rect 12194 9818 12200 9820
rect 12256 9818 12280 9820
rect 12336 9818 12360 9820
rect 12416 9818 12440 9820
rect 12496 9818 12502 9820
rect 12256 9766 12258 9818
rect 12438 9766 12440 9818
rect 12194 9764 12200 9766
rect 12256 9764 12280 9766
rect 12336 9764 12360 9766
rect 12416 9764 12440 9766
rect 12496 9764 12502 9766
rect 12194 9744 12502 9764
rect 12544 9722 12572 10220
rect 12716 10202 12768 10208
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 11796 9444 11848 9450
rect 11796 9386 11848 9392
rect 11886 9344 11942 9353
rect 11942 9302 12020 9330
rect 11886 9279 11942 9288
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11888 9036 11940 9042
rect 11888 8978 11940 8984
rect 11796 8968 11848 8974
rect 11716 8928 11796 8956
rect 11716 8566 11744 8928
rect 11796 8910 11848 8916
rect 11794 8800 11850 8809
rect 11794 8735 11850 8744
rect 11808 8634 11836 8735
rect 11796 8628 11848 8634
rect 11796 8570 11848 8576
rect 11704 8560 11756 8566
rect 11704 8502 11756 8508
rect 11518 8463 11574 8472
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11518 7848 11574 7857
rect 11518 7783 11574 7792
rect 11532 7274 11560 7783
rect 11520 7268 11572 7274
rect 11520 7210 11572 7216
rect 11520 6860 11572 6866
rect 11520 6802 11572 6808
rect 11532 6497 11560 6802
rect 11624 6798 11652 8434
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 11716 6644 11744 8230
rect 11808 7886 11836 8366
rect 11900 8129 11928 8978
rect 11992 8401 12020 9302
rect 12084 8974 12112 9454
rect 12452 9217 12480 9590
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 12438 9208 12494 9217
rect 12438 9143 12494 9152
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 12176 8820 12204 8910
rect 12084 8792 12204 8820
rect 11978 8392 12034 8401
rect 11978 8327 12034 8336
rect 11886 8120 11942 8129
rect 11886 8055 11942 8064
rect 11796 7880 11848 7886
rect 11796 7822 11848 7828
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11808 6866 11836 7686
rect 11900 7002 11928 7686
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11992 7177 12020 7346
rect 11978 7168 12034 7177
rect 11978 7103 12034 7112
rect 11888 6996 11940 7002
rect 11888 6938 11940 6944
rect 11796 6860 11848 6866
rect 11796 6802 11848 6808
rect 11888 6860 11940 6866
rect 11888 6802 11940 6808
rect 11624 6616 11744 6644
rect 11796 6656 11848 6662
rect 11518 6488 11574 6497
rect 11518 6423 11574 6432
rect 11520 6384 11572 6390
rect 11520 6326 11572 6332
rect 11532 6168 11560 6326
rect 11624 6322 11652 6616
rect 11796 6598 11848 6604
rect 11702 6488 11758 6497
rect 11702 6423 11758 6432
rect 11716 6322 11744 6423
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11704 6316 11756 6322
rect 11704 6258 11756 6264
rect 11612 6180 11664 6186
rect 11532 6140 11612 6168
rect 11612 6122 11664 6128
rect 11428 6112 11480 6118
rect 11716 6066 11744 6258
rect 11428 6054 11480 6060
rect 11624 6038 11744 6066
rect 11624 5710 11652 6038
rect 11808 5914 11836 6598
rect 11900 6066 11928 6802
rect 12084 6712 12112 8792
rect 12194 8732 12502 8752
rect 12194 8730 12200 8732
rect 12256 8730 12280 8732
rect 12336 8730 12360 8732
rect 12416 8730 12440 8732
rect 12496 8730 12502 8732
rect 12256 8678 12258 8730
rect 12438 8678 12440 8730
rect 12194 8676 12200 8678
rect 12256 8676 12280 8678
rect 12336 8676 12360 8678
rect 12416 8676 12440 8678
rect 12496 8676 12502 8678
rect 12194 8656 12502 8676
rect 12164 8560 12216 8566
rect 12162 8528 12164 8537
rect 12544 8537 12572 9522
rect 12216 8528 12218 8537
rect 12530 8528 12586 8537
rect 12162 8463 12218 8472
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12348 8492 12400 8498
rect 12530 8463 12586 8472
rect 12348 8434 12400 8440
rect 12268 8090 12296 8434
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12360 7954 12388 8434
rect 12636 8430 12664 10066
rect 12728 9042 12756 10202
rect 12820 9926 12848 11086
rect 12898 11047 12954 11056
rect 12912 11014 12940 11047
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 13004 10810 13032 11290
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 12898 10704 12954 10713
rect 12954 10662 13032 10690
rect 12898 10639 12954 10648
rect 12898 10568 12954 10577
rect 12898 10503 12954 10512
rect 12808 9920 12860 9926
rect 12808 9862 12860 9868
rect 12820 9194 12848 9862
rect 12912 9518 12940 10503
rect 13004 9586 13032 10662
rect 13096 10130 13124 11494
rect 13188 11150 13216 13126
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13176 11144 13228 11150
rect 13176 11086 13228 11092
rect 13188 10810 13216 11086
rect 13176 10804 13228 10810
rect 13176 10746 13228 10752
rect 13084 10124 13136 10130
rect 13084 10066 13136 10072
rect 13188 10062 13216 10746
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13280 9761 13308 12174
rect 13372 12170 13400 16546
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13544 12436 13596 12442
rect 13544 12378 13596 12384
rect 13452 12368 13504 12374
rect 13452 12310 13504 12316
rect 13360 12164 13412 12170
rect 13360 12106 13412 12112
rect 13372 11762 13400 12106
rect 13464 12102 13492 12310
rect 13556 12220 13584 12378
rect 13648 12322 13676 14282
rect 13832 12442 13860 15914
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 13648 12294 13768 12322
rect 13556 12192 13676 12220
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13372 11257 13400 11494
rect 13358 11248 13414 11257
rect 13464 11218 13492 12038
rect 13542 11384 13598 11393
rect 13542 11319 13544 11328
rect 13596 11319 13598 11328
rect 13544 11290 13596 11296
rect 13358 11183 13414 11192
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 13372 10742 13400 10950
rect 13450 10840 13506 10849
rect 13450 10775 13506 10784
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13372 9994 13400 10678
rect 13464 10674 13492 10775
rect 13452 10668 13504 10674
rect 13452 10610 13504 10616
rect 13452 10532 13504 10538
rect 13452 10474 13504 10480
rect 13464 10033 13492 10474
rect 13450 10024 13506 10033
rect 13360 9988 13412 9994
rect 13450 9959 13506 9968
rect 13360 9930 13412 9936
rect 13372 9897 13400 9930
rect 13358 9888 13414 9897
rect 13358 9823 13414 9832
rect 13266 9752 13322 9761
rect 13266 9687 13322 9696
rect 13360 9716 13412 9722
rect 13174 9616 13230 9625
rect 12992 9580 13044 9586
rect 13174 9551 13230 9560
rect 12992 9522 13044 9528
rect 12900 9512 12952 9518
rect 12900 9454 12952 9460
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13096 9353 13124 9454
rect 13188 9382 13216 9551
rect 13176 9376 13228 9382
rect 13082 9344 13138 9353
rect 13176 9318 13228 9324
rect 13082 9279 13138 9288
rect 12820 9166 13032 9194
rect 12900 9104 12952 9110
rect 12898 9072 12900 9081
rect 12952 9072 12954 9081
rect 12716 9036 12768 9042
rect 12898 9007 12954 9016
rect 12716 8978 12768 8984
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12820 8809 12848 8910
rect 12806 8800 12862 8809
rect 12806 8735 12862 8744
rect 12806 8664 12862 8673
rect 12806 8599 12862 8608
rect 12716 8492 12768 8498
rect 12716 8434 12768 8440
rect 12624 8424 12676 8430
rect 12728 8401 12756 8434
rect 12624 8366 12676 8372
rect 12714 8392 12770 8401
rect 12714 8327 12770 8336
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12544 8129 12572 8230
rect 12530 8120 12586 8129
rect 12530 8055 12586 8064
rect 12164 7948 12216 7954
rect 12164 7890 12216 7896
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 12176 7732 12204 7890
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12176 7704 12572 7732
rect 12194 7644 12502 7664
rect 12194 7642 12200 7644
rect 12256 7642 12280 7644
rect 12336 7642 12360 7644
rect 12416 7642 12440 7644
rect 12496 7642 12502 7644
rect 12256 7590 12258 7642
rect 12438 7590 12440 7642
rect 12194 7588 12200 7590
rect 12256 7588 12280 7590
rect 12336 7588 12360 7590
rect 12416 7588 12440 7590
rect 12496 7588 12502 7590
rect 12194 7568 12502 7588
rect 12256 7472 12308 7478
rect 12256 7414 12308 7420
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 11992 6684 12112 6712
rect 11992 6497 12020 6684
rect 12176 6644 12204 6938
rect 12268 6934 12296 7414
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12348 7268 12400 7274
rect 12348 7210 12400 7216
rect 12256 6928 12308 6934
rect 12256 6870 12308 6876
rect 12360 6780 12388 7210
rect 12452 7177 12480 7346
rect 12544 7206 12572 7704
rect 12636 7274 12664 7754
rect 12716 7404 12768 7410
rect 12820 7392 12848 8599
rect 13004 8566 13032 9166
rect 13280 9042 13308 9687
rect 13360 9658 13412 9664
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13174 8936 13230 8945
rect 13084 8900 13136 8906
rect 13372 8922 13400 9658
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13464 9353 13492 9522
rect 13450 9344 13506 9353
rect 13450 9279 13506 9288
rect 13174 8871 13230 8880
rect 13280 8894 13400 8922
rect 13084 8842 13136 8848
rect 13096 8673 13124 8842
rect 13082 8664 13138 8673
rect 13188 8634 13216 8871
rect 13082 8599 13138 8608
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 12992 8560 13044 8566
rect 13044 8520 13124 8548
rect 12992 8502 13044 8508
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 12900 8288 12952 8294
rect 12900 8230 12952 8236
rect 12768 7364 12848 7392
rect 12716 7346 12768 7352
rect 12714 7304 12770 7313
rect 12624 7268 12676 7274
rect 12714 7239 12716 7248
rect 12624 7210 12676 7216
rect 12768 7239 12770 7248
rect 12716 7210 12768 7216
rect 12532 7200 12584 7206
rect 12438 7168 12494 7177
rect 12808 7200 12860 7206
rect 12532 7142 12584 7148
rect 12622 7168 12678 7177
rect 12438 7103 12494 7112
rect 12808 7142 12860 7148
rect 12622 7103 12678 7112
rect 12530 7032 12586 7041
rect 12530 6967 12586 6976
rect 12440 6792 12492 6798
rect 12360 6752 12440 6780
rect 12440 6734 12492 6740
rect 12084 6616 12204 6644
rect 11978 6488 12034 6497
rect 11978 6423 12034 6432
rect 12084 6254 12112 6616
rect 12194 6556 12502 6576
rect 12194 6554 12200 6556
rect 12256 6554 12280 6556
rect 12336 6554 12360 6556
rect 12416 6554 12440 6556
rect 12496 6554 12502 6556
rect 12256 6502 12258 6554
rect 12438 6502 12440 6554
rect 12194 6500 12200 6502
rect 12256 6500 12280 6502
rect 12336 6500 12360 6502
rect 12416 6500 12440 6502
rect 12496 6500 12502 6502
rect 12194 6480 12502 6500
rect 12544 6440 12572 6967
rect 12452 6412 12572 6440
rect 12164 6384 12216 6390
rect 12164 6326 12216 6332
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 11900 6038 12112 6066
rect 11796 5908 11848 5914
rect 11796 5850 11848 5856
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11428 5568 11480 5574
rect 11428 5510 11480 5516
rect 11520 5568 11572 5574
rect 11520 5510 11572 5516
rect 11440 5001 11468 5510
rect 11426 4992 11482 5001
rect 11426 4927 11482 4936
rect 11428 4752 11480 4758
rect 11428 4694 11480 4700
rect 11440 3670 11468 4694
rect 11428 3664 11480 3670
rect 11428 3606 11480 3612
rect 11532 3534 11560 5510
rect 11610 5400 11666 5409
rect 11610 5335 11666 5344
rect 11624 5234 11652 5335
rect 11612 5228 11664 5234
rect 11612 5170 11664 5176
rect 11610 4856 11666 4865
rect 11610 4791 11612 4800
rect 11664 4791 11666 4800
rect 11612 4762 11664 4768
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11624 4264 11652 4558
rect 11716 4486 11744 5782
rect 11794 5672 11850 5681
rect 12084 5642 12112 6038
rect 12176 5846 12204 6326
rect 12256 6248 12308 6254
rect 12308 6208 12388 6236
rect 12256 6190 12308 6196
rect 12164 5840 12216 5846
rect 12164 5782 12216 5788
rect 12360 5681 12388 6208
rect 12452 5914 12480 6412
rect 12636 6236 12664 7103
rect 12716 6860 12768 6866
rect 12716 6802 12768 6808
rect 12544 6208 12664 6236
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12544 5710 12572 6208
rect 12624 5840 12676 5846
rect 12624 5782 12676 5788
rect 12532 5704 12584 5710
rect 12346 5672 12402 5681
rect 11794 5607 11850 5616
rect 12072 5636 12124 5642
rect 11808 5574 11836 5607
rect 12532 5646 12584 5652
rect 12346 5607 12402 5616
rect 12072 5578 12124 5584
rect 11796 5568 11848 5574
rect 11796 5510 11848 5516
rect 11980 5568 12032 5574
rect 11980 5510 12032 5516
rect 11992 5370 12020 5510
rect 11980 5364 12032 5370
rect 12084 5352 12112 5578
rect 12636 5574 12664 5782
rect 12728 5778 12756 6802
rect 12820 6254 12848 7142
rect 12912 6866 12940 8230
rect 13004 7750 13032 8366
rect 12992 7744 13044 7750
rect 12990 7712 12992 7721
rect 13044 7712 13046 7721
rect 12990 7647 13046 7656
rect 13096 7585 13124 8520
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13188 8401 13216 8434
rect 13174 8392 13230 8401
rect 13174 8327 13230 8336
rect 13174 8256 13230 8265
rect 13174 8191 13230 8200
rect 13082 7576 13138 7585
rect 13082 7511 13138 7520
rect 12992 7472 13044 7478
rect 13188 7460 13216 8191
rect 13280 7750 13308 8894
rect 13360 8560 13412 8566
rect 13360 8502 13412 8508
rect 13372 8401 13400 8502
rect 13358 8392 13414 8401
rect 13358 8327 13414 8336
rect 13360 8084 13412 8090
rect 13360 8026 13412 8032
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13280 7546 13308 7686
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 12992 7414 13044 7420
rect 13096 7432 13216 7460
rect 12900 6860 12952 6866
rect 12900 6802 12952 6808
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12912 6254 12940 6326
rect 12808 6248 12860 6254
rect 12808 6190 12860 6196
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12900 6112 12952 6118
rect 12806 6080 12862 6089
rect 12900 6054 12952 6060
rect 12806 6015 12862 6024
rect 12820 5846 12848 6015
rect 12912 5914 12940 6054
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 12808 5840 12860 5846
rect 12808 5782 12860 5788
rect 12898 5808 12954 5817
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12532 5568 12584 5574
rect 12532 5510 12584 5516
rect 12624 5568 12676 5574
rect 12624 5510 12676 5516
rect 12194 5468 12502 5488
rect 12194 5466 12200 5468
rect 12256 5466 12280 5468
rect 12336 5466 12360 5468
rect 12416 5466 12440 5468
rect 12496 5466 12502 5468
rect 12256 5414 12258 5466
rect 12438 5414 12440 5466
rect 12194 5412 12200 5414
rect 12256 5412 12280 5414
rect 12336 5412 12360 5414
rect 12416 5412 12440 5414
rect 12496 5412 12502 5414
rect 12194 5392 12502 5412
rect 12084 5324 12204 5352
rect 11980 5306 12032 5312
rect 11796 5296 11848 5302
rect 11796 5238 11848 5244
rect 11886 5264 11942 5273
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11624 4236 11744 4264
rect 11610 4176 11666 4185
rect 11610 4111 11612 4120
rect 11664 4111 11666 4120
rect 11612 4082 11664 4088
rect 11716 3584 11744 4236
rect 11808 4154 11836 5238
rect 11942 5222 12112 5250
rect 11886 5199 11942 5208
rect 11980 5092 12032 5098
rect 11980 5034 12032 5040
rect 11992 5001 12020 5034
rect 11978 4992 12034 5001
rect 11978 4927 12034 4936
rect 11888 4684 11940 4690
rect 11940 4644 12020 4672
rect 11888 4626 11940 4632
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11900 4321 11928 4422
rect 11886 4312 11942 4321
rect 11886 4247 11942 4256
rect 11808 4126 11928 4154
rect 11796 4072 11848 4078
rect 11796 4014 11848 4020
rect 11624 3556 11744 3584
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11428 3392 11480 3398
rect 11428 3334 11480 3340
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11256 2604 11376 2632
rect 11256 2553 11284 2604
rect 11112 2468 11192 2496
rect 11242 2544 11298 2553
rect 11242 2479 11298 2488
rect 11336 2508 11388 2514
rect 11060 2450 11112 2456
rect 11336 2450 11388 2456
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10980 2106 11008 2246
rect 10968 2100 11020 2106
rect 10968 2042 11020 2048
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 11060 1760 11112 1766
rect 11060 1702 11112 1708
rect 10876 808 10928 814
rect 9182 734 9260 762
rect 9126 711 9182 720
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 9770 640 9826 649
rect 9770 575 9826 584
rect 9784 270 9812 575
rect 9772 264 9824 270
rect 9772 206 9824 212
rect 10046 0 10102 800
rect 10414 0 10470 800
rect 10690 0 10746 800
rect 11072 800 11100 1702
rect 11164 1601 11192 2042
rect 11150 1592 11206 1601
rect 11150 1527 11206 1536
rect 11256 1222 11284 2382
rect 11348 2009 11376 2450
rect 11334 2000 11390 2009
rect 11440 1970 11468 3334
rect 11532 2446 11560 3334
rect 11520 2440 11572 2446
rect 11520 2382 11572 2388
rect 11520 2304 11572 2310
rect 11518 2272 11520 2281
rect 11572 2272 11574 2281
rect 11518 2207 11574 2216
rect 11518 2136 11574 2145
rect 11518 2071 11574 2080
rect 11532 1970 11560 2071
rect 11624 2038 11652 3556
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 11716 3097 11744 3402
rect 11808 3369 11836 4014
rect 11794 3360 11850 3369
rect 11794 3295 11850 3304
rect 11794 3224 11850 3233
rect 11794 3159 11796 3168
rect 11848 3159 11850 3168
rect 11796 3130 11848 3136
rect 11702 3088 11758 3097
rect 11702 3023 11758 3032
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11612 2032 11664 2038
rect 11612 1974 11664 1980
rect 11334 1935 11390 1944
rect 11428 1964 11480 1970
rect 11428 1906 11480 1912
rect 11520 1964 11572 1970
rect 11520 1906 11572 1912
rect 11716 1834 11744 2926
rect 11796 2576 11848 2582
rect 11796 2518 11848 2524
rect 11704 1828 11756 1834
rect 11704 1770 11756 1776
rect 11428 1692 11480 1698
rect 11428 1634 11480 1640
rect 11440 1601 11468 1634
rect 11426 1592 11482 1601
rect 11426 1527 11482 1536
rect 11244 1216 11296 1222
rect 11244 1158 11296 1164
rect 11440 800 11468 1527
rect 11808 1358 11836 2518
rect 11900 2446 11928 4126
rect 11992 3534 12020 4644
rect 12084 4622 12112 5222
rect 12176 5166 12204 5324
rect 12544 5302 12572 5510
rect 12820 5352 12848 5782
rect 13004 5760 13032 7414
rect 13096 6730 13124 7432
rect 13372 7392 13400 8026
rect 13464 7834 13492 9279
rect 13556 8906 13584 11290
rect 13648 11014 13676 12192
rect 13636 11008 13688 11014
rect 13636 10950 13688 10956
rect 13636 10464 13688 10470
rect 13636 10406 13688 10412
rect 13648 10130 13676 10406
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13636 9920 13688 9926
rect 13636 9862 13688 9868
rect 13648 9110 13676 9862
rect 13740 9382 13768 12294
rect 13832 11937 13860 12378
rect 13818 11928 13874 11937
rect 13924 11898 13952 17818
rect 14016 17066 14044 19200
rect 14384 17954 14412 19200
rect 14384 17926 14504 17954
rect 14004 17060 14056 17066
rect 14004 17002 14056 17008
rect 14068 16892 14376 16912
rect 14068 16890 14074 16892
rect 14130 16890 14154 16892
rect 14210 16890 14234 16892
rect 14290 16890 14314 16892
rect 14370 16890 14376 16892
rect 14130 16838 14132 16890
rect 14312 16838 14314 16890
rect 14068 16836 14074 16838
rect 14130 16836 14154 16838
rect 14210 16836 14234 16838
rect 14290 16836 14314 16838
rect 14370 16836 14376 16838
rect 14068 16816 14376 16836
rect 14068 15804 14376 15824
rect 14068 15802 14074 15804
rect 14130 15802 14154 15804
rect 14210 15802 14234 15804
rect 14290 15802 14314 15804
rect 14370 15802 14376 15804
rect 14130 15750 14132 15802
rect 14312 15750 14314 15802
rect 14068 15748 14074 15750
rect 14130 15748 14154 15750
rect 14210 15748 14234 15750
rect 14290 15748 14314 15750
rect 14370 15748 14376 15750
rect 14068 15728 14376 15748
rect 14068 14716 14376 14736
rect 14068 14714 14074 14716
rect 14130 14714 14154 14716
rect 14210 14714 14234 14716
rect 14290 14714 14314 14716
rect 14370 14714 14376 14716
rect 14130 14662 14132 14714
rect 14312 14662 14314 14714
rect 14068 14660 14074 14662
rect 14130 14660 14154 14662
rect 14210 14660 14234 14662
rect 14290 14660 14314 14662
rect 14370 14660 14376 14662
rect 14068 14640 14376 14660
rect 14068 13628 14376 13648
rect 14068 13626 14074 13628
rect 14130 13626 14154 13628
rect 14210 13626 14234 13628
rect 14290 13626 14314 13628
rect 14370 13626 14376 13628
rect 14130 13574 14132 13626
rect 14312 13574 14314 13626
rect 14068 13572 14074 13574
rect 14130 13572 14154 13574
rect 14210 13572 14234 13574
rect 14290 13572 14314 13574
rect 14370 13572 14376 13574
rect 14068 13552 14376 13572
rect 14068 12540 14376 12560
rect 14068 12538 14074 12540
rect 14130 12538 14154 12540
rect 14210 12538 14234 12540
rect 14290 12538 14314 12540
rect 14370 12538 14376 12540
rect 14130 12486 14132 12538
rect 14312 12486 14314 12538
rect 14068 12484 14074 12486
rect 14130 12484 14154 12486
rect 14210 12484 14234 12486
rect 14290 12484 14314 12486
rect 14370 12484 14376 12486
rect 14068 12464 14376 12484
rect 14476 12424 14504 17926
rect 14556 15632 14608 15638
rect 14556 15574 14608 15580
rect 14384 12396 14504 12424
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13818 11863 13874 11872
rect 13912 11892 13964 11898
rect 13912 11834 13964 11840
rect 13818 11792 13874 11801
rect 13818 11727 13874 11736
rect 13832 10266 13860 11727
rect 13912 11688 13964 11694
rect 14016 11676 14044 12038
rect 13964 11648 14044 11676
rect 13912 11630 13964 11636
rect 13924 11150 13952 11630
rect 14108 11626 14136 12242
rect 14384 12186 14412 12396
rect 14462 12336 14518 12345
rect 14462 12271 14464 12280
rect 14516 12271 14518 12280
rect 14464 12242 14516 12248
rect 14384 12158 14504 12186
rect 14568 12170 14596 15574
rect 14648 14612 14700 14618
rect 14648 14554 14700 14560
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14278 12064 14334 12073
rect 14200 11665 14228 12038
rect 14278 11999 14334 12008
rect 14186 11656 14242 11665
rect 14096 11620 14148 11626
rect 14292 11626 14320 11999
rect 14186 11591 14242 11600
rect 14280 11620 14332 11626
rect 14096 11562 14148 11568
rect 14280 11562 14332 11568
rect 14068 11452 14376 11472
rect 14068 11450 14074 11452
rect 14130 11450 14154 11452
rect 14210 11450 14234 11452
rect 14290 11450 14314 11452
rect 14370 11450 14376 11452
rect 14130 11398 14132 11450
rect 14312 11398 14314 11450
rect 14068 11396 14074 11398
rect 14130 11396 14154 11398
rect 14210 11396 14234 11398
rect 14290 11396 14314 11398
rect 14370 11396 14376 11398
rect 14068 11376 14376 11396
rect 14372 11280 14424 11286
rect 14278 11248 14334 11257
rect 14004 11212 14056 11218
rect 14372 11222 14424 11228
rect 14278 11183 14334 11192
rect 14004 11154 14056 11160
rect 13912 11144 13964 11150
rect 13912 11086 13964 11092
rect 14016 10810 14044 11154
rect 14096 11076 14148 11082
rect 14096 11018 14148 11024
rect 14108 10985 14136 11018
rect 14188 11008 14240 11014
rect 14094 10976 14150 10985
rect 14188 10950 14240 10956
rect 14094 10911 14150 10920
rect 14108 10810 14136 10911
rect 14004 10804 14056 10810
rect 13924 10764 14004 10792
rect 13820 10260 13872 10266
rect 13820 10202 13872 10208
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13728 9376 13780 9382
rect 13832 9353 13860 9998
rect 13728 9318 13780 9324
rect 13818 9344 13874 9353
rect 13818 9279 13874 9288
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 13924 8956 13952 10764
rect 14004 10746 14056 10752
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14108 10606 14136 10746
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14200 10538 14228 10950
rect 14292 10810 14320 11183
rect 14280 10804 14332 10810
rect 14280 10746 14332 10752
rect 14384 10742 14412 11222
rect 14372 10736 14424 10742
rect 14372 10678 14424 10684
rect 14188 10532 14240 10538
rect 14188 10474 14240 10480
rect 14068 10364 14376 10384
rect 14068 10362 14074 10364
rect 14130 10362 14154 10364
rect 14210 10362 14234 10364
rect 14290 10362 14314 10364
rect 14370 10362 14376 10364
rect 14130 10310 14132 10362
rect 14312 10310 14314 10362
rect 14068 10308 14074 10310
rect 14130 10308 14154 10310
rect 14210 10308 14234 10310
rect 14290 10308 14314 10310
rect 14370 10308 14376 10310
rect 14068 10288 14376 10308
rect 14476 10248 14504 12158
rect 14556 12164 14608 12170
rect 14556 12106 14608 12112
rect 14554 11928 14610 11937
rect 14554 11863 14556 11872
rect 14608 11863 14610 11872
rect 14556 11834 14608 11840
rect 14568 11354 14596 11834
rect 14556 11348 14608 11354
rect 14556 11290 14608 11296
rect 14568 10713 14596 11290
rect 14660 11234 14688 14554
rect 14752 11898 14780 19200
rect 15120 15910 15148 19200
rect 15488 17882 15516 19200
rect 15476 17876 15528 17882
rect 15476 17818 15528 17824
rect 15474 17776 15530 17785
rect 15474 17711 15530 17720
rect 15488 16574 15516 17711
rect 15396 16546 15516 16574
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 14922 14512 14978 14521
rect 14922 14447 14978 14456
rect 14832 13252 14884 13258
rect 14832 13194 14884 13200
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14752 11393 14780 11834
rect 14738 11384 14794 11393
rect 14738 11319 14794 11328
rect 14660 11206 14780 11234
rect 14648 11144 14700 11150
rect 14648 11086 14700 11092
rect 14554 10704 14610 10713
rect 14554 10639 14610 10648
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14292 10220 14504 10248
rect 14188 10192 14240 10198
rect 14186 10160 14188 10169
rect 14292 10180 14320 10220
rect 14240 10160 14320 10180
rect 14242 10152 14320 10160
rect 14568 10112 14596 10542
rect 14186 10095 14242 10104
rect 14476 10084 14596 10112
rect 14096 9920 14148 9926
rect 14094 9888 14096 9897
rect 14188 9920 14240 9926
rect 14148 9888 14150 9897
rect 14188 9862 14240 9868
rect 14094 9823 14150 9832
rect 14200 9722 14228 9862
rect 14188 9716 14240 9722
rect 14188 9658 14240 9664
rect 14476 9450 14504 10084
rect 14556 9988 14608 9994
rect 14556 9930 14608 9936
rect 14568 9761 14596 9930
rect 14554 9752 14610 9761
rect 14554 9687 14610 9696
rect 14660 9586 14688 11086
rect 14752 11014 14780 11206
rect 14740 11008 14792 11014
rect 14740 10950 14792 10956
rect 14752 10470 14780 10950
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 9722 14780 10406
rect 14844 9722 14872 13194
rect 14936 11150 14964 14447
rect 15108 11688 15160 11694
rect 15108 11630 15160 11636
rect 15016 11552 15068 11558
rect 15016 11494 15068 11500
rect 14924 11144 14976 11150
rect 14924 11086 14976 11092
rect 14922 10976 14978 10985
rect 14922 10911 14978 10920
rect 14740 9716 14792 9722
rect 14740 9658 14792 9664
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14648 9580 14700 9586
rect 14648 9522 14700 9528
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14068 9276 14376 9296
rect 14068 9274 14074 9276
rect 14130 9274 14154 9276
rect 14210 9274 14234 9276
rect 14290 9274 14314 9276
rect 14370 9274 14376 9276
rect 14130 9222 14132 9274
rect 14312 9222 14314 9274
rect 14068 9220 14074 9222
rect 14130 9220 14154 9222
rect 14210 9220 14234 9222
rect 14290 9220 14314 9222
rect 14370 9220 14376 9222
rect 14068 9200 14376 9220
rect 14462 9208 14518 9217
rect 14568 9178 14596 9454
rect 14462 9143 14518 9152
rect 14556 9172 14608 9178
rect 14476 9110 14504 9143
rect 14556 9114 14608 9120
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14556 9036 14608 9042
rect 14556 8978 14608 8984
rect 13924 8928 14044 8956
rect 13544 8900 13596 8906
rect 13544 8842 13596 8848
rect 13556 8430 13584 8842
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13542 8120 13598 8129
rect 13542 8055 13598 8064
rect 13556 7954 13584 8055
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13464 7806 13584 7834
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13188 7364 13400 7392
rect 13084 6724 13136 6730
rect 13084 6666 13136 6672
rect 13096 6497 13124 6666
rect 13082 6488 13138 6497
rect 13082 6423 13138 6432
rect 13084 6248 13136 6254
rect 13188 6236 13216 7364
rect 13358 7032 13414 7041
rect 13358 6967 13414 6976
rect 13268 6928 13320 6934
rect 13268 6870 13320 6876
rect 13280 6474 13308 6870
rect 13372 6866 13400 6967
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13280 6446 13400 6474
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13136 6208 13216 6236
rect 13084 6190 13136 6196
rect 12954 5752 13032 5760
rect 12898 5743 12900 5752
rect 12952 5732 13032 5752
rect 12900 5714 12952 5720
rect 12992 5568 13044 5574
rect 13096 5545 13124 6190
rect 13176 6112 13228 6118
rect 13280 6089 13308 6326
rect 13176 6054 13228 6060
rect 13266 6080 13322 6089
rect 13188 5896 13216 6054
rect 13266 6015 13322 6024
rect 13372 5930 13400 6446
rect 13464 6236 13492 7686
rect 13556 7410 13584 7806
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13648 7002 13676 8366
rect 13832 8294 13860 8774
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 13740 8266 13860 8294
rect 13740 7818 13768 8266
rect 13818 8120 13874 8129
rect 13818 8055 13874 8064
rect 13832 7818 13860 8055
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13820 7812 13872 7818
rect 13820 7754 13872 7760
rect 13924 7750 13952 8570
rect 14016 8430 14044 8928
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14004 8424 14056 8430
rect 14004 8366 14056 8372
rect 14068 8188 14376 8208
rect 14068 8186 14074 8188
rect 14130 8186 14154 8188
rect 14210 8186 14234 8188
rect 14290 8186 14314 8188
rect 14370 8186 14376 8188
rect 14130 8134 14132 8186
rect 14312 8134 14314 8186
rect 14068 8132 14074 8134
rect 14130 8132 14154 8134
rect 14210 8132 14234 8134
rect 14290 8132 14314 8134
rect 14370 8132 14376 8134
rect 14068 8112 14376 8132
rect 14004 8016 14056 8022
rect 14056 7976 14136 8004
rect 14004 7958 14056 7964
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13726 7576 13782 7585
rect 14016 7528 14044 7822
rect 14108 7818 14136 7976
rect 14096 7812 14148 7818
rect 14096 7754 14148 7760
rect 14476 7750 14504 8570
rect 14568 8498 14596 8978
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14568 8129 14596 8298
rect 14554 8120 14610 8129
rect 14554 8055 14610 8064
rect 14660 7818 14688 9522
rect 14752 8634 14780 9658
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 14844 9450 14872 9522
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 14844 9110 14872 9386
rect 14832 9104 14884 9110
rect 14832 9046 14884 9052
rect 14844 8809 14872 9046
rect 14830 8800 14886 8809
rect 14830 8735 14886 8744
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14648 7812 14700 7818
rect 14648 7754 14700 7760
rect 14464 7744 14516 7750
rect 14464 7686 14516 7692
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 13726 7511 13728 7520
rect 13780 7511 13782 7520
rect 13728 7482 13780 7488
rect 13832 7500 14044 7528
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13740 7002 13768 7278
rect 13636 6996 13688 7002
rect 13636 6938 13688 6944
rect 13728 6996 13780 7002
rect 13728 6938 13780 6944
rect 13634 6896 13690 6905
rect 13634 6831 13690 6840
rect 13544 6656 13596 6662
rect 13544 6598 13596 6604
rect 13556 6458 13584 6598
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13464 6208 13584 6236
rect 13450 6080 13506 6089
rect 13450 6015 13506 6024
rect 13177 5868 13216 5896
rect 13280 5902 13400 5930
rect 13177 5760 13205 5868
rect 13280 5846 13308 5902
rect 13268 5840 13320 5846
rect 13268 5782 13320 5788
rect 13358 5808 13414 5817
rect 13177 5732 13216 5760
rect 13358 5743 13414 5752
rect 12992 5510 13044 5516
rect 13082 5536 13138 5545
rect 12728 5324 12848 5352
rect 12900 5364 12952 5370
rect 12532 5296 12584 5302
rect 12254 5264 12310 5273
rect 12254 5199 12256 5208
rect 12308 5199 12310 5208
rect 12438 5264 12494 5273
rect 12532 5238 12584 5244
rect 12438 5199 12494 5208
rect 12256 5170 12308 5176
rect 12164 5160 12216 5166
rect 12164 5102 12216 5108
rect 12348 5092 12400 5098
rect 12348 5034 12400 5040
rect 12256 5024 12308 5030
rect 12256 4966 12308 4972
rect 12268 4729 12296 4966
rect 12254 4720 12310 4729
rect 12360 4706 12388 5034
rect 12452 4826 12480 5199
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12622 4992 12678 5001
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12544 4706 12572 4966
rect 12622 4927 12678 4936
rect 12360 4678 12572 4706
rect 12254 4655 12310 4664
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12084 4264 12112 4422
rect 12194 4380 12502 4400
rect 12194 4378 12200 4380
rect 12256 4378 12280 4380
rect 12336 4378 12360 4380
rect 12416 4378 12440 4380
rect 12496 4378 12502 4380
rect 12256 4326 12258 4378
rect 12438 4326 12440 4378
rect 12194 4324 12200 4326
rect 12256 4324 12280 4326
rect 12336 4324 12360 4326
rect 12416 4324 12440 4326
rect 12496 4324 12502 4326
rect 12194 4304 12502 4324
rect 12084 4236 12296 4264
rect 12072 4072 12124 4078
rect 12072 4014 12124 4020
rect 11980 3528 12032 3534
rect 11980 3470 12032 3476
rect 11980 3392 12032 3398
rect 11980 3334 12032 3340
rect 11992 3194 12020 3334
rect 11980 3188 12032 3194
rect 11980 3130 12032 3136
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 12084 2106 12112 4014
rect 12268 3670 12296 4236
rect 12346 4176 12402 4185
rect 12346 4111 12402 4120
rect 12256 3664 12308 3670
rect 12256 3606 12308 3612
rect 12360 3602 12388 4111
rect 12440 4072 12492 4078
rect 12438 4040 12440 4049
rect 12492 4040 12494 4049
rect 12438 3975 12494 3984
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12348 3596 12400 3602
rect 12348 3538 12400 3544
rect 12452 3380 12480 3878
rect 12544 3738 12572 4422
rect 12636 4282 12664 4927
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12532 3732 12584 3738
rect 12532 3674 12584 3680
rect 12728 3584 12756 5324
rect 12900 5306 12952 5312
rect 12808 5228 12860 5234
rect 12808 5170 12860 5176
rect 12820 4010 12848 5170
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12912 3738 12940 5306
rect 13004 4690 13032 5510
rect 13082 5471 13138 5480
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 13096 4486 13124 5238
rect 13084 4480 13136 4486
rect 13084 4422 13136 4428
rect 13084 4276 13136 4282
rect 13084 4218 13136 4224
rect 12990 4040 13046 4049
rect 12990 3975 13046 3984
rect 12808 3732 12860 3738
rect 12808 3674 12860 3680
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12636 3556 12756 3584
rect 12452 3352 12572 3380
rect 12194 3292 12502 3312
rect 12194 3290 12200 3292
rect 12256 3290 12280 3292
rect 12336 3290 12360 3292
rect 12416 3290 12440 3292
rect 12496 3290 12502 3292
rect 12256 3238 12258 3290
rect 12438 3238 12440 3290
rect 12194 3236 12200 3238
rect 12256 3236 12280 3238
rect 12336 3236 12360 3238
rect 12416 3236 12440 3238
rect 12496 3236 12502 3238
rect 12194 3216 12502 3236
rect 12164 3120 12216 3126
rect 12162 3088 12164 3097
rect 12256 3120 12308 3126
rect 12216 3088 12218 3097
rect 12256 3062 12308 3068
rect 12438 3088 12494 3097
rect 12162 3023 12218 3032
rect 12268 2990 12296 3062
rect 12438 3023 12494 3032
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 12452 2292 12480 3023
rect 12544 2446 12572 3352
rect 12636 3126 12664 3556
rect 12714 3496 12770 3505
rect 12714 3431 12770 3440
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12728 2650 12756 3431
rect 12820 3058 12848 3674
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12900 2508 12952 2514
rect 12900 2450 12952 2456
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 12452 2264 12572 2292
rect 12194 2204 12502 2224
rect 12194 2202 12200 2204
rect 12256 2202 12280 2204
rect 12336 2202 12360 2204
rect 12416 2202 12440 2204
rect 12496 2202 12502 2204
rect 12256 2150 12258 2202
rect 12438 2150 12440 2202
rect 12194 2148 12200 2150
rect 12256 2148 12280 2150
rect 12336 2148 12360 2150
rect 12416 2148 12440 2150
rect 12496 2148 12502 2150
rect 12194 2128 12502 2148
rect 12072 2100 12124 2106
rect 12544 2088 12572 2264
rect 12636 2106 12664 2314
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 12072 2042 12124 2048
rect 12452 2060 12572 2088
rect 12624 2100 12676 2106
rect 12070 2000 12126 2009
rect 12070 1935 12126 1944
rect 11886 1456 11942 1465
rect 11886 1391 11942 1400
rect 11796 1352 11848 1358
rect 11796 1294 11848 1300
rect 11900 1204 11928 1391
rect 11808 1176 11928 1204
rect 11520 1148 11572 1154
rect 11520 1090 11572 1096
rect 10876 750 10928 756
rect 11058 0 11114 800
rect 11426 0 11482 800
rect 11532 746 11560 1090
rect 11808 800 11836 1176
rect 12084 800 12112 1935
rect 12452 800 12480 2060
rect 12624 2042 12676 2048
rect 12820 800 12848 2246
rect 12912 1737 12940 2450
rect 12898 1728 12954 1737
rect 12898 1663 12954 1672
rect 13004 882 13032 3975
rect 13096 3505 13124 4218
rect 13082 3496 13138 3505
rect 13082 3431 13138 3440
rect 13084 3392 13136 3398
rect 13084 3334 13136 3340
rect 13096 3074 13124 3334
rect 13188 3194 13216 5732
rect 13372 5284 13400 5743
rect 13280 5256 13400 5284
rect 13280 4622 13308 5256
rect 13360 5024 13412 5030
rect 13360 4966 13412 4972
rect 13268 4616 13320 4622
rect 13268 4558 13320 4564
rect 13268 4480 13320 4486
rect 13266 4448 13268 4457
rect 13320 4448 13322 4457
rect 13266 4383 13322 4392
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13280 3534 13308 3878
rect 13268 3528 13320 3534
rect 13268 3470 13320 3476
rect 13372 3482 13400 4966
rect 13464 3738 13492 6015
rect 13556 5710 13584 6208
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13648 5234 13676 6831
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13740 5370 13768 6734
rect 13832 6254 13860 7500
rect 14372 7404 14424 7410
rect 14372 7346 14424 7352
rect 14004 7268 14056 7274
rect 13924 7228 14004 7256
rect 13924 6662 13952 7228
rect 14004 7210 14056 7216
rect 14384 7188 14412 7346
rect 14476 7313 14504 7686
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14462 7304 14518 7313
rect 14462 7239 14518 7248
rect 14384 7160 14504 7188
rect 14068 7100 14376 7120
rect 14068 7098 14074 7100
rect 14130 7098 14154 7100
rect 14210 7098 14234 7100
rect 14290 7098 14314 7100
rect 14370 7098 14376 7100
rect 14130 7046 14132 7098
rect 14312 7046 14314 7098
rect 14068 7044 14074 7046
rect 14130 7044 14154 7046
rect 14210 7044 14234 7046
rect 14290 7044 14314 7046
rect 14370 7044 14376 7046
rect 14068 7024 14376 7044
rect 14280 6928 14332 6934
rect 14280 6870 14332 6876
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 14096 6656 14148 6662
rect 14096 6598 14148 6604
rect 14188 6656 14240 6662
rect 14188 6598 14240 6604
rect 14002 6488 14058 6497
rect 14108 6458 14136 6598
rect 14002 6423 14004 6432
rect 14056 6423 14058 6432
rect 14096 6452 14148 6458
rect 14004 6394 14056 6400
rect 14096 6394 14148 6400
rect 13912 6316 13964 6322
rect 13912 6258 13964 6264
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5953 13860 6054
rect 13818 5944 13874 5953
rect 13818 5879 13874 5888
rect 13728 5364 13780 5370
rect 13924 5352 13952 6258
rect 14200 6186 14228 6598
rect 14292 6186 14320 6870
rect 14476 6497 14504 7160
rect 14568 6798 14596 7346
rect 14648 6860 14700 6866
rect 14648 6802 14700 6808
rect 14556 6792 14608 6798
rect 14660 6769 14688 6802
rect 14556 6734 14608 6740
rect 14646 6760 14702 6769
rect 14646 6695 14702 6704
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14462 6488 14518 6497
rect 14462 6423 14518 6432
rect 14568 6372 14596 6598
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14476 6361 14596 6372
rect 14462 6352 14596 6361
rect 14518 6344 14596 6352
rect 14660 6304 14688 6394
rect 14462 6287 14518 6296
rect 14568 6276 14688 6304
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 14280 6180 14332 6186
rect 14280 6122 14332 6128
rect 14068 6012 14376 6032
rect 14068 6010 14074 6012
rect 14130 6010 14154 6012
rect 14210 6010 14234 6012
rect 14290 6010 14314 6012
rect 14370 6010 14376 6012
rect 14130 5958 14132 6010
rect 14312 5958 14314 6010
rect 14068 5956 14074 5958
rect 14130 5956 14154 5958
rect 14210 5956 14234 5958
rect 14290 5956 14314 5958
rect 14370 5956 14376 5958
rect 14068 5936 14376 5956
rect 14004 5840 14056 5846
rect 14004 5782 14056 5788
rect 13728 5306 13780 5312
rect 13832 5324 13952 5352
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13542 4856 13598 4865
rect 13542 4791 13598 4800
rect 13556 4214 13584 4791
rect 13636 4752 13688 4758
rect 13636 4694 13688 4700
rect 13544 4208 13596 4214
rect 13648 4185 13676 4694
rect 13544 4150 13596 4156
rect 13634 4176 13690 4185
rect 13634 4111 13690 4120
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13464 3641 13492 3674
rect 13556 3670 13584 4014
rect 13740 3992 13768 5170
rect 13832 5030 13860 5324
rect 14016 5302 14044 5782
rect 14186 5672 14242 5681
rect 14096 5636 14148 5642
rect 14186 5607 14242 5616
rect 14096 5578 14148 5584
rect 14004 5296 14056 5302
rect 14004 5238 14056 5244
rect 14108 5137 14136 5578
rect 14200 5166 14228 5607
rect 14278 5536 14334 5545
rect 14278 5471 14334 5480
rect 14292 5234 14320 5471
rect 14370 5400 14426 5409
rect 14370 5335 14426 5344
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 14188 5160 14240 5166
rect 14094 5128 14150 5137
rect 14188 5102 14240 5108
rect 14278 5128 14334 5137
rect 14094 5063 14150 5072
rect 14278 5063 14280 5072
rect 14332 5063 14334 5072
rect 14280 5034 14332 5040
rect 13820 5024 13872 5030
rect 14384 5012 14412 5335
rect 14476 5137 14504 6190
rect 14462 5128 14518 5137
rect 14462 5063 14518 5072
rect 14384 4984 14504 5012
rect 13820 4966 13872 4972
rect 14068 4924 14376 4944
rect 14068 4922 14074 4924
rect 14130 4922 14154 4924
rect 14210 4922 14234 4924
rect 14290 4922 14314 4924
rect 14370 4922 14376 4924
rect 14130 4870 14132 4922
rect 14312 4870 14314 4922
rect 14068 4868 14074 4870
rect 14130 4868 14154 4870
rect 14210 4868 14234 4870
rect 14290 4868 14314 4870
rect 14370 4868 14376 4870
rect 14068 4848 14376 4868
rect 14370 4720 14426 4729
rect 14370 4655 14426 4664
rect 14188 4616 14240 4622
rect 14188 4558 14240 4564
rect 14200 4282 14228 4558
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 14188 4276 14240 4282
rect 14188 4218 14240 4224
rect 14108 4049 14136 4218
rect 14278 4176 14334 4185
rect 14278 4111 14280 4120
rect 14332 4111 14334 4120
rect 14280 4082 14332 4088
rect 14384 4078 14412 4655
rect 14476 4282 14504 4984
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14372 4072 14424 4078
rect 14094 4040 14150 4049
rect 14004 4004 14056 4010
rect 13648 3964 13768 3992
rect 13924 3964 14004 3992
rect 13544 3664 13596 3670
rect 13450 3632 13506 3641
rect 13544 3606 13596 3612
rect 13450 3567 13506 3576
rect 13544 3528 13596 3534
rect 13542 3496 13544 3505
rect 13596 3496 13598 3505
rect 13372 3454 13492 3482
rect 13268 3392 13320 3398
rect 13320 3352 13400 3380
rect 13268 3334 13320 3340
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13268 3188 13320 3194
rect 13268 3130 13320 3136
rect 13280 3074 13308 3130
rect 13096 3046 13308 3074
rect 13176 2916 13228 2922
rect 13176 2858 13228 2864
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 13096 2446 13124 2790
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13188 1578 13216 2858
rect 13268 2508 13320 2514
rect 13268 2450 13320 2456
rect 13280 1970 13308 2450
rect 13268 1964 13320 1970
rect 13268 1906 13320 1912
rect 13096 1550 13216 1578
rect 13096 1154 13124 1550
rect 13174 1320 13230 1329
rect 13174 1255 13230 1264
rect 13084 1148 13136 1154
rect 13084 1090 13136 1096
rect 12992 876 13044 882
rect 12992 818 13044 824
rect 13188 800 13216 1255
rect 13372 1193 13400 3352
rect 13464 3058 13492 3454
rect 13542 3431 13598 3440
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13452 2916 13504 2922
rect 13452 2858 13504 2864
rect 13464 1494 13492 2858
rect 13452 1488 13504 1494
rect 13452 1430 13504 1436
rect 13358 1184 13414 1193
rect 13358 1119 13414 1128
rect 13464 800 13492 1430
rect 11520 740 11572 746
rect 11520 682 11572 688
rect 11794 0 11850 800
rect 12070 0 12126 800
rect 12438 0 12494 800
rect 12806 0 12862 800
rect 13174 0 13230 800
rect 13450 0 13506 800
rect 13556 105 13584 3334
rect 13648 3074 13676 3964
rect 13924 3924 13952 3964
rect 14372 4014 14424 4020
rect 14094 3975 14150 3984
rect 14004 3946 14056 3952
rect 13726 3904 13782 3913
rect 13726 3839 13782 3848
rect 13832 3896 13952 3924
rect 13740 3602 13768 3839
rect 13728 3596 13780 3602
rect 13728 3538 13780 3544
rect 13648 3046 13768 3074
rect 13636 2984 13688 2990
rect 13636 2926 13688 2932
rect 13542 96 13598 105
rect 13648 66 13676 2926
rect 13740 1630 13768 3046
rect 13832 2990 13860 3896
rect 14068 3836 14376 3856
rect 14068 3834 14074 3836
rect 14130 3834 14154 3836
rect 14210 3834 14234 3836
rect 14290 3834 14314 3836
rect 14370 3834 14376 3836
rect 14130 3782 14132 3834
rect 14312 3782 14314 3834
rect 14068 3780 14074 3782
rect 14130 3780 14154 3782
rect 14210 3780 14234 3782
rect 14290 3780 14314 3782
rect 14370 3780 14376 3782
rect 14068 3760 14376 3780
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 13820 2984 13872 2990
rect 13820 2926 13872 2932
rect 13818 2816 13874 2825
rect 13818 2751 13874 2760
rect 13728 1624 13780 1630
rect 13728 1566 13780 1572
rect 13832 800 13860 2751
rect 13924 2650 13952 3470
rect 14464 3188 14516 3194
rect 14568 3176 14596 6276
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 14660 5302 14688 6122
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14660 4826 14688 4966
rect 14648 4820 14700 4826
rect 14648 4762 14700 4768
rect 14752 4264 14780 7686
rect 14844 6730 14872 8434
rect 14936 7546 14964 10911
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 14936 6769 14964 7482
rect 15028 7410 15056 11494
rect 15120 11121 15148 11630
rect 15106 11112 15162 11121
rect 15106 11047 15162 11056
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15120 10810 15148 10950
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15120 9722 15148 10746
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 15120 8673 15148 9658
rect 15106 8664 15162 8673
rect 15212 8634 15240 15302
rect 15290 13968 15346 13977
rect 15290 13903 15346 13912
rect 15304 9382 15332 13903
rect 15396 11694 15424 16546
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15396 11354 15424 11494
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15384 11144 15436 11150
rect 15384 11086 15436 11092
rect 15292 9376 15344 9382
rect 15292 9318 15344 9324
rect 15292 9104 15344 9110
rect 15292 9046 15344 9052
rect 15106 8599 15162 8608
rect 15200 8628 15252 8634
rect 15120 8514 15148 8599
rect 15200 8570 15252 8576
rect 15120 8486 15240 8514
rect 15106 8120 15162 8129
rect 15106 8055 15162 8064
rect 15120 7954 15148 8055
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 15212 7818 15240 8486
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 14922 6760 14978 6769
rect 14832 6724 14884 6730
rect 14922 6695 14978 6704
rect 14832 6666 14884 6672
rect 14844 6361 14872 6666
rect 14924 6656 14976 6662
rect 14924 6598 14976 6604
rect 14936 6390 14964 6598
rect 14924 6384 14976 6390
rect 14830 6352 14886 6361
rect 14924 6326 14976 6332
rect 14830 6287 14886 6296
rect 14832 6248 14884 6254
rect 14830 6216 14832 6225
rect 14884 6216 14886 6225
rect 14830 6151 14886 6160
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14936 5953 14964 6054
rect 14922 5944 14978 5953
rect 14922 5879 14924 5888
rect 14976 5879 14978 5888
rect 14924 5850 14976 5856
rect 14832 5840 14884 5846
rect 14830 5808 14832 5817
rect 14884 5808 14886 5817
rect 14830 5743 14886 5752
rect 14922 5672 14978 5681
rect 14832 5636 14884 5642
rect 14922 5607 14978 5616
rect 14832 5578 14884 5584
rect 14844 5545 14872 5578
rect 14830 5536 14886 5545
rect 14830 5471 14886 5480
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14844 4826 14872 5170
rect 14936 4826 14964 5607
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14924 4820 14976 4826
rect 14924 4762 14976 4768
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 14660 4236 14780 4264
rect 14660 3942 14688 4236
rect 14832 4208 14884 4214
rect 14752 4168 14832 4196
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14648 3460 14700 3466
rect 14648 3402 14700 3408
rect 14516 3148 14596 3176
rect 14464 3130 14516 3136
rect 14464 2984 14516 2990
rect 14516 2944 14596 2972
rect 14464 2926 14516 2932
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 14068 2748 14376 2768
rect 14068 2746 14074 2748
rect 14130 2746 14154 2748
rect 14210 2746 14234 2748
rect 14290 2746 14314 2748
rect 14370 2746 14376 2748
rect 14130 2694 14132 2746
rect 14312 2694 14314 2746
rect 14068 2692 14074 2694
rect 14130 2692 14154 2694
rect 14210 2692 14234 2694
rect 14290 2692 14314 2694
rect 14370 2692 14376 2694
rect 14068 2672 14376 2692
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 14096 2576 14148 2582
rect 14096 2518 14148 2524
rect 14108 1057 14136 2518
rect 14280 2372 14332 2378
rect 14280 2314 14332 2320
rect 14094 1048 14150 1057
rect 14094 983 14150 992
rect 14186 912 14242 921
rect 14292 898 14320 2314
rect 14476 1986 14504 2790
rect 14242 870 14320 898
rect 14384 1958 14504 1986
rect 14186 847 14242 856
rect 14200 800 14228 847
rect 13542 31 13598 40
rect 13636 60 13688 66
rect 13636 2 13688 8
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14384 134 14412 1958
rect 14568 1850 14596 2944
rect 14476 1822 14596 1850
rect 14476 1222 14504 1822
rect 14660 1290 14688 3402
rect 14752 2553 14780 4168
rect 14832 4150 14884 4156
rect 14936 4146 14964 4626
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 14936 4049 14964 4082
rect 14922 4040 14978 4049
rect 14832 4004 14884 4010
rect 14922 3975 14978 3984
rect 14832 3946 14884 3952
rect 14844 3233 14872 3946
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14830 3224 14886 3233
rect 14830 3159 14886 3168
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14738 2544 14794 2553
rect 14738 2479 14794 2488
rect 14740 2372 14792 2378
rect 14740 2314 14792 2320
rect 14648 1284 14700 1290
rect 14648 1226 14700 1232
rect 14464 1216 14516 1222
rect 14752 1170 14780 2314
rect 14464 1158 14516 1164
rect 14568 1142 14780 1170
rect 14568 800 14596 1142
rect 14844 800 14872 2994
rect 14936 1902 14964 3878
rect 15028 2106 15056 7142
rect 15120 6746 15148 7754
rect 15304 7750 15332 9046
rect 15396 8514 15424 11086
rect 15488 9178 15516 13806
rect 15580 12434 15608 15506
rect 15580 12406 15700 12434
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15580 11354 15608 11494
rect 15568 11348 15620 11354
rect 15568 11290 15620 11296
rect 15568 11076 15620 11082
rect 15568 11018 15620 11024
rect 15476 9172 15528 9178
rect 15476 9114 15528 9120
rect 15580 8634 15608 11018
rect 15672 10690 15700 12406
rect 15764 11082 15792 15846
rect 15856 12986 15884 19200
rect 16118 17912 16174 17921
rect 16118 17847 16174 17856
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15672 10662 15792 10690
rect 15658 10568 15714 10577
rect 15658 10503 15714 10512
rect 15672 10266 15700 10503
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15672 8906 15700 10202
rect 15660 8900 15712 8906
rect 15660 8842 15712 8848
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15396 8486 15608 8514
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 15474 7984 15530 7993
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15200 7472 15252 7478
rect 15198 7440 15200 7449
rect 15252 7440 15254 7449
rect 15198 7375 15254 7384
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 15212 6866 15240 7210
rect 15200 6860 15252 6866
rect 15200 6802 15252 6808
rect 15120 6718 15240 6746
rect 15108 6656 15160 6662
rect 15108 6598 15160 6604
rect 15120 5273 15148 6598
rect 15106 5264 15162 5273
rect 15106 5199 15162 5208
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 15120 4622 15148 4762
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 15016 2100 15068 2106
rect 15016 2042 15068 2048
rect 14924 1896 14976 1902
rect 14924 1838 14976 1844
rect 15120 1018 15148 3334
rect 15212 3194 15240 6718
rect 15304 5370 15332 7278
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15304 4826 15332 5034
rect 15292 4820 15344 4826
rect 15292 4762 15344 4768
rect 15396 4729 15424 7958
rect 15474 7919 15476 7928
rect 15528 7919 15530 7928
rect 15476 7890 15528 7896
rect 15474 7712 15530 7721
rect 15474 7647 15530 7656
rect 15488 5370 15516 7647
rect 15580 7002 15608 8486
rect 15660 8424 15712 8430
rect 15660 8366 15712 8372
rect 15672 7886 15700 8366
rect 15660 7880 15712 7886
rect 15660 7822 15712 7828
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15566 6488 15622 6497
rect 15566 6423 15622 6432
rect 15476 5364 15528 5370
rect 15476 5306 15528 5312
rect 15580 5302 15608 6423
rect 15672 6186 15700 7686
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15658 6080 15714 6089
rect 15658 6015 15714 6024
rect 15568 5296 15620 5302
rect 15474 5264 15530 5273
rect 15568 5238 15620 5244
rect 15474 5199 15530 5208
rect 15488 5166 15516 5199
rect 15476 5160 15528 5166
rect 15476 5102 15528 5108
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15476 4752 15528 4758
rect 15382 4720 15438 4729
rect 15476 4694 15528 4700
rect 15382 4655 15438 4664
rect 15384 4616 15436 4622
rect 15290 4584 15346 4593
rect 15384 4558 15436 4564
rect 15290 4519 15292 4528
rect 15344 4519 15346 4528
rect 15292 4490 15344 4496
rect 15396 3738 15424 4558
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15304 3534 15332 3674
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15396 2990 15424 3130
rect 15384 2984 15436 2990
rect 15212 2944 15384 2972
rect 15108 1012 15160 1018
rect 15108 954 15160 960
rect 15212 800 15240 2944
rect 15384 2926 15436 2932
rect 15488 2774 15516 4694
rect 15580 3534 15608 4966
rect 15672 4690 15700 6015
rect 15764 5778 15792 10662
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15856 5710 15884 11290
rect 15948 7857 15976 11630
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 15934 7848 15990 7857
rect 15934 7783 15990 7792
rect 16040 6322 16068 11562
rect 16132 9217 16160 17847
rect 16224 12918 16252 19200
rect 16394 18320 16450 18329
rect 16394 18255 16450 18264
rect 16212 12912 16264 12918
rect 16212 12854 16264 12860
rect 16224 11937 16252 12854
rect 16210 11928 16266 11937
rect 16210 11863 16266 11872
rect 16212 11824 16264 11830
rect 16212 11766 16264 11772
rect 16224 10810 16252 11766
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16118 9208 16174 9217
rect 16118 9143 16174 9152
rect 16120 9104 16172 9110
rect 16120 9046 16172 9052
rect 16132 8090 16160 9046
rect 16224 8838 16252 10746
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16210 8528 16266 8537
rect 16210 8463 16266 8472
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 16028 6316 16080 6322
rect 16028 6258 16080 6264
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15752 5636 15804 5642
rect 15752 5578 15804 5584
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15764 4570 15792 5578
rect 15672 4542 15792 4570
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15396 2746 15516 2774
rect 14372 128 14424 134
rect 14372 70 14424 76
rect 14554 0 14610 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15396 202 15424 2746
rect 15672 2582 15700 4542
rect 15752 4480 15804 4486
rect 15752 4422 15804 4428
rect 15660 2576 15712 2582
rect 15660 2518 15712 2524
rect 15568 2508 15620 2514
rect 15568 2450 15620 2456
rect 15580 800 15608 2450
rect 15764 2446 15792 4422
rect 15856 3058 15884 5646
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15948 2922 15976 6054
rect 16040 5642 16068 6122
rect 16028 5636 16080 5642
rect 16028 5578 16080 5584
rect 16132 5234 16160 7754
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 15936 2916 15988 2922
rect 15936 2858 15988 2864
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 15936 2372 15988 2378
rect 15936 2314 15988 2320
rect 15948 800 15976 2314
rect 16224 800 16252 8463
rect 16316 5846 16344 11698
rect 16408 9489 16436 18255
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 16394 9480 16450 9489
rect 16394 9415 16450 9424
rect 16500 9081 16528 12106
rect 16592 11286 16620 19200
rect 16960 12374 16988 19200
rect 16948 12368 17000 12374
rect 16948 12310 17000 12316
rect 16672 12096 16724 12102
rect 16672 12038 16724 12044
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16592 9110 16620 10474
rect 16580 9104 16632 9110
rect 16486 9072 16542 9081
rect 16580 9046 16632 9052
rect 16486 9007 16542 9016
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16304 5840 16356 5846
rect 16304 5782 16356 5788
rect 16316 4185 16344 5782
rect 16408 5030 16436 8774
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16500 4486 16528 9007
rect 16578 8392 16634 8401
rect 16578 8327 16634 8336
rect 16592 5914 16620 8327
rect 16580 5908 16632 5914
rect 16580 5850 16632 5856
rect 16488 4480 16540 4486
rect 16488 4422 16540 4428
rect 16592 4298 16620 5850
rect 16500 4270 16620 4298
rect 16302 4176 16358 4185
rect 16302 4111 16358 4120
rect 16316 1562 16344 4111
rect 16500 2310 16528 4270
rect 16684 3194 16712 12038
rect 16764 8288 16816 8294
rect 16764 8230 16816 8236
rect 16776 5574 16804 8230
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16672 3188 16724 3194
rect 16672 3130 16724 3136
rect 16948 3120 17000 3126
rect 16948 3062 17000 3068
rect 16580 2984 16632 2990
rect 16580 2926 16632 2932
rect 16488 2304 16540 2310
rect 16488 2246 16540 2252
rect 16304 1556 16356 1562
rect 16304 1498 16356 1504
rect 16592 800 16620 2926
rect 16960 800 16988 3062
rect 15384 196 15436 202
rect 15384 138 15436 144
rect 15566 0 15622 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16946 0 17002 800
<< via2 >>
rect 1398 17856 1454 17912
rect 570 15816 626 15872
rect 202 15680 258 15736
rect 1490 15544 1546 15600
rect 1030 7928 1086 7984
rect 1582 14592 1638 14648
rect 1674 14320 1730 14376
rect 1306 13912 1362 13968
rect 1306 11736 1362 11792
rect 1398 9424 1454 9480
rect 1214 2080 1270 2136
rect 386 992 442 1048
rect 1582 13368 1638 13424
rect 2134 16496 2190 16552
rect 1950 14476 2006 14512
rect 1950 14456 1952 14476
rect 1952 14456 2004 14476
rect 2004 14456 2006 14476
rect 1766 12552 1822 12608
rect 1582 11892 1638 11928
rect 1582 11872 1584 11892
rect 1584 11872 1636 11892
rect 1636 11872 1638 11892
rect 1674 11328 1730 11384
rect 2226 15408 2282 15464
rect 1858 11056 1914 11112
rect 2134 12824 2190 12880
rect 2134 12688 2190 12744
rect 1674 9036 1730 9072
rect 1674 9016 1676 9036
rect 1676 9016 1728 9036
rect 1728 9016 1730 9036
rect 2594 17720 2650 17776
rect 2226 12416 2282 12472
rect 2226 12144 2282 12200
rect 2226 11056 2282 11112
rect 2134 10512 2190 10568
rect 1858 8880 1914 8936
rect 2134 9424 2190 9480
rect 2318 9968 2374 10024
rect 1766 6840 1822 6896
rect 1582 4684 1638 4720
rect 1582 4664 1584 4684
rect 1584 4664 1636 4684
rect 1636 4664 1638 4684
rect 1674 3984 1730 4040
rect 4066 19352 4122 19408
rect 2830 16890 2886 16892
rect 2910 16890 2966 16892
rect 2990 16890 3046 16892
rect 3070 16890 3126 16892
rect 2830 16838 2876 16890
rect 2876 16838 2886 16890
rect 2910 16838 2940 16890
rect 2940 16838 2952 16890
rect 2952 16838 2966 16890
rect 2990 16838 3004 16890
rect 3004 16838 3016 16890
rect 3016 16838 3046 16890
rect 3070 16838 3080 16890
rect 3080 16838 3126 16890
rect 2830 16836 2886 16838
rect 2910 16836 2966 16838
rect 2990 16836 3046 16838
rect 3070 16836 3126 16838
rect 2830 15802 2886 15804
rect 2910 15802 2966 15804
rect 2990 15802 3046 15804
rect 3070 15802 3126 15804
rect 2830 15750 2876 15802
rect 2876 15750 2886 15802
rect 2910 15750 2940 15802
rect 2940 15750 2952 15802
rect 2952 15750 2966 15802
rect 2990 15750 3004 15802
rect 3004 15750 3016 15802
rect 3016 15750 3046 15802
rect 3070 15750 3080 15802
rect 3080 15750 3126 15802
rect 2830 15748 2886 15750
rect 2910 15748 2966 15750
rect 2990 15748 3046 15750
rect 3070 15748 3126 15750
rect 2830 14714 2886 14716
rect 2910 14714 2966 14716
rect 2990 14714 3046 14716
rect 3070 14714 3126 14716
rect 2830 14662 2876 14714
rect 2876 14662 2886 14714
rect 2910 14662 2940 14714
rect 2940 14662 2952 14714
rect 2952 14662 2966 14714
rect 2990 14662 3004 14714
rect 3004 14662 3016 14714
rect 3016 14662 3046 14714
rect 3070 14662 3080 14714
rect 3080 14662 3126 14714
rect 2830 14660 2886 14662
rect 2910 14660 2966 14662
rect 2990 14660 3046 14662
rect 3070 14660 3126 14662
rect 3054 14320 3110 14376
rect 2830 13626 2886 13628
rect 2910 13626 2966 13628
rect 2990 13626 3046 13628
rect 3070 13626 3126 13628
rect 2830 13574 2876 13626
rect 2876 13574 2886 13626
rect 2910 13574 2940 13626
rect 2940 13574 2952 13626
rect 2952 13574 2966 13626
rect 2990 13574 3004 13626
rect 3004 13574 3016 13626
rect 3016 13574 3046 13626
rect 3070 13574 3080 13626
rect 3080 13574 3126 13626
rect 2830 13572 2886 13574
rect 2910 13572 2966 13574
rect 2990 13572 3046 13574
rect 3070 13572 3126 13574
rect 3422 16360 3478 16416
rect 3330 14592 3386 14648
rect 3330 14048 3386 14104
rect 3790 16088 3846 16144
rect 3514 15136 3570 15192
rect 3698 15020 3754 15056
rect 3698 15000 3700 15020
rect 3700 15000 3752 15020
rect 3752 15000 3754 15020
rect 3974 18400 4030 18456
rect 3882 14864 3938 14920
rect 3606 14728 3662 14784
rect 3514 14184 3570 14240
rect 3514 13948 3516 13968
rect 3516 13948 3568 13968
rect 3568 13948 3570 13968
rect 3514 13912 3570 13948
rect 2778 12688 2834 12744
rect 3330 13368 3386 13424
rect 2830 12538 2886 12540
rect 2910 12538 2966 12540
rect 2990 12538 3046 12540
rect 3070 12538 3126 12540
rect 2830 12486 2876 12538
rect 2876 12486 2886 12538
rect 2910 12486 2940 12538
rect 2940 12486 2952 12538
rect 2952 12486 2966 12538
rect 2990 12486 3004 12538
rect 3004 12486 3016 12538
rect 3016 12486 3046 12538
rect 3070 12486 3080 12538
rect 3080 12486 3126 12538
rect 2830 12484 2886 12486
rect 2910 12484 2966 12486
rect 2990 12484 3046 12486
rect 3070 12484 3126 12486
rect 2778 12144 2834 12200
rect 2686 11892 2742 11928
rect 2686 11872 2688 11892
rect 2688 11872 2740 11892
rect 2740 11872 2742 11892
rect 2830 11450 2886 11452
rect 2910 11450 2966 11452
rect 2990 11450 3046 11452
rect 3070 11450 3126 11452
rect 2830 11398 2876 11450
rect 2876 11398 2886 11450
rect 2910 11398 2940 11450
rect 2940 11398 2952 11450
rect 2952 11398 2966 11450
rect 2990 11398 3004 11450
rect 3004 11398 3016 11450
rect 3016 11398 3046 11450
rect 3070 11398 3080 11450
rect 3080 11398 3126 11450
rect 2830 11396 2886 11398
rect 2910 11396 2966 11398
rect 2990 11396 3046 11398
rect 3070 11396 3126 11398
rect 2594 10784 2650 10840
rect 2778 10784 2834 10840
rect 2830 10362 2886 10364
rect 2910 10362 2966 10364
rect 2990 10362 3046 10364
rect 3070 10362 3126 10364
rect 2830 10310 2876 10362
rect 2876 10310 2886 10362
rect 2910 10310 2940 10362
rect 2940 10310 2952 10362
rect 2952 10310 2966 10362
rect 2990 10310 3004 10362
rect 3004 10310 3016 10362
rect 3016 10310 3046 10362
rect 3070 10310 3080 10362
rect 3080 10310 3126 10362
rect 2830 10308 2886 10310
rect 2910 10308 2966 10310
rect 2990 10308 3046 10310
rect 3070 10308 3126 10310
rect 2594 9832 2650 9888
rect 2962 9580 3018 9616
rect 2962 9560 2964 9580
rect 2964 9560 3016 9580
rect 3016 9560 3018 9580
rect 2318 8472 2374 8528
rect 2226 6568 2282 6624
rect 2134 5480 2190 5536
rect 2410 6704 2466 6760
rect 2318 5616 2374 5672
rect 2226 4392 2282 4448
rect 2134 2760 2190 2816
rect 2042 2488 2098 2544
rect 1858 2216 1914 2272
rect 1950 1672 2006 1728
rect 1214 40 1270 96
rect 2594 6568 2650 6624
rect 2502 4392 2558 4448
rect 2830 9274 2886 9276
rect 2910 9274 2966 9276
rect 2990 9274 3046 9276
rect 3070 9274 3126 9276
rect 2830 9222 2876 9274
rect 2876 9222 2886 9274
rect 2910 9222 2940 9274
rect 2940 9222 2952 9274
rect 2952 9222 2966 9274
rect 2990 9222 3004 9274
rect 3004 9222 3016 9274
rect 3016 9222 3046 9274
rect 3070 9222 3080 9274
rect 3080 9222 3126 9274
rect 2830 9220 2886 9222
rect 2910 9220 2966 9222
rect 2990 9220 3046 9222
rect 3070 9220 3126 9222
rect 3330 11328 3386 11384
rect 3330 10648 3386 10704
rect 3606 13232 3662 13288
rect 3882 14184 3938 14240
rect 3790 13776 3846 13832
rect 3790 13640 3846 13696
rect 3698 12416 3754 12472
rect 3698 12280 3754 12336
rect 3514 11192 3570 11248
rect 2830 8186 2886 8188
rect 2910 8186 2966 8188
rect 2990 8186 3046 8188
rect 3070 8186 3126 8188
rect 2830 8134 2876 8186
rect 2876 8134 2886 8186
rect 2910 8134 2940 8186
rect 2940 8134 2952 8186
rect 2952 8134 2966 8186
rect 2990 8134 3004 8186
rect 3004 8134 3016 8186
rect 3016 8134 3046 8186
rect 3070 8134 3080 8186
rect 3080 8134 3126 8186
rect 2830 8132 2886 8134
rect 2910 8132 2966 8134
rect 2990 8132 3046 8134
rect 3070 8132 3126 8134
rect 3146 7384 3202 7440
rect 3054 7268 3110 7304
rect 3054 7248 3056 7268
rect 3056 7248 3108 7268
rect 3108 7248 3110 7268
rect 2830 7098 2886 7100
rect 2910 7098 2966 7100
rect 2990 7098 3046 7100
rect 3070 7098 3126 7100
rect 2830 7046 2876 7098
rect 2876 7046 2886 7098
rect 2910 7046 2940 7098
rect 2940 7046 2952 7098
rect 2952 7046 2966 7098
rect 2990 7046 3004 7098
rect 3004 7046 3016 7098
rect 3016 7046 3046 7098
rect 3070 7046 3080 7098
rect 3080 7046 3126 7098
rect 2830 7044 2886 7046
rect 2910 7044 2966 7046
rect 2990 7044 3046 7046
rect 3070 7044 3126 7046
rect 2830 6010 2886 6012
rect 2910 6010 2966 6012
rect 2990 6010 3046 6012
rect 3070 6010 3126 6012
rect 2830 5958 2876 6010
rect 2876 5958 2886 6010
rect 2910 5958 2940 6010
rect 2940 5958 2952 6010
rect 2952 5958 2966 6010
rect 2990 5958 3004 6010
rect 3004 5958 3016 6010
rect 3016 5958 3046 6010
rect 3070 5958 3080 6010
rect 3080 5958 3126 6010
rect 2830 5956 2886 5958
rect 2910 5956 2966 5958
rect 2990 5956 3046 5958
rect 3070 5956 3126 5958
rect 2830 4922 2886 4924
rect 2910 4922 2966 4924
rect 2990 4922 3046 4924
rect 3070 4922 3126 4924
rect 2830 4870 2876 4922
rect 2876 4870 2886 4922
rect 2910 4870 2940 4922
rect 2940 4870 2952 4922
rect 2952 4870 2966 4922
rect 2990 4870 3004 4922
rect 3004 4870 3016 4922
rect 3016 4870 3046 4922
rect 3070 4870 3080 4922
rect 3080 4870 3126 4922
rect 2830 4868 2886 4870
rect 2910 4868 2966 4870
rect 2990 4868 3046 4870
rect 3070 4868 3126 4870
rect 2962 4664 3018 4720
rect 2830 3834 2886 3836
rect 2910 3834 2966 3836
rect 2990 3834 3046 3836
rect 3070 3834 3126 3836
rect 2830 3782 2876 3834
rect 2876 3782 2886 3834
rect 2910 3782 2940 3834
rect 2940 3782 2952 3834
rect 2952 3782 2966 3834
rect 2990 3782 3004 3834
rect 3004 3782 3016 3834
rect 3016 3782 3046 3834
rect 3070 3782 3080 3834
rect 3080 3782 3126 3834
rect 2830 3780 2886 3782
rect 2910 3780 2966 3782
rect 2990 3780 3046 3782
rect 3070 3780 3126 3782
rect 2318 2896 2374 2952
rect 2318 2796 2320 2816
rect 2320 2796 2372 2816
rect 2372 2796 2374 2816
rect 2318 2760 2374 2796
rect 2318 2508 2374 2544
rect 2318 2488 2320 2508
rect 2320 2488 2372 2508
rect 2372 2488 2374 2508
rect 2594 3304 2650 3360
rect 2778 3168 2834 3224
rect 4158 14220 4160 14240
rect 4160 14220 4212 14240
rect 4212 14220 4214 14240
rect 4158 14184 4214 14220
rect 4158 13948 4160 13968
rect 4160 13948 4212 13968
rect 4212 13948 4214 13968
rect 4158 13912 4214 13948
rect 4158 13504 4214 13560
rect 3882 11056 3938 11112
rect 4066 11464 4122 11520
rect 3974 10648 4030 10704
rect 3974 10104 4030 10160
rect 3882 9152 3938 9208
rect 3330 6432 3386 6488
rect 3238 4428 3240 4448
rect 3240 4428 3292 4448
rect 3292 4428 3294 4448
rect 3238 4392 3294 4428
rect 3238 3576 3294 3632
rect 2830 2746 2886 2748
rect 2910 2746 2966 2748
rect 2990 2746 3046 2748
rect 3070 2746 3126 2748
rect 2830 2694 2876 2746
rect 2876 2694 2886 2746
rect 2910 2694 2940 2746
rect 2940 2694 2952 2746
rect 2952 2694 2966 2746
rect 2990 2694 3004 2746
rect 3004 2694 3016 2746
rect 3016 2694 3046 2746
rect 3070 2694 3080 2746
rect 3080 2694 3126 2746
rect 2830 2692 2886 2694
rect 2910 2692 2966 2694
rect 2990 2692 3046 2694
rect 3070 2692 3126 2694
rect 3606 8200 3662 8256
rect 3606 7656 3662 7712
rect 3790 6976 3846 7032
rect 5170 17992 5226 18048
rect 4704 17434 4760 17436
rect 4784 17434 4840 17436
rect 4864 17434 4920 17436
rect 4944 17434 5000 17436
rect 4704 17382 4750 17434
rect 4750 17382 4760 17434
rect 4784 17382 4814 17434
rect 4814 17382 4826 17434
rect 4826 17382 4840 17434
rect 4864 17382 4878 17434
rect 4878 17382 4890 17434
rect 4890 17382 4920 17434
rect 4944 17382 4954 17434
rect 4954 17382 5000 17434
rect 4704 17380 4760 17382
rect 4784 17380 4840 17382
rect 4864 17380 4920 17382
rect 4944 17380 5000 17382
rect 4704 16346 4760 16348
rect 4784 16346 4840 16348
rect 4864 16346 4920 16348
rect 4944 16346 5000 16348
rect 4704 16294 4750 16346
rect 4750 16294 4760 16346
rect 4784 16294 4814 16346
rect 4814 16294 4826 16346
rect 4826 16294 4840 16346
rect 4864 16294 4878 16346
rect 4878 16294 4890 16346
rect 4890 16294 4920 16346
rect 4944 16294 4954 16346
rect 4954 16294 5000 16346
rect 4704 16292 4760 16294
rect 4784 16292 4840 16294
rect 4864 16292 4920 16294
rect 4944 16292 5000 16294
rect 4704 15258 4760 15260
rect 4784 15258 4840 15260
rect 4864 15258 4920 15260
rect 4944 15258 5000 15260
rect 4704 15206 4750 15258
rect 4750 15206 4760 15258
rect 4784 15206 4814 15258
rect 4814 15206 4826 15258
rect 4826 15206 4840 15258
rect 4864 15206 4878 15258
rect 4878 15206 4890 15258
rect 4890 15206 4920 15258
rect 4944 15206 4954 15258
rect 4954 15206 5000 15258
rect 4704 15204 4760 15206
rect 4784 15204 4840 15206
rect 4864 15204 4920 15206
rect 4944 15204 5000 15206
rect 4704 14170 4760 14172
rect 4784 14170 4840 14172
rect 4864 14170 4920 14172
rect 4944 14170 5000 14172
rect 4704 14118 4750 14170
rect 4750 14118 4760 14170
rect 4784 14118 4814 14170
rect 4814 14118 4826 14170
rect 4826 14118 4840 14170
rect 4864 14118 4878 14170
rect 4878 14118 4890 14170
rect 4890 14118 4920 14170
rect 4944 14118 4954 14170
rect 4954 14118 5000 14170
rect 4704 14116 4760 14118
rect 4784 14116 4840 14118
rect 4864 14116 4920 14118
rect 4944 14116 5000 14118
rect 4342 10240 4398 10296
rect 3974 8336 4030 8392
rect 3698 5344 3754 5400
rect 3790 5244 3792 5264
rect 3792 5244 3844 5264
rect 3844 5244 3846 5264
rect 3790 5208 3846 5244
rect 3698 5072 3754 5128
rect 3606 3440 3662 3496
rect 3514 1400 3570 1456
rect 3422 448 3478 504
rect 3974 3304 4030 3360
rect 4704 13082 4760 13084
rect 4784 13082 4840 13084
rect 4864 13082 4920 13084
rect 4944 13082 5000 13084
rect 4704 13030 4750 13082
rect 4750 13030 4760 13082
rect 4784 13030 4814 13082
rect 4814 13030 4826 13082
rect 4826 13030 4840 13082
rect 4864 13030 4878 13082
rect 4878 13030 4890 13082
rect 4890 13030 4920 13082
rect 4944 13030 4954 13082
rect 4954 13030 5000 13082
rect 4704 13028 4760 13030
rect 4784 13028 4840 13030
rect 4864 13028 4920 13030
rect 4944 13028 5000 13030
rect 5354 17448 5410 17504
rect 5262 17312 5318 17368
rect 5170 14048 5226 14104
rect 5354 17040 5410 17096
rect 5354 15408 5410 15464
rect 5630 15408 5686 15464
rect 5630 15136 5686 15192
rect 5630 14728 5686 14784
rect 6090 15680 6146 15736
rect 5906 15408 5962 15464
rect 5814 14592 5870 14648
rect 5538 14356 5540 14376
rect 5540 14356 5592 14376
rect 5592 14356 5594 14376
rect 5538 14320 5594 14356
rect 5446 13932 5502 13968
rect 5446 13912 5448 13932
rect 5448 13912 5500 13932
rect 5500 13912 5502 13932
rect 5354 13776 5410 13832
rect 5446 13232 5502 13288
rect 4986 12144 5042 12200
rect 5078 12008 5134 12064
rect 4704 11994 4760 11996
rect 4784 11994 4840 11996
rect 4864 11994 4920 11996
rect 4944 11994 5000 11996
rect 4704 11942 4750 11994
rect 4750 11942 4760 11994
rect 4784 11942 4814 11994
rect 4814 11942 4826 11994
rect 4826 11942 4840 11994
rect 4864 11942 4878 11994
rect 4878 11942 4890 11994
rect 4890 11942 4920 11994
rect 4944 11942 4954 11994
rect 4954 11942 5000 11994
rect 4704 11940 4760 11942
rect 4784 11940 4840 11942
rect 4864 11940 4920 11942
rect 4944 11940 5000 11942
rect 4618 11348 4674 11384
rect 4618 11328 4620 11348
rect 4620 11328 4672 11348
rect 4672 11328 4674 11348
rect 5354 12008 5410 12064
rect 5262 11872 5318 11928
rect 4802 11192 4858 11248
rect 5262 11600 5318 11656
rect 4704 10906 4760 10908
rect 4784 10906 4840 10908
rect 4864 10906 4920 10908
rect 4944 10906 5000 10908
rect 4704 10854 4750 10906
rect 4750 10854 4760 10906
rect 4784 10854 4814 10906
rect 4814 10854 4826 10906
rect 4826 10854 4840 10906
rect 4864 10854 4878 10906
rect 4878 10854 4890 10906
rect 4890 10854 4920 10906
rect 4944 10854 4954 10906
rect 4954 10854 5000 10906
rect 4704 10852 4760 10854
rect 4784 10852 4840 10854
rect 4864 10852 4920 10854
rect 4944 10852 5000 10854
rect 4802 10240 4858 10296
rect 4704 9818 4760 9820
rect 4784 9818 4840 9820
rect 4864 9818 4920 9820
rect 4944 9818 5000 9820
rect 4704 9766 4750 9818
rect 4750 9766 4760 9818
rect 4784 9766 4814 9818
rect 4814 9766 4826 9818
rect 4826 9766 4840 9818
rect 4864 9766 4878 9818
rect 4878 9766 4890 9818
rect 4890 9766 4920 9818
rect 4944 9766 4954 9818
rect 4954 9766 5000 9818
rect 4704 9764 4760 9766
rect 4784 9764 4840 9766
rect 4864 9764 4920 9766
rect 4944 9764 5000 9766
rect 5078 9696 5134 9752
rect 4704 8730 4760 8732
rect 4784 8730 4840 8732
rect 4864 8730 4920 8732
rect 4944 8730 5000 8732
rect 4704 8678 4750 8730
rect 4750 8678 4760 8730
rect 4784 8678 4814 8730
rect 4814 8678 4826 8730
rect 4826 8678 4840 8730
rect 4864 8678 4878 8730
rect 4878 8678 4890 8730
rect 4890 8678 4920 8730
rect 4944 8678 4954 8730
rect 4954 8678 5000 8730
rect 4704 8676 4760 8678
rect 4784 8676 4840 8678
rect 4864 8676 4920 8678
rect 4944 8676 5000 8678
rect 4704 7642 4760 7644
rect 4784 7642 4840 7644
rect 4864 7642 4920 7644
rect 4944 7642 5000 7644
rect 4704 7590 4750 7642
rect 4750 7590 4760 7642
rect 4784 7590 4814 7642
rect 4814 7590 4826 7642
rect 4826 7590 4840 7642
rect 4864 7590 4878 7642
rect 4878 7590 4890 7642
rect 4890 7590 4920 7642
rect 4944 7590 4954 7642
rect 4954 7590 5000 7642
rect 4704 7588 4760 7590
rect 4784 7588 4840 7590
rect 4864 7588 4920 7590
rect 4944 7588 5000 7590
rect 4526 6976 4582 7032
rect 4434 6840 4490 6896
rect 4704 6554 4760 6556
rect 4784 6554 4840 6556
rect 4864 6554 4920 6556
rect 4944 6554 5000 6556
rect 4704 6502 4750 6554
rect 4750 6502 4760 6554
rect 4784 6502 4814 6554
rect 4814 6502 4826 6554
rect 4826 6502 4840 6554
rect 4864 6502 4878 6554
rect 4878 6502 4890 6554
rect 4890 6502 4920 6554
rect 4944 6502 4954 6554
rect 4954 6502 5000 6554
rect 4704 6500 4760 6502
rect 4784 6500 4840 6502
rect 4864 6500 4920 6502
rect 4944 6500 5000 6502
rect 4158 4120 4214 4176
rect 4250 3168 4306 3224
rect 3974 2352 4030 2408
rect 4894 6296 4950 6352
rect 4618 5888 4674 5944
rect 4894 5752 4950 5808
rect 5078 5752 5134 5808
rect 5630 13504 5686 13560
rect 6090 14728 6146 14784
rect 5998 13776 6054 13832
rect 5906 13640 5962 13696
rect 5722 13368 5778 13424
rect 5538 12552 5594 12608
rect 5538 12280 5594 12336
rect 5446 11600 5502 11656
rect 5906 12960 5962 13016
rect 5814 12416 5870 12472
rect 5722 12044 5724 12064
rect 5724 12044 5776 12064
rect 5776 12044 5778 12064
rect 5722 12008 5778 12044
rect 5630 11056 5686 11112
rect 5630 10804 5686 10840
rect 5630 10784 5632 10804
rect 5632 10784 5684 10804
rect 5684 10784 5686 10804
rect 5538 9424 5594 9480
rect 5446 9152 5502 9208
rect 5814 11328 5870 11384
rect 5998 12280 6054 12336
rect 6182 13776 6238 13832
rect 6578 16890 6634 16892
rect 6658 16890 6714 16892
rect 6738 16890 6794 16892
rect 6818 16890 6874 16892
rect 6578 16838 6624 16890
rect 6624 16838 6634 16890
rect 6658 16838 6688 16890
rect 6688 16838 6700 16890
rect 6700 16838 6714 16890
rect 6738 16838 6752 16890
rect 6752 16838 6764 16890
rect 6764 16838 6794 16890
rect 6818 16838 6828 16890
rect 6828 16838 6874 16890
rect 6578 16836 6634 16838
rect 6658 16836 6714 16838
rect 6738 16836 6794 16838
rect 6818 16836 6874 16838
rect 7010 15952 7066 16008
rect 6578 15802 6634 15804
rect 6658 15802 6714 15804
rect 6738 15802 6794 15804
rect 6818 15802 6874 15804
rect 6578 15750 6624 15802
rect 6624 15750 6634 15802
rect 6658 15750 6688 15802
rect 6688 15750 6700 15802
rect 6700 15750 6714 15802
rect 6738 15750 6752 15802
rect 6752 15750 6764 15802
rect 6764 15750 6794 15802
rect 6818 15750 6828 15802
rect 6828 15750 6874 15802
rect 6578 15748 6634 15750
rect 6658 15748 6714 15750
rect 6738 15748 6794 15750
rect 6818 15748 6874 15750
rect 6578 14714 6634 14716
rect 6658 14714 6714 14716
rect 6738 14714 6794 14716
rect 6818 14714 6874 14716
rect 6578 14662 6624 14714
rect 6624 14662 6634 14714
rect 6658 14662 6688 14714
rect 6688 14662 6700 14714
rect 6700 14662 6714 14714
rect 6738 14662 6752 14714
rect 6752 14662 6764 14714
rect 6764 14662 6794 14714
rect 6818 14662 6828 14714
rect 6828 14662 6874 14714
rect 6578 14660 6634 14662
rect 6658 14660 6714 14662
rect 6738 14660 6794 14662
rect 6818 14660 6874 14662
rect 6734 14320 6790 14376
rect 6642 14184 6698 14240
rect 6918 14320 6974 14376
rect 6826 14184 6882 14240
rect 6578 13626 6634 13628
rect 6658 13626 6714 13628
rect 6738 13626 6794 13628
rect 6818 13626 6874 13628
rect 6578 13574 6624 13626
rect 6624 13574 6634 13626
rect 6658 13574 6688 13626
rect 6688 13574 6700 13626
rect 6700 13574 6714 13626
rect 6738 13574 6752 13626
rect 6752 13574 6764 13626
rect 6764 13574 6794 13626
rect 6818 13574 6828 13626
rect 6828 13574 6874 13626
rect 6578 13572 6634 13574
rect 6658 13572 6714 13574
rect 6738 13572 6794 13574
rect 6818 13572 6874 13574
rect 7010 13912 7066 13968
rect 7562 17720 7618 17776
rect 7562 17176 7618 17232
rect 7378 15000 7434 15056
rect 6366 12688 6422 12744
rect 6090 11464 6146 11520
rect 6090 11056 6146 11112
rect 5998 10920 6054 10976
rect 5814 8880 5870 8936
rect 5538 8336 5594 8392
rect 5354 6024 5410 6080
rect 4704 5466 4760 5468
rect 4784 5466 4840 5468
rect 4864 5466 4920 5468
rect 4944 5466 5000 5468
rect 4704 5414 4750 5466
rect 4750 5414 4760 5466
rect 4784 5414 4814 5466
rect 4814 5414 4826 5466
rect 4826 5414 4840 5466
rect 4864 5414 4878 5466
rect 4878 5414 4890 5466
rect 4890 5414 4920 5466
rect 4944 5414 4954 5466
rect 4954 5414 5000 5466
rect 4704 5412 4760 5414
rect 4784 5412 4840 5414
rect 4864 5412 4920 5414
rect 4944 5412 5000 5414
rect 4704 4378 4760 4380
rect 4784 4378 4840 4380
rect 4864 4378 4920 4380
rect 4944 4378 5000 4380
rect 4704 4326 4750 4378
rect 4750 4326 4760 4378
rect 4784 4326 4814 4378
rect 4814 4326 4826 4378
rect 4826 4326 4840 4378
rect 4864 4326 4878 4378
rect 4878 4326 4890 4378
rect 4890 4326 4920 4378
rect 4944 4326 4954 4378
rect 4954 4326 5000 4378
rect 4704 4324 4760 4326
rect 4784 4324 4840 4326
rect 4864 4324 4920 4326
rect 4944 4324 5000 4326
rect 5170 4528 5226 4584
rect 4704 3290 4760 3292
rect 4784 3290 4840 3292
rect 4864 3290 4920 3292
rect 4944 3290 5000 3292
rect 4704 3238 4750 3290
rect 4750 3238 4760 3290
rect 4784 3238 4814 3290
rect 4814 3238 4826 3290
rect 4826 3238 4840 3290
rect 4864 3238 4878 3290
rect 4878 3238 4890 3290
rect 4890 3238 4920 3290
rect 4944 3238 4954 3290
rect 4954 3238 5000 3290
rect 4704 3236 4760 3238
rect 4784 3236 4840 3238
rect 4864 3236 4920 3238
rect 4944 3236 5000 3238
rect 4710 2760 4766 2816
rect 4526 2644 4582 2680
rect 4526 2624 4528 2644
rect 4528 2624 4580 2644
rect 4580 2624 4582 2644
rect 4526 2080 4582 2136
rect 4704 2202 4760 2204
rect 4784 2202 4840 2204
rect 4864 2202 4920 2204
rect 4944 2202 5000 2204
rect 4704 2150 4750 2202
rect 4750 2150 4760 2202
rect 4784 2150 4814 2202
rect 4814 2150 4826 2202
rect 4826 2150 4840 2202
rect 4864 2150 4878 2202
rect 4878 2150 4890 2202
rect 4890 2150 4920 2202
rect 4944 2150 4954 2202
rect 4954 2150 5000 2202
rect 4704 2148 4760 2150
rect 4784 2148 4840 2150
rect 4864 2148 4920 2150
rect 4944 2148 5000 2150
rect 5262 4392 5318 4448
rect 5814 8064 5870 8120
rect 5630 7948 5686 7984
rect 5630 7928 5632 7948
rect 5632 7928 5684 7948
rect 5684 7928 5686 7948
rect 5538 5616 5594 5672
rect 5630 3440 5686 3496
rect 5538 2760 5594 2816
rect 5446 2488 5502 2544
rect 5906 7792 5962 7848
rect 5998 7656 6054 7712
rect 6366 12008 6422 12064
rect 6918 13368 6974 13424
rect 7102 13524 7158 13560
rect 7102 13504 7104 13524
rect 7104 13504 7156 13524
rect 7156 13504 7158 13524
rect 6578 12538 6634 12540
rect 6658 12538 6714 12540
rect 6738 12538 6794 12540
rect 6818 12538 6874 12540
rect 6578 12486 6624 12538
rect 6624 12486 6634 12538
rect 6658 12486 6688 12538
rect 6688 12486 6700 12538
rect 6700 12486 6714 12538
rect 6738 12486 6752 12538
rect 6752 12486 6764 12538
rect 6764 12486 6794 12538
rect 6818 12486 6828 12538
rect 6828 12486 6874 12538
rect 6578 12484 6634 12486
rect 6658 12484 6714 12486
rect 6738 12484 6794 12486
rect 6818 12484 6874 12486
rect 6274 9832 6330 9888
rect 6826 12008 6882 12064
rect 6578 11450 6634 11452
rect 6658 11450 6714 11452
rect 6738 11450 6794 11452
rect 6818 11450 6874 11452
rect 6578 11398 6624 11450
rect 6624 11398 6634 11450
rect 6658 11398 6688 11450
rect 6688 11398 6700 11450
rect 6700 11398 6714 11450
rect 6738 11398 6752 11450
rect 6752 11398 6764 11450
rect 6764 11398 6794 11450
rect 6818 11398 6828 11450
rect 6828 11398 6874 11450
rect 6578 11396 6634 11398
rect 6658 11396 6714 11398
rect 6738 11396 6794 11398
rect 6818 11396 6874 11398
rect 6826 10784 6882 10840
rect 7194 12824 7250 12880
rect 7194 12708 7250 12744
rect 7194 12688 7196 12708
rect 7196 12688 7248 12708
rect 7248 12688 7250 12708
rect 7102 12144 7158 12200
rect 6578 10362 6634 10364
rect 6658 10362 6714 10364
rect 6738 10362 6794 10364
rect 6818 10362 6874 10364
rect 6578 10310 6624 10362
rect 6624 10310 6634 10362
rect 6658 10310 6688 10362
rect 6688 10310 6700 10362
rect 6700 10310 6714 10362
rect 6738 10310 6752 10362
rect 6752 10310 6764 10362
rect 6764 10310 6794 10362
rect 6818 10310 6828 10362
rect 6828 10310 6874 10362
rect 6578 10308 6634 10310
rect 6658 10308 6714 10310
rect 6738 10308 6794 10310
rect 6818 10308 6874 10310
rect 7194 11736 7250 11792
rect 7746 15700 7802 15736
rect 7746 15680 7748 15700
rect 7748 15680 7800 15700
rect 7800 15680 7802 15700
rect 7838 15272 7894 15328
rect 7838 15136 7894 15192
rect 7746 14728 7802 14784
rect 7838 14592 7894 14648
rect 8022 14592 8078 14648
rect 7102 10376 7158 10432
rect 7010 10240 7066 10296
rect 6918 9424 6974 9480
rect 6578 9274 6634 9276
rect 6658 9274 6714 9276
rect 6738 9274 6794 9276
rect 6818 9274 6874 9276
rect 6578 9222 6624 9274
rect 6624 9222 6634 9274
rect 6658 9222 6688 9274
rect 6688 9222 6700 9274
rect 6700 9222 6714 9274
rect 6738 9222 6752 9274
rect 6752 9222 6764 9274
rect 6764 9222 6794 9274
rect 6818 9222 6828 9274
rect 6828 9222 6874 9274
rect 6578 9220 6634 9222
rect 6658 9220 6714 9222
rect 6738 9220 6794 9222
rect 6818 9220 6874 9222
rect 6578 8186 6634 8188
rect 6658 8186 6714 8188
rect 6738 8186 6794 8188
rect 6818 8186 6874 8188
rect 6578 8134 6624 8186
rect 6624 8134 6634 8186
rect 6658 8134 6688 8186
rect 6688 8134 6700 8186
rect 6700 8134 6714 8186
rect 6738 8134 6752 8186
rect 6752 8134 6764 8186
rect 6764 8134 6794 8186
rect 6818 8134 6828 8186
rect 6828 8134 6874 8186
rect 6578 8132 6634 8134
rect 6658 8132 6714 8134
rect 6738 8132 6794 8134
rect 6818 8132 6874 8134
rect 6090 6840 6146 6896
rect 7010 8900 7066 8936
rect 7010 8880 7012 8900
rect 7012 8880 7064 8900
rect 7064 8880 7066 8900
rect 6458 7248 6514 7304
rect 6918 7248 6974 7304
rect 6578 7098 6634 7100
rect 6658 7098 6714 7100
rect 6738 7098 6794 7100
rect 6818 7098 6874 7100
rect 6578 7046 6624 7098
rect 6624 7046 6634 7098
rect 6658 7046 6688 7098
rect 6688 7046 6700 7098
rect 6700 7046 6714 7098
rect 6738 7046 6752 7098
rect 6752 7046 6764 7098
rect 6764 7046 6794 7098
rect 6818 7046 6828 7098
rect 6828 7046 6874 7098
rect 6578 7044 6634 7046
rect 6658 7044 6714 7046
rect 6738 7044 6794 7046
rect 6818 7044 6874 7046
rect 5814 3304 5870 3360
rect 5906 3168 5962 3224
rect 6578 6010 6634 6012
rect 6658 6010 6714 6012
rect 6738 6010 6794 6012
rect 6818 6010 6874 6012
rect 6578 5958 6624 6010
rect 6624 5958 6634 6010
rect 6658 5958 6688 6010
rect 6688 5958 6700 6010
rect 6700 5958 6714 6010
rect 6738 5958 6752 6010
rect 6752 5958 6764 6010
rect 6764 5958 6794 6010
rect 6818 5958 6828 6010
rect 6828 5958 6874 6010
rect 6578 5956 6634 5958
rect 6658 5956 6714 5958
rect 6738 5956 6794 5958
rect 6818 5956 6874 5958
rect 6090 2760 6146 2816
rect 5906 2624 5962 2680
rect 5814 2488 5870 2544
rect 6090 2216 6146 2272
rect 7746 14048 7802 14104
rect 7746 13640 7802 13696
rect 7286 9288 7342 9344
rect 7470 8880 7526 8936
rect 7286 7656 7342 7712
rect 7286 7112 7342 7168
rect 7102 6996 7158 7032
rect 7102 6976 7104 6996
rect 7104 6976 7156 6996
rect 7156 6976 7158 6996
rect 6918 5208 6974 5264
rect 6578 4922 6634 4924
rect 6658 4922 6714 4924
rect 6738 4922 6794 4924
rect 6818 4922 6874 4924
rect 6578 4870 6624 4922
rect 6624 4870 6634 4922
rect 6658 4870 6688 4922
rect 6688 4870 6700 4922
rect 6700 4870 6714 4922
rect 6738 4870 6752 4922
rect 6752 4870 6764 4922
rect 6764 4870 6794 4922
rect 6818 4870 6828 4922
rect 6828 4870 6874 4922
rect 6578 4868 6634 4870
rect 6658 4868 6714 4870
rect 6738 4868 6794 4870
rect 6818 4868 6874 4870
rect 7102 5072 7158 5128
rect 7102 4800 7158 4856
rect 6550 4020 6552 4040
rect 6552 4020 6604 4040
rect 6604 4020 6606 4040
rect 6550 3984 6606 4020
rect 7010 4120 7066 4176
rect 6826 3984 6882 4040
rect 6578 3834 6634 3836
rect 6658 3834 6714 3836
rect 6738 3834 6794 3836
rect 6818 3834 6874 3836
rect 6578 3782 6624 3834
rect 6624 3782 6634 3834
rect 6658 3782 6688 3834
rect 6688 3782 6700 3834
rect 6700 3782 6714 3834
rect 6738 3782 6752 3834
rect 6752 3782 6764 3834
rect 6764 3782 6794 3834
rect 6818 3782 6828 3834
rect 6828 3782 6874 3834
rect 6578 3780 6634 3782
rect 6658 3780 6714 3782
rect 6738 3780 6794 3782
rect 6818 3780 6874 3782
rect 6366 3032 6422 3088
rect 6274 2896 6330 2952
rect 6578 2746 6634 2748
rect 6658 2746 6714 2748
rect 6738 2746 6794 2748
rect 6818 2746 6874 2748
rect 6578 2694 6624 2746
rect 6624 2694 6634 2746
rect 6658 2694 6688 2746
rect 6688 2694 6700 2746
rect 6700 2694 6714 2746
rect 6738 2694 6752 2746
rect 6752 2694 6764 2746
rect 6764 2694 6794 2746
rect 6818 2694 6828 2746
rect 6828 2694 6874 2746
rect 6578 2692 6634 2694
rect 6658 2692 6714 2694
rect 6738 2692 6794 2694
rect 6818 2692 6874 2694
rect 6826 2524 6828 2544
rect 6828 2524 6880 2544
rect 6880 2524 6882 2544
rect 6826 2488 6882 2524
rect 7470 6296 7526 6352
rect 7746 11328 7802 11384
rect 8022 12960 8078 13016
rect 8022 12280 8078 12336
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8498 17434
rect 8498 17382 8508 17434
rect 8532 17382 8562 17434
rect 8562 17382 8574 17434
rect 8574 17382 8588 17434
rect 8612 17382 8626 17434
rect 8626 17382 8638 17434
rect 8638 17382 8668 17434
rect 8692 17382 8702 17434
rect 8702 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8498 16346
rect 8498 16294 8508 16346
rect 8532 16294 8562 16346
rect 8562 16294 8574 16346
rect 8574 16294 8588 16346
rect 8612 16294 8626 16346
rect 8626 16294 8638 16346
rect 8638 16294 8668 16346
rect 8692 16294 8702 16346
rect 8702 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8498 15258
rect 8498 15206 8508 15258
rect 8532 15206 8562 15258
rect 8562 15206 8574 15258
rect 8574 15206 8588 15258
rect 8612 15206 8626 15258
rect 8626 15206 8638 15258
rect 8638 15206 8668 15258
rect 8692 15206 8702 15258
rect 8702 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8498 14170
rect 8498 14118 8508 14170
rect 8532 14118 8562 14170
rect 8562 14118 8574 14170
rect 8574 14118 8588 14170
rect 8612 14118 8626 14170
rect 8626 14118 8638 14170
rect 8638 14118 8668 14170
rect 8692 14118 8702 14170
rect 8702 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8498 13082
rect 8498 13030 8508 13082
rect 8532 13030 8562 13082
rect 8562 13030 8574 13082
rect 8574 13030 8588 13082
rect 8612 13030 8626 13082
rect 8626 13030 8638 13082
rect 8638 13030 8668 13082
rect 8692 13030 8702 13082
rect 8702 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 8206 12416 8262 12472
rect 8114 11772 8116 11792
rect 8116 11772 8168 11792
rect 8168 11772 8170 11792
rect 8114 11736 8170 11772
rect 8758 12280 8814 12336
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8498 11994
rect 8498 11942 8508 11994
rect 8532 11942 8562 11994
rect 8562 11942 8574 11994
rect 8574 11942 8588 11994
rect 8612 11942 8626 11994
rect 8626 11942 8638 11994
rect 8638 11942 8668 11994
rect 8692 11942 8702 11994
rect 8702 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 8114 11328 8170 11384
rect 7930 10548 7932 10568
rect 7932 10548 7984 10568
rect 7984 10548 7986 10568
rect 7930 10512 7986 10548
rect 7930 9832 7986 9888
rect 8114 10920 8170 10976
rect 8114 10784 8170 10840
rect 8114 9696 8170 9752
rect 7930 7248 7986 7304
rect 7378 5908 7434 5944
rect 7378 5888 7380 5908
rect 7380 5888 7432 5908
rect 7432 5888 7434 5908
rect 7286 4936 7342 4992
rect 7010 1808 7066 1864
rect 7470 4936 7526 4992
rect 7470 3984 7526 4040
rect 7378 3712 7434 3768
rect 7378 3304 7434 3360
rect 7470 3188 7526 3224
rect 7746 4156 7748 4176
rect 7748 4156 7800 4176
rect 7800 4156 7802 4176
rect 7746 4120 7802 4156
rect 7746 3984 7802 4040
rect 7470 3168 7472 3188
rect 7472 3168 7524 3188
rect 7524 3168 7526 3188
rect 7470 2896 7526 2952
rect 7470 2624 7526 2680
rect 8574 11736 8630 11792
rect 9402 14864 9458 14920
rect 9402 14320 9458 14376
rect 9034 12280 9090 12336
rect 9402 14068 9458 14104
rect 9402 14048 9404 14068
rect 9404 14048 9456 14068
rect 9456 14048 9458 14068
rect 9678 17856 9734 17912
rect 9862 17856 9918 17912
rect 9862 16632 9918 16688
rect 9586 15000 9642 15056
rect 9678 14592 9734 14648
rect 10326 16890 10382 16892
rect 10406 16890 10462 16892
rect 10486 16890 10542 16892
rect 10566 16890 10622 16892
rect 10326 16838 10372 16890
rect 10372 16838 10382 16890
rect 10406 16838 10436 16890
rect 10436 16838 10448 16890
rect 10448 16838 10462 16890
rect 10486 16838 10500 16890
rect 10500 16838 10512 16890
rect 10512 16838 10542 16890
rect 10566 16838 10576 16890
rect 10576 16838 10622 16890
rect 10326 16836 10382 16838
rect 10406 16836 10462 16838
rect 10486 16836 10542 16838
rect 10566 16836 10622 16838
rect 10326 15802 10382 15804
rect 10406 15802 10462 15804
rect 10486 15802 10542 15804
rect 10566 15802 10622 15804
rect 10326 15750 10372 15802
rect 10372 15750 10382 15802
rect 10406 15750 10436 15802
rect 10436 15750 10448 15802
rect 10448 15750 10462 15802
rect 10486 15750 10500 15802
rect 10500 15750 10512 15802
rect 10512 15750 10542 15802
rect 10566 15750 10576 15802
rect 10576 15750 10622 15802
rect 10326 15748 10382 15750
rect 10406 15748 10462 15750
rect 10486 15748 10542 15750
rect 10566 15748 10622 15750
rect 9770 13812 9772 13832
rect 9772 13812 9824 13832
rect 9824 13812 9826 13832
rect 9770 13776 9826 13812
rect 10326 14714 10382 14716
rect 10406 14714 10462 14716
rect 10486 14714 10542 14716
rect 10566 14714 10622 14716
rect 10326 14662 10372 14714
rect 10372 14662 10382 14714
rect 10406 14662 10436 14714
rect 10436 14662 10448 14714
rect 10448 14662 10462 14714
rect 10486 14662 10500 14714
rect 10500 14662 10512 14714
rect 10512 14662 10542 14714
rect 10566 14662 10576 14714
rect 10576 14662 10622 14714
rect 10326 14660 10382 14662
rect 10406 14660 10462 14662
rect 10486 14660 10542 14662
rect 10566 14660 10622 14662
rect 9402 13268 9404 13288
rect 9404 13268 9456 13288
rect 9456 13268 9458 13288
rect 9402 13232 9458 13268
rect 10138 13524 10194 13560
rect 10138 13504 10140 13524
rect 10140 13504 10192 13524
rect 10192 13504 10194 13524
rect 10326 13626 10382 13628
rect 10406 13626 10462 13628
rect 10486 13626 10542 13628
rect 10566 13626 10622 13628
rect 10326 13574 10372 13626
rect 10372 13574 10382 13626
rect 10406 13574 10436 13626
rect 10436 13574 10448 13626
rect 10448 13574 10462 13626
rect 10486 13574 10500 13626
rect 10500 13574 10512 13626
rect 10512 13574 10542 13626
rect 10566 13574 10576 13626
rect 10576 13574 10622 13626
rect 10326 13572 10382 13574
rect 10406 13572 10462 13574
rect 10486 13572 10542 13574
rect 10566 13572 10622 13574
rect 10966 16496 11022 16552
rect 11058 15952 11114 16008
rect 9954 13232 10010 13288
rect 10230 13232 10286 13288
rect 11058 15000 11114 15056
rect 12200 17434 12256 17436
rect 12280 17434 12336 17436
rect 12360 17434 12416 17436
rect 12440 17434 12496 17436
rect 12200 17382 12246 17434
rect 12246 17382 12256 17434
rect 12280 17382 12310 17434
rect 12310 17382 12322 17434
rect 12322 17382 12336 17434
rect 12360 17382 12374 17434
rect 12374 17382 12386 17434
rect 12386 17382 12416 17434
rect 12440 17382 12450 17434
rect 12450 17382 12496 17434
rect 12200 17380 12256 17382
rect 12280 17380 12336 17382
rect 12360 17380 12416 17382
rect 12440 17380 12496 17382
rect 12200 16346 12256 16348
rect 12280 16346 12336 16348
rect 12360 16346 12416 16348
rect 12440 16346 12496 16348
rect 12200 16294 12246 16346
rect 12246 16294 12256 16346
rect 12280 16294 12310 16346
rect 12310 16294 12322 16346
rect 12322 16294 12336 16346
rect 12360 16294 12374 16346
rect 12374 16294 12386 16346
rect 12386 16294 12416 16346
rect 12440 16294 12450 16346
rect 12450 16294 12496 16346
rect 12200 16292 12256 16294
rect 12280 16292 12336 16294
rect 12360 16292 12416 16294
rect 12440 16292 12496 16294
rect 12530 15544 12586 15600
rect 12200 15258 12256 15260
rect 12280 15258 12336 15260
rect 12360 15258 12416 15260
rect 12440 15258 12496 15260
rect 12200 15206 12246 15258
rect 12246 15206 12256 15258
rect 12280 15206 12310 15258
rect 12310 15206 12322 15258
rect 12322 15206 12336 15258
rect 12360 15206 12374 15258
rect 12374 15206 12386 15258
rect 12386 15206 12416 15258
rect 12440 15206 12450 15258
rect 12450 15206 12496 15258
rect 12200 15204 12256 15206
rect 12280 15204 12336 15206
rect 12360 15204 12416 15206
rect 12440 15204 12496 15206
rect 9678 12144 9734 12200
rect 9126 11872 9182 11928
rect 8942 11736 8998 11792
rect 9218 11736 9274 11792
rect 9310 11600 9366 11656
rect 9034 11464 9090 11520
rect 9402 11192 9458 11248
rect 8574 11056 8630 11112
rect 8758 11056 8814 11112
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8498 10906
rect 8498 10854 8508 10906
rect 8532 10854 8562 10906
rect 8562 10854 8574 10906
rect 8574 10854 8588 10906
rect 8612 10854 8626 10906
rect 8626 10854 8638 10906
rect 8638 10854 8668 10906
rect 8692 10854 8702 10906
rect 8702 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 8390 10512 8446 10568
rect 8942 10920 8998 10976
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8498 9818
rect 8498 9766 8508 9818
rect 8532 9766 8562 9818
rect 8562 9766 8574 9818
rect 8574 9766 8588 9818
rect 8612 9766 8626 9818
rect 8626 9766 8638 9818
rect 8638 9766 8668 9818
rect 8692 9766 8702 9818
rect 8702 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 8850 9696 8906 9752
rect 9034 9716 9090 9752
rect 9034 9696 9036 9716
rect 9036 9696 9088 9716
rect 9088 9696 9090 9716
rect 9034 9560 9090 9616
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8498 8730
rect 8498 8678 8508 8730
rect 8532 8678 8562 8730
rect 8562 8678 8574 8730
rect 8574 8678 8588 8730
rect 8612 8678 8626 8730
rect 8626 8678 8638 8730
rect 8638 8678 8668 8730
rect 8692 8678 8702 8730
rect 8702 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8498 7642
rect 8498 7590 8508 7642
rect 8532 7590 8562 7642
rect 8562 7590 8574 7642
rect 8574 7590 8588 7642
rect 8612 7590 8626 7642
rect 8626 7590 8638 7642
rect 8638 7590 8668 7642
rect 8692 7590 8702 7642
rect 8702 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8298 7248 8354 7304
rect 8114 6024 8170 6080
rect 8298 6840 8354 6896
rect 8850 6840 8906 6896
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8498 6554
rect 8498 6502 8508 6554
rect 8532 6502 8562 6554
rect 8562 6502 8574 6554
rect 8574 6502 8588 6554
rect 8612 6502 8626 6554
rect 8626 6502 8638 6554
rect 8638 6502 8668 6554
rect 8692 6502 8702 6554
rect 8702 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 9034 8744 9090 8800
rect 8298 6160 8354 6216
rect 9126 6976 9182 7032
rect 8850 6160 8906 6216
rect 8022 4936 8078 4992
rect 8022 4392 8078 4448
rect 7930 2252 7932 2272
rect 7932 2252 7984 2272
rect 7984 2252 7986 2272
rect 7930 2216 7986 2252
rect 8206 4256 8262 4312
rect 8114 3984 8170 4040
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8498 5466
rect 8498 5414 8508 5466
rect 8532 5414 8562 5466
rect 8562 5414 8574 5466
rect 8574 5414 8588 5466
rect 8612 5414 8626 5466
rect 8626 5414 8638 5466
rect 8638 5414 8668 5466
rect 8692 5414 8702 5466
rect 8702 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 9586 11192 9642 11248
rect 9310 10104 9366 10160
rect 9402 9968 9458 10024
rect 9586 9696 9642 9752
rect 9862 12416 9918 12472
rect 9678 8744 9734 8800
rect 10326 12538 10382 12540
rect 10406 12538 10462 12540
rect 10486 12538 10542 12540
rect 10566 12538 10622 12540
rect 10326 12486 10372 12538
rect 10372 12486 10382 12538
rect 10406 12486 10436 12538
rect 10436 12486 10448 12538
rect 10448 12486 10462 12538
rect 10486 12486 10500 12538
rect 10500 12486 10512 12538
rect 10512 12486 10542 12538
rect 10566 12486 10576 12538
rect 10576 12486 10622 12538
rect 10326 12484 10382 12486
rect 10406 12484 10462 12486
rect 10486 12484 10542 12486
rect 10566 12484 10622 12486
rect 10046 12280 10102 12336
rect 9954 11328 10010 11384
rect 10230 11736 10286 11792
rect 10598 12008 10654 12064
rect 10138 11464 10194 11520
rect 10138 10548 10140 10568
rect 10140 10548 10192 10568
rect 10192 10548 10194 10568
rect 10138 10512 10194 10548
rect 9862 9560 9918 9616
rect 10138 10412 10140 10432
rect 10140 10412 10192 10432
rect 10192 10412 10194 10432
rect 10138 10376 10194 10412
rect 10138 10260 10194 10296
rect 10138 10240 10140 10260
rect 10140 10240 10192 10260
rect 10192 10240 10194 10260
rect 9862 8336 9918 8392
rect 10326 11450 10382 11452
rect 10406 11450 10462 11452
rect 10486 11450 10542 11452
rect 10566 11450 10622 11452
rect 10326 11398 10372 11450
rect 10372 11398 10382 11450
rect 10406 11398 10436 11450
rect 10436 11398 10448 11450
rect 10448 11398 10462 11450
rect 10486 11398 10500 11450
rect 10500 11398 10512 11450
rect 10512 11398 10542 11450
rect 10566 11398 10576 11450
rect 10576 11398 10622 11450
rect 10326 11396 10382 11398
rect 10406 11396 10462 11398
rect 10486 11396 10542 11398
rect 10566 11396 10622 11398
rect 10322 11212 10378 11248
rect 10322 11192 10324 11212
rect 10324 11192 10376 11212
rect 10376 11192 10378 11212
rect 10598 11192 10654 11248
rect 11058 12824 11114 12880
rect 10966 12280 11022 12336
rect 10326 10362 10382 10364
rect 10406 10362 10462 10364
rect 10486 10362 10542 10364
rect 10566 10362 10622 10364
rect 10326 10310 10372 10362
rect 10372 10310 10382 10362
rect 10406 10310 10436 10362
rect 10436 10310 10448 10362
rect 10448 10310 10462 10362
rect 10486 10310 10500 10362
rect 10500 10310 10512 10362
rect 10512 10310 10542 10362
rect 10566 10310 10576 10362
rect 10576 10310 10622 10362
rect 10326 10308 10382 10310
rect 10406 10308 10462 10310
rect 10486 10308 10542 10310
rect 10566 10308 10622 10310
rect 10782 10240 10838 10296
rect 10690 9968 10746 10024
rect 10598 9560 10654 9616
rect 10230 9424 10286 9480
rect 10690 9424 10746 9480
rect 10326 9274 10382 9276
rect 10406 9274 10462 9276
rect 10486 9274 10542 9276
rect 10566 9274 10622 9276
rect 10326 9222 10372 9274
rect 10372 9222 10382 9274
rect 10406 9222 10436 9274
rect 10436 9222 10448 9274
rect 10448 9222 10462 9274
rect 10486 9222 10500 9274
rect 10500 9222 10512 9274
rect 10512 9222 10542 9274
rect 10566 9222 10576 9274
rect 10576 9222 10622 9274
rect 10326 9220 10382 9222
rect 10406 9220 10462 9222
rect 10486 9220 10542 9222
rect 10566 9220 10622 9222
rect 10046 9016 10102 9072
rect 10046 8608 10102 8664
rect 10138 8336 10194 8392
rect 10046 8200 10102 8256
rect 9954 8064 10010 8120
rect 9494 6976 9550 7032
rect 9402 6160 9458 6216
rect 8482 4800 8538 4856
rect 8942 4392 8998 4448
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8498 4378
rect 8498 4326 8508 4378
rect 8532 4326 8562 4378
rect 8562 4326 8574 4378
rect 8574 4326 8588 4378
rect 8612 4326 8626 4378
rect 8626 4326 8638 4378
rect 8638 4326 8668 4378
rect 8692 4326 8702 4378
rect 8702 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8114 3032 8170 3088
rect 9218 5616 9274 5672
rect 9218 4664 9274 4720
rect 8758 3612 8760 3632
rect 8760 3612 8812 3632
rect 8812 3612 8814 3632
rect 8758 3576 8814 3612
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8498 3290
rect 8498 3238 8508 3290
rect 8532 3238 8562 3290
rect 8562 3238 8574 3290
rect 8574 3238 8588 3290
rect 8612 3238 8626 3290
rect 8626 3238 8638 3290
rect 8638 3238 8668 3290
rect 8692 3238 8702 3290
rect 8702 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 7654 1400 7710 1456
rect 8298 2624 8354 2680
rect 8390 2488 8446 2544
rect 8758 2916 8814 2952
rect 8758 2896 8760 2916
rect 8760 2896 8812 2916
rect 8812 2896 8814 2916
rect 8758 2644 8814 2680
rect 8758 2624 8760 2644
rect 8760 2624 8812 2644
rect 8812 2624 8814 2644
rect 9218 3032 9274 3088
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8498 2202
rect 8498 2150 8508 2202
rect 8532 2150 8562 2202
rect 8562 2150 8574 2202
rect 8574 2150 8588 2202
rect 8612 2150 8626 2202
rect 8626 2150 8638 2202
rect 8638 2150 8668 2202
rect 8692 2150 8702 2202
rect 8702 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 9126 2352 9182 2408
rect 9402 4256 9458 4312
rect 9402 3712 9458 3768
rect 9678 7928 9734 7984
rect 10326 8186 10382 8188
rect 10406 8186 10462 8188
rect 10486 8186 10542 8188
rect 10566 8186 10622 8188
rect 10326 8134 10372 8186
rect 10372 8134 10382 8186
rect 10406 8134 10436 8186
rect 10436 8134 10448 8186
rect 10448 8134 10462 8186
rect 10486 8134 10500 8186
rect 10500 8134 10512 8186
rect 10512 8134 10542 8186
rect 10566 8134 10576 8186
rect 10576 8134 10622 8186
rect 10326 8132 10382 8134
rect 10406 8132 10462 8134
rect 10486 8132 10542 8134
rect 10566 8132 10622 8134
rect 10782 8336 10838 8392
rect 10138 7112 10194 7168
rect 10046 6976 10102 7032
rect 10690 7656 10746 7712
rect 10326 7098 10382 7100
rect 10406 7098 10462 7100
rect 10486 7098 10542 7100
rect 10566 7098 10622 7100
rect 10326 7046 10372 7098
rect 10372 7046 10382 7098
rect 10406 7046 10436 7098
rect 10436 7046 10448 7098
rect 10448 7046 10462 7098
rect 10486 7046 10500 7098
rect 10500 7046 10512 7098
rect 10512 7046 10542 7098
rect 10566 7046 10576 7098
rect 10576 7046 10622 7098
rect 10326 7044 10382 7046
rect 10406 7044 10462 7046
rect 10486 7044 10542 7046
rect 10566 7044 10622 7046
rect 10782 6996 10838 7032
rect 10782 6976 10784 6996
rect 10784 6976 10836 6996
rect 10836 6976 10838 6996
rect 9954 6024 10010 6080
rect 9954 5480 10010 5536
rect 9862 4936 9918 4992
rect 9770 4800 9826 4856
rect 9586 4020 9588 4040
rect 9588 4020 9640 4040
rect 9640 4020 9642 4040
rect 9586 3984 9642 4020
rect 9678 3712 9734 3768
rect 9310 2488 9366 2544
rect 9954 4256 10010 4312
rect 9862 3612 9864 3632
rect 9864 3612 9916 3632
rect 9916 3612 9918 3632
rect 9862 3576 9918 3612
rect 10966 10376 11022 10432
rect 10966 9832 11022 9888
rect 10966 9152 11022 9208
rect 11242 12824 11298 12880
rect 11150 12144 11206 12200
rect 11242 10648 11298 10704
rect 11150 9868 11152 9888
rect 11152 9868 11204 9888
rect 11204 9868 11206 9888
rect 11150 9832 11206 9868
rect 11150 9560 11206 9616
rect 11242 9424 11298 9480
rect 11242 7792 11298 7848
rect 11150 7404 11206 7440
rect 11150 7384 11152 7404
rect 11152 7384 11204 7404
rect 11204 7384 11206 7404
rect 11058 7248 11114 7304
rect 11426 13096 11482 13152
rect 12200 14170 12256 14172
rect 12280 14170 12336 14172
rect 12360 14170 12416 14172
rect 12440 14170 12496 14172
rect 12200 14118 12246 14170
rect 12246 14118 12256 14170
rect 12280 14118 12310 14170
rect 12310 14118 12322 14170
rect 12322 14118 12336 14170
rect 12360 14118 12374 14170
rect 12374 14118 12386 14170
rect 12386 14118 12416 14170
rect 12440 14118 12450 14170
rect 12450 14118 12496 14170
rect 12200 14116 12256 14118
rect 12280 14116 12336 14118
rect 12360 14116 12416 14118
rect 12440 14116 12496 14118
rect 12070 13504 12126 13560
rect 12070 13368 12126 13424
rect 11886 12688 11942 12744
rect 11518 11736 11574 11792
rect 11518 11056 11574 11112
rect 11794 12044 11796 12064
rect 11796 12044 11848 12064
rect 11848 12044 11850 12064
rect 11794 12008 11850 12044
rect 11702 10784 11758 10840
rect 10138 5888 10194 5944
rect 10326 6010 10382 6012
rect 10406 6010 10462 6012
rect 10486 6010 10542 6012
rect 10566 6010 10622 6012
rect 10326 5958 10372 6010
rect 10372 5958 10382 6010
rect 10406 5958 10436 6010
rect 10436 5958 10448 6010
rect 10448 5958 10462 6010
rect 10486 5958 10500 6010
rect 10500 5958 10512 6010
rect 10512 5958 10542 6010
rect 10566 5958 10576 6010
rect 10576 5958 10622 6010
rect 10326 5956 10382 5958
rect 10406 5956 10462 5958
rect 10486 5956 10542 5958
rect 10566 5956 10622 5958
rect 10782 6060 10784 6080
rect 10784 6060 10836 6080
rect 10836 6060 10838 6080
rect 10782 6024 10838 6060
rect 10782 5888 10838 5944
rect 10690 5616 10746 5672
rect 10322 5244 10324 5264
rect 10324 5244 10376 5264
rect 10376 5244 10378 5264
rect 10322 5208 10378 5244
rect 10598 5480 10654 5536
rect 10414 5072 10470 5128
rect 10326 4922 10382 4924
rect 10406 4922 10462 4924
rect 10486 4922 10542 4924
rect 10566 4922 10622 4924
rect 10326 4870 10372 4922
rect 10372 4870 10382 4922
rect 10406 4870 10436 4922
rect 10436 4870 10448 4922
rect 10448 4870 10462 4922
rect 10486 4870 10500 4922
rect 10500 4870 10512 4922
rect 10512 4870 10542 4922
rect 10566 4870 10576 4922
rect 10576 4870 10622 4922
rect 10326 4868 10382 4870
rect 10406 4868 10462 4870
rect 10486 4868 10542 4870
rect 10566 4868 10622 4870
rect 11334 7112 11390 7168
rect 11242 6704 11298 6760
rect 11150 6432 11206 6488
rect 11058 6024 11114 6080
rect 11058 5888 11114 5944
rect 11242 5616 11298 5672
rect 11242 5344 11298 5400
rect 10966 4936 11022 4992
rect 10874 4800 10930 4856
rect 10230 4256 10286 4312
rect 11242 4528 11298 4584
rect 10322 3984 10378 4040
rect 10874 3984 10930 4040
rect 10326 3834 10382 3836
rect 10406 3834 10462 3836
rect 10486 3834 10542 3836
rect 10566 3834 10622 3836
rect 10326 3782 10372 3834
rect 10372 3782 10382 3834
rect 10406 3782 10436 3834
rect 10436 3782 10448 3834
rect 10448 3782 10462 3834
rect 10486 3782 10500 3834
rect 10500 3782 10512 3834
rect 10512 3782 10542 3834
rect 10566 3782 10576 3834
rect 10576 3782 10622 3834
rect 10326 3780 10382 3782
rect 10406 3780 10462 3782
rect 10486 3780 10542 3782
rect 10566 3780 10622 3782
rect 10230 3576 10286 3632
rect 10506 3440 10562 3496
rect 10414 3032 10470 3088
rect 10690 3032 10746 3088
rect 10138 2896 10194 2952
rect 10598 2932 10600 2952
rect 10600 2932 10652 2952
rect 10652 2932 10654 2952
rect 10598 2896 10654 2932
rect 10046 2508 10102 2544
rect 10046 2488 10048 2508
rect 10048 2488 10100 2508
rect 10100 2488 10102 2508
rect 9586 1400 9642 1456
rect 9218 1264 9274 1320
rect 6734 176 6790 232
rect 9126 720 9182 776
rect 10326 2746 10382 2748
rect 10406 2746 10462 2748
rect 10486 2746 10542 2748
rect 10566 2746 10622 2748
rect 10326 2694 10372 2746
rect 10372 2694 10382 2746
rect 10406 2694 10436 2746
rect 10436 2694 10448 2746
rect 10448 2694 10462 2746
rect 10486 2694 10500 2746
rect 10500 2694 10512 2746
rect 10512 2694 10542 2746
rect 10566 2694 10576 2746
rect 10576 2694 10622 2746
rect 10326 2692 10382 2694
rect 10406 2692 10462 2694
rect 10486 2692 10542 2694
rect 10566 2692 10622 2694
rect 10322 2488 10378 2544
rect 10782 2760 10838 2816
rect 10966 3168 11022 3224
rect 11058 2624 11114 2680
rect 11242 3168 11298 3224
rect 11610 9832 11666 9888
rect 11518 9288 11574 9344
rect 11518 8472 11574 8528
rect 11978 12436 12034 12472
rect 11978 12416 11980 12436
rect 11980 12416 12032 12436
rect 12032 12416 12034 12436
rect 11978 11636 11980 11656
rect 11980 11636 12032 11656
rect 12032 11636 12034 11656
rect 11978 11600 12034 11636
rect 11978 11348 12034 11384
rect 11978 11328 11980 11348
rect 11980 11328 12032 11348
rect 12032 11328 12034 11348
rect 11978 11192 12034 11248
rect 11886 9968 11942 10024
rect 12200 13082 12256 13084
rect 12280 13082 12336 13084
rect 12360 13082 12416 13084
rect 12440 13082 12496 13084
rect 12200 13030 12246 13082
rect 12246 13030 12256 13082
rect 12280 13030 12310 13082
rect 12310 13030 12322 13082
rect 12322 13030 12336 13082
rect 12360 13030 12374 13082
rect 12374 13030 12386 13082
rect 12386 13030 12416 13082
rect 12440 13030 12450 13082
rect 12450 13030 12496 13082
rect 12200 13028 12256 13030
rect 12280 13028 12336 13030
rect 12360 13028 12416 13030
rect 12440 13028 12496 13030
rect 12530 12824 12586 12880
rect 12714 13232 12770 13288
rect 12200 11994 12256 11996
rect 12280 11994 12336 11996
rect 12360 11994 12416 11996
rect 12440 11994 12496 11996
rect 12200 11942 12246 11994
rect 12246 11942 12256 11994
rect 12280 11942 12310 11994
rect 12310 11942 12322 11994
rect 12322 11942 12336 11994
rect 12360 11942 12374 11994
rect 12374 11942 12386 11994
rect 12386 11942 12416 11994
rect 12440 11942 12450 11994
rect 12450 11942 12496 11994
rect 12200 11940 12256 11942
rect 12280 11940 12336 11942
rect 12360 11940 12416 11942
rect 12440 11940 12496 11942
rect 12162 11600 12218 11656
rect 12622 12044 12624 12064
rect 12624 12044 12676 12064
rect 12676 12044 12678 12064
rect 12622 12008 12678 12044
rect 12622 11328 12678 11384
rect 12898 12416 12954 12472
rect 12898 12144 12954 12200
rect 12200 10906 12256 10908
rect 12280 10906 12336 10908
rect 12360 10906 12416 10908
rect 12440 10906 12496 10908
rect 12200 10854 12246 10906
rect 12246 10854 12256 10906
rect 12280 10854 12310 10906
rect 12310 10854 12322 10906
rect 12322 10854 12336 10906
rect 12360 10854 12374 10906
rect 12374 10854 12386 10906
rect 12386 10854 12416 10906
rect 12440 10854 12450 10906
rect 12450 10854 12496 10906
rect 12200 10852 12256 10854
rect 12280 10852 12336 10854
rect 12360 10852 12416 10854
rect 12440 10852 12496 10854
rect 12438 10668 12494 10704
rect 12438 10648 12440 10668
rect 12440 10648 12492 10668
rect 12492 10648 12494 10668
rect 12806 11328 12862 11384
rect 11978 9832 12034 9888
rect 12200 9818 12256 9820
rect 12280 9818 12336 9820
rect 12360 9818 12416 9820
rect 12440 9818 12496 9820
rect 12200 9766 12246 9818
rect 12246 9766 12256 9818
rect 12280 9766 12310 9818
rect 12310 9766 12322 9818
rect 12322 9766 12336 9818
rect 12360 9766 12374 9818
rect 12374 9766 12386 9818
rect 12386 9766 12416 9818
rect 12440 9766 12450 9818
rect 12450 9766 12496 9818
rect 12200 9764 12256 9766
rect 12280 9764 12336 9766
rect 12360 9764 12416 9766
rect 12440 9764 12496 9766
rect 11886 9288 11942 9344
rect 11794 8744 11850 8800
rect 11518 7792 11574 7848
rect 12438 9152 12494 9208
rect 11978 8336 12034 8392
rect 11886 8064 11942 8120
rect 11978 7112 12034 7168
rect 11518 6432 11574 6488
rect 11702 6432 11758 6488
rect 12200 8730 12256 8732
rect 12280 8730 12336 8732
rect 12360 8730 12416 8732
rect 12440 8730 12496 8732
rect 12200 8678 12246 8730
rect 12246 8678 12256 8730
rect 12280 8678 12310 8730
rect 12310 8678 12322 8730
rect 12322 8678 12336 8730
rect 12360 8678 12374 8730
rect 12374 8678 12386 8730
rect 12386 8678 12416 8730
rect 12440 8678 12450 8730
rect 12450 8678 12496 8730
rect 12200 8676 12256 8678
rect 12280 8676 12336 8678
rect 12360 8676 12416 8678
rect 12440 8676 12496 8678
rect 12162 8508 12164 8528
rect 12164 8508 12216 8528
rect 12216 8508 12218 8528
rect 12162 8472 12218 8508
rect 12530 8472 12586 8528
rect 12898 11056 12954 11112
rect 12898 10648 12954 10704
rect 12898 10512 12954 10568
rect 13358 11192 13414 11248
rect 13542 11348 13598 11384
rect 13542 11328 13544 11348
rect 13544 11328 13596 11348
rect 13596 11328 13598 11348
rect 13450 10784 13506 10840
rect 13450 9968 13506 10024
rect 13358 9832 13414 9888
rect 13266 9696 13322 9752
rect 13174 9560 13230 9616
rect 13082 9288 13138 9344
rect 12898 9052 12900 9072
rect 12900 9052 12952 9072
rect 12952 9052 12954 9072
rect 12898 9016 12954 9052
rect 12806 8744 12862 8800
rect 12806 8608 12862 8664
rect 12714 8336 12770 8392
rect 12530 8064 12586 8120
rect 12200 7642 12256 7644
rect 12280 7642 12336 7644
rect 12360 7642 12416 7644
rect 12440 7642 12496 7644
rect 12200 7590 12246 7642
rect 12246 7590 12256 7642
rect 12280 7590 12310 7642
rect 12310 7590 12322 7642
rect 12322 7590 12336 7642
rect 12360 7590 12374 7642
rect 12374 7590 12386 7642
rect 12386 7590 12416 7642
rect 12440 7590 12450 7642
rect 12450 7590 12496 7642
rect 12200 7588 12256 7590
rect 12280 7588 12336 7590
rect 12360 7588 12416 7590
rect 12440 7588 12496 7590
rect 13174 8880 13230 8936
rect 13450 9288 13506 9344
rect 13082 8608 13138 8664
rect 12714 7268 12770 7304
rect 12714 7248 12716 7268
rect 12716 7248 12768 7268
rect 12768 7248 12770 7268
rect 12438 7112 12494 7168
rect 12622 7112 12678 7168
rect 12530 6976 12586 7032
rect 11978 6432 12034 6488
rect 12200 6554 12256 6556
rect 12280 6554 12336 6556
rect 12360 6554 12416 6556
rect 12440 6554 12496 6556
rect 12200 6502 12246 6554
rect 12246 6502 12256 6554
rect 12280 6502 12310 6554
rect 12310 6502 12322 6554
rect 12322 6502 12336 6554
rect 12360 6502 12374 6554
rect 12374 6502 12386 6554
rect 12386 6502 12416 6554
rect 12440 6502 12450 6554
rect 12450 6502 12496 6554
rect 12200 6500 12256 6502
rect 12280 6500 12336 6502
rect 12360 6500 12416 6502
rect 12440 6500 12496 6502
rect 11426 4936 11482 4992
rect 11610 5344 11666 5400
rect 11610 4820 11666 4856
rect 11610 4800 11612 4820
rect 11612 4800 11664 4820
rect 11664 4800 11666 4820
rect 11794 5616 11850 5672
rect 12346 5616 12402 5672
rect 12990 7692 12992 7712
rect 12992 7692 13044 7712
rect 13044 7692 13046 7712
rect 12990 7656 13046 7692
rect 13174 8336 13230 8392
rect 13174 8200 13230 8256
rect 13082 7520 13138 7576
rect 13358 8336 13414 8392
rect 12806 6024 12862 6080
rect 12200 5466 12256 5468
rect 12280 5466 12336 5468
rect 12360 5466 12416 5468
rect 12440 5466 12496 5468
rect 12200 5414 12246 5466
rect 12246 5414 12256 5466
rect 12280 5414 12310 5466
rect 12310 5414 12322 5466
rect 12322 5414 12336 5466
rect 12360 5414 12374 5466
rect 12374 5414 12386 5466
rect 12386 5414 12416 5466
rect 12440 5414 12450 5466
rect 12450 5414 12496 5466
rect 12200 5412 12256 5414
rect 12280 5412 12336 5414
rect 12360 5412 12416 5414
rect 12440 5412 12496 5414
rect 11610 4140 11666 4176
rect 11610 4120 11612 4140
rect 11612 4120 11664 4140
rect 11664 4120 11666 4140
rect 11886 5208 11942 5264
rect 11978 4936 12034 4992
rect 11886 4256 11942 4312
rect 11242 2488 11298 2544
rect 9770 584 9826 640
rect 11150 1536 11206 1592
rect 11334 1944 11390 2000
rect 11518 2252 11520 2272
rect 11520 2252 11572 2272
rect 11572 2252 11574 2272
rect 11518 2216 11574 2252
rect 11518 2080 11574 2136
rect 11794 3304 11850 3360
rect 11794 3188 11850 3224
rect 11794 3168 11796 3188
rect 11796 3168 11848 3188
rect 11848 3168 11850 3188
rect 11702 3032 11758 3088
rect 11426 1536 11482 1592
rect 12898 5772 12954 5808
rect 12898 5752 12900 5772
rect 12900 5752 12952 5772
rect 12952 5752 12954 5772
rect 13818 11872 13874 11928
rect 14074 16890 14130 16892
rect 14154 16890 14210 16892
rect 14234 16890 14290 16892
rect 14314 16890 14370 16892
rect 14074 16838 14120 16890
rect 14120 16838 14130 16890
rect 14154 16838 14184 16890
rect 14184 16838 14196 16890
rect 14196 16838 14210 16890
rect 14234 16838 14248 16890
rect 14248 16838 14260 16890
rect 14260 16838 14290 16890
rect 14314 16838 14324 16890
rect 14324 16838 14370 16890
rect 14074 16836 14130 16838
rect 14154 16836 14210 16838
rect 14234 16836 14290 16838
rect 14314 16836 14370 16838
rect 14074 15802 14130 15804
rect 14154 15802 14210 15804
rect 14234 15802 14290 15804
rect 14314 15802 14370 15804
rect 14074 15750 14120 15802
rect 14120 15750 14130 15802
rect 14154 15750 14184 15802
rect 14184 15750 14196 15802
rect 14196 15750 14210 15802
rect 14234 15750 14248 15802
rect 14248 15750 14260 15802
rect 14260 15750 14290 15802
rect 14314 15750 14324 15802
rect 14324 15750 14370 15802
rect 14074 15748 14130 15750
rect 14154 15748 14210 15750
rect 14234 15748 14290 15750
rect 14314 15748 14370 15750
rect 14074 14714 14130 14716
rect 14154 14714 14210 14716
rect 14234 14714 14290 14716
rect 14314 14714 14370 14716
rect 14074 14662 14120 14714
rect 14120 14662 14130 14714
rect 14154 14662 14184 14714
rect 14184 14662 14196 14714
rect 14196 14662 14210 14714
rect 14234 14662 14248 14714
rect 14248 14662 14260 14714
rect 14260 14662 14290 14714
rect 14314 14662 14324 14714
rect 14324 14662 14370 14714
rect 14074 14660 14130 14662
rect 14154 14660 14210 14662
rect 14234 14660 14290 14662
rect 14314 14660 14370 14662
rect 14074 13626 14130 13628
rect 14154 13626 14210 13628
rect 14234 13626 14290 13628
rect 14314 13626 14370 13628
rect 14074 13574 14120 13626
rect 14120 13574 14130 13626
rect 14154 13574 14184 13626
rect 14184 13574 14196 13626
rect 14196 13574 14210 13626
rect 14234 13574 14248 13626
rect 14248 13574 14260 13626
rect 14260 13574 14290 13626
rect 14314 13574 14324 13626
rect 14324 13574 14370 13626
rect 14074 13572 14130 13574
rect 14154 13572 14210 13574
rect 14234 13572 14290 13574
rect 14314 13572 14370 13574
rect 14074 12538 14130 12540
rect 14154 12538 14210 12540
rect 14234 12538 14290 12540
rect 14314 12538 14370 12540
rect 14074 12486 14120 12538
rect 14120 12486 14130 12538
rect 14154 12486 14184 12538
rect 14184 12486 14196 12538
rect 14196 12486 14210 12538
rect 14234 12486 14248 12538
rect 14248 12486 14260 12538
rect 14260 12486 14290 12538
rect 14314 12486 14324 12538
rect 14324 12486 14370 12538
rect 14074 12484 14130 12486
rect 14154 12484 14210 12486
rect 14234 12484 14290 12486
rect 14314 12484 14370 12486
rect 13818 11736 13874 11792
rect 14462 12300 14518 12336
rect 14462 12280 14464 12300
rect 14464 12280 14516 12300
rect 14516 12280 14518 12300
rect 14278 12008 14334 12064
rect 14186 11600 14242 11656
rect 14074 11450 14130 11452
rect 14154 11450 14210 11452
rect 14234 11450 14290 11452
rect 14314 11450 14370 11452
rect 14074 11398 14120 11450
rect 14120 11398 14130 11450
rect 14154 11398 14184 11450
rect 14184 11398 14196 11450
rect 14196 11398 14210 11450
rect 14234 11398 14248 11450
rect 14248 11398 14260 11450
rect 14260 11398 14290 11450
rect 14314 11398 14324 11450
rect 14324 11398 14370 11450
rect 14074 11396 14130 11398
rect 14154 11396 14210 11398
rect 14234 11396 14290 11398
rect 14314 11396 14370 11398
rect 14278 11192 14334 11248
rect 14094 10920 14150 10976
rect 13818 9288 13874 9344
rect 14074 10362 14130 10364
rect 14154 10362 14210 10364
rect 14234 10362 14290 10364
rect 14314 10362 14370 10364
rect 14074 10310 14120 10362
rect 14120 10310 14130 10362
rect 14154 10310 14184 10362
rect 14184 10310 14196 10362
rect 14196 10310 14210 10362
rect 14234 10310 14248 10362
rect 14248 10310 14260 10362
rect 14260 10310 14290 10362
rect 14314 10310 14324 10362
rect 14324 10310 14370 10362
rect 14074 10308 14130 10310
rect 14154 10308 14210 10310
rect 14234 10308 14290 10310
rect 14314 10308 14370 10310
rect 14554 11892 14610 11928
rect 14554 11872 14556 11892
rect 14556 11872 14608 11892
rect 14608 11872 14610 11892
rect 15474 17720 15530 17776
rect 14922 14456 14978 14512
rect 14738 11328 14794 11384
rect 14554 10648 14610 10704
rect 14186 10140 14188 10160
rect 14188 10140 14240 10160
rect 14240 10140 14242 10160
rect 14186 10104 14242 10140
rect 14094 9868 14096 9888
rect 14096 9868 14148 9888
rect 14148 9868 14150 9888
rect 14094 9832 14150 9868
rect 14554 9696 14610 9752
rect 14922 10920 14978 10976
rect 14074 9274 14130 9276
rect 14154 9274 14210 9276
rect 14234 9274 14290 9276
rect 14314 9274 14370 9276
rect 14074 9222 14120 9274
rect 14120 9222 14130 9274
rect 14154 9222 14184 9274
rect 14184 9222 14196 9274
rect 14196 9222 14210 9274
rect 14234 9222 14248 9274
rect 14248 9222 14260 9274
rect 14260 9222 14290 9274
rect 14314 9222 14324 9274
rect 14324 9222 14370 9274
rect 14074 9220 14130 9222
rect 14154 9220 14210 9222
rect 14234 9220 14290 9222
rect 14314 9220 14370 9222
rect 14462 9152 14518 9208
rect 13542 8064 13598 8120
rect 13082 6432 13138 6488
rect 13358 6976 13414 7032
rect 13266 6024 13322 6080
rect 13818 8064 13874 8120
rect 14074 8186 14130 8188
rect 14154 8186 14210 8188
rect 14234 8186 14290 8188
rect 14314 8186 14370 8188
rect 14074 8134 14120 8186
rect 14120 8134 14130 8186
rect 14154 8134 14184 8186
rect 14184 8134 14196 8186
rect 14196 8134 14210 8186
rect 14234 8134 14248 8186
rect 14248 8134 14260 8186
rect 14260 8134 14290 8186
rect 14314 8134 14324 8186
rect 14324 8134 14370 8186
rect 14074 8132 14130 8134
rect 14154 8132 14210 8134
rect 14234 8132 14290 8134
rect 14314 8132 14370 8134
rect 13726 7540 13782 7576
rect 13726 7520 13728 7540
rect 13728 7520 13780 7540
rect 13780 7520 13782 7540
rect 14554 8064 14610 8120
rect 14830 8744 14886 8800
rect 13634 6840 13690 6896
rect 13450 6024 13506 6080
rect 13358 5752 13414 5808
rect 12254 5228 12310 5264
rect 12254 5208 12256 5228
rect 12256 5208 12308 5228
rect 12308 5208 12310 5228
rect 12438 5208 12494 5264
rect 12254 4664 12310 4720
rect 12622 4936 12678 4992
rect 12200 4378 12256 4380
rect 12280 4378 12336 4380
rect 12360 4378 12416 4380
rect 12440 4378 12496 4380
rect 12200 4326 12246 4378
rect 12246 4326 12256 4378
rect 12280 4326 12310 4378
rect 12310 4326 12322 4378
rect 12322 4326 12336 4378
rect 12360 4326 12374 4378
rect 12374 4326 12386 4378
rect 12386 4326 12416 4378
rect 12440 4326 12450 4378
rect 12450 4326 12496 4378
rect 12200 4324 12256 4326
rect 12280 4324 12336 4326
rect 12360 4324 12416 4326
rect 12440 4324 12496 4326
rect 12346 4120 12402 4176
rect 12438 4020 12440 4040
rect 12440 4020 12492 4040
rect 12492 4020 12494 4040
rect 12438 3984 12494 4020
rect 13082 5480 13138 5536
rect 12990 3984 13046 4040
rect 12200 3290 12256 3292
rect 12280 3290 12336 3292
rect 12360 3290 12416 3292
rect 12440 3290 12496 3292
rect 12200 3238 12246 3290
rect 12246 3238 12256 3290
rect 12280 3238 12310 3290
rect 12310 3238 12322 3290
rect 12322 3238 12336 3290
rect 12360 3238 12374 3290
rect 12374 3238 12386 3290
rect 12386 3238 12416 3290
rect 12440 3238 12450 3290
rect 12450 3238 12496 3290
rect 12200 3236 12256 3238
rect 12280 3236 12336 3238
rect 12360 3236 12416 3238
rect 12440 3236 12496 3238
rect 12162 3068 12164 3088
rect 12164 3068 12216 3088
rect 12216 3068 12218 3088
rect 12162 3032 12218 3068
rect 12438 3032 12494 3088
rect 12714 3440 12770 3496
rect 12200 2202 12256 2204
rect 12280 2202 12336 2204
rect 12360 2202 12416 2204
rect 12440 2202 12496 2204
rect 12200 2150 12246 2202
rect 12246 2150 12256 2202
rect 12280 2150 12310 2202
rect 12310 2150 12322 2202
rect 12322 2150 12336 2202
rect 12360 2150 12374 2202
rect 12374 2150 12386 2202
rect 12386 2150 12416 2202
rect 12440 2150 12450 2202
rect 12450 2150 12496 2202
rect 12200 2148 12256 2150
rect 12280 2148 12336 2150
rect 12360 2148 12416 2150
rect 12440 2148 12496 2150
rect 12070 1944 12126 2000
rect 11886 1400 11942 1456
rect 12898 1672 12954 1728
rect 13082 3440 13138 3496
rect 13266 4428 13268 4448
rect 13268 4428 13320 4448
rect 13320 4428 13322 4448
rect 13266 4392 13322 4428
rect 14462 7248 14518 7304
rect 14074 7098 14130 7100
rect 14154 7098 14210 7100
rect 14234 7098 14290 7100
rect 14314 7098 14370 7100
rect 14074 7046 14120 7098
rect 14120 7046 14130 7098
rect 14154 7046 14184 7098
rect 14184 7046 14196 7098
rect 14196 7046 14210 7098
rect 14234 7046 14248 7098
rect 14248 7046 14260 7098
rect 14260 7046 14290 7098
rect 14314 7046 14324 7098
rect 14324 7046 14370 7098
rect 14074 7044 14130 7046
rect 14154 7044 14210 7046
rect 14234 7044 14290 7046
rect 14314 7044 14370 7046
rect 14002 6452 14058 6488
rect 14002 6432 14004 6452
rect 14004 6432 14056 6452
rect 14056 6432 14058 6452
rect 13818 5888 13874 5944
rect 14646 6704 14702 6760
rect 14462 6432 14518 6488
rect 14462 6296 14518 6352
rect 14074 6010 14130 6012
rect 14154 6010 14210 6012
rect 14234 6010 14290 6012
rect 14314 6010 14370 6012
rect 14074 5958 14120 6010
rect 14120 5958 14130 6010
rect 14154 5958 14184 6010
rect 14184 5958 14196 6010
rect 14196 5958 14210 6010
rect 14234 5958 14248 6010
rect 14248 5958 14260 6010
rect 14260 5958 14290 6010
rect 14314 5958 14324 6010
rect 14324 5958 14370 6010
rect 14074 5956 14130 5958
rect 14154 5956 14210 5958
rect 14234 5956 14290 5958
rect 14314 5956 14370 5958
rect 13542 4800 13598 4856
rect 13634 4120 13690 4176
rect 14186 5616 14242 5672
rect 14278 5480 14334 5536
rect 14370 5344 14426 5400
rect 14094 5072 14150 5128
rect 14278 5092 14334 5128
rect 14278 5072 14280 5092
rect 14280 5072 14332 5092
rect 14332 5072 14334 5092
rect 14462 5072 14518 5128
rect 14074 4922 14130 4924
rect 14154 4922 14210 4924
rect 14234 4922 14290 4924
rect 14314 4922 14370 4924
rect 14074 4870 14120 4922
rect 14120 4870 14130 4922
rect 14154 4870 14184 4922
rect 14184 4870 14196 4922
rect 14196 4870 14210 4922
rect 14234 4870 14248 4922
rect 14248 4870 14260 4922
rect 14260 4870 14290 4922
rect 14314 4870 14324 4922
rect 14324 4870 14370 4922
rect 14074 4868 14130 4870
rect 14154 4868 14210 4870
rect 14234 4868 14290 4870
rect 14314 4868 14370 4870
rect 14370 4664 14426 4720
rect 14278 4140 14334 4176
rect 14278 4120 14280 4140
rect 14280 4120 14332 4140
rect 14332 4120 14334 4140
rect 13450 3576 13506 3632
rect 13174 1264 13230 1320
rect 13542 3476 13544 3496
rect 13544 3476 13596 3496
rect 13596 3476 13598 3496
rect 13542 3440 13598 3476
rect 13358 1128 13414 1184
rect 14094 3984 14150 4040
rect 13726 3848 13782 3904
rect 13542 40 13598 96
rect 14074 3834 14130 3836
rect 14154 3834 14210 3836
rect 14234 3834 14290 3836
rect 14314 3834 14370 3836
rect 14074 3782 14120 3834
rect 14120 3782 14130 3834
rect 14154 3782 14184 3834
rect 14184 3782 14196 3834
rect 14196 3782 14210 3834
rect 14234 3782 14248 3834
rect 14248 3782 14260 3834
rect 14260 3782 14290 3834
rect 14314 3782 14324 3834
rect 14324 3782 14370 3834
rect 14074 3780 14130 3782
rect 14154 3780 14210 3782
rect 14234 3780 14290 3782
rect 14314 3780 14370 3782
rect 13818 2760 13874 2816
rect 15106 11056 15162 11112
rect 15106 8608 15162 8664
rect 15290 13912 15346 13968
rect 15106 8064 15162 8120
rect 14922 6704 14978 6760
rect 14830 6296 14886 6352
rect 14830 6196 14832 6216
rect 14832 6196 14884 6216
rect 14884 6196 14886 6216
rect 14830 6160 14886 6196
rect 14922 5908 14978 5944
rect 14922 5888 14924 5908
rect 14924 5888 14976 5908
rect 14976 5888 14978 5908
rect 14830 5788 14832 5808
rect 14832 5788 14884 5808
rect 14884 5788 14886 5808
rect 14830 5752 14886 5788
rect 14922 5616 14978 5672
rect 14830 5480 14886 5536
rect 14074 2746 14130 2748
rect 14154 2746 14210 2748
rect 14234 2746 14290 2748
rect 14314 2746 14370 2748
rect 14074 2694 14120 2746
rect 14120 2694 14130 2746
rect 14154 2694 14184 2746
rect 14184 2694 14196 2746
rect 14196 2694 14210 2746
rect 14234 2694 14248 2746
rect 14248 2694 14260 2746
rect 14260 2694 14290 2746
rect 14314 2694 14324 2746
rect 14324 2694 14370 2746
rect 14074 2692 14130 2694
rect 14154 2692 14210 2694
rect 14234 2692 14290 2694
rect 14314 2692 14370 2694
rect 14094 992 14150 1048
rect 14186 856 14242 912
rect 14922 3984 14978 4040
rect 14830 3168 14886 3224
rect 14738 2488 14794 2544
rect 16118 17856 16174 17912
rect 15658 10512 15714 10568
rect 15198 7420 15200 7440
rect 15200 7420 15252 7440
rect 15252 7420 15254 7440
rect 15198 7384 15254 7420
rect 15106 5208 15162 5264
rect 15474 7948 15530 7984
rect 15474 7928 15476 7948
rect 15476 7928 15528 7948
rect 15528 7928 15530 7948
rect 15474 7656 15530 7712
rect 15566 6432 15622 6488
rect 15658 6024 15714 6080
rect 15474 5208 15530 5264
rect 15382 4664 15438 4720
rect 15290 4548 15346 4584
rect 15290 4528 15292 4548
rect 15292 4528 15344 4548
rect 15344 4528 15346 4548
rect 15934 7792 15990 7848
rect 16394 18264 16450 18320
rect 16210 11872 16266 11928
rect 16118 9152 16174 9208
rect 16210 8472 16266 8528
rect 16394 9424 16450 9480
rect 16486 9016 16542 9072
rect 16578 8336 16634 8392
rect 16302 4120 16358 4176
<< metal3 >>
rect 0 19410 800 19440
rect 4061 19410 4127 19413
rect 0 19408 4127 19410
rect 0 19352 4066 19408
rect 4122 19352 4127 19408
rect 0 19350 4127 19352
rect 0 19320 800 19350
rect 4061 19347 4127 19350
rect 0 18458 800 18488
rect 3969 18458 4035 18461
rect 0 18456 4035 18458
rect 0 18400 3974 18456
rect 4030 18400 4035 18456
rect 0 18398 4035 18400
rect 0 18368 800 18398
rect 3969 18395 4035 18398
rect 4102 18260 4108 18324
rect 4172 18322 4178 18324
rect 16389 18322 16455 18325
rect 4172 18320 16455 18322
rect 4172 18264 16394 18320
rect 16450 18264 16455 18320
rect 4172 18262 16455 18264
rect 4172 18260 4178 18262
rect 16389 18259 16455 18262
rect 5165 18050 5231 18053
rect 10726 18050 10732 18052
rect 5165 18048 10732 18050
rect 5165 17992 5170 18048
rect 5226 17992 10732 18048
rect 5165 17990 10732 17992
rect 5165 17987 5231 17990
rect 10726 17988 10732 17990
rect 10796 17988 10802 18052
rect 1393 17914 1459 17917
rect 9673 17914 9739 17917
rect 1393 17912 9739 17914
rect 1393 17856 1398 17912
rect 1454 17856 9678 17912
rect 9734 17856 9739 17912
rect 1393 17854 9739 17856
rect 1393 17851 1459 17854
rect 9673 17851 9739 17854
rect 9857 17914 9923 17917
rect 16113 17914 16179 17917
rect 9857 17912 16179 17914
rect 9857 17856 9862 17912
rect 9918 17856 16118 17912
rect 16174 17856 16179 17912
rect 9857 17854 16179 17856
rect 9857 17851 9923 17854
rect 16113 17851 16179 17854
rect 2589 17778 2655 17781
rect 7557 17778 7623 17781
rect 15469 17778 15535 17781
rect 2589 17776 2790 17778
rect 2589 17720 2594 17776
rect 2650 17720 2790 17776
rect 2589 17718 2790 17720
rect 2589 17715 2655 17718
rect 2730 17642 2790 17718
rect 7557 17776 15535 17778
rect 7557 17720 7562 17776
rect 7618 17720 15474 17776
rect 15530 17720 15535 17776
rect 7557 17718 15535 17720
rect 7557 17715 7623 17718
rect 15469 17715 15535 17718
rect 12566 17642 12572 17644
rect 2730 17582 12572 17642
rect 12566 17580 12572 17582
rect 12636 17580 12642 17644
rect 5349 17506 5415 17509
rect 7782 17506 7788 17508
rect 5349 17504 7788 17506
rect 5349 17448 5354 17504
rect 5410 17448 7788 17504
rect 5349 17446 7788 17448
rect 5349 17443 5415 17446
rect 7782 17444 7788 17446
rect 7852 17444 7858 17508
rect 4692 17440 5012 17441
rect 0 17280 800 17400
rect 4692 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5012 17440
rect 4692 17375 5012 17376
rect 8440 17440 8760 17441
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 17375 8760 17376
rect 12188 17440 12508 17441
rect 12188 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12508 17440
rect 12188 17375 12508 17376
rect 5257 17370 5323 17373
rect 5257 17368 7804 17370
rect 5257 17312 5262 17368
rect 5318 17312 7804 17368
rect 5257 17310 7804 17312
rect 5257 17307 5323 17310
rect 2630 17172 2636 17236
rect 2700 17234 2706 17236
rect 7557 17234 7623 17237
rect 2700 17232 7623 17234
rect 2700 17176 7562 17232
rect 7618 17176 7623 17232
rect 2700 17174 7623 17176
rect 7744 17234 7804 17310
rect 13302 17234 13308 17236
rect 7744 17174 13308 17234
rect 2700 17172 2706 17174
rect 7557 17171 7623 17174
rect 13302 17172 13308 17174
rect 13372 17172 13378 17236
rect 5349 17098 5415 17101
rect 13118 17098 13124 17100
rect 5349 17096 13124 17098
rect 5349 17040 5354 17096
rect 5410 17040 13124 17096
rect 5349 17038 13124 17040
rect 5349 17035 5415 17038
rect 13118 17036 13124 17038
rect 13188 17036 13194 17100
rect 2818 16896 3138 16897
rect 2818 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3138 16896
rect 2818 16831 3138 16832
rect 6566 16896 6886 16897
rect 6566 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6886 16896
rect 6566 16831 6886 16832
rect 10314 16896 10634 16897
rect 10314 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10634 16896
rect 10314 16831 10634 16832
rect 14062 16896 14382 16897
rect 14062 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14382 16896
rect 14062 16831 14382 16832
rect 4286 16628 4292 16692
rect 4356 16690 4362 16692
rect 9857 16690 9923 16693
rect 4356 16688 9923 16690
rect 4356 16632 9862 16688
rect 9918 16632 9923 16688
rect 4356 16630 9923 16632
rect 4356 16628 4362 16630
rect 9857 16627 9923 16630
rect 16400 16600 17200 16720
rect 2129 16554 2195 16557
rect 10961 16554 11027 16557
rect 2129 16552 11027 16554
rect 2129 16496 2134 16552
rect 2190 16496 10966 16552
rect 11022 16496 11027 16552
rect 2129 16494 11027 16496
rect 2129 16491 2195 16494
rect 10961 16491 11027 16494
rect 0 16418 800 16448
rect 3417 16418 3483 16421
rect 0 16416 3483 16418
rect 0 16360 3422 16416
rect 3478 16360 3483 16416
rect 0 16358 3483 16360
rect 0 16328 800 16358
rect 3417 16355 3483 16358
rect 4692 16352 5012 16353
rect 4692 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5012 16352
rect 4692 16287 5012 16288
rect 8440 16352 8760 16353
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 16287 8760 16288
rect 12188 16352 12508 16353
rect 12188 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12508 16352
rect 12188 16287 12508 16288
rect 3785 16146 3851 16149
rect 9070 16146 9076 16148
rect 3785 16144 9076 16146
rect 3785 16088 3790 16144
rect 3846 16088 9076 16144
rect 3785 16086 9076 16088
rect 3785 16083 3851 16086
rect 9070 16084 9076 16086
rect 9140 16084 9146 16148
rect 7005 16012 7071 16013
rect 7005 16010 7052 16012
rect 6924 16008 7052 16010
rect 7116 16010 7122 16012
rect 11053 16010 11119 16013
rect 7116 16008 11119 16010
rect 6924 15952 7010 16008
rect 7116 15952 11058 16008
rect 11114 15952 11119 16008
rect 6924 15950 7052 15952
rect 7005 15948 7052 15950
rect 7116 15950 11119 15952
rect 7116 15948 7122 15950
rect 7005 15947 7071 15948
rect 11053 15947 11119 15950
rect 565 15874 631 15877
rect 1158 15874 1164 15876
rect 565 15872 1164 15874
rect 565 15816 570 15872
rect 626 15816 1164 15872
rect 565 15814 1164 15816
rect 565 15811 631 15814
rect 1158 15812 1164 15814
rect 1228 15812 1234 15876
rect 2818 15808 3138 15809
rect 2818 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3138 15808
rect 2818 15743 3138 15744
rect 6566 15808 6886 15809
rect 6566 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6886 15808
rect 6566 15743 6886 15744
rect 10314 15808 10634 15809
rect 10314 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10634 15808
rect 10314 15743 10634 15744
rect 14062 15808 14382 15809
rect 14062 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14382 15808
rect 14062 15743 14382 15744
rect 197 15738 263 15741
rect 1342 15738 1348 15740
rect 197 15736 1348 15738
rect 197 15680 202 15736
rect 258 15680 1348 15736
rect 197 15678 1348 15680
rect 197 15675 263 15678
rect 1342 15676 1348 15678
rect 1412 15676 1418 15740
rect 4470 15676 4476 15740
rect 4540 15738 4546 15740
rect 6085 15738 6151 15741
rect 4540 15736 6151 15738
rect 4540 15680 6090 15736
rect 6146 15680 6151 15736
rect 4540 15678 6151 15680
rect 4540 15676 4546 15678
rect 6085 15675 6151 15678
rect 7741 15738 7807 15741
rect 9806 15738 9812 15740
rect 7741 15736 9812 15738
rect 7741 15680 7746 15736
rect 7802 15680 9812 15736
rect 7741 15678 9812 15680
rect 7741 15675 7807 15678
rect 9806 15676 9812 15678
rect 9876 15676 9882 15740
rect 1485 15602 1551 15605
rect 12525 15602 12591 15605
rect 1485 15600 12591 15602
rect 1485 15544 1490 15600
rect 1546 15544 12530 15600
rect 12586 15544 12591 15600
rect 1485 15542 12591 15544
rect 1485 15539 1551 15542
rect 12525 15539 12591 15542
rect 0 15466 800 15496
rect 2221 15466 2287 15469
rect 5349 15468 5415 15469
rect 0 15464 2287 15466
rect 0 15408 2226 15464
rect 2282 15408 2287 15464
rect 0 15406 2287 15408
rect 0 15376 800 15406
rect 2221 15403 2287 15406
rect 3558 15406 5274 15466
rect 3558 15197 3618 15406
rect 5214 15330 5274 15406
rect 5349 15464 5396 15468
rect 5460 15466 5466 15468
rect 5625 15466 5691 15469
rect 5460 15464 5691 15466
rect 5349 15408 5354 15464
rect 5460 15408 5630 15464
rect 5686 15408 5691 15464
rect 5349 15404 5396 15408
rect 5460 15406 5691 15408
rect 5460 15404 5466 15406
rect 5349 15403 5415 15404
rect 5625 15403 5691 15406
rect 5901 15466 5967 15469
rect 11462 15466 11468 15468
rect 5901 15464 11468 15466
rect 5901 15408 5906 15464
rect 5962 15408 11468 15464
rect 5901 15406 11468 15408
rect 5901 15403 5967 15406
rect 11462 15404 11468 15406
rect 11532 15404 11538 15468
rect 7833 15330 7899 15333
rect 5214 15328 7899 15330
rect 5214 15272 7838 15328
rect 7894 15272 7899 15328
rect 5214 15270 7899 15272
rect 7833 15267 7899 15270
rect 4692 15264 5012 15265
rect 4692 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5012 15264
rect 4692 15199 5012 15200
rect 8440 15264 8760 15265
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 15199 8760 15200
rect 12188 15264 12508 15265
rect 12188 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12508 15264
rect 12188 15199 12508 15200
rect 3509 15192 3618 15197
rect 3509 15136 3514 15192
rect 3570 15136 3618 15192
rect 3509 15134 3618 15136
rect 5625 15194 5691 15197
rect 7833 15194 7899 15197
rect 5625 15192 7899 15194
rect 5625 15136 5630 15192
rect 5686 15136 7838 15192
rect 7894 15136 7899 15192
rect 5625 15134 7899 15136
rect 3509 15131 3575 15134
rect 5625 15131 5691 15134
rect 7833 15131 7899 15134
rect 3693 15058 3759 15061
rect 7373 15058 7439 15061
rect 3693 15056 7439 15058
rect 3693 15000 3698 15056
rect 3754 15000 7378 15056
rect 7434 15000 7439 15056
rect 3693 14998 7439 15000
rect 3693 14995 3759 14998
rect 7373 14995 7439 14998
rect 7966 14996 7972 15060
rect 8036 15058 8042 15060
rect 9581 15058 9647 15061
rect 8036 15056 9647 15058
rect 8036 15000 9586 15056
rect 9642 15000 9647 15056
rect 8036 14998 9647 15000
rect 8036 14996 8042 14998
rect 9581 14995 9647 14998
rect 11053 15058 11119 15061
rect 13854 15058 13860 15060
rect 11053 15056 13860 15058
rect 11053 15000 11058 15056
rect 11114 15000 13860 15056
rect 11053 14998 13860 15000
rect 11053 14995 11119 14998
rect 13854 14996 13860 14998
rect 13924 14996 13930 15060
rect 3877 14922 3943 14925
rect 9397 14922 9463 14925
rect 3877 14920 9463 14922
rect 3877 14864 3882 14920
rect 3938 14864 9402 14920
rect 9458 14864 9463 14920
rect 3877 14862 9463 14864
rect 3877 14859 3943 14862
rect 9397 14859 9463 14862
rect 3601 14786 3667 14789
rect 5625 14786 5691 14789
rect 3601 14784 5691 14786
rect 3601 14728 3606 14784
rect 3662 14728 5630 14784
rect 5686 14728 5691 14784
rect 3601 14726 5691 14728
rect 3601 14723 3667 14726
rect 5625 14723 5691 14726
rect 5758 14724 5764 14788
rect 5828 14786 5834 14788
rect 6085 14786 6151 14789
rect 5828 14784 6151 14786
rect 5828 14728 6090 14784
rect 6146 14728 6151 14784
rect 5828 14726 6151 14728
rect 5828 14724 5834 14726
rect 6085 14723 6151 14726
rect 7741 14786 7807 14789
rect 9254 14786 9260 14788
rect 7741 14784 9260 14786
rect 7741 14728 7746 14784
rect 7802 14728 9260 14784
rect 7741 14726 9260 14728
rect 7741 14723 7807 14726
rect 9254 14724 9260 14726
rect 9324 14724 9330 14788
rect 2818 14720 3138 14721
rect 2818 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3138 14720
rect 2818 14655 3138 14656
rect 6566 14720 6886 14721
rect 6566 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6886 14720
rect 6566 14655 6886 14656
rect 10314 14720 10634 14721
rect 10314 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10634 14720
rect 10314 14655 10634 14656
rect 14062 14720 14382 14721
rect 14062 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14382 14720
rect 14062 14655 14382 14656
rect 974 14588 980 14652
rect 1044 14650 1050 14652
rect 1577 14650 1643 14653
rect 1044 14648 1643 14650
rect 1044 14592 1582 14648
rect 1638 14592 1643 14648
rect 1044 14590 1643 14592
rect 1044 14588 1050 14590
rect 1577 14587 1643 14590
rect 3325 14652 3391 14653
rect 3325 14648 3372 14652
rect 3436 14650 3442 14652
rect 5809 14650 5875 14653
rect 3436 14648 5875 14650
rect 3325 14592 3330 14648
rect 3436 14592 5814 14648
rect 5870 14592 5875 14648
rect 3325 14588 3372 14592
rect 3436 14590 5875 14592
rect 3436 14588 3442 14590
rect 3325 14587 3391 14588
rect 5809 14587 5875 14590
rect 7833 14650 7899 14653
rect 8017 14650 8083 14653
rect 9673 14650 9739 14653
rect 7833 14648 9739 14650
rect 7833 14592 7838 14648
rect 7894 14592 8022 14648
rect 8078 14592 9678 14648
rect 9734 14592 9739 14648
rect 7833 14590 9739 14592
rect 7833 14587 7899 14590
rect 8017 14587 8083 14590
rect 9673 14587 9739 14590
rect 1710 14452 1716 14516
rect 1780 14514 1786 14516
rect 1945 14514 2011 14517
rect 14917 14514 14983 14517
rect 1780 14512 2011 14514
rect 1780 14456 1950 14512
rect 2006 14456 2011 14512
rect 1780 14454 2011 14456
rect 1780 14452 1786 14454
rect 1945 14451 2011 14454
rect 2730 14512 14983 14514
rect 2730 14456 14922 14512
rect 14978 14456 14983 14512
rect 2730 14454 14983 14456
rect 0 14378 800 14408
rect 1669 14378 1735 14381
rect 0 14376 1735 14378
rect 0 14320 1674 14376
rect 1730 14320 1735 14376
rect 0 14318 1735 14320
rect 0 14288 800 14318
rect 1669 14315 1735 14318
rect 1526 14180 1532 14244
rect 1596 14242 1602 14244
rect 2730 14242 2790 14454
rect 14917 14451 14983 14454
rect 3049 14378 3115 14381
rect 4102 14378 4108 14380
rect 3049 14376 4108 14378
rect 3049 14320 3054 14376
rect 3110 14320 4108 14376
rect 3049 14318 4108 14320
rect 3049 14315 3115 14318
rect 4102 14316 4108 14318
rect 4172 14316 4178 14380
rect 5533 14378 5599 14381
rect 6729 14378 6795 14381
rect 4478 14318 5458 14378
rect 1596 14182 2790 14242
rect 3509 14242 3575 14245
rect 3877 14242 3943 14245
rect 3509 14240 3943 14242
rect 3509 14184 3514 14240
rect 3570 14184 3882 14240
rect 3938 14184 3943 14240
rect 3509 14182 3943 14184
rect 1596 14180 1602 14182
rect 3509 14179 3575 14182
rect 3877 14179 3943 14182
rect 4153 14242 4219 14245
rect 4478 14242 4538 14318
rect 4153 14240 4538 14242
rect 4153 14184 4158 14240
rect 4214 14184 4538 14240
rect 4153 14182 4538 14184
rect 5398 14242 5458 14318
rect 5533 14376 6795 14378
rect 5533 14320 5538 14376
rect 5594 14320 6734 14376
rect 6790 14320 6795 14376
rect 5533 14318 6795 14320
rect 5533 14315 5599 14318
rect 6729 14315 6795 14318
rect 6913 14378 6979 14381
rect 9397 14378 9463 14381
rect 6913 14376 9463 14378
rect 6913 14320 6918 14376
rect 6974 14320 9402 14376
rect 9458 14320 9463 14376
rect 6913 14318 9463 14320
rect 6913 14315 6979 14318
rect 9397 14315 9463 14318
rect 6637 14242 6703 14245
rect 5398 14240 6703 14242
rect 5398 14184 6642 14240
rect 6698 14184 6703 14240
rect 5398 14182 6703 14184
rect 4153 14179 4219 14182
rect 6637 14179 6703 14182
rect 6821 14242 6887 14245
rect 7598 14242 7604 14244
rect 6821 14240 7604 14242
rect 6821 14184 6826 14240
rect 6882 14184 7604 14240
rect 6821 14182 7604 14184
rect 6821 14179 6887 14182
rect 7598 14180 7604 14182
rect 7668 14180 7674 14244
rect 4692 14176 5012 14177
rect 4692 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5012 14176
rect 4692 14111 5012 14112
rect 8440 14176 8760 14177
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 14111 8760 14112
rect 12188 14176 12508 14177
rect 12188 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12508 14176
rect 12188 14111 12508 14112
rect 3325 14106 3391 14109
rect 3918 14106 3924 14108
rect 3325 14104 3924 14106
rect 3325 14048 3330 14104
rect 3386 14048 3924 14104
rect 3325 14046 3924 14048
rect 3325 14043 3391 14046
rect 3918 14044 3924 14046
rect 3988 14044 3994 14108
rect 5165 14106 5231 14109
rect 7741 14106 7807 14109
rect 5165 14104 7807 14106
rect 5165 14048 5170 14104
rect 5226 14048 7746 14104
rect 7802 14048 7807 14104
rect 5165 14046 7807 14048
rect 5165 14043 5231 14046
rect 7741 14043 7807 14046
rect 9254 14044 9260 14108
rect 9324 14106 9330 14108
rect 9397 14106 9463 14109
rect 9324 14104 9463 14106
rect 9324 14048 9402 14104
rect 9458 14048 9463 14104
rect 9324 14046 9463 14048
rect 9324 14044 9330 14046
rect 9397 14043 9463 14046
rect 1301 13970 1367 13973
rect 3509 13970 3575 13973
rect 1301 13968 3575 13970
rect 1301 13912 1306 13968
rect 1362 13912 3514 13968
rect 3570 13912 3575 13968
rect 1301 13910 3575 13912
rect 1301 13907 1367 13910
rect 3509 13907 3575 13910
rect 4153 13970 4219 13973
rect 5441 13970 5507 13973
rect 4153 13968 5507 13970
rect 4153 13912 4158 13968
rect 4214 13912 5446 13968
rect 5502 13912 5507 13968
rect 4153 13910 5507 13912
rect 4153 13907 4219 13910
rect 5441 13907 5507 13910
rect 7005 13970 7071 13973
rect 15285 13970 15351 13973
rect 7005 13968 15351 13970
rect 7005 13912 7010 13968
rect 7066 13912 15290 13968
rect 15346 13912 15351 13968
rect 7005 13910 15351 13912
rect 7005 13907 7071 13910
rect 15285 13907 15351 13910
rect 3785 13836 3851 13837
rect 3734 13834 3740 13836
rect 3694 13774 3740 13834
rect 3804 13832 3851 13836
rect 3846 13776 3851 13832
rect 3734 13772 3740 13774
rect 3804 13772 3851 13776
rect 4102 13772 4108 13836
rect 4172 13834 4178 13836
rect 5349 13834 5415 13837
rect 4172 13832 5415 13834
rect 4172 13776 5354 13832
rect 5410 13776 5415 13832
rect 4172 13774 5415 13776
rect 4172 13772 4178 13774
rect 3785 13771 3851 13772
rect 5349 13771 5415 13774
rect 5574 13772 5580 13836
rect 5644 13834 5650 13836
rect 5993 13834 6059 13837
rect 5644 13832 6059 13834
rect 5644 13776 5998 13832
rect 6054 13776 6059 13832
rect 5644 13774 6059 13776
rect 5644 13772 5650 13774
rect 5993 13771 6059 13774
rect 6177 13834 6243 13837
rect 9622 13834 9628 13836
rect 6177 13832 9628 13834
rect 6177 13776 6182 13832
rect 6238 13776 9628 13832
rect 6177 13774 9628 13776
rect 6177 13771 6243 13774
rect 9622 13772 9628 13774
rect 9692 13772 9698 13836
rect 9765 13834 9831 13837
rect 11094 13834 11100 13836
rect 9765 13832 11100 13834
rect 9765 13776 9770 13832
rect 9826 13776 11100 13832
rect 9765 13774 11100 13776
rect 9765 13771 9831 13774
rect 11094 13772 11100 13774
rect 11164 13772 11170 13836
rect 3785 13698 3851 13701
rect 5901 13698 5967 13701
rect 3785 13696 5967 13698
rect 3785 13640 3790 13696
rect 3846 13640 5906 13696
rect 5962 13640 5967 13696
rect 3785 13638 5967 13640
rect 3785 13635 3851 13638
rect 5901 13635 5967 13638
rect 7741 13698 7807 13701
rect 7741 13696 9690 13698
rect 7741 13640 7746 13696
rect 7802 13640 9690 13696
rect 7741 13638 9690 13640
rect 7741 13635 7807 13638
rect 2818 13632 3138 13633
rect 2818 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3138 13632
rect 2818 13567 3138 13568
rect 6566 13632 6886 13633
rect 6566 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6886 13632
rect 6566 13567 6886 13568
rect 4153 13562 4219 13565
rect 5625 13562 5691 13565
rect 4153 13560 5691 13562
rect 4153 13504 4158 13560
rect 4214 13504 5630 13560
rect 5686 13504 5691 13560
rect 4153 13502 5691 13504
rect 4153 13499 4219 13502
rect 5625 13499 5691 13502
rect 7097 13562 7163 13565
rect 9438 13562 9444 13564
rect 7097 13560 9444 13562
rect 7097 13504 7102 13560
rect 7158 13504 9444 13560
rect 7097 13502 9444 13504
rect 7097 13499 7163 13502
rect 9438 13500 9444 13502
rect 9508 13500 9514 13564
rect 9630 13562 9690 13638
rect 10314 13632 10634 13633
rect 10314 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10634 13632
rect 10314 13567 10634 13568
rect 14062 13632 14382 13633
rect 14062 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14382 13632
rect 14062 13567 14382 13568
rect 10133 13564 10199 13565
rect 10133 13562 10180 13564
rect 9630 13560 10180 13562
rect 9630 13504 10138 13560
rect 9630 13502 10180 13504
rect 10133 13500 10180 13502
rect 10244 13500 10250 13564
rect 12065 13562 12131 13565
rect 13670 13562 13676 13564
rect 12065 13560 13676 13562
rect 12065 13504 12070 13560
rect 12126 13504 13676 13560
rect 12065 13502 13676 13504
rect 10133 13499 10199 13500
rect 12065 13499 12131 13502
rect 13670 13500 13676 13502
rect 13740 13500 13746 13564
rect 0 13426 800 13456
rect 1577 13426 1643 13429
rect 0 13424 1643 13426
rect 0 13368 1582 13424
rect 1638 13368 1643 13424
rect 0 13366 1643 13368
rect 0 13336 800 13366
rect 1577 13363 1643 13366
rect 3325 13426 3391 13429
rect 4286 13426 4292 13428
rect 3325 13424 4292 13426
rect 3325 13368 3330 13424
rect 3386 13368 4292 13424
rect 3325 13366 4292 13368
rect 3325 13363 3391 13366
rect 4286 13364 4292 13366
rect 4356 13364 4362 13428
rect 5717 13426 5783 13429
rect 4478 13424 5783 13426
rect 4478 13368 5722 13424
rect 5778 13368 5783 13424
rect 4478 13366 5783 13368
rect 3601 13290 3667 13293
rect 4478 13290 4538 13366
rect 5717 13363 5783 13366
rect 6913 13426 6979 13429
rect 12065 13426 12131 13429
rect 6913 13424 12131 13426
rect 6913 13368 6918 13424
rect 6974 13368 12070 13424
rect 12126 13368 12131 13424
rect 6913 13366 12131 13368
rect 6913 13363 6979 13366
rect 12065 13363 12131 13366
rect 3601 13288 4538 13290
rect 3601 13232 3606 13288
rect 3662 13232 4538 13288
rect 3601 13230 4538 13232
rect 5441 13290 5507 13293
rect 9397 13290 9463 13293
rect 9949 13292 10015 13293
rect 9949 13290 9996 13292
rect 5441 13288 9322 13290
rect 5441 13232 5446 13288
rect 5502 13232 9322 13288
rect 5441 13230 9322 13232
rect 3601 13227 3667 13230
rect 5441 13227 5507 13230
rect 9262 13154 9322 13230
rect 9397 13288 9996 13290
rect 9397 13232 9402 13288
rect 9458 13232 9954 13288
rect 9397 13230 9996 13232
rect 9397 13227 9463 13230
rect 9949 13228 9996 13230
rect 10060 13228 10066 13292
rect 10225 13290 10291 13293
rect 12709 13290 12775 13293
rect 10225 13288 12775 13290
rect 10225 13232 10230 13288
rect 10286 13232 12714 13288
rect 12770 13232 12775 13288
rect 10225 13230 12775 13232
rect 9949 13227 10015 13228
rect 10225 13227 10291 13230
rect 12709 13227 12775 13230
rect 11421 13154 11487 13157
rect 9262 13152 11487 13154
rect 9262 13096 11426 13152
rect 11482 13096 11487 13152
rect 9262 13094 11487 13096
rect 11421 13091 11487 13094
rect 4692 13088 5012 13089
rect 4692 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5012 13088
rect 4692 13023 5012 13024
rect 8440 13088 8760 13089
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 13023 8760 13024
rect 12188 13088 12508 13089
rect 12188 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12508 13088
rect 12188 13023 12508 13024
rect 5390 12956 5396 13020
rect 5460 13018 5466 13020
rect 5901 13018 5967 13021
rect 5460 13016 5967 13018
rect 5460 12960 5906 13016
rect 5962 12960 5967 13016
rect 5460 12958 5967 12960
rect 5460 12956 5466 12958
rect 5901 12955 5967 12958
rect 7230 12956 7236 13020
rect 7300 13018 7306 13020
rect 8017 13018 8083 13021
rect 7300 13016 8083 13018
rect 7300 12960 8022 13016
rect 8078 12960 8083 13016
rect 7300 12958 8083 12960
rect 7300 12956 7306 12958
rect 8017 12955 8083 12958
rect 9438 12956 9444 13020
rect 9508 13018 9514 13020
rect 12014 13018 12020 13020
rect 9508 12958 12020 13018
rect 9508 12956 9514 12958
rect 12014 12956 12020 12958
rect 12084 12956 12090 13020
rect 2129 12882 2195 12885
rect 7189 12882 7255 12885
rect 11053 12882 11119 12885
rect 2129 12880 7114 12882
rect 2129 12824 2134 12880
rect 2190 12824 7114 12880
rect 2129 12822 7114 12824
rect 2129 12819 2195 12822
rect 2129 12746 2195 12749
rect 2773 12746 2839 12749
rect 2129 12744 2839 12746
rect 2129 12688 2134 12744
rect 2190 12688 2778 12744
rect 2834 12688 2839 12744
rect 2129 12686 2839 12688
rect 2129 12683 2195 12686
rect 2773 12683 2839 12686
rect 5390 12684 5396 12748
rect 5460 12746 5466 12748
rect 6361 12746 6427 12749
rect 5460 12744 6427 12746
rect 5460 12688 6366 12744
rect 6422 12688 6427 12744
rect 5460 12686 6427 12688
rect 5460 12684 5466 12686
rect 6361 12683 6427 12686
rect 1761 12610 1827 12613
rect 2446 12610 2452 12612
rect 1761 12608 2452 12610
rect 1761 12552 1766 12608
rect 1822 12552 2452 12608
rect 1761 12550 2452 12552
rect 1761 12547 1827 12550
rect 2446 12548 2452 12550
rect 2516 12548 2522 12612
rect 5206 12548 5212 12612
rect 5276 12610 5282 12612
rect 5533 12610 5599 12613
rect 5276 12608 5599 12610
rect 5276 12552 5538 12608
rect 5594 12552 5599 12608
rect 5276 12550 5599 12552
rect 7054 12610 7114 12822
rect 7189 12880 11119 12882
rect 7189 12824 7194 12880
rect 7250 12824 11058 12880
rect 11114 12824 11119 12880
rect 7189 12822 11119 12824
rect 7189 12819 7255 12822
rect 11053 12819 11119 12822
rect 11237 12884 11303 12885
rect 11237 12880 11284 12884
rect 11348 12882 11354 12884
rect 12525 12882 12591 12885
rect 12934 12882 12940 12884
rect 11237 12824 11242 12880
rect 11237 12820 11284 12824
rect 11348 12822 11394 12882
rect 12525 12880 12940 12882
rect 12525 12824 12530 12880
rect 12586 12824 12940 12880
rect 12525 12822 12940 12824
rect 11348 12820 11354 12822
rect 11237 12819 11303 12820
rect 12525 12819 12591 12822
rect 12934 12820 12940 12822
rect 13004 12820 13010 12884
rect 7189 12746 7255 12749
rect 11881 12746 11947 12749
rect 7189 12744 11947 12746
rect 7189 12688 7194 12744
rect 7250 12688 11886 12744
rect 11942 12688 11947 12744
rect 7189 12686 11947 12688
rect 7189 12683 7255 12686
rect 11881 12683 11947 12686
rect 8150 12610 8156 12612
rect 7054 12550 8156 12610
rect 5276 12548 5282 12550
rect 5533 12547 5599 12550
rect 8150 12548 8156 12550
rect 8220 12610 8226 12612
rect 8220 12550 10242 12610
rect 8220 12548 8226 12550
rect 2818 12544 3138 12545
rect 0 12474 800 12504
rect 2818 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3138 12544
rect 2818 12479 3138 12480
rect 6566 12544 6886 12545
rect 6566 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6886 12544
rect 6566 12479 6886 12480
rect 2221 12474 2287 12477
rect 0 12472 2287 12474
rect 0 12416 2226 12472
rect 2282 12416 2287 12472
rect 0 12414 2287 12416
rect 0 12384 800 12414
rect 2221 12411 2287 12414
rect 3550 12412 3556 12476
rect 3620 12474 3626 12476
rect 3693 12474 3759 12477
rect 5809 12474 5875 12477
rect 3620 12472 3759 12474
rect 3620 12416 3698 12472
rect 3754 12416 3759 12472
rect 3620 12414 3759 12416
rect 3620 12412 3626 12414
rect 3693 12411 3759 12414
rect 4110 12472 5875 12474
rect 4110 12416 5814 12472
rect 5870 12416 5875 12472
rect 4110 12414 5875 12416
rect 3693 12338 3759 12341
rect 4110 12338 4170 12414
rect 5809 12411 5875 12414
rect 8201 12474 8267 12477
rect 9857 12474 9923 12477
rect 8201 12472 9923 12474
rect 8201 12416 8206 12472
rect 8262 12416 9862 12472
rect 9918 12416 9923 12472
rect 8201 12414 9923 12416
rect 8201 12411 8267 12414
rect 9857 12411 9923 12414
rect 10182 12372 10242 12550
rect 10314 12544 10634 12545
rect 10314 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10634 12544
rect 10314 12479 10634 12480
rect 14062 12544 14382 12545
rect 14062 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14382 12544
rect 14062 12479 14382 12480
rect 10726 12412 10732 12476
rect 10796 12474 10802 12476
rect 11973 12474 12039 12477
rect 10796 12472 12039 12474
rect 10796 12416 11978 12472
rect 12034 12416 12039 12472
rect 10796 12414 12039 12416
rect 10796 12412 10802 12414
rect 11973 12411 12039 12414
rect 12893 12474 12959 12477
rect 13486 12474 13492 12476
rect 12893 12472 13492 12474
rect 12893 12416 12898 12472
rect 12954 12416 13492 12472
rect 12893 12414 13492 12416
rect 12893 12411 12959 12414
rect 13486 12412 13492 12414
rect 13556 12412 13562 12476
rect 3693 12336 4170 12338
rect 3693 12280 3698 12336
rect 3754 12280 4170 12336
rect 3693 12278 4170 12280
rect 3693 12275 3759 12278
rect 5206 12276 5212 12340
rect 5276 12338 5282 12340
rect 5533 12338 5599 12341
rect 5276 12336 5599 12338
rect 5276 12280 5538 12336
rect 5594 12280 5599 12336
rect 5276 12278 5599 12280
rect 5276 12276 5282 12278
rect 5533 12275 5599 12278
rect 5993 12338 6059 12341
rect 5993 12336 7298 12338
rect 5993 12280 5998 12336
rect 6054 12280 7298 12336
rect 5993 12278 7298 12280
rect 5993 12275 6059 12278
rect 2221 12202 2287 12205
rect 2773 12202 2839 12205
rect 2221 12200 2839 12202
rect 2221 12144 2226 12200
rect 2282 12144 2778 12200
rect 2834 12144 2839 12200
rect 2221 12142 2839 12144
rect 2221 12139 2287 12142
rect 2773 12139 2839 12142
rect 4981 12202 5047 12205
rect 7097 12202 7163 12205
rect 4981 12200 7163 12202
rect 4981 12144 4986 12200
rect 5042 12144 7102 12200
rect 7158 12144 7163 12200
rect 4981 12142 7163 12144
rect 7238 12202 7298 12278
rect 7782 12276 7788 12340
rect 7852 12338 7858 12340
rect 8017 12338 8083 12341
rect 7852 12336 8083 12338
rect 7852 12280 8022 12336
rect 8078 12280 8083 12336
rect 7852 12278 8083 12280
rect 7852 12276 7858 12278
rect 8017 12275 8083 12278
rect 8753 12338 8819 12341
rect 9029 12340 9095 12341
rect 8886 12338 8892 12340
rect 8753 12336 8892 12338
rect 8753 12280 8758 12336
rect 8814 12280 8892 12336
rect 8753 12278 8892 12280
rect 8753 12275 8819 12278
rect 8886 12276 8892 12278
rect 8956 12276 8962 12340
rect 9029 12336 9076 12340
rect 9140 12338 9146 12340
rect 9029 12280 9034 12336
rect 9029 12276 9076 12280
rect 9140 12278 9186 12338
rect 9140 12276 9146 12278
rect 9254 12276 9260 12340
rect 9324 12338 9330 12340
rect 10041 12338 10107 12341
rect 9324 12336 10107 12338
rect 9324 12280 10046 12336
rect 10102 12280 10107 12336
rect 10182 12338 10288 12372
rect 10961 12338 11027 12341
rect 10182 12336 11027 12338
rect 10182 12312 10966 12336
rect 9324 12278 10107 12280
rect 10228 12280 10966 12312
rect 11022 12280 11027 12336
rect 10228 12278 11027 12280
rect 9324 12276 9330 12278
rect 9029 12275 9095 12276
rect 10041 12275 10107 12278
rect 10961 12275 11027 12278
rect 13854 12276 13860 12340
rect 13924 12338 13930 12340
rect 14457 12338 14523 12341
rect 13924 12336 14523 12338
rect 13924 12280 14462 12336
rect 14518 12280 14523 12336
rect 13924 12278 14523 12280
rect 13924 12276 13930 12278
rect 14457 12275 14523 12278
rect 9673 12202 9739 12205
rect 11145 12202 11211 12205
rect 7238 12142 9460 12202
rect 4981 12139 5047 12142
rect 7097 12139 7163 12142
rect 790 12004 796 12068
rect 860 12066 866 12068
rect 1158 12066 1164 12068
rect 860 12006 1164 12066
rect 860 12004 866 12006
rect 1158 12004 1164 12006
rect 1228 12004 1234 12068
rect 5073 12066 5139 12069
rect 5349 12066 5415 12069
rect 5717 12068 5783 12069
rect 5717 12066 5764 12068
rect 5073 12064 5415 12066
rect 5073 12008 5078 12064
rect 5134 12008 5354 12064
rect 5410 12008 5415 12064
rect 5073 12006 5415 12008
rect 5672 12064 5764 12066
rect 5672 12008 5722 12064
rect 5672 12006 5764 12008
rect 5073 12003 5139 12006
rect 5349 12003 5415 12006
rect 5717 12004 5764 12006
rect 5828 12004 5834 12068
rect 6361 12066 6427 12069
rect 6821 12066 6887 12069
rect 6361 12064 6887 12066
rect 6361 12008 6366 12064
rect 6422 12008 6826 12064
rect 6882 12008 6887 12064
rect 6361 12006 6887 12008
rect 5717 12003 5783 12004
rect 6361 12003 6427 12006
rect 6821 12003 6887 12006
rect 4692 12000 5012 12001
rect 4692 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5012 12000
rect 4692 11935 5012 11936
rect 8440 12000 8760 12001
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 11935 8760 11936
rect 1158 11868 1164 11932
rect 1228 11930 1234 11932
rect 1577 11930 1643 11933
rect 2681 11932 2747 11933
rect 2630 11930 2636 11932
rect 1228 11928 1643 11930
rect 1228 11872 1582 11928
rect 1638 11872 1643 11928
rect 1228 11870 1643 11872
rect 2590 11870 2636 11930
rect 2700 11928 2747 11932
rect 2742 11872 2747 11928
rect 1228 11868 1234 11870
rect 1577 11867 1643 11870
rect 2630 11868 2636 11870
rect 2700 11868 2747 11872
rect 2681 11867 2747 11868
rect 5257 11930 5323 11933
rect 7414 11930 7420 11932
rect 5257 11928 7420 11930
rect 5257 11872 5262 11928
rect 5318 11872 7420 11928
rect 5257 11870 7420 11872
rect 5257 11867 5323 11870
rect 7414 11868 7420 11870
rect 7484 11868 7490 11932
rect 9121 11930 9187 11933
rect 9254 11930 9260 11932
rect 9121 11928 9260 11930
rect 9121 11872 9126 11928
rect 9182 11872 9260 11928
rect 9121 11870 9260 11872
rect 9121 11867 9187 11870
rect 9254 11868 9260 11870
rect 9324 11868 9330 11932
rect 9400 11930 9460 12142
rect 9673 12200 11211 12202
rect 9673 12144 9678 12200
rect 9734 12144 11150 12200
rect 11206 12144 11211 12200
rect 9673 12142 11211 12144
rect 9673 12139 9739 12142
rect 11145 12139 11211 12142
rect 11646 12140 11652 12204
rect 11716 12202 11722 12204
rect 12893 12202 12959 12205
rect 11716 12200 12959 12202
rect 11716 12144 12898 12200
rect 12954 12144 12959 12200
rect 11716 12142 12959 12144
rect 11716 12140 11722 12142
rect 12893 12139 12959 12142
rect 9622 12004 9628 12068
rect 9692 12066 9698 12068
rect 10593 12066 10659 12069
rect 9692 12064 10659 12066
rect 9692 12008 10598 12064
rect 10654 12008 10659 12064
rect 9692 12006 10659 12008
rect 9692 12004 9698 12006
rect 10593 12003 10659 12006
rect 11278 12004 11284 12068
rect 11348 12066 11354 12068
rect 11789 12066 11855 12069
rect 11348 12064 11855 12066
rect 11348 12008 11794 12064
rect 11850 12008 11855 12064
rect 11348 12006 11855 12008
rect 11348 12004 11354 12006
rect 11789 12003 11855 12006
rect 12617 12066 12683 12069
rect 14273 12066 14339 12069
rect 12617 12064 14339 12066
rect 12617 12008 12622 12064
rect 12678 12008 14278 12064
rect 14334 12008 14339 12064
rect 12617 12006 14339 12008
rect 12617 12003 12683 12006
rect 14273 12003 14339 12006
rect 12188 12000 12508 12001
rect 12188 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12508 12000
rect 12188 11935 12508 11936
rect 13813 11932 13879 11933
rect 9400 11870 10932 11930
rect 1301 11794 1367 11797
rect 7189 11794 7255 11797
rect 1301 11792 7255 11794
rect 1301 11736 1306 11792
rect 1362 11736 7194 11792
rect 7250 11736 7255 11792
rect 1301 11734 7255 11736
rect 1301 11731 1367 11734
rect 7189 11731 7255 11734
rect 7782 11732 7788 11796
rect 7852 11794 7858 11796
rect 8109 11794 8175 11797
rect 7852 11792 8175 11794
rect 7852 11736 8114 11792
rect 8170 11736 8175 11792
rect 7852 11734 8175 11736
rect 7852 11732 7858 11734
rect 8109 11731 8175 11734
rect 8569 11794 8635 11797
rect 8937 11794 9003 11797
rect 8569 11792 9003 11794
rect 8569 11736 8574 11792
rect 8630 11736 8942 11792
rect 8998 11736 9003 11792
rect 8569 11734 9003 11736
rect 8569 11731 8635 11734
rect 8937 11731 9003 11734
rect 9213 11796 9279 11797
rect 9213 11792 9260 11796
rect 9324 11794 9330 11796
rect 9213 11736 9218 11792
rect 9213 11732 9260 11736
rect 9324 11734 9370 11794
rect 9324 11732 9330 11734
rect 9806 11732 9812 11796
rect 9876 11794 9882 11796
rect 10225 11794 10291 11797
rect 9876 11792 10291 11794
rect 9876 11736 10230 11792
rect 10286 11736 10291 11792
rect 9876 11734 10291 11736
rect 9876 11732 9882 11734
rect 9213 11731 9279 11732
rect 10225 11731 10291 11734
rect 3550 11596 3556 11660
rect 3620 11658 3626 11660
rect 5257 11658 5323 11661
rect 3620 11656 5323 11658
rect 3620 11600 5262 11656
rect 5318 11600 5323 11656
rect 3620 11598 5323 11600
rect 3620 11596 3626 11598
rect 5257 11595 5323 11598
rect 5441 11658 5507 11661
rect 9305 11658 9371 11661
rect 5441 11656 9371 11658
rect 5441 11600 5446 11656
rect 5502 11600 9310 11656
rect 9366 11600 9371 11656
rect 5441 11598 9371 11600
rect 5441 11595 5507 11598
rect 9305 11595 9371 11598
rect 9446 11598 10794 11658
rect 4061 11522 4127 11525
rect 6085 11522 6151 11525
rect 4061 11520 6151 11522
rect 4061 11464 4066 11520
rect 4122 11464 6090 11520
rect 6146 11464 6151 11520
rect 4061 11462 6151 11464
rect 4061 11459 4127 11462
rect 6085 11459 6151 11462
rect 7598 11460 7604 11524
rect 7668 11522 7674 11524
rect 9029 11522 9095 11525
rect 7668 11520 9095 11522
rect 7668 11464 9034 11520
rect 9090 11464 9095 11520
rect 7668 11462 9095 11464
rect 7668 11460 7674 11462
rect 9029 11459 9095 11462
rect 2818 11456 3138 11457
rect 0 11386 800 11416
rect 2818 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3138 11456
rect 2818 11391 3138 11392
rect 6566 11456 6886 11457
rect 6566 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6886 11456
rect 6566 11391 6886 11392
rect 1669 11386 1735 11389
rect 0 11384 1735 11386
rect 0 11328 1674 11384
rect 1730 11328 1735 11384
rect 0 11326 1735 11328
rect 0 11296 800 11326
rect 1669 11323 1735 11326
rect 3325 11386 3391 11389
rect 3325 11384 3572 11386
rect 3325 11328 3330 11384
rect 3386 11328 3572 11384
rect 3325 11326 3572 11328
rect 3325 11323 3391 11326
rect 3512 11253 3572 11326
rect 4470 11324 4476 11388
rect 4540 11386 4546 11388
rect 4613 11386 4679 11389
rect 4540 11384 4679 11386
rect 4540 11328 4618 11384
rect 4674 11328 4679 11384
rect 4540 11326 4679 11328
rect 4540 11324 4546 11326
rect 4613 11323 4679 11326
rect 5809 11386 5875 11389
rect 6310 11386 6316 11388
rect 5809 11384 6316 11386
rect 5809 11328 5814 11384
rect 5870 11328 6316 11384
rect 5809 11326 6316 11328
rect 5809 11323 5875 11326
rect 6310 11324 6316 11326
rect 6380 11324 6386 11388
rect 7741 11386 7807 11389
rect 8109 11386 8175 11389
rect 9446 11386 9506 11598
rect 9622 11460 9628 11524
rect 9692 11522 9698 11524
rect 10133 11522 10199 11525
rect 9692 11520 10199 11522
rect 9692 11464 10138 11520
rect 10194 11464 10199 11520
rect 9692 11462 10199 11464
rect 9692 11460 9698 11462
rect 10133 11459 10199 11462
rect 10314 11456 10634 11457
rect 10314 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10634 11456
rect 10314 11391 10634 11392
rect 7741 11384 9506 11386
rect 7741 11328 7746 11384
rect 7802 11328 8114 11384
rect 8170 11328 9506 11384
rect 7741 11326 9506 11328
rect 9949 11388 10015 11389
rect 9949 11384 9996 11388
rect 10060 11386 10066 11388
rect 9949 11328 9954 11384
rect 7741 11323 7807 11326
rect 8109 11323 8175 11326
rect 9949 11324 9996 11328
rect 10060 11326 10106 11386
rect 10060 11324 10066 11326
rect 9949 11323 10015 11324
rect 3509 11248 3575 11253
rect 3509 11192 3514 11248
rect 3570 11192 3575 11248
rect 3509 11187 3575 11192
rect 4797 11250 4863 11253
rect 7966 11250 7972 11252
rect 4797 11248 7972 11250
rect 4797 11192 4802 11248
rect 4858 11192 7972 11248
rect 4797 11190 7972 11192
rect 4797 11187 4863 11190
rect 7966 11188 7972 11190
rect 8036 11188 8042 11252
rect 9397 11250 9463 11253
rect 9581 11250 9647 11253
rect 9397 11248 9647 11250
rect 9397 11192 9402 11248
rect 9458 11192 9586 11248
rect 9642 11192 9647 11248
rect 9397 11190 9647 11192
rect 9397 11187 9463 11190
rect 9581 11187 9647 11190
rect 9990 11188 9996 11252
rect 10060 11250 10066 11252
rect 10317 11250 10383 11253
rect 10060 11248 10383 11250
rect 10060 11192 10322 11248
rect 10378 11192 10383 11248
rect 10060 11190 10383 11192
rect 10060 11188 10066 11190
rect 10317 11187 10383 11190
rect 10593 11250 10659 11253
rect 10734 11250 10794 11598
rect 10872 11522 10932 11870
rect 13813 11928 13860 11932
rect 13924 11930 13930 11932
rect 14549 11930 14615 11933
rect 16205 11930 16271 11933
rect 13813 11872 13818 11928
rect 13813 11868 13860 11872
rect 13924 11870 13970 11930
rect 14549 11928 16271 11930
rect 14549 11872 14554 11928
rect 14610 11872 16210 11928
rect 16266 11872 16271 11928
rect 14549 11870 16271 11872
rect 13924 11868 13930 11870
rect 13813 11867 13879 11868
rect 14549 11867 14615 11870
rect 16205 11867 16271 11870
rect 11513 11794 11579 11797
rect 13813 11794 13879 11797
rect 11513 11792 13879 11794
rect 11513 11736 11518 11792
rect 11574 11736 13818 11792
rect 13874 11736 13879 11792
rect 11513 11734 13879 11736
rect 11513 11731 11579 11734
rect 13813 11731 13879 11734
rect 11973 11658 12039 11661
rect 12157 11658 12223 11661
rect 11973 11656 12223 11658
rect 11973 11600 11978 11656
rect 12034 11600 12162 11656
rect 12218 11600 12223 11656
rect 11973 11598 12223 11600
rect 11973 11595 12039 11598
rect 12157 11595 12223 11598
rect 12750 11596 12756 11660
rect 12820 11658 12826 11660
rect 14181 11658 14247 11661
rect 12820 11656 14247 11658
rect 12820 11600 14186 11656
rect 14242 11600 14247 11656
rect 12820 11598 14247 11600
rect 12820 11596 12826 11598
rect 14181 11595 14247 11598
rect 10872 11462 13876 11522
rect 11830 11324 11836 11388
rect 11900 11386 11906 11388
rect 11973 11386 12039 11389
rect 11900 11384 12039 11386
rect 11900 11328 11978 11384
rect 12034 11328 12039 11384
rect 11900 11326 12039 11328
rect 11900 11324 11906 11326
rect 11973 11323 12039 11326
rect 12617 11386 12683 11389
rect 12801 11386 12867 11389
rect 13537 11388 13603 11389
rect 12617 11384 12867 11386
rect 12617 11328 12622 11384
rect 12678 11328 12806 11384
rect 12862 11328 12867 11384
rect 12617 11326 12867 11328
rect 12617 11323 12683 11326
rect 12801 11323 12867 11326
rect 13486 11324 13492 11388
rect 13556 11386 13603 11388
rect 13556 11384 13648 11386
rect 13598 11328 13648 11384
rect 13556 11326 13648 11328
rect 13556 11324 13603 11326
rect 13537 11323 13603 11324
rect 10593 11248 10794 11250
rect 10593 11192 10598 11248
rect 10654 11192 10794 11248
rect 10593 11190 10794 11192
rect 10593 11187 10659 11190
rect 11462 11188 11468 11252
rect 11532 11250 11538 11252
rect 11973 11250 12039 11253
rect 13353 11250 13419 11253
rect 11532 11248 12039 11250
rect 11532 11192 11978 11248
rect 12034 11192 12039 11248
rect 11532 11190 12039 11192
rect 11532 11188 11538 11190
rect 11973 11187 12039 11190
rect 12896 11248 13419 11250
rect 12896 11192 13358 11248
rect 13414 11192 13419 11248
rect 12896 11190 13419 11192
rect 13816 11250 13876 11462
rect 14062 11456 14382 11457
rect 14062 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14382 11456
rect 14062 11391 14382 11392
rect 14733 11388 14799 11389
rect 14733 11384 14780 11388
rect 14844 11386 14850 11388
rect 14733 11328 14738 11384
rect 14733 11324 14780 11328
rect 14844 11326 14890 11386
rect 14844 11324 14850 11326
rect 14733 11323 14799 11324
rect 14273 11250 14339 11253
rect 13816 11248 14339 11250
rect 13816 11192 14278 11248
rect 14334 11192 14339 11248
rect 13816 11190 14339 11192
rect 12896 11117 12956 11190
rect 13353 11187 13419 11190
rect 14273 11187 14339 11190
rect 1853 11116 1919 11117
rect 1853 11112 1900 11116
rect 1964 11114 1970 11116
rect 2221 11114 2287 11117
rect 3877 11114 3943 11117
rect 5625 11114 5691 11117
rect 1853 11056 1858 11112
rect 1853 11052 1900 11056
rect 1964 11054 2010 11114
rect 2221 11112 5691 11114
rect 2221 11056 2226 11112
rect 2282 11056 3882 11112
rect 3938 11056 5630 11112
rect 5686 11056 5691 11112
rect 2221 11054 5691 11056
rect 1964 11052 1970 11054
rect 1853 11051 1919 11052
rect 2221 11051 2287 11054
rect 3877 11051 3943 11054
rect 5625 11051 5691 11054
rect 6085 11114 6151 11117
rect 8569 11114 8635 11117
rect 6085 11112 8635 11114
rect 6085 11056 6090 11112
rect 6146 11056 8574 11112
rect 8630 11056 8635 11112
rect 6085 11054 8635 11056
rect 6085 11051 6151 11054
rect 8569 11051 8635 11054
rect 8753 11114 8819 11117
rect 10910 11114 10916 11116
rect 8753 11112 10916 11114
rect 8753 11056 8758 11112
rect 8814 11056 10916 11112
rect 8753 11054 10916 11056
rect 8753 11051 8819 11054
rect 10910 11052 10916 11054
rect 10980 11052 10986 11116
rect 11513 11114 11579 11117
rect 12566 11114 12572 11116
rect 11513 11112 12572 11114
rect 11513 11056 11518 11112
rect 11574 11056 12572 11112
rect 11513 11054 12572 11056
rect 11513 11051 11579 11054
rect 12566 11052 12572 11054
rect 12636 11052 12642 11116
rect 12893 11112 12959 11117
rect 15101 11114 15167 11117
rect 12893 11056 12898 11112
rect 12954 11056 12959 11112
rect 12893 11051 12959 11056
rect 14920 11112 15167 11114
rect 14920 11056 15106 11112
rect 15162 11056 15167 11112
rect 14920 11054 15167 11056
rect 14920 10981 14980 11054
rect 15101 11051 15167 11054
rect 5993 10978 6059 10981
rect 8109 10978 8175 10981
rect 5993 10976 8175 10978
rect 5993 10920 5998 10976
rect 6054 10920 8114 10976
rect 8170 10920 8175 10976
rect 5993 10918 8175 10920
rect 5993 10915 6059 10918
rect 8109 10915 8175 10918
rect 8937 10978 9003 10981
rect 8937 10976 12128 10978
rect 8937 10920 8942 10976
rect 8998 10920 12128 10976
rect 8937 10918 12128 10920
rect 8937 10915 9003 10918
rect 4692 10912 5012 10913
rect 4692 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5012 10912
rect 4692 10847 5012 10848
rect 8440 10912 8760 10913
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 10847 8760 10848
rect 2589 10842 2655 10845
rect 2773 10842 2839 10845
rect 3366 10842 3372 10844
rect 2589 10840 3372 10842
rect 2589 10784 2594 10840
rect 2650 10784 2778 10840
rect 2834 10784 3372 10840
rect 2589 10782 3372 10784
rect 2589 10779 2655 10782
rect 2773 10779 2839 10782
rect 3366 10780 3372 10782
rect 3436 10780 3442 10844
rect 5625 10842 5691 10845
rect 6821 10842 6887 10845
rect 5625 10840 6887 10842
rect 5625 10784 5630 10840
rect 5686 10784 6826 10840
rect 6882 10784 6887 10840
rect 5625 10782 6887 10784
rect 5625 10779 5691 10782
rect 6821 10779 6887 10782
rect 7414 10780 7420 10844
rect 7484 10842 7490 10844
rect 8109 10842 8175 10845
rect 7484 10840 8175 10842
rect 7484 10784 8114 10840
rect 8170 10784 8175 10840
rect 7484 10782 8175 10784
rect 7484 10780 7490 10782
rect 8109 10779 8175 10782
rect 9438 10780 9444 10844
rect 9508 10842 9514 10844
rect 11697 10842 11763 10845
rect 9508 10840 11763 10842
rect 9508 10784 11702 10840
rect 11758 10784 11763 10840
rect 9508 10782 11763 10784
rect 9508 10780 9514 10782
rect 11697 10779 11763 10782
rect 3325 10706 3391 10709
rect 3969 10706 4035 10709
rect 11237 10706 11303 10709
rect 3325 10704 3848 10706
rect 3325 10648 3330 10704
rect 3386 10648 3848 10704
rect 3325 10646 3848 10648
rect 3325 10643 3391 10646
rect 2129 10570 2195 10573
rect 3788 10570 3848 10646
rect 3969 10704 11303 10706
rect 3969 10648 3974 10704
rect 4030 10648 11242 10704
rect 11298 10648 11303 10704
rect 3969 10646 11303 10648
rect 12068 10706 12128 10918
rect 13854 10916 13860 10980
rect 13924 10978 13930 10980
rect 14089 10978 14155 10981
rect 13924 10976 14155 10978
rect 13924 10920 14094 10976
rect 14150 10920 14155 10976
rect 13924 10918 14155 10920
rect 13924 10916 13930 10918
rect 14089 10915 14155 10918
rect 14917 10976 14983 10981
rect 14917 10920 14922 10976
rect 14978 10920 14983 10976
rect 14917 10915 14983 10920
rect 12188 10912 12508 10913
rect 12188 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12508 10912
rect 12188 10847 12508 10848
rect 13118 10780 13124 10844
rect 13188 10842 13194 10844
rect 13445 10842 13511 10845
rect 14590 10842 14596 10844
rect 13188 10840 14596 10842
rect 13188 10784 13450 10840
rect 13506 10784 14596 10840
rect 13188 10782 14596 10784
rect 13188 10780 13194 10782
rect 13445 10779 13511 10782
rect 14590 10780 14596 10782
rect 14660 10780 14666 10844
rect 12433 10706 12499 10709
rect 12893 10706 12959 10709
rect 12068 10704 12680 10706
rect 12068 10648 12438 10704
rect 12494 10648 12680 10704
rect 12068 10646 12680 10648
rect 3969 10643 4035 10646
rect 11237 10643 11303 10646
rect 12433 10643 12499 10646
rect 7925 10570 7991 10573
rect 2129 10568 3388 10570
rect 2129 10512 2134 10568
rect 2190 10512 3388 10568
rect 2129 10510 3388 10512
rect 3788 10568 7991 10570
rect 3788 10512 7930 10568
rect 7986 10512 7991 10568
rect 3788 10510 7991 10512
rect 2129 10507 2195 10510
rect 0 10434 800 10464
rect 3328 10434 3388 10510
rect 7925 10507 7991 10510
rect 8385 10570 8451 10573
rect 9070 10570 9076 10572
rect 8385 10568 9076 10570
rect 8385 10512 8390 10568
rect 8446 10512 9076 10568
rect 8385 10510 9076 10512
rect 8385 10507 8451 10510
rect 9070 10508 9076 10510
rect 9140 10570 9146 10572
rect 9990 10570 9996 10572
rect 9140 10510 9996 10570
rect 9140 10508 9146 10510
rect 9990 10508 9996 10510
rect 10060 10508 10066 10572
rect 10133 10570 10199 10573
rect 11646 10570 11652 10572
rect 10133 10568 11652 10570
rect 10133 10512 10138 10568
rect 10194 10512 11652 10568
rect 10133 10510 11652 10512
rect 10133 10507 10199 10510
rect 11646 10508 11652 10510
rect 11716 10508 11722 10572
rect 12620 10570 12680 10646
rect 12893 10704 13140 10706
rect 12893 10648 12898 10704
rect 12954 10648 13140 10704
rect 12893 10646 13140 10648
rect 12893 10643 12959 10646
rect 12893 10570 12959 10573
rect 12620 10568 12959 10570
rect 12620 10512 12898 10568
rect 12954 10512 12959 10568
rect 12620 10510 12959 10512
rect 13080 10570 13140 10646
rect 13670 10644 13676 10708
rect 13740 10706 13746 10708
rect 14549 10706 14615 10709
rect 13740 10704 14615 10706
rect 13740 10648 14554 10704
rect 14610 10648 14615 10704
rect 13740 10646 14615 10648
rect 13740 10644 13746 10646
rect 14549 10643 14615 10646
rect 13486 10570 13492 10572
rect 13080 10510 13492 10570
rect 12893 10507 12959 10510
rect 13486 10508 13492 10510
rect 13556 10508 13562 10572
rect 15653 10570 15719 10573
rect 13862 10568 15719 10570
rect 13862 10512 15658 10568
rect 15714 10512 15719 10568
rect 13862 10510 15719 10512
rect 7097 10434 7163 10437
rect 10133 10434 10199 10437
rect 0 10374 1410 10434
rect 3328 10374 4170 10434
rect 0 10344 800 10374
rect 1350 10162 1410 10374
rect 2818 10368 3138 10369
rect 2818 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3138 10368
rect 2818 10303 3138 10304
rect 3969 10162 4035 10165
rect 1350 10160 4035 10162
rect 1350 10104 3974 10160
rect 4030 10104 4035 10160
rect 1350 10102 4035 10104
rect 4110 10162 4170 10374
rect 7097 10432 10199 10434
rect 7097 10376 7102 10432
rect 7158 10376 10138 10432
rect 10194 10376 10199 10432
rect 7097 10374 10199 10376
rect 7097 10371 7163 10374
rect 10133 10371 10199 10374
rect 10961 10434 11027 10437
rect 13862 10434 13922 10510
rect 15653 10507 15719 10510
rect 10961 10432 13922 10434
rect 10961 10376 10966 10432
rect 11022 10376 13922 10432
rect 10961 10374 13922 10376
rect 10961 10371 11027 10374
rect 6566 10368 6886 10369
rect 6566 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6886 10368
rect 6566 10303 6886 10304
rect 10314 10368 10634 10369
rect 10314 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10634 10368
rect 10314 10303 10634 10304
rect 14062 10368 14382 10369
rect 14062 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14382 10368
rect 14062 10303 14382 10304
rect 4337 10298 4403 10301
rect 4797 10298 4863 10301
rect 4337 10296 4863 10298
rect 4337 10240 4342 10296
rect 4398 10240 4802 10296
rect 4858 10240 4863 10296
rect 4337 10238 4863 10240
rect 4337 10235 4403 10238
rect 4797 10235 4863 10238
rect 7005 10298 7071 10301
rect 10133 10298 10199 10301
rect 7005 10296 10199 10298
rect 7005 10240 7010 10296
rect 7066 10240 10138 10296
rect 10194 10240 10199 10296
rect 7005 10238 10199 10240
rect 7005 10235 7071 10238
rect 10133 10235 10199 10238
rect 10777 10298 10843 10301
rect 13854 10298 13860 10300
rect 10777 10296 13860 10298
rect 10777 10240 10782 10296
rect 10838 10240 13860 10296
rect 10777 10238 13860 10240
rect 10777 10235 10843 10238
rect 13854 10236 13860 10238
rect 13924 10236 13930 10300
rect 8886 10162 8892 10164
rect 4110 10102 8892 10162
rect 3969 10099 4035 10102
rect 8886 10100 8892 10102
rect 8956 10100 8962 10164
rect 9305 10162 9371 10165
rect 12750 10162 12756 10164
rect 9305 10160 12756 10162
rect 9305 10104 9310 10160
rect 9366 10104 12756 10160
rect 9305 10102 12756 10104
rect 9305 10099 9371 10102
rect 12750 10100 12756 10102
rect 12820 10100 12826 10164
rect 14181 10162 14247 10165
rect 13264 10160 14247 10162
rect 13264 10104 14186 10160
rect 14242 10104 14247 10160
rect 13264 10102 14247 10104
rect 2313 10026 2379 10029
rect 9397 10026 9463 10029
rect 2313 10024 9463 10026
rect 2313 9968 2318 10024
rect 2374 9968 9402 10024
rect 9458 9968 9463 10024
rect 2313 9966 9463 9968
rect 2313 9963 2379 9966
rect 9397 9963 9463 9966
rect 10685 10026 10751 10029
rect 11881 10026 11947 10029
rect 13264 10026 13324 10102
rect 14181 10099 14247 10102
rect 10685 10024 13324 10026
rect 10685 9968 10690 10024
rect 10746 9968 11886 10024
rect 11942 9968 13324 10024
rect 10685 9966 13324 9968
rect 13445 10026 13511 10029
rect 16400 10026 17200 10056
rect 13445 10024 17200 10026
rect 13445 9968 13450 10024
rect 13506 9968 17200 10024
rect 13445 9966 17200 9968
rect 10685 9963 10751 9966
rect 11881 9963 11947 9966
rect 13445 9963 13511 9966
rect 16400 9936 17200 9966
rect 2589 9890 2655 9893
rect 4102 9890 4108 9892
rect 2589 9888 4108 9890
rect 2589 9832 2594 9888
rect 2650 9832 4108 9888
rect 2589 9830 4108 9832
rect 2589 9827 2655 9830
rect 4102 9828 4108 9830
rect 4172 9890 4178 9892
rect 4470 9890 4476 9892
rect 4172 9830 4476 9890
rect 4172 9828 4178 9830
rect 4470 9828 4476 9830
rect 4540 9828 4546 9892
rect 6269 9890 6335 9893
rect 7925 9890 7991 9893
rect 6269 9888 7991 9890
rect 6269 9832 6274 9888
rect 6330 9832 7930 9888
rect 7986 9832 7991 9888
rect 6269 9830 7991 9832
rect 6269 9827 6335 9830
rect 7925 9827 7991 9830
rect 10174 9828 10180 9892
rect 10244 9890 10250 9892
rect 10961 9890 11027 9893
rect 11145 9892 11211 9893
rect 10244 9888 11027 9890
rect 10244 9832 10966 9888
rect 11022 9832 11027 9888
rect 10244 9830 11027 9832
rect 10244 9828 10250 9830
rect 10961 9827 11027 9830
rect 11094 9828 11100 9892
rect 11164 9890 11211 9892
rect 11605 9890 11671 9893
rect 11973 9890 12039 9893
rect 11164 9888 12039 9890
rect 11206 9832 11610 9888
rect 11666 9832 11978 9888
rect 12034 9832 12039 9888
rect 11164 9830 12039 9832
rect 11164 9828 11211 9830
rect 11145 9827 11211 9828
rect 11605 9827 11671 9830
rect 11973 9827 12039 9830
rect 13353 9890 13419 9893
rect 13486 9890 13492 9892
rect 13353 9888 13492 9890
rect 13353 9832 13358 9888
rect 13414 9832 13492 9888
rect 13353 9830 13492 9832
rect 13353 9827 13419 9830
rect 13486 9828 13492 9830
rect 13556 9828 13562 9892
rect 13854 9828 13860 9892
rect 13924 9890 13930 9892
rect 14089 9890 14155 9893
rect 13924 9888 14155 9890
rect 13924 9832 14094 9888
rect 14150 9832 14155 9888
rect 13924 9830 14155 9832
rect 13924 9828 13930 9830
rect 14089 9827 14155 9830
rect 4692 9824 5012 9825
rect 4692 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5012 9824
rect 4692 9759 5012 9760
rect 8440 9824 8760 9825
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 9759 8760 9760
rect 12188 9824 12508 9825
rect 12188 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12508 9824
rect 12188 9759 12508 9760
rect 5073 9754 5139 9757
rect 8109 9754 8175 9757
rect 5073 9752 8175 9754
rect 5073 9696 5078 9752
rect 5134 9696 8114 9752
rect 8170 9696 8175 9752
rect 5073 9694 8175 9696
rect 5073 9691 5139 9694
rect 8109 9691 8175 9694
rect 8845 9754 8911 9757
rect 9029 9754 9095 9757
rect 8845 9752 9095 9754
rect 8845 9696 8850 9752
rect 8906 9696 9034 9752
rect 9090 9696 9095 9752
rect 8845 9694 9095 9696
rect 8845 9691 8911 9694
rect 9029 9691 9095 9694
rect 9581 9754 9647 9757
rect 13118 9754 13124 9756
rect 9581 9752 12128 9754
rect 9581 9696 9586 9752
rect 9642 9696 12128 9752
rect 9581 9694 12128 9696
rect 9581 9691 9647 9694
rect 2957 9618 3023 9621
rect 7414 9618 7420 9620
rect 2957 9616 7420 9618
rect 2957 9560 2962 9616
rect 3018 9560 7420 9616
rect 2957 9558 7420 9560
rect 2957 9555 3023 9558
rect 7414 9556 7420 9558
rect 7484 9618 7490 9620
rect 9029 9618 9095 9621
rect 7484 9616 9095 9618
rect 7484 9560 9034 9616
rect 9090 9560 9095 9616
rect 7484 9558 9095 9560
rect 7484 9556 7490 9558
rect 9029 9555 9095 9558
rect 9857 9618 9923 9621
rect 10593 9618 10659 9621
rect 9857 9616 10659 9618
rect 9857 9560 9862 9616
rect 9918 9560 10598 9616
rect 10654 9560 10659 9616
rect 9857 9558 10659 9560
rect 9857 9555 9923 9558
rect 10593 9555 10659 9558
rect 10910 9556 10916 9620
rect 10980 9618 10986 9620
rect 11145 9618 11211 9621
rect 10980 9616 11211 9618
rect 10980 9560 11150 9616
rect 11206 9560 11211 9616
rect 10980 9558 11211 9560
rect 12068 9618 12128 9694
rect 12988 9694 13124 9754
rect 12988 9618 13048 9694
rect 13118 9692 13124 9694
rect 13188 9692 13194 9756
rect 13261 9754 13327 9757
rect 14549 9754 14615 9757
rect 13261 9752 14615 9754
rect 13261 9696 13266 9752
rect 13322 9696 14554 9752
rect 14610 9696 14615 9752
rect 13261 9694 14615 9696
rect 13261 9691 13327 9694
rect 14549 9691 14615 9694
rect 12068 9558 13048 9618
rect 13169 9618 13235 9621
rect 13302 9618 13308 9620
rect 13169 9616 13308 9618
rect 13169 9560 13174 9616
rect 13230 9560 13308 9616
rect 13169 9558 13308 9560
rect 10980 9556 10986 9558
rect 11145 9555 11211 9558
rect 13169 9555 13235 9558
rect 13302 9556 13308 9558
rect 13372 9556 13378 9620
rect 0 9482 800 9512
rect 1393 9482 1459 9485
rect 0 9480 1459 9482
rect 0 9424 1398 9480
rect 1454 9424 1459 9480
rect 0 9422 1459 9424
rect 0 9392 800 9422
rect 1393 9419 1459 9422
rect 2129 9482 2195 9485
rect 5533 9482 5599 9485
rect 2129 9480 5599 9482
rect 2129 9424 2134 9480
rect 2190 9424 5538 9480
rect 5594 9424 5599 9480
rect 2129 9422 5599 9424
rect 2129 9419 2195 9422
rect 5533 9419 5599 9422
rect 6913 9482 6979 9485
rect 10225 9482 10291 9485
rect 10685 9482 10751 9485
rect 6913 9480 10751 9482
rect 6913 9424 6918 9480
rect 6974 9424 10230 9480
rect 10286 9424 10690 9480
rect 10746 9424 10751 9480
rect 6913 9422 10751 9424
rect 6913 9419 6979 9422
rect 10225 9419 10291 9422
rect 10685 9419 10751 9422
rect 11237 9482 11303 9485
rect 16389 9482 16455 9485
rect 11237 9480 16455 9482
rect 11237 9424 11242 9480
rect 11298 9424 16394 9480
rect 16450 9424 16455 9480
rect 11237 9422 16455 9424
rect 11237 9419 11303 9422
rect 16389 9419 16455 9422
rect 7281 9348 7347 9349
rect 7230 9284 7236 9348
rect 7300 9346 7347 9348
rect 11513 9346 11579 9349
rect 11881 9346 11947 9349
rect 7300 9344 7392 9346
rect 7342 9288 7392 9344
rect 7300 9286 7392 9288
rect 11513 9344 11947 9346
rect 11513 9288 11518 9344
rect 11574 9288 11886 9344
rect 11942 9288 11947 9344
rect 11513 9286 11947 9288
rect 7300 9284 7347 9286
rect 7281 9283 7347 9284
rect 11513 9283 11579 9286
rect 11881 9283 11947 9286
rect 12014 9284 12020 9348
rect 12084 9346 12090 9348
rect 13077 9346 13143 9349
rect 12084 9344 13143 9346
rect 12084 9288 13082 9344
rect 13138 9288 13143 9344
rect 12084 9286 13143 9288
rect 12084 9284 12090 9286
rect 13077 9283 13143 9286
rect 13445 9346 13511 9349
rect 13813 9346 13879 9349
rect 13445 9344 13879 9346
rect 13445 9288 13450 9344
rect 13506 9288 13818 9344
rect 13874 9288 13879 9344
rect 13445 9286 13879 9288
rect 13445 9283 13511 9286
rect 13813 9283 13879 9286
rect 2818 9280 3138 9281
rect 2818 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3138 9280
rect 2818 9215 3138 9216
rect 6566 9280 6886 9281
rect 6566 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6886 9280
rect 6566 9215 6886 9216
rect 10314 9280 10634 9281
rect 10314 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10634 9280
rect 10314 9215 10634 9216
rect 14062 9280 14382 9281
rect 14062 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14382 9280
rect 14062 9215 14382 9216
rect 3877 9210 3943 9213
rect 5441 9210 5507 9213
rect 3877 9208 5507 9210
rect 3877 9152 3882 9208
rect 3938 9152 5446 9208
rect 5502 9152 5507 9208
rect 3877 9150 5507 9152
rect 3877 9147 3943 9150
rect 5441 9147 5507 9150
rect 7230 9148 7236 9212
rect 7300 9210 7306 9212
rect 10961 9210 11027 9213
rect 12433 9210 12499 9213
rect 7300 9150 10242 9210
rect 7300 9148 7306 9150
rect 1669 9074 1735 9077
rect 10041 9074 10107 9077
rect 1669 9072 10107 9074
rect 1669 9016 1674 9072
rect 1730 9016 10046 9072
rect 10102 9016 10107 9072
rect 1669 9014 10107 9016
rect 10182 9074 10242 9150
rect 10961 9208 12499 9210
rect 10961 9152 10966 9208
rect 11022 9152 12438 9208
rect 12494 9152 12499 9208
rect 10961 9150 12499 9152
rect 10961 9147 11027 9150
rect 12433 9147 12499 9150
rect 12566 9148 12572 9212
rect 12636 9210 12642 9212
rect 14457 9210 14523 9213
rect 16113 9210 16179 9213
rect 12636 9150 13140 9210
rect 12636 9148 12642 9150
rect 12893 9074 12959 9077
rect 10182 9072 12959 9074
rect 10182 9016 12898 9072
rect 12954 9016 12959 9072
rect 10182 9014 12959 9016
rect 13080 9074 13140 9150
rect 14457 9208 16179 9210
rect 14457 9152 14462 9208
rect 14518 9152 16118 9208
rect 16174 9152 16179 9208
rect 14457 9150 16179 9152
rect 14457 9147 14523 9150
rect 16113 9147 16179 9150
rect 16481 9074 16547 9077
rect 13080 9072 16547 9074
rect 13080 9016 16486 9072
rect 16542 9016 16547 9072
rect 13080 9014 16547 9016
rect 1669 9011 1735 9014
rect 10041 9011 10107 9014
rect 12893 9011 12959 9014
rect 16481 9011 16547 9014
rect 1853 8938 1919 8941
rect 5809 8938 5875 8941
rect 1853 8936 5875 8938
rect 1853 8880 1858 8936
rect 1914 8880 5814 8936
rect 5870 8880 5875 8936
rect 1853 8878 5875 8880
rect 1853 8875 1919 8878
rect 5809 8875 5875 8878
rect 6310 8876 6316 8940
rect 6380 8938 6386 8940
rect 7005 8938 7071 8941
rect 6380 8936 7071 8938
rect 6380 8880 7010 8936
rect 7066 8880 7071 8936
rect 6380 8878 7071 8880
rect 6380 8876 6386 8878
rect 7005 8875 7071 8878
rect 7465 8938 7531 8941
rect 13169 8938 13235 8941
rect 7465 8936 13235 8938
rect 7465 8880 7470 8936
rect 7526 8880 13174 8936
rect 13230 8880 13235 8936
rect 7465 8878 13235 8880
rect 7465 8875 7531 8878
rect 13169 8875 13235 8878
rect 9029 8802 9095 8805
rect 9673 8802 9739 8805
rect 11789 8804 11855 8805
rect 9806 8802 9812 8804
rect 9029 8800 9812 8802
rect 9029 8744 9034 8800
rect 9090 8744 9678 8800
rect 9734 8744 9812 8800
rect 9029 8742 9812 8744
rect 9029 8739 9095 8742
rect 9673 8739 9739 8742
rect 9806 8740 9812 8742
rect 9876 8740 9882 8804
rect 11789 8802 11836 8804
rect 11744 8800 11836 8802
rect 11744 8744 11794 8800
rect 11744 8742 11836 8744
rect 11789 8740 11836 8742
rect 11900 8740 11906 8804
rect 12801 8802 12867 8805
rect 14825 8802 14891 8805
rect 12801 8800 14891 8802
rect 12801 8744 12806 8800
rect 12862 8744 14830 8800
rect 14886 8744 14891 8800
rect 12801 8742 14891 8744
rect 11789 8739 11855 8740
rect 12801 8739 12867 8742
rect 14825 8739 14891 8742
rect 4692 8736 5012 8737
rect 4692 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5012 8736
rect 4692 8671 5012 8672
rect 8440 8736 8760 8737
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 8671 8760 8672
rect 12188 8736 12508 8737
rect 12188 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12508 8736
rect 12188 8671 12508 8672
rect 10041 8666 10107 8669
rect 12801 8666 12867 8669
rect 12934 8666 12940 8668
rect 10041 8664 11852 8666
rect 10041 8608 10046 8664
rect 10102 8608 11852 8664
rect 10041 8606 11852 8608
rect 10041 8603 10107 8606
rect 2313 8530 2379 8533
rect 11513 8530 11579 8533
rect 2313 8528 11579 8530
rect 2313 8472 2318 8528
rect 2374 8472 11518 8528
rect 11574 8472 11579 8528
rect 2313 8470 11579 8472
rect 11792 8530 11852 8606
rect 12801 8664 12940 8666
rect 12801 8608 12806 8664
rect 12862 8608 12940 8664
rect 12801 8606 12940 8608
rect 12801 8603 12867 8606
rect 12934 8604 12940 8606
rect 13004 8604 13010 8668
rect 13077 8666 13143 8669
rect 15101 8666 15167 8669
rect 13077 8664 15167 8666
rect 13077 8608 13082 8664
rect 13138 8608 15106 8664
rect 15162 8608 15167 8664
rect 13077 8606 15167 8608
rect 13077 8603 13143 8606
rect 15101 8603 15167 8606
rect 12157 8530 12223 8533
rect 11792 8528 12223 8530
rect 11792 8472 12162 8528
rect 12218 8472 12223 8528
rect 11792 8470 12223 8472
rect 2313 8467 2379 8470
rect 11513 8467 11579 8470
rect 12157 8467 12223 8470
rect 12525 8530 12591 8533
rect 16205 8530 16271 8533
rect 12525 8528 16271 8530
rect 12525 8472 12530 8528
rect 12586 8472 16210 8528
rect 16266 8472 16271 8528
rect 12525 8470 16271 8472
rect 12525 8467 12591 8470
rect 16205 8467 16271 8470
rect 0 8394 800 8424
rect 3969 8394 4035 8397
rect 5533 8396 5599 8397
rect 5533 8394 5580 8396
rect 0 8392 4035 8394
rect 0 8336 3974 8392
rect 4030 8336 4035 8392
rect 0 8334 4035 8336
rect 5488 8392 5580 8394
rect 5488 8336 5538 8392
rect 5488 8334 5580 8336
rect 0 8304 800 8334
rect 3969 8331 4035 8334
rect 5533 8332 5580 8334
rect 5644 8332 5650 8396
rect 6310 8332 6316 8396
rect 6380 8394 6386 8396
rect 9857 8394 9923 8397
rect 6380 8392 9923 8394
rect 6380 8336 9862 8392
rect 9918 8336 9923 8392
rect 6380 8334 9923 8336
rect 6380 8332 6386 8334
rect 5533 8331 5599 8332
rect 9857 8331 9923 8334
rect 10133 8394 10199 8397
rect 10777 8394 10843 8397
rect 10133 8392 10843 8394
rect 10133 8336 10138 8392
rect 10194 8336 10782 8392
rect 10838 8336 10843 8392
rect 10133 8334 10843 8336
rect 10133 8331 10199 8334
rect 10777 8331 10843 8334
rect 11830 8332 11836 8396
rect 11900 8394 11906 8396
rect 11973 8394 12039 8397
rect 12709 8394 12775 8397
rect 13169 8396 13235 8397
rect 11900 8392 12775 8394
rect 11900 8336 11978 8392
rect 12034 8336 12714 8392
rect 12770 8336 12775 8392
rect 11900 8334 12775 8336
rect 11900 8332 11906 8334
rect 11973 8331 12039 8334
rect 12709 8331 12775 8334
rect 13118 8332 13124 8396
rect 13188 8394 13235 8396
rect 13353 8394 13419 8397
rect 13670 8394 13676 8396
rect 13188 8392 13280 8394
rect 13230 8336 13280 8392
rect 13188 8334 13280 8336
rect 13353 8392 13676 8394
rect 13353 8336 13358 8392
rect 13414 8336 13676 8392
rect 13353 8334 13676 8336
rect 13188 8332 13235 8334
rect 13169 8331 13235 8332
rect 13353 8331 13419 8334
rect 13670 8332 13676 8334
rect 13740 8332 13746 8396
rect 16573 8394 16639 8397
rect 13816 8392 16639 8394
rect 13816 8336 16578 8392
rect 16634 8336 16639 8392
rect 13816 8334 16639 8336
rect 3601 8258 3667 8261
rect 3918 8258 3924 8260
rect 3601 8256 3924 8258
rect 3601 8200 3606 8256
rect 3662 8200 3924 8256
rect 3601 8198 3924 8200
rect 3601 8195 3667 8198
rect 3918 8196 3924 8198
rect 3988 8196 3994 8260
rect 5214 8198 6378 8258
rect 2818 8192 3138 8193
rect 2818 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3138 8192
rect 2818 8127 3138 8128
rect 3734 8060 3740 8124
rect 3804 8122 3810 8124
rect 5214 8122 5274 8198
rect 3804 8062 5274 8122
rect 3804 8060 3810 8062
rect 5390 8060 5396 8124
rect 5460 8122 5466 8124
rect 5809 8122 5875 8125
rect 5460 8120 5875 8122
rect 5460 8064 5814 8120
rect 5870 8064 5875 8120
rect 5460 8062 5875 8064
rect 5460 8060 5466 8062
rect 5809 8059 5875 8062
rect 1025 7986 1091 7989
rect 5625 7986 5691 7989
rect 1025 7984 5691 7986
rect 1025 7928 1030 7984
rect 1086 7928 5630 7984
rect 5686 7928 5691 7984
rect 1025 7926 5691 7928
rect 6318 7986 6378 8198
rect 7966 8196 7972 8260
rect 8036 8258 8042 8260
rect 10041 8258 10107 8261
rect 8036 8256 10107 8258
rect 8036 8200 10046 8256
rect 10102 8200 10107 8256
rect 8036 8198 10107 8200
rect 10780 8258 10840 8331
rect 11278 8258 11284 8260
rect 10780 8198 11284 8258
rect 8036 8196 8042 8198
rect 10041 8195 10107 8198
rect 11278 8196 11284 8198
rect 11348 8258 11354 8260
rect 12934 8258 12940 8260
rect 11348 8198 12940 8258
rect 11348 8196 11354 8198
rect 12934 8196 12940 8198
rect 13004 8196 13010 8260
rect 13169 8258 13235 8261
rect 13356 8258 13416 8331
rect 13169 8256 13416 8258
rect 13169 8200 13174 8256
rect 13230 8200 13416 8256
rect 13169 8198 13416 8200
rect 6566 8192 6886 8193
rect 6566 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6886 8192
rect 6566 8127 6886 8128
rect 10314 8192 10634 8193
rect 10314 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10634 8192
rect 10314 8127 10634 8128
rect 8150 8060 8156 8124
rect 8220 8122 8226 8124
rect 9254 8122 9260 8124
rect 8220 8062 9260 8122
rect 8220 8060 8226 8062
rect 9254 8060 9260 8062
rect 9324 8060 9330 8124
rect 9949 8122 10015 8125
rect 9492 8120 10015 8122
rect 9492 8064 9954 8120
rect 10010 8064 10015 8120
rect 9492 8062 10015 8064
rect 9492 7986 9552 8062
rect 9949 8059 10015 8062
rect 11881 8122 11947 8125
rect 12525 8124 12591 8125
rect 12014 8122 12020 8124
rect 11881 8120 12020 8122
rect 11881 8064 11886 8120
rect 11942 8064 12020 8120
rect 11881 8062 12020 8064
rect 11881 8059 11947 8062
rect 12014 8060 12020 8062
rect 12084 8060 12090 8124
rect 12525 8120 12572 8124
rect 12636 8122 12642 8124
rect 12942 8122 13002 8196
rect 13169 8195 13235 8198
rect 13816 8125 13876 8334
rect 16573 8331 16639 8334
rect 14062 8192 14382 8193
rect 14062 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14382 8192
rect 14062 8127 14382 8128
rect 13537 8122 13603 8125
rect 12525 8064 12530 8120
rect 12525 8060 12572 8064
rect 12636 8062 12682 8122
rect 12942 8120 13603 8122
rect 12942 8064 13542 8120
rect 13598 8064 13603 8120
rect 12942 8062 13603 8064
rect 12636 8060 12642 8062
rect 12525 8059 12591 8060
rect 13537 8059 13603 8062
rect 13813 8120 13879 8125
rect 13813 8064 13818 8120
rect 13874 8064 13879 8120
rect 13813 8059 13879 8064
rect 14549 8122 14615 8125
rect 14958 8122 14964 8124
rect 14549 8120 14964 8122
rect 14549 8064 14554 8120
rect 14610 8064 14964 8120
rect 14549 8062 14964 8064
rect 14549 8059 14615 8062
rect 14958 8060 14964 8062
rect 15028 8060 15034 8124
rect 15101 8122 15167 8125
rect 15326 8122 15332 8124
rect 15101 8120 15332 8122
rect 15101 8064 15106 8120
rect 15162 8064 15332 8120
rect 15101 8062 15332 8064
rect 15101 8059 15167 8062
rect 15326 8060 15332 8062
rect 15396 8060 15402 8124
rect 6318 7926 9552 7986
rect 9673 7986 9739 7989
rect 15469 7986 15535 7989
rect 9673 7984 15535 7986
rect 9673 7928 9678 7984
rect 9734 7928 15474 7984
rect 15530 7928 15535 7984
rect 9673 7926 15535 7928
rect 1025 7923 1091 7926
rect 5625 7923 5691 7926
rect 9673 7923 9739 7926
rect 15469 7923 15535 7926
rect 1342 7788 1348 7852
rect 1412 7850 1418 7852
rect 5390 7850 5396 7852
rect 1412 7790 5396 7850
rect 1412 7788 1418 7790
rect 5390 7788 5396 7790
rect 5460 7788 5466 7852
rect 5901 7850 5967 7853
rect 11237 7850 11303 7853
rect 5901 7848 11303 7850
rect 5901 7792 5906 7848
rect 5962 7792 11242 7848
rect 11298 7792 11303 7848
rect 5901 7790 11303 7792
rect 5901 7787 5967 7790
rect 11237 7787 11303 7790
rect 11513 7850 11579 7853
rect 15929 7850 15995 7853
rect 11513 7848 15995 7850
rect 11513 7792 11518 7848
rect 11574 7792 15934 7848
rect 15990 7792 15995 7848
rect 11513 7790 15995 7792
rect 11513 7787 11579 7790
rect 15929 7787 15995 7790
rect 3601 7716 3667 7717
rect 3550 7714 3556 7716
rect 3510 7654 3556 7714
rect 3620 7712 3667 7716
rect 3662 7656 3667 7712
rect 3550 7652 3556 7654
rect 3620 7652 3667 7656
rect 3601 7651 3667 7652
rect 5993 7714 6059 7717
rect 7281 7714 7347 7717
rect 5993 7712 7347 7714
rect 5993 7656 5998 7712
rect 6054 7656 7286 7712
rect 7342 7656 7347 7712
rect 5993 7654 7347 7656
rect 5993 7651 6059 7654
rect 7281 7651 7347 7654
rect 9806 7652 9812 7716
rect 9876 7714 9882 7716
rect 10685 7714 10751 7717
rect 9876 7712 10751 7714
rect 9876 7656 10690 7712
rect 10746 7656 10751 7712
rect 9876 7654 10751 7656
rect 9876 7652 9882 7654
rect 10685 7651 10751 7654
rect 12985 7714 13051 7717
rect 15469 7714 15535 7717
rect 12985 7712 15535 7714
rect 12985 7656 12990 7712
rect 13046 7656 15474 7712
rect 15530 7656 15535 7712
rect 12985 7654 15535 7656
rect 12985 7651 13051 7654
rect 15469 7651 15535 7654
rect 4692 7648 5012 7649
rect 4692 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5012 7648
rect 4692 7583 5012 7584
rect 8440 7648 8760 7649
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 7583 8760 7584
rect 12188 7648 12508 7649
rect 12188 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12508 7648
rect 12188 7583 12508 7584
rect 8886 7516 8892 7580
rect 8956 7578 8962 7580
rect 13077 7578 13143 7581
rect 13721 7580 13787 7581
rect 13302 7578 13308 7580
rect 8956 7518 12036 7578
rect 8956 7516 8962 7518
rect 0 7442 800 7472
rect 3141 7442 3207 7445
rect 0 7440 3207 7442
rect 0 7384 3146 7440
rect 3202 7384 3207 7440
rect 0 7382 3207 7384
rect 0 7352 800 7382
rect 3141 7379 3207 7382
rect 5942 7380 5948 7444
rect 6012 7442 6018 7444
rect 11145 7442 11211 7445
rect 6012 7440 11211 7442
rect 6012 7384 11150 7440
rect 11206 7384 11211 7440
rect 6012 7382 11211 7384
rect 11976 7442 12036 7518
rect 13077 7576 13308 7578
rect 13077 7520 13082 7576
rect 13138 7520 13308 7576
rect 13077 7518 13308 7520
rect 13077 7515 13143 7518
rect 13302 7516 13308 7518
rect 13372 7516 13378 7580
rect 13670 7516 13676 7580
rect 13740 7578 13787 7580
rect 13740 7576 13832 7578
rect 13782 7520 13832 7576
rect 13740 7518 13832 7520
rect 13740 7516 13787 7518
rect 13721 7515 13787 7516
rect 15193 7442 15259 7445
rect 11976 7440 15259 7442
rect 11976 7384 15198 7440
rect 15254 7384 15259 7440
rect 11976 7382 15259 7384
rect 6012 7380 6018 7382
rect 11145 7379 11211 7382
rect 15193 7379 15259 7382
rect 3049 7306 3115 7309
rect 6453 7306 6519 7309
rect 3049 7304 6519 7306
rect 3049 7248 3054 7304
rect 3110 7248 6458 7304
rect 6514 7248 6519 7304
rect 3049 7246 6519 7248
rect 3049 7243 3115 7246
rect 6453 7243 6519 7246
rect 6913 7306 6979 7309
rect 7925 7306 7991 7309
rect 6913 7304 7991 7306
rect 6913 7248 6918 7304
rect 6974 7248 7930 7304
rect 7986 7248 7991 7304
rect 6913 7246 7991 7248
rect 6913 7243 6979 7246
rect 7925 7243 7991 7246
rect 8293 7306 8359 7309
rect 11053 7306 11119 7309
rect 8293 7304 11119 7306
rect 8293 7248 8298 7304
rect 8354 7248 11058 7304
rect 11114 7248 11119 7304
rect 8293 7246 11119 7248
rect 8293 7243 8359 7246
rect 11053 7243 11119 7246
rect 11462 7244 11468 7308
rect 11532 7306 11538 7308
rect 12566 7306 12572 7308
rect 11532 7246 12572 7306
rect 11532 7244 11538 7246
rect 12566 7244 12572 7246
rect 12636 7306 12642 7308
rect 12709 7306 12775 7309
rect 12636 7304 12775 7306
rect 12636 7248 12714 7304
rect 12770 7248 12775 7304
rect 12636 7246 12775 7248
rect 12636 7244 12642 7246
rect 12709 7243 12775 7246
rect 13118 7244 13124 7308
rect 13188 7306 13194 7308
rect 14457 7306 14523 7309
rect 13188 7304 14523 7306
rect 13188 7248 14462 7304
rect 14518 7248 14523 7304
rect 13188 7246 14523 7248
rect 13188 7244 13194 7246
rect 14457 7243 14523 7246
rect 7281 7170 7347 7173
rect 10133 7170 10199 7173
rect 7281 7168 10199 7170
rect 7281 7112 7286 7168
rect 7342 7112 10138 7168
rect 10194 7112 10199 7168
rect 7281 7110 10199 7112
rect 7281 7107 7347 7110
rect 10133 7107 10199 7110
rect 11329 7170 11395 7173
rect 11973 7170 12039 7173
rect 11329 7168 12039 7170
rect 11329 7112 11334 7168
rect 11390 7112 11978 7168
rect 12034 7112 12039 7168
rect 11329 7110 12039 7112
rect 11329 7107 11395 7110
rect 11973 7107 12039 7110
rect 12433 7170 12499 7173
rect 12617 7170 12683 7173
rect 12433 7168 12683 7170
rect 12433 7112 12438 7168
rect 12494 7112 12622 7168
rect 12678 7112 12683 7168
rect 12433 7110 12683 7112
rect 12433 7107 12499 7110
rect 12617 7107 12683 7110
rect 2818 7104 3138 7105
rect 2818 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3138 7104
rect 2818 7039 3138 7040
rect 6566 7104 6886 7105
rect 6566 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6886 7104
rect 6566 7039 6886 7040
rect 10314 7104 10634 7105
rect 10314 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10634 7104
rect 10314 7039 10634 7040
rect 14062 7104 14382 7105
rect 14062 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14382 7104
rect 14062 7039 14382 7040
rect 3785 7036 3851 7037
rect 3734 6972 3740 7036
rect 3804 7034 3851 7036
rect 4521 7034 4587 7037
rect 7097 7034 7163 7037
rect 9121 7034 9187 7037
rect 3804 7032 3896 7034
rect 3846 6976 3896 7032
rect 3804 6974 3896 6976
rect 4521 7032 6332 7034
rect 4521 6976 4526 7032
rect 4582 6976 6332 7032
rect 4521 6974 6332 6976
rect 3804 6972 3851 6974
rect 3785 6971 3851 6972
rect 4521 6971 4587 6974
rect 1761 6900 1827 6901
rect 1710 6898 1716 6900
rect 1670 6838 1716 6898
rect 1780 6896 1827 6900
rect 4429 6900 4495 6901
rect 4429 6898 4476 6900
rect 1822 6840 1827 6896
rect 1710 6836 1716 6838
rect 1780 6836 1827 6840
rect 4384 6896 4476 6898
rect 4384 6840 4434 6896
rect 4384 6838 4476 6840
rect 1761 6835 1827 6836
rect 4429 6836 4476 6838
rect 4540 6836 4546 6900
rect 5758 6836 5764 6900
rect 5828 6898 5834 6900
rect 6085 6898 6151 6901
rect 5828 6896 6151 6898
rect 5828 6840 6090 6896
rect 6146 6840 6151 6896
rect 5828 6838 6151 6840
rect 6272 6898 6332 6974
rect 7097 7032 9187 7034
rect 7097 6976 7102 7032
rect 7158 6976 9126 7032
rect 9182 6976 9187 7032
rect 7097 6974 9187 6976
rect 7097 6971 7163 6974
rect 9121 6971 9187 6974
rect 9489 7034 9555 7037
rect 10041 7034 10107 7037
rect 9489 7032 10107 7034
rect 9489 6976 9494 7032
rect 9550 6976 10046 7032
rect 10102 6976 10107 7032
rect 9489 6974 10107 6976
rect 9489 6971 9555 6974
rect 10041 6971 10107 6974
rect 10777 7034 10843 7037
rect 12525 7034 12591 7037
rect 12750 7034 12756 7036
rect 10777 7032 12220 7034
rect 10777 6976 10782 7032
rect 10838 6976 12220 7032
rect 10777 6974 12220 6976
rect 10777 6971 10843 6974
rect 8293 6898 8359 6901
rect 6272 6896 8359 6898
rect 6272 6840 8298 6896
rect 8354 6840 8359 6896
rect 6272 6838 8359 6840
rect 5828 6836 5834 6838
rect 4429 6835 4495 6836
rect 6085 6835 6151 6838
rect 8293 6835 8359 6838
rect 8845 6898 8911 6901
rect 12014 6898 12020 6900
rect 8845 6896 12020 6898
rect 8845 6840 8850 6896
rect 8906 6840 12020 6896
rect 8845 6838 12020 6840
rect 8845 6835 8911 6838
rect 12014 6836 12020 6838
rect 12084 6836 12090 6900
rect 12160 6898 12220 6974
rect 12525 7032 12756 7034
rect 12525 6976 12530 7032
rect 12586 6976 12756 7032
rect 12525 6974 12756 6976
rect 12525 6971 12591 6974
rect 12750 6972 12756 6974
rect 12820 6972 12826 7036
rect 13353 7034 13419 7037
rect 13486 7034 13492 7036
rect 13353 7032 13492 7034
rect 13353 6976 13358 7032
rect 13414 6976 13492 7032
rect 13353 6974 13492 6976
rect 13353 6971 13419 6974
rect 13486 6972 13492 6974
rect 13556 6972 13562 7036
rect 13629 6898 13695 6901
rect 14958 6898 14964 6900
rect 12160 6896 14964 6898
rect 12160 6840 13634 6896
rect 13690 6840 14964 6896
rect 12160 6838 14964 6840
rect 13629 6835 13695 6838
rect 14958 6836 14964 6838
rect 15028 6836 15034 6900
rect 2405 6762 2471 6765
rect 11237 6762 11303 6765
rect 14641 6762 14707 6765
rect 2405 6760 14707 6762
rect 2405 6704 2410 6760
rect 2466 6704 11242 6760
rect 11298 6704 14646 6760
rect 14702 6704 14707 6760
rect 2405 6702 14707 6704
rect 2405 6699 2471 6702
rect 11237 6699 11303 6702
rect 14641 6699 14707 6702
rect 14917 6764 14983 6765
rect 14917 6760 14964 6764
rect 15028 6762 15034 6764
rect 14917 6704 14922 6760
rect 14917 6700 14964 6704
rect 15028 6702 15074 6762
rect 15028 6700 15034 6702
rect 14917 6699 14983 6700
rect 2221 6626 2287 6629
rect 2589 6626 2655 6629
rect 2221 6624 2655 6626
rect 2221 6568 2226 6624
rect 2282 6568 2594 6624
rect 2650 6568 2655 6624
rect 2221 6566 2655 6568
rect 2221 6563 2287 6566
rect 2589 6563 2655 6566
rect 12750 6564 12756 6628
rect 12820 6626 12826 6628
rect 13854 6626 13860 6628
rect 12820 6566 13860 6626
rect 12820 6564 12826 6566
rect 13854 6564 13860 6566
rect 13924 6626 13930 6628
rect 15510 6626 15516 6628
rect 13924 6566 15516 6626
rect 13924 6564 13930 6566
rect 15510 6564 15516 6566
rect 15580 6564 15586 6628
rect 4692 6560 5012 6561
rect 0 6490 800 6520
rect 4692 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5012 6560
rect 4692 6495 5012 6496
rect 8440 6560 8760 6561
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 6495 8760 6496
rect 12188 6560 12508 6561
rect 12188 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12508 6560
rect 12188 6495 12508 6496
rect 3325 6490 3391 6493
rect 11145 6492 11211 6493
rect 10910 6490 10916 6492
rect 0 6488 3391 6490
rect 0 6432 3330 6488
rect 3386 6432 3391 6488
rect 0 6430 3391 6432
rect 0 6400 800 6430
rect 3325 6427 3391 6430
rect 9032 6430 10916 6490
rect 4889 6354 4955 6357
rect 7465 6354 7531 6357
rect 4889 6352 7531 6354
rect 4889 6296 4894 6352
rect 4950 6296 7470 6352
rect 7526 6296 7531 6352
rect 4889 6294 7531 6296
rect 4889 6291 4955 6294
rect 7465 6291 7531 6294
rect 790 6156 796 6220
rect 860 6218 866 6220
rect 8293 6218 8359 6221
rect 860 6216 8359 6218
rect 860 6160 8298 6216
rect 8354 6160 8359 6216
rect 860 6158 8359 6160
rect 860 6156 866 6158
rect 8293 6155 8359 6158
rect 8845 6218 8911 6221
rect 9032 6218 9092 6430
rect 10910 6428 10916 6430
rect 10980 6428 10986 6492
rect 11094 6490 11100 6492
rect 11054 6430 11100 6490
rect 11164 6488 11211 6492
rect 11206 6432 11211 6488
rect 11094 6428 11100 6430
rect 11164 6428 11211 6432
rect 11278 6428 11284 6492
rect 11348 6490 11354 6492
rect 11513 6490 11579 6493
rect 11348 6488 11579 6490
rect 11348 6432 11518 6488
rect 11574 6432 11579 6488
rect 11348 6430 11579 6432
rect 11348 6428 11354 6430
rect 11145 6427 11211 6428
rect 11513 6427 11579 6430
rect 11697 6490 11763 6493
rect 11973 6490 12039 6493
rect 11697 6488 12039 6490
rect 11697 6432 11702 6488
rect 11758 6432 11978 6488
rect 12034 6432 12039 6488
rect 11697 6430 12039 6432
rect 11697 6427 11763 6430
rect 11973 6427 12039 6430
rect 12750 6428 12756 6492
rect 12820 6490 12826 6492
rect 13077 6490 13143 6493
rect 12820 6488 13143 6490
rect 12820 6432 13082 6488
rect 13138 6432 13143 6488
rect 12820 6430 13143 6432
rect 12820 6428 12826 6430
rect 13077 6427 13143 6430
rect 13854 6428 13860 6492
rect 13924 6490 13930 6492
rect 13997 6490 14063 6493
rect 13924 6488 14063 6490
rect 13924 6432 14002 6488
rect 14058 6432 14063 6488
rect 13924 6430 14063 6432
rect 13924 6428 13930 6430
rect 13997 6427 14063 6430
rect 14457 6490 14523 6493
rect 15561 6490 15627 6493
rect 14457 6488 15627 6490
rect 14457 6432 14462 6488
rect 14518 6432 15566 6488
rect 15622 6432 15627 6488
rect 14457 6430 15627 6432
rect 14457 6427 14523 6430
rect 15561 6427 15627 6430
rect 9990 6292 9996 6356
rect 10060 6354 10066 6356
rect 14457 6354 14523 6357
rect 10060 6352 14523 6354
rect 10060 6296 14462 6352
rect 14518 6296 14523 6352
rect 10060 6294 14523 6296
rect 10060 6292 10066 6294
rect 14457 6291 14523 6294
rect 14825 6354 14891 6357
rect 14825 6352 15716 6354
rect 14825 6296 14830 6352
rect 14886 6296 15716 6352
rect 14825 6294 15716 6296
rect 14825 6291 14891 6294
rect 8845 6216 9092 6218
rect 8845 6160 8850 6216
rect 8906 6160 9092 6216
rect 8845 6158 9092 6160
rect 9397 6218 9463 6221
rect 14825 6218 14891 6221
rect 9397 6216 14891 6218
rect 9397 6160 9402 6216
rect 9458 6160 14830 6216
rect 14886 6160 14891 6216
rect 9397 6158 14891 6160
rect 8845 6155 8911 6158
rect 9397 6155 9463 6158
rect 14825 6155 14891 6158
rect 15656 6085 15716 6294
rect 5349 6082 5415 6085
rect 5574 6082 5580 6084
rect 5349 6080 5580 6082
rect 5349 6024 5354 6080
rect 5410 6024 5580 6080
rect 5349 6022 5580 6024
rect 5349 6019 5415 6022
rect 5574 6020 5580 6022
rect 5644 6020 5650 6084
rect 8109 6082 8175 6085
rect 9949 6082 10015 6085
rect 8109 6080 10015 6082
rect 8109 6024 8114 6080
rect 8170 6024 9954 6080
rect 10010 6024 10015 6080
rect 8109 6022 10015 6024
rect 8109 6019 8175 6022
rect 9949 6019 10015 6022
rect 10777 6082 10843 6085
rect 11053 6084 11119 6085
rect 10910 6082 10916 6084
rect 10777 6080 10916 6082
rect 10777 6024 10782 6080
rect 10838 6024 10916 6080
rect 10777 6022 10916 6024
rect 10777 6019 10843 6022
rect 10910 6020 10916 6022
rect 10980 6020 10986 6084
rect 11053 6080 11100 6084
rect 11164 6082 11170 6084
rect 11053 6024 11058 6080
rect 11053 6020 11100 6024
rect 11164 6022 11210 6082
rect 11164 6020 11170 6022
rect 11278 6020 11284 6084
rect 11348 6082 11354 6084
rect 12801 6082 12867 6085
rect 11348 6080 12867 6082
rect 11348 6024 12806 6080
rect 12862 6024 12867 6080
rect 11348 6022 12867 6024
rect 11348 6020 11354 6022
rect 11053 6019 11119 6020
rect 12801 6019 12867 6022
rect 13261 6082 13327 6085
rect 13445 6082 13511 6085
rect 13261 6080 13511 6082
rect 13261 6024 13266 6080
rect 13322 6024 13450 6080
rect 13506 6024 13511 6080
rect 13261 6022 13511 6024
rect 13261 6019 13327 6022
rect 13445 6019 13511 6022
rect 15653 6080 15719 6085
rect 15653 6024 15658 6080
rect 15714 6024 15719 6080
rect 15653 6019 15719 6024
rect 2818 6016 3138 6017
rect 2818 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3138 6016
rect 2818 5951 3138 5952
rect 6566 6016 6886 6017
rect 6566 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6886 6016
rect 6566 5951 6886 5952
rect 10314 6016 10634 6017
rect 10314 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10634 6016
rect 10314 5951 10634 5952
rect 14062 6016 14382 6017
rect 14062 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14382 6016
rect 14062 5951 14382 5952
rect 4470 5884 4476 5948
rect 4540 5946 4546 5948
rect 4613 5946 4679 5949
rect 4540 5944 4679 5946
rect 4540 5888 4618 5944
rect 4674 5888 4679 5944
rect 4540 5886 4679 5888
rect 4540 5884 4546 5886
rect 4613 5883 4679 5886
rect 7373 5946 7439 5949
rect 7782 5946 7788 5948
rect 7373 5944 7788 5946
rect 7373 5888 7378 5944
rect 7434 5888 7788 5944
rect 7373 5886 7788 5888
rect 7373 5883 7439 5886
rect 7782 5884 7788 5886
rect 7852 5884 7858 5948
rect 7966 5884 7972 5948
rect 8036 5946 8042 5948
rect 10133 5946 10199 5949
rect 8036 5944 10199 5946
rect 8036 5888 10138 5944
rect 10194 5888 10199 5944
rect 8036 5886 10199 5888
rect 8036 5884 8042 5886
rect 10133 5883 10199 5886
rect 10777 5946 10843 5949
rect 11053 5946 11119 5949
rect 13813 5946 13879 5949
rect 10777 5944 13879 5946
rect 10777 5888 10782 5944
rect 10838 5888 11058 5944
rect 11114 5888 13818 5944
rect 13874 5888 13879 5944
rect 10777 5886 13879 5888
rect 10777 5883 10843 5886
rect 11053 5883 11119 5886
rect 13813 5883 13879 5886
rect 14774 5884 14780 5948
rect 14844 5946 14850 5948
rect 14917 5946 14983 5949
rect 14844 5944 15026 5946
rect 14844 5888 14922 5944
rect 14978 5888 15026 5944
rect 14844 5886 15026 5888
rect 14844 5884 14850 5886
rect 14917 5883 15026 5886
rect 1342 5748 1348 5812
rect 1412 5810 1418 5812
rect 4889 5810 4955 5813
rect 1412 5808 4955 5810
rect 1412 5752 4894 5808
rect 4950 5752 4955 5808
rect 1412 5750 4955 5752
rect 1412 5748 1418 5750
rect 4889 5747 4955 5750
rect 5073 5810 5139 5813
rect 12893 5810 12959 5813
rect 13353 5812 13419 5813
rect 5073 5808 12959 5810
rect 5073 5752 5078 5808
rect 5134 5752 12898 5808
rect 12954 5752 12959 5808
rect 5073 5750 12959 5752
rect 5073 5747 5139 5750
rect 12893 5747 12959 5750
rect 13302 5748 13308 5812
rect 13372 5810 13419 5812
rect 14825 5810 14891 5813
rect 13372 5808 14891 5810
rect 13414 5752 14830 5808
rect 14886 5752 14891 5808
rect 13372 5750 14891 5752
rect 13372 5748 13419 5750
rect 13353 5747 13419 5748
rect 14825 5747 14891 5750
rect 14966 5677 15026 5883
rect 2313 5676 2379 5677
rect 2262 5674 2268 5676
rect 2222 5614 2268 5674
rect 2332 5672 2379 5676
rect 5533 5674 5599 5677
rect 2374 5616 2379 5672
rect 2262 5612 2268 5614
rect 2332 5612 2379 5616
rect 2313 5611 2379 5612
rect 2730 5672 5599 5674
rect 2730 5616 5538 5672
rect 5594 5616 5599 5672
rect 2730 5614 5599 5616
rect 2129 5538 2195 5541
rect 2730 5538 2790 5614
rect 5533 5611 5599 5614
rect 6126 5612 6132 5676
rect 6196 5674 6202 5676
rect 9213 5674 9279 5677
rect 6196 5672 9279 5674
rect 6196 5616 9218 5672
rect 9274 5616 9279 5672
rect 6196 5614 9279 5616
rect 6196 5612 6202 5614
rect 9213 5611 9279 5614
rect 9622 5612 9628 5676
rect 9692 5674 9698 5676
rect 10174 5674 10180 5676
rect 9692 5614 10180 5674
rect 9692 5612 9698 5614
rect 10174 5612 10180 5614
rect 10244 5612 10250 5676
rect 10685 5674 10751 5677
rect 11237 5674 11303 5677
rect 10685 5672 11303 5674
rect 10685 5616 10690 5672
rect 10746 5616 11242 5672
rect 11298 5616 11303 5672
rect 10685 5614 11303 5616
rect 10685 5611 10751 5614
rect 11237 5611 11303 5614
rect 11789 5674 11855 5677
rect 12341 5674 12407 5677
rect 14181 5674 14247 5677
rect 11789 5672 14247 5674
rect 11789 5616 11794 5672
rect 11850 5616 12346 5672
rect 12402 5616 14186 5672
rect 14242 5616 14247 5672
rect 11789 5614 14247 5616
rect 11789 5611 11855 5614
rect 12341 5611 12407 5614
rect 14181 5611 14247 5614
rect 14917 5672 15026 5677
rect 14917 5616 14922 5672
rect 14978 5616 15026 5672
rect 14917 5614 15026 5616
rect 14917 5611 14983 5614
rect 2129 5536 2790 5538
rect 2129 5480 2134 5536
rect 2190 5480 2790 5536
rect 2129 5478 2790 5480
rect 9949 5538 10015 5541
rect 10593 5538 10659 5541
rect 10726 5538 10732 5540
rect 9949 5536 10732 5538
rect 9949 5480 9954 5536
rect 10010 5480 10598 5536
rect 10654 5480 10732 5536
rect 9949 5478 10732 5480
rect 2129 5475 2195 5478
rect 9949 5475 10015 5478
rect 10593 5475 10659 5478
rect 10726 5476 10732 5478
rect 10796 5476 10802 5540
rect 13077 5538 13143 5541
rect 13302 5538 13308 5540
rect 11102 5478 12128 5538
rect 4692 5472 5012 5473
rect 0 5402 800 5432
rect 4692 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5012 5472
rect 4692 5407 5012 5408
rect 8440 5472 8760 5473
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 5407 8760 5408
rect 3693 5402 3759 5405
rect 0 5400 3759 5402
rect 0 5344 3698 5400
rect 3754 5344 3759 5400
rect 0 5342 3759 5344
rect 0 5312 800 5342
rect 3693 5339 3759 5342
rect 5206 5340 5212 5404
rect 5276 5402 5282 5404
rect 11102 5402 11162 5478
rect 5276 5342 7114 5402
rect 5276 5340 5282 5342
rect 3785 5266 3851 5269
rect 6913 5266 6979 5269
rect 3785 5264 6979 5266
rect 3785 5208 3790 5264
rect 3846 5208 6918 5264
rect 6974 5208 6979 5264
rect 3785 5206 6979 5208
rect 7054 5266 7114 5342
rect 8848 5342 11162 5402
rect 11237 5400 11303 5405
rect 11605 5404 11671 5405
rect 11605 5402 11652 5404
rect 11237 5344 11242 5400
rect 11298 5344 11303 5400
rect 8848 5266 8908 5342
rect 11237 5339 11303 5344
rect 11560 5400 11652 5402
rect 11560 5344 11610 5400
rect 11560 5342 11652 5344
rect 11605 5340 11652 5342
rect 11716 5340 11722 5404
rect 11605 5339 11671 5340
rect 7054 5206 8908 5266
rect 10317 5266 10383 5269
rect 10317 5264 10656 5266
rect 10317 5208 10322 5264
rect 10378 5208 10656 5264
rect 10317 5206 10656 5208
rect 3785 5203 3851 5206
rect 6913 5203 6979 5206
rect 10317 5203 10383 5206
rect 3693 5130 3759 5133
rect 7097 5130 7163 5133
rect 3693 5128 9920 5130
rect 3693 5072 3698 5128
rect 3754 5072 7102 5128
rect 7158 5072 9920 5128
rect 3693 5070 9920 5072
rect 3693 5067 3759 5070
rect 7097 5067 7163 5070
rect 9860 4997 9920 5070
rect 10174 5068 10180 5132
rect 10244 5130 10250 5132
rect 10409 5130 10475 5133
rect 10244 5128 10475 5130
rect 10244 5072 10414 5128
rect 10470 5072 10475 5128
rect 10244 5070 10475 5072
rect 10596 5130 10656 5206
rect 10726 5204 10732 5268
rect 10796 5266 10802 5268
rect 11094 5266 11100 5268
rect 10796 5206 11100 5266
rect 10796 5204 10802 5206
rect 11094 5204 11100 5206
rect 11164 5204 11170 5268
rect 11240 5266 11300 5339
rect 12068 5300 12128 5478
rect 13077 5536 13308 5538
rect 13077 5480 13082 5536
rect 13138 5480 13308 5536
rect 13077 5478 13308 5480
rect 13077 5475 13143 5478
rect 13302 5476 13308 5478
rect 13372 5476 13378 5540
rect 13670 5476 13676 5540
rect 13740 5538 13746 5540
rect 14273 5538 14339 5541
rect 14825 5540 14891 5541
rect 13740 5536 14339 5538
rect 13740 5480 14278 5536
rect 14334 5480 14339 5536
rect 13740 5478 14339 5480
rect 13740 5476 13746 5478
rect 14273 5475 14339 5478
rect 14774 5476 14780 5540
rect 14844 5538 14891 5540
rect 14844 5536 14936 5538
rect 14886 5480 14936 5536
rect 14844 5478 14936 5480
rect 14844 5476 14891 5478
rect 14825 5475 14891 5476
rect 12188 5472 12508 5473
rect 12188 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12508 5472
rect 12188 5407 12508 5408
rect 12750 5340 12756 5404
rect 12820 5402 12826 5404
rect 14365 5402 14431 5405
rect 12820 5400 14431 5402
rect 12820 5344 14370 5400
rect 14426 5344 14431 5400
rect 12820 5342 14431 5344
rect 12820 5340 12826 5342
rect 14365 5339 14431 5342
rect 12068 5269 12266 5300
rect 11881 5266 11947 5269
rect 11240 5264 11947 5266
rect 11240 5208 11886 5264
rect 11942 5208 11947 5264
rect 12068 5264 12315 5269
rect 12068 5240 12254 5264
rect 11240 5206 11947 5208
rect 12206 5208 12254 5240
rect 12310 5208 12315 5264
rect 12206 5206 12315 5208
rect 11881 5203 11947 5206
rect 12249 5203 12315 5206
rect 12433 5266 12499 5269
rect 15101 5266 15167 5269
rect 12433 5264 15167 5266
rect 12433 5208 12438 5264
rect 12494 5208 15106 5264
rect 15162 5208 15167 5264
rect 12433 5206 15167 5208
rect 12433 5203 12499 5206
rect 15101 5203 15167 5206
rect 15469 5268 15535 5269
rect 15469 5264 15516 5268
rect 15580 5266 15586 5268
rect 15469 5208 15474 5264
rect 15469 5204 15516 5208
rect 15580 5206 15626 5266
rect 15580 5204 15586 5206
rect 15469 5203 15535 5204
rect 14089 5130 14155 5133
rect 14273 5130 14339 5133
rect 10596 5128 14339 5130
rect 10596 5072 14094 5128
rect 14150 5072 14278 5128
rect 14334 5072 14339 5128
rect 10596 5070 14339 5072
rect 10244 5068 10250 5070
rect 10409 5067 10475 5070
rect 14089 5067 14155 5070
rect 14273 5067 14339 5070
rect 14457 5130 14523 5133
rect 15142 5130 15148 5132
rect 14457 5128 15148 5130
rect 14457 5072 14462 5128
rect 14518 5072 15148 5128
rect 14457 5070 15148 5072
rect 14457 5067 14523 5070
rect 15142 5068 15148 5070
rect 15212 5068 15218 5132
rect 7281 4994 7347 4997
rect 7465 4994 7531 4997
rect 7281 4992 7531 4994
rect 7281 4936 7286 4992
rect 7342 4936 7470 4992
rect 7526 4936 7531 4992
rect 7281 4934 7531 4936
rect 7281 4931 7347 4934
rect 7465 4931 7531 4934
rect 8017 4994 8083 4997
rect 9622 4994 9628 4996
rect 8017 4992 9628 4994
rect 8017 4936 8022 4992
rect 8078 4936 9628 4992
rect 8017 4934 9628 4936
rect 8017 4931 8083 4934
rect 9622 4932 9628 4934
rect 9692 4932 9698 4996
rect 9857 4992 9923 4997
rect 9857 4936 9862 4992
rect 9918 4936 9923 4992
rect 9857 4931 9923 4936
rect 10961 4994 11027 4997
rect 11094 4994 11100 4996
rect 10961 4992 11100 4994
rect 10961 4936 10966 4992
rect 11022 4936 11100 4992
rect 10961 4934 11100 4936
rect 10961 4931 11027 4934
rect 11094 4932 11100 4934
rect 11164 4932 11170 4996
rect 11421 4994 11487 4997
rect 11973 4994 12039 4997
rect 12617 4994 12683 4997
rect 13486 4994 13492 4996
rect 11421 4992 11898 4994
rect 11421 4936 11426 4992
rect 11482 4936 11898 4992
rect 11421 4934 11898 4936
rect 11421 4931 11487 4934
rect 2818 4928 3138 4929
rect 2818 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3138 4928
rect 2818 4863 3138 4864
rect 6566 4928 6886 4929
rect 6566 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6886 4928
rect 6566 4863 6886 4864
rect 10314 4928 10634 4929
rect 10314 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10634 4928
rect 10314 4863 10634 4864
rect 7097 4858 7163 4861
rect 8477 4858 8543 4861
rect 7097 4856 8543 4858
rect 7097 4800 7102 4856
rect 7158 4800 8482 4856
rect 8538 4800 8543 4856
rect 7097 4798 8543 4800
rect 7097 4795 7163 4798
rect 8477 4795 8543 4798
rect 9622 4796 9628 4860
rect 9692 4858 9698 4860
rect 9765 4858 9831 4861
rect 9692 4856 9831 4858
rect 9692 4800 9770 4856
rect 9826 4800 9831 4856
rect 9692 4798 9831 4800
rect 9692 4796 9698 4798
rect 9765 4795 9831 4798
rect 10869 4858 10935 4861
rect 11605 4858 11671 4861
rect 10869 4856 11671 4858
rect 10869 4800 10874 4856
rect 10930 4800 11610 4856
rect 11666 4800 11671 4856
rect 10869 4798 11671 4800
rect 11838 4858 11898 4934
rect 11973 4992 13492 4994
rect 11973 4936 11978 4992
rect 12034 4936 12622 4992
rect 12678 4936 13492 4992
rect 11973 4934 13492 4936
rect 11973 4931 12039 4934
rect 12617 4931 12683 4934
rect 13486 4932 13492 4934
rect 13556 4932 13562 4996
rect 14062 4928 14382 4929
rect 14062 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14382 4928
rect 14062 4863 14382 4864
rect 13537 4858 13603 4861
rect 11838 4856 13603 4858
rect 11838 4800 13542 4856
rect 13598 4800 13603 4856
rect 11838 4798 13603 4800
rect 10869 4795 10935 4798
rect 11605 4795 11671 4798
rect 13537 4795 13603 4798
rect 974 4660 980 4724
rect 1044 4722 1050 4724
rect 1577 4722 1643 4725
rect 1044 4720 1643 4722
rect 1044 4664 1582 4720
rect 1638 4664 1643 4720
rect 1044 4662 1643 4664
rect 1044 4660 1050 4662
rect 1577 4659 1643 4662
rect 2957 4722 3023 4725
rect 9213 4722 9279 4725
rect 12249 4722 12315 4725
rect 2957 4720 12315 4722
rect 2957 4664 2962 4720
rect 3018 4664 9218 4720
rect 9274 4664 12254 4720
rect 12310 4664 12315 4720
rect 2957 4662 12315 4664
rect 2957 4659 3023 4662
rect 9213 4659 9279 4662
rect 12249 4659 12315 4662
rect 14365 4722 14431 4725
rect 15377 4722 15443 4725
rect 14365 4720 15443 4722
rect 14365 4664 14370 4720
rect 14426 4664 15382 4720
rect 15438 4664 15443 4720
rect 14365 4662 15443 4664
rect 14365 4659 14431 4662
rect 15377 4659 15443 4662
rect 5165 4586 5231 4589
rect 10174 4586 10180 4588
rect 5165 4584 10180 4586
rect 5165 4528 5170 4584
rect 5226 4528 10180 4584
rect 5165 4526 10180 4528
rect 5165 4523 5231 4526
rect 10174 4524 10180 4526
rect 10244 4524 10250 4588
rect 11237 4586 11303 4589
rect 11462 4586 11468 4588
rect 11237 4584 11468 4586
rect 11237 4528 11242 4584
rect 11298 4528 11468 4584
rect 11237 4526 11468 4528
rect 11237 4523 11303 4526
rect 11462 4524 11468 4526
rect 11532 4524 11538 4588
rect 15285 4586 15351 4589
rect 12068 4584 15351 4586
rect 12068 4528 15290 4584
rect 15346 4528 15351 4584
rect 12068 4526 15351 4528
rect 0 4450 800 4480
rect 2221 4450 2287 4453
rect 0 4448 2287 4450
rect 0 4392 2226 4448
rect 2282 4392 2287 4448
rect 0 4390 2287 4392
rect 0 4360 800 4390
rect 2221 4387 2287 4390
rect 2497 4450 2563 4453
rect 3233 4450 3299 4453
rect 3366 4450 3372 4452
rect 2497 4448 3372 4450
rect 2497 4392 2502 4448
rect 2558 4392 3238 4448
rect 3294 4392 3372 4448
rect 2497 4390 3372 4392
rect 2497 4387 2563 4390
rect 3233 4387 3299 4390
rect 3366 4388 3372 4390
rect 3436 4388 3442 4452
rect 5257 4450 5323 4453
rect 8017 4450 8083 4453
rect 5257 4448 8083 4450
rect 5257 4392 5262 4448
rect 5318 4392 8022 4448
rect 8078 4392 8083 4448
rect 5257 4390 8083 4392
rect 5257 4387 5323 4390
rect 8017 4387 8083 4390
rect 8937 4450 9003 4453
rect 12068 4450 12128 4526
rect 15285 4523 15351 4526
rect 8937 4448 12128 4450
rect 8937 4392 8942 4448
rect 8998 4392 12128 4448
rect 8937 4390 12128 4392
rect 8937 4387 9003 4390
rect 12750 4388 12756 4452
rect 12820 4450 12826 4452
rect 13261 4450 13327 4453
rect 12820 4448 13327 4450
rect 12820 4392 13266 4448
rect 13322 4392 13327 4448
rect 12820 4390 13327 4392
rect 12820 4388 12826 4390
rect 13261 4387 13327 4390
rect 4692 4384 5012 4385
rect 4692 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5012 4384
rect 4692 4319 5012 4320
rect 8440 4384 8760 4385
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 4319 8760 4320
rect 12188 4384 12508 4385
rect 12188 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12508 4384
rect 12188 4319 12508 4320
rect 7598 4252 7604 4316
rect 7668 4314 7674 4316
rect 8201 4314 8267 4317
rect 7668 4312 8267 4314
rect 7668 4256 8206 4312
rect 8262 4256 8267 4312
rect 7668 4254 8267 4256
rect 7668 4252 7674 4254
rect 8201 4251 8267 4254
rect 9397 4314 9463 4317
rect 9949 4314 10015 4317
rect 9397 4312 10015 4314
rect 9397 4256 9402 4312
rect 9458 4256 9954 4312
rect 10010 4256 10015 4312
rect 9397 4254 10015 4256
rect 9397 4251 9463 4254
rect 9949 4251 10015 4254
rect 10225 4314 10291 4317
rect 11881 4314 11947 4317
rect 15326 4314 15332 4316
rect 10225 4312 11947 4314
rect 10225 4256 10230 4312
rect 10286 4256 11886 4312
rect 11942 4256 11947 4312
rect 10225 4254 11947 4256
rect 10225 4251 10291 4254
rect 11881 4251 11947 4254
rect 12712 4254 15332 4314
rect 4153 4178 4219 4181
rect 7005 4178 7071 4181
rect 4153 4176 7071 4178
rect 4153 4120 4158 4176
rect 4214 4120 7010 4176
rect 7066 4120 7071 4176
rect 4153 4118 7071 4120
rect 4153 4115 4219 4118
rect 7005 4115 7071 4118
rect 7741 4178 7807 4181
rect 10910 4178 10916 4180
rect 7741 4176 10916 4178
rect 7741 4120 7746 4176
rect 7802 4120 10916 4176
rect 7741 4118 10916 4120
rect 7741 4115 7807 4118
rect 10910 4116 10916 4118
rect 10980 4116 10986 4180
rect 11462 4116 11468 4180
rect 11532 4178 11538 4180
rect 11605 4178 11671 4181
rect 11532 4176 11671 4178
rect 11532 4120 11610 4176
rect 11666 4120 11671 4176
rect 11532 4118 11671 4120
rect 11532 4116 11538 4118
rect 11605 4115 11671 4118
rect 12341 4178 12407 4181
rect 12566 4178 12572 4180
rect 12341 4176 12572 4178
rect 12341 4120 12346 4176
rect 12402 4120 12572 4176
rect 12341 4118 12572 4120
rect 12341 4115 12407 4118
rect 12566 4116 12572 4118
rect 12636 4116 12642 4180
rect 1526 3980 1532 4044
rect 1596 4042 1602 4044
rect 1669 4042 1735 4045
rect 1596 4040 1735 4042
rect 1596 3984 1674 4040
rect 1730 3984 1735 4040
rect 1596 3982 1735 3984
rect 1596 3980 1602 3982
rect 1669 3979 1735 3982
rect 5390 3980 5396 4044
rect 5460 4042 5466 4044
rect 6545 4042 6611 4045
rect 5460 4040 6611 4042
rect 5460 3984 6550 4040
rect 6606 3984 6611 4040
rect 5460 3982 6611 3984
rect 5460 3980 5466 3982
rect 6545 3979 6611 3982
rect 6821 4042 6887 4045
rect 7046 4042 7052 4044
rect 6821 4040 7052 4042
rect 6821 3984 6826 4040
rect 6882 3984 7052 4040
rect 6821 3982 7052 3984
rect 6821 3979 6887 3982
rect 7046 3980 7052 3982
rect 7116 3980 7122 4044
rect 7465 4042 7531 4045
rect 7741 4042 7807 4045
rect 7465 4040 7807 4042
rect 7465 3984 7470 4040
rect 7526 3984 7746 4040
rect 7802 3984 7807 4040
rect 7465 3982 7807 3984
rect 7465 3979 7531 3982
rect 7741 3979 7807 3982
rect 8109 4042 8175 4045
rect 9581 4042 9647 4045
rect 8109 4040 9647 4042
rect 8109 3984 8114 4040
rect 8170 3984 9586 4040
rect 9642 3984 9647 4040
rect 8109 3982 9647 3984
rect 8109 3979 8175 3982
rect 9581 3979 9647 3982
rect 10317 4042 10383 4045
rect 10869 4042 10935 4045
rect 12433 4042 12499 4045
rect 12712 4042 12772 4254
rect 15326 4252 15332 4254
rect 15396 4252 15402 4316
rect 13302 4116 13308 4180
rect 13372 4178 13378 4180
rect 13629 4178 13695 4181
rect 13372 4176 13695 4178
rect 13372 4120 13634 4176
rect 13690 4120 13695 4176
rect 13372 4118 13695 4120
rect 13372 4116 13378 4118
rect 13629 4115 13695 4118
rect 14273 4178 14339 4181
rect 16297 4178 16363 4181
rect 14273 4176 16363 4178
rect 14273 4120 14278 4176
rect 14334 4120 16302 4176
rect 16358 4120 16363 4176
rect 14273 4118 16363 4120
rect 14273 4115 14339 4118
rect 16297 4115 16363 4118
rect 10317 4040 10794 4042
rect 10317 3984 10322 4040
rect 10378 3984 10794 4040
rect 10317 3982 10794 3984
rect 10317 3979 10383 3982
rect 10734 3906 10794 3982
rect 10869 4040 12772 4042
rect 10869 3984 10874 4040
rect 10930 3984 12438 4040
rect 12494 3984 12772 4040
rect 10869 3982 12772 3984
rect 12985 4042 13051 4045
rect 14089 4042 14155 4045
rect 14917 4044 14983 4045
rect 14917 4042 14964 4044
rect 12985 4040 14155 4042
rect 12985 3984 12990 4040
rect 13046 3984 14094 4040
rect 14150 3984 14155 4040
rect 12985 3982 14155 3984
rect 14872 4040 14964 4042
rect 14872 3984 14922 4040
rect 14872 3982 14964 3984
rect 10869 3979 10935 3982
rect 12433 3979 12499 3982
rect 12985 3979 13051 3982
rect 14089 3979 14155 3982
rect 14917 3980 14964 3982
rect 15028 3980 15034 4044
rect 14917 3979 14983 3980
rect 13721 3906 13787 3909
rect 10734 3904 13787 3906
rect 10734 3848 13726 3904
rect 13782 3848 13787 3904
rect 10734 3846 13787 3848
rect 13721 3843 13787 3846
rect 2818 3840 3138 3841
rect 2818 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3138 3840
rect 2818 3775 3138 3776
rect 6566 3840 6886 3841
rect 6566 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6886 3840
rect 6566 3775 6886 3776
rect 10314 3840 10634 3841
rect 10314 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10634 3840
rect 10314 3775 10634 3776
rect 14062 3840 14382 3841
rect 14062 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14382 3840
rect 14062 3775 14382 3776
rect 7373 3770 7439 3773
rect 8150 3770 8156 3772
rect 7373 3768 8156 3770
rect 7373 3712 7378 3768
rect 7434 3712 8156 3768
rect 7373 3710 8156 3712
rect 7373 3707 7439 3710
rect 8150 3708 8156 3710
rect 8220 3770 8226 3772
rect 9397 3770 9463 3773
rect 8220 3768 9463 3770
rect 8220 3712 9402 3768
rect 9458 3712 9463 3768
rect 8220 3710 9463 3712
rect 8220 3708 8226 3710
rect 9397 3707 9463 3710
rect 9673 3770 9739 3773
rect 9990 3770 9996 3772
rect 9673 3768 9996 3770
rect 9673 3712 9678 3768
rect 9734 3712 9996 3768
rect 9673 3710 9996 3712
rect 9673 3707 9739 3710
rect 9990 3708 9996 3710
rect 10060 3708 10066 3772
rect 12014 3708 12020 3772
rect 12084 3770 12090 3772
rect 12084 3710 13876 3770
rect 12084 3708 12090 3710
rect 3233 3634 3299 3637
rect 8753 3634 8819 3637
rect 3233 3632 8819 3634
rect 3233 3576 3238 3632
rect 3294 3576 8758 3632
rect 8814 3576 8819 3632
rect 3233 3574 8819 3576
rect 3233 3571 3299 3574
rect 8753 3571 8819 3574
rect 9254 3572 9260 3636
rect 9324 3634 9330 3636
rect 9857 3634 9923 3637
rect 9324 3632 9923 3634
rect 9324 3576 9862 3632
rect 9918 3576 9923 3632
rect 9324 3574 9923 3576
rect 9324 3572 9330 3574
rect 9857 3571 9923 3574
rect 10225 3634 10291 3637
rect 13445 3634 13511 3637
rect 10225 3632 13511 3634
rect 10225 3576 10230 3632
rect 10286 3576 13450 3632
rect 13506 3576 13511 3632
rect 10225 3574 13511 3576
rect 10225 3571 10291 3574
rect 13445 3571 13511 3574
rect 0 3498 800 3528
rect 3601 3498 3667 3501
rect 0 3496 3667 3498
rect 0 3440 3606 3496
rect 3662 3440 3667 3496
rect 0 3438 3667 3440
rect 0 3408 800 3438
rect 3601 3435 3667 3438
rect 5625 3498 5691 3501
rect 10501 3498 10567 3501
rect 11462 3498 11468 3500
rect 5625 3496 10196 3498
rect 5625 3440 5630 3496
rect 5686 3440 10196 3496
rect 5625 3438 10196 3440
rect 5625 3435 5691 3438
rect 2589 3362 2655 3365
rect 3969 3362 4035 3365
rect 2589 3360 4035 3362
rect 2589 3304 2594 3360
rect 2650 3304 3974 3360
rect 4030 3304 4035 3360
rect 2589 3302 4035 3304
rect 2589 3299 2655 3302
rect 3969 3299 4035 3302
rect 5809 3362 5875 3365
rect 7373 3362 7439 3365
rect 5809 3360 7439 3362
rect 5809 3304 5814 3360
rect 5870 3304 7378 3360
rect 7434 3304 7439 3360
rect 5809 3302 7439 3304
rect 10136 3362 10196 3438
rect 10501 3496 11468 3498
rect 10501 3440 10506 3496
rect 10562 3440 11468 3496
rect 10501 3438 11468 3440
rect 10501 3435 10567 3438
rect 11462 3436 11468 3438
rect 11532 3436 11538 3500
rect 11646 3436 11652 3500
rect 11716 3498 11722 3500
rect 12709 3498 12775 3501
rect 11716 3496 12775 3498
rect 11716 3440 12714 3496
rect 12770 3440 12775 3496
rect 11716 3438 12775 3440
rect 11716 3436 11722 3438
rect 12709 3435 12775 3438
rect 13077 3498 13143 3501
rect 13537 3498 13603 3501
rect 13077 3496 13603 3498
rect 13077 3440 13082 3496
rect 13138 3440 13542 3496
rect 13598 3440 13603 3496
rect 13077 3438 13603 3440
rect 13077 3435 13143 3438
rect 13537 3435 13603 3438
rect 11789 3362 11855 3365
rect 10136 3360 11855 3362
rect 10136 3304 11794 3360
rect 11850 3304 11855 3360
rect 10136 3302 11855 3304
rect 13816 3362 13876 3710
rect 16400 3362 17200 3392
rect 13816 3302 17200 3362
rect 5809 3299 5875 3302
rect 7373 3299 7439 3302
rect 11789 3299 11855 3302
rect 4692 3296 5012 3297
rect 4692 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5012 3296
rect 4692 3231 5012 3232
rect 8440 3296 8760 3297
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 3231 8760 3232
rect 12188 3296 12508 3297
rect 12188 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12508 3296
rect 16400 3272 17200 3302
rect 12188 3231 12508 3232
rect 2773 3226 2839 3229
rect 4245 3226 4311 3229
rect 5901 3228 5967 3229
rect 5901 3226 5948 3228
rect 2773 3224 4311 3226
rect 2773 3168 2778 3224
rect 2834 3168 4250 3224
rect 4306 3168 4311 3224
rect 2773 3166 4311 3168
rect 5856 3224 5948 3226
rect 5856 3168 5906 3224
rect 5856 3166 5948 3168
rect 2773 3163 2839 3166
rect 4245 3163 4311 3166
rect 5901 3164 5948 3166
rect 6012 3164 6018 3228
rect 7230 3164 7236 3228
rect 7300 3226 7306 3228
rect 7465 3226 7531 3229
rect 7300 3224 7531 3226
rect 7300 3168 7470 3224
rect 7526 3168 7531 3224
rect 7300 3166 7531 3168
rect 7300 3164 7306 3166
rect 5901 3163 5967 3164
rect 7465 3163 7531 3166
rect 9990 3164 9996 3228
rect 10060 3226 10066 3228
rect 10961 3226 11027 3229
rect 10060 3224 11027 3226
rect 10060 3168 10966 3224
rect 11022 3168 11027 3224
rect 10060 3166 11027 3168
rect 10060 3164 10066 3166
rect 10961 3163 11027 3166
rect 11237 3224 11303 3229
rect 11237 3168 11242 3224
rect 11298 3168 11303 3224
rect 11237 3163 11303 3168
rect 11462 3164 11468 3228
rect 11532 3226 11538 3228
rect 11789 3226 11855 3229
rect 13486 3226 13492 3228
rect 11532 3224 11855 3226
rect 11532 3168 11794 3224
rect 11850 3168 11855 3224
rect 11532 3166 11855 3168
rect 11532 3164 11538 3166
rect 11789 3163 11855 3166
rect 13172 3166 13492 3226
rect 2446 3028 2452 3092
rect 2516 3090 2522 3092
rect 6361 3090 6427 3093
rect 2516 3088 6427 3090
rect 2516 3032 6366 3088
rect 6422 3032 6427 3088
rect 2516 3030 6427 3032
rect 2516 3028 2522 3030
rect 6361 3027 6427 3030
rect 8109 3090 8175 3093
rect 9213 3090 9279 3093
rect 10409 3090 10475 3093
rect 8109 3088 9092 3090
rect 8109 3032 8114 3088
rect 8170 3032 9092 3088
rect 8109 3030 9092 3032
rect 8109 3027 8175 3030
rect 2313 2954 2379 2957
rect 6269 2954 6335 2957
rect 7465 2954 7531 2957
rect 2313 2952 7531 2954
rect 2313 2896 2318 2952
rect 2374 2896 6274 2952
rect 6330 2896 7470 2952
rect 7526 2896 7531 2952
rect 2313 2894 7531 2896
rect 2313 2891 2379 2894
rect 6269 2891 6335 2894
rect 7465 2891 7531 2894
rect 8753 2954 8819 2957
rect 8886 2954 8892 2956
rect 8753 2952 8892 2954
rect 8753 2896 8758 2952
rect 8814 2896 8892 2952
rect 8753 2894 8892 2896
rect 8753 2891 8819 2894
rect 8886 2892 8892 2894
rect 8956 2892 8962 2956
rect 9032 2954 9092 3030
rect 9213 3088 10475 3090
rect 9213 3032 9218 3088
rect 9274 3032 10414 3088
rect 10470 3032 10475 3088
rect 9213 3030 10475 3032
rect 9213 3027 9279 3030
rect 10409 3027 10475 3030
rect 10685 3090 10751 3093
rect 11240 3090 11300 3163
rect 10685 3088 11300 3090
rect 10685 3032 10690 3088
rect 10746 3032 11300 3088
rect 10685 3030 11300 3032
rect 11697 3090 11763 3093
rect 12157 3090 12223 3093
rect 11697 3088 12223 3090
rect 11697 3032 11702 3088
rect 11758 3032 12162 3088
rect 12218 3032 12223 3088
rect 11697 3030 12223 3032
rect 10685 3027 10751 3030
rect 11697 3027 11763 3030
rect 12157 3027 12223 3030
rect 12433 3090 12499 3093
rect 12934 3090 12940 3092
rect 12433 3088 12940 3090
rect 12433 3032 12438 3088
rect 12494 3032 12940 3088
rect 12433 3030 12940 3032
rect 12433 3027 12499 3030
rect 12934 3028 12940 3030
rect 13004 3028 13010 3092
rect 9622 2954 9628 2956
rect 9032 2894 9628 2954
rect 9622 2892 9628 2894
rect 9692 2954 9698 2956
rect 10133 2954 10199 2957
rect 9692 2952 10199 2954
rect 9692 2896 10138 2952
rect 10194 2896 10199 2952
rect 9692 2894 10199 2896
rect 9692 2892 9698 2894
rect 10133 2891 10199 2894
rect 10593 2954 10659 2957
rect 10593 2952 11208 2954
rect 10593 2896 10598 2952
rect 10654 2896 11208 2952
rect 10593 2894 11208 2896
rect 10593 2891 10659 2894
rect 2129 2818 2195 2821
rect 2313 2818 2379 2821
rect 2129 2816 2379 2818
rect 2129 2760 2134 2816
rect 2190 2760 2318 2816
rect 2374 2760 2379 2816
rect 2129 2758 2379 2760
rect 2129 2755 2195 2758
rect 2313 2755 2379 2758
rect 4470 2756 4476 2820
rect 4540 2818 4546 2820
rect 4705 2818 4771 2821
rect 4540 2816 4771 2818
rect 4540 2760 4710 2816
rect 4766 2760 4771 2816
rect 4540 2758 4771 2760
rect 4540 2756 4546 2758
rect 4705 2755 4771 2758
rect 5533 2818 5599 2821
rect 6085 2818 6151 2821
rect 10777 2820 10843 2821
rect 5533 2816 6151 2818
rect 5533 2760 5538 2816
rect 5594 2760 6090 2816
rect 6146 2760 6151 2816
rect 5533 2758 6151 2760
rect 5533 2755 5599 2758
rect 6085 2755 6151 2758
rect 7414 2756 7420 2820
rect 7484 2818 7490 2820
rect 9990 2818 9996 2820
rect 7484 2758 9996 2818
rect 7484 2756 7490 2758
rect 9990 2756 9996 2758
rect 10060 2756 10066 2820
rect 10726 2756 10732 2820
rect 10796 2818 10843 2820
rect 11148 2818 11208 2894
rect 13172 2818 13232 3166
rect 13486 3164 13492 3166
rect 13556 3226 13562 3228
rect 14825 3226 14891 3229
rect 13556 3224 14891 3226
rect 13556 3168 14830 3224
rect 14886 3168 14891 3224
rect 13556 3166 14891 3168
rect 13556 3164 13562 3166
rect 14825 3163 14891 3166
rect 15142 3090 15148 3092
rect 10796 2816 10888 2818
rect 10838 2760 10888 2816
rect 10796 2758 10888 2760
rect 11148 2758 13232 2818
rect 13310 3030 15148 3090
rect 10796 2756 10843 2758
rect 10777 2755 10843 2756
rect 2818 2752 3138 2753
rect 2818 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3138 2752
rect 2818 2687 3138 2688
rect 6566 2752 6886 2753
rect 6566 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6886 2752
rect 6566 2687 6886 2688
rect 10314 2752 10634 2753
rect 10314 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10634 2752
rect 10314 2687 10634 2688
rect 1894 2620 1900 2684
rect 1964 2682 1970 2684
rect 4521 2682 4587 2685
rect 5206 2682 5212 2684
rect 1964 2622 2698 2682
rect 1964 2620 1970 2622
rect 1342 2484 1348 2548
rect 1412 2546 1418 2548
rect 2037 2546 2103 2549
rect 2313 2548 2379 2549
rect 1412 2544 2103 2546
rect 1412 2488 2042 2544
rect 2098 2488 2103 2544
rect 1412 2486 2103 2488
rect 1412 2484 1418 2486
rect 2037 2483 2103 2486
rect 2262 2484 2268 2548
rect 2332 2546 2379 2548
rect 2638 2546 2698 2622
rect 4521 2680 5212 2682
rect 4521 2624 4526 2680
rect 4582 2624 5212 2680
rect 4521 2622 5212 2624
rect 4521 2619 4587 2622
rect 5206 2620 5212 2622
rect 5276 2620 5282 2684
rect 5901 2682 5967 2685
rect 6310 2682 6316 2684
rect 5901 2680 6316 2682
rect 5901 2624 5906 2680
rect 5962 2624 6316 2680
rect 5901 2622 6316 2624
rect 5901 2619 5967 2622
rect 6310 2620 6316 2622
rect 6380 2620 6386 2684
rect 7465 2682 7531 2685
rect 8293 2682 8359 2685
rect 7465 2680 8359 2682
rect 7465 2624 7470 2680
rect 7526 2624 8298 2680
rect 8354 2624 8359 2680
rect 7465 2622 8359 2624
rect 7465 2619 7531 2622
rect 8293 2619 8359 2622
rect 8753 2682 8819 2685
rect 9070 2682 9076 2684
rect 8753 2680 9076 2682
rect 8753 2624 8758 2680
rect 8814 2624 9076 2680
rect 8753 2622 9076 2624
rect 8753 2619 8819 2622
rect 9070 2620 9076 2622
rect 9140 2620 9146 2684
rect 11053 2682 11119 2685
rect 13310 2682 13370 3030
rect 15142 3028 15148 3030
rect 15212 3028 15218 3092
rect 14590 2954 14596 2956
rect 13862 2894 14596 2954
rect 13862 2821 13922 2894
rect 14590 2892 14596 2894
rect 14660 2892 14666 2956
rect 13813 2816 13922 2821
rect 13813 2760 13818 2816
rect 13874 2760 13922 2816
rect 13813 2758 13922 2760
rect 13813 2755 13879 2758
rect 14062 2752 14382 2753
rect 14062 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14382 2752
rect 14062 2687 14382 2688
rect 11053 2680 13370 2682
rect 11053 2624 11058 2680
rect 11114 2624 13370 2680
rect 11053 2622 13370 2624
rect 11053 2619 11119 2622
rect 5441 2546 5507 2549
rect 5809 2548 5875 2549
rect 2332 2544 2424 2546
rect 2374 2488 2424 2544
rect 2332 2486 2424 2488
rect 2638 2544 5507 2546
rect 2638 2488 5446 2544
rect 5502 2488 5507 2544
rect 2638 2486 5507 2488
rect 2332 2484 2379 2486
rect 2313 2483 2379 2484
rect 5441 2483 5507 2486
rect 5758 2484 5764 2548
rect 5828 2546 5875 2548
rect 6821 2546 6887 2549
rect 7230 2546 7236 2548
rect 5828 2544 5920 2546
rect 5870 2488 5920 2544
rect 5828 2486 5920 2488
rect 6821 2544 7236 2546
rect 6821 2488 6826 2544
rect 6882 2488 7236 2544
rect 6821 2486 7236 2488
rect 5828 2484 5875 2486
rect 5809 2483 5875 2484
rect 6821 2483 6887 2486
rect 7230 2484 7236 2486
rect 7300 2484 7306 2548
rect 8385 2546 8451 2549
rect 9305 2548 9371 2549
rect 9254 2546 9260 2548
rect 8385 2544 9260 2546
rect 9324 2546 9371 2548
rect 9324 2544 9416 2546
rect 8385 2488 8390 2544
rect 8446 2488 9260 2544
rect 9366 2488 9416 2544
rect 8385 2486 9260 2488
rect 8385 2483 8451 2486
rect 9254 2484 9260 2486
rect 9324 2486 9416 2488
rect 9324 2484 9371 2486
rect 9806 2484 9812 2548
rect 9876 2546 9882 2548
rect 10041 2546 10107 2549
rect 9876 2544 10107 2546
rect 9876 2488 10046 2544
rect 10102 2488 10107 2544
rect 9876 2486 10107 2488
rect 9876 2484 9882 2486
rect 9305 2483 9371 2484
rect 10041 2483 10107 2486
rect 10317 2546 10383 2549
rect 11237 2546 11303 2549
rect 10317 2544 11303 2546
rect 10317 2488 10322 2544
rect 10378 2488 11242 2544
rect 11298 2488 11303 2544
rect 10317 2486 11303 2488
rect 10317 2483 10383 2486
rect 11237 2483 11303 2486
rect 11462 2484 11468 2548
rect 11532 2546 11538 2548
rect 14733 2546 14799 2549
rect 11532 2544 14799 2546
rect 11532 2488 14738 2544
rect 14794 2488 14799 2544
rect 11532 2486 14799 2488
rect 11532 2484 11538 2486
rect 14733 2483 14799 2486
rect 0 2410 800 2440
rect 3969 2410 4035 2413
rect 9121 2410 9187 2413
rect 13854 2410 13860 2412
rect 0 2408 4035 2410
rect 0 2352 3974 2408
rect 4030 2352 4035 2408
rect 0 2350 4035 2352
rect 0 2320 800 2350
rect 3969 2347 4035 2350
rect 4478 2350 8954 2410
rect 1853 2274 1919 2277
rect 4478 2274 4538 2350
rect 1853 2272 4538 2274
rect 1853 2216 1858 2272
rect 1914 2216 4538 2272
rect 1853 2214 4538 2216
rect 1853 2211 1919 2214
rect 5574 2212 5580 2276
rect 5644 2274 5650 2276
rect 6085 2274 6151 2277
rect 7925 2276 7991 2277
rect 7925 2274 7972 2276
rect 5644 2272 6151 2274
rect 5644 2216 6090 2272
rect 6146 2216 6151 2272
rect 5644 2214 6151 2216
rect 7880 2272 7972 2274
rect 7880 2216 7930 2272
rect 7880 2214 7972 2216
rect 5644 2212 5650 2214
rect 6085 2211 6151 2214
rect 7925 2212 7972 2214
rect 8036 2212 8042 2276
rect 8894 2274 8954 2350
rect 9121 2408 13860 2410
rect 9121 2352 9126 2408
rect 9182 2352 13860 2408
rect 9121 2350 13860 2352
rect 9121 2347 9187 2350
rect 13854 2348 13860 2350
rect 13924 2348 13930 2412
rect 11513 2274 11579 2277
rect 8894 2272 11579 2274
rect 8894 2216 11518 2272
rect 11574 2216 11579 2272
rect 8894 2214 11579 2216
rect 7925 2211 7991 2212
rect 11513 2211 11579 2214
rect 4692 2208 5012 2209
rect 4692 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5012 2208
rect 4692 2143 5012 2144
rect 8440 2208 8760 2209
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2143 8760 2144
rect 12188 2208 12508 2209
rect 12188 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12508 2208
rect 12188 2143 12508 2144
rect 1209 2138 1275 2141
rect 4521 2138 4587 2141
rect 1209 2136 4587 2138
rect 1209 2080 1214 2136
rect 1270 2080 4526 2136
rect 4582 2080 4587 2136
rect 1209 2078 4587 2080
rect 1209 2075 1275 2078
rect 4521 2075 4587 2078
rect 10910 2076 10916 2140
rect 10980 2138 10986 2140
rect 11513 2138 11579 2141
rect 10980 2136 11579 2138
rect 10980 2080 11518 2136
rect 11574 2080 11579 2136
rect 10980 2078 11579 2080
rect 10980 2076 10986 2078
rect 11513 2075 11579 2078
rect 7782 1940 7788 2004
rect 7852 2002 7858 2004
rect 11329 2002 11395 2005
rect 7852 2000 11395 2002
rect 7852 1944 11334 2000
rect 11390 1944 11395 2000
rect 7852 1942 11395 1944
rect 7852 1940 7858 1942
rect 11329 1939 11395 1942
rect 11830 1940 11836 2004
rect 11900 2002 11906 2004
rect 12065 2002 12131 2005
rect 11900 2000 12131 2002
rect 11900 1944 12070 2000
rect 12126 1944 12131 2000
rect 11900 1942 12131 1944
rect 11900 1940 11906 1942
rect 12065 1939 12131 1942
rect 7005 1866 7071 1869
rect 11462 1866 11468 1868
rect 7005 1864 11468 1866
rect 7005 1808 7010 1864
rect 7066 1808 11468 1864
rect 7005 1806 11468 1808
rect 7005 1803 7071 1806
rect 11462 1804 11468 1806
rect 11532 1804 11538 1868
rect 1945 1730 2011 1733
rect 1945 1728 2790 1730
rect 1945 1672 1950 1728
rect 2006 1672 2790 1728
rect 1945 1670 2790 1672
rect 1945 1667 2011 1670
rect 2730 1594 2790 1670
rect 7598 1668 7604 1732
rect 7668 1730 7674 1732
rect 12893 1730 12959 1733
rect 7668 1728 12959 1730
rect 7668 1672 12898 1728
rect 12954 1672 12959 1728
rect 7668 1670 12959 1672
rect 7668 1668 7674 1670
rect 12893 1667 12959 1670
rect 11145 1594 11211 1597
rect 2730 1592 11211 1594
rect 2730 1536 11150 1592
rect 11206 1536 11211 1592
rect 2730 1534 11211 1536
rect 11145 1531 11211 1534
rect 11421 1594 11487 1597
rect 12934 1594 12940 1596
rect 11421 1592 12940 1594
rect 11421 1536 11426 1592
rect 11482 1536 12940 1592
rect 11421 1534 12940 1536
rect 11421 1531 11487 1534
rect 12934 1532 12940 1534
rect 13004 1532 13010 1596
rect 0 1458 800 1488
rect 3509 1458 3575 1461
rect 0 1456 3575 1458
rect 0 1400 3514 1456
rect 3570 1400 3575 1456
rect 0 1398 3575 1400
rect 0 1368 800 1398
rect 3509 1395 3575 1398
rect 7649 1458 7715 1461
rect 9581 1458 9647 1461
rect 7649 1456 9647 1458
rect 7649 1400 7654 1456
rect 7710 1400 9586 1456
rect 9642 1400 9647 1456
rect 7649 1398 9647 1400
rect 7649 1395 7715 1398
rect 9581 1395 9647 1398
rect 11881 1458 11947 1461
rect 13670 1458 13676 1460
rect 11881 1456 13676 1458
rect 11881 1400 11886 1456
rect 11942 1400 13676 1456
rect 11881 1398 13676 1400
rect 11881 1395 11947 1398
rect 13670 1396 13676 1398
rect 13740 1396 13746 1460
rect 1158 1260 1164 1324
rect 1228 1322 1234 1324
rect 9213 1322 9279 1325
rect 1228 1320 9279 1322
rect 1228 1264 9218 1320
rect 9274 1264 9279 1320
rect 1228 1262 9279 1264
rect 1228 1260 1234 1262
rect 9213 1259 9279 1262
rect 13169 1322 13235 1325
rect 14774 1322 14780 1324
rect 13169 1320 14780 1322
rect 13169 1264 13174 1320
rect 13230 1264 14780 1320
rect 13169 1262 14780 1264
rect 13169 1259 13235 1262
rect 14774 1260 14780 1262
rect 14844 1260 14850 1324
rect 3366 1124 3372 1188
rect 3436 1186 3442 1188
rect 13353 1186 13419 1189
rect 3436 1184 13419 1186
rect 3436 1128 13358 1184
rect 13414 1128 13419 1184
rect 3436 1126 13419 1128
rect 3436 1124 3442 1126
rect 13353 1123 13419 1126
rect 381 1050 447 1053
rect 14089 1050 14155 1053
rect 381 1048 14155 1050
rect 381 992 386 1048
rect 442 992 14094 1048
rect 14150 992 14155 1048
rect 381 990 14155 992
rect 381 987 447 990
rect 14089 987 14155 990
rect 7046 852 7052 916
rect 7116 914 7122 916
rect 14181 914 14247 917
rect 7116 912 14247 914
rect 7116 856 14186 912
rect 14242 856 14247 912
rect 7116 854 14247 856
rect 7116 852 7122 854
rect 14181 851 14247 854
rect 6126 716 6132 780
rect 6196 778 6202 780
rect 9121 778 9187 781
rect 6196 776 9187 778
rect 6196 720 9126 776
rect 9182 720 9187 776
rect 6196 718 9187 720
rect 6196 716 6202 718
rect 9121 715 9187 718
rect 9765 642 9831 645
rect 13302 642 13308 644
rect 9765 640 13308 642
rect 9765 584 9770 640
rect 9826 584 13308 640
rect 9765 582 13308 584
rect 9765 579 9831 582
rect 13302 580 13308 582
rect 13372 580 13378 644
rect 0 506 800 536
rect 3417 506 3483 509
rect 0 504 3483 506
rect 0 448 3422 504
rect 3478 448 3483 504
rect 0 446 3483 448
rect 0 416 800 446
rect 3417 443 3483 446
rect 6729 234 6795 237
rect 12750 234 12756 236
rect 6729 232 12756 234
rect 6729 176 6734 232
rect 6790 176 12756 232
rect 6729 174 12756 176
rect 6729 171 6795 174
rect 12750 172 12756 174
rect 12820 172 12826 236
rect 1209 98 1275 101
rect 13537 98 13603 101
rect 1209 96 13603 98
rect 1209 40 1214 96
rect 1270 40 13542 96
rect 13598 40 13603 96
rect 1209 38 13603 40
rect 1209 35 1275 38
rect 13537 35 13603 38
<< via3 >>
rect 4108 18260 4172 18324
rect 10732 17988 10796 18052
rect 12572 17580 12636 17644
rect 7788 17444 7852 17508
rect 4700 17436 4764 17440
rect 4700 17380 4704 17436
rect 4704 17380 4760 17436
rect 4760 17380 4764 17436
rect 4700 17376 4764 17380
rect 4780 17436 4844 17440
rect 4780 17380 4784 17436
rect 4784 17380 4840 17436
rect 4840 17380 4844 17436
rect 4780 17376 4844 17380
rect 4860 17436 4924 17440
rect 4860 17380 4864 17436
rect 4864 17380 4920 17436
rect 4920 17380 4924 17436
rect 4860 17376 4924 17380
rect 4940 17436 5004 17440
rect 4940 17380 4944 17436
rect 4944 17380 5000 17436
rect 5000 17380 5004 17436
rect 4940 17376 5004 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 12196 17436 12260 17440
rect 12196 17380 12200 17436
rect 12200 17380 12256 17436
rect 12256 17380 12260 17436
rect 12196 17376 12260 17380
rect 12276 17436 12340 17440
rect 12276 17380 12280 17436
rect 12280 17380 12336 17436
rect 12336 17380 12340 17436
rect 12276 17376 12340 17380
rect 12356 17436 12420 17440
rect 12356 17380 12360 17436
rect 12360 17380 12416 17436
rect 12416 17380 12420 17436
rect 12356 17376 12420 17380
rect 12436 17436 12500 17440
rect 12436 17380 12440 17436
rect 12440 17380 12496 17436
rect 12496 17380 12500 17436
rect 12436 17376 12500 17380
rect 2636 17172 2700 17236
rect 13308 17172 13372 17236
rect 13124 17036 13188 17100
rect 2826 16892 2890 16896
rect 2826 16836 2830 16892
rect 2830 16836 2886 16892
rect 2886 16836 2890 16892
rect 2826 16832 2890 16836
rect 2906 16892 2970 16896
rect 2906 16836 2910 16892
rect 2910 16836 2966 16892
rect 2966 16836 2970 16892
rect 2906 16832 2970 16836
rect 2986 16892 3050 16896
rect 2986 16836 2990 16892
rect 2990 16836 3046 16892
rect 3046 16836 3050 16892
rect 2986 16832 3050 16836
rect 3066 16892 3130 16896
rect 3066 16836 3070 16892
rect 3070 16836 3126 16892
rect 3126 16836 3130 16892
rect 3066 16832 3130 16836
rect 6574 16892 6638 16896
rect 6574 16836 6578 16892
rect 6578 16836 6634 16892
rect 6634 16836 6638 16892
rect 6574 16832 6638 16836
rect 6654 16892 6718 16896
rect 6654 16836 6658 16892
rect 6658 16836 6714 16892
rect 6714 16836 6718 16892
rect 6654 16832 6718 16836
rect 6734 16892 6798 16896
rect 6734 16836 6738 16892
rect 6738 16836 6794 16892
rect 6794 16836 6798 16892
rect 6734 16832 6798 16836
rect 6814 16892 6878 16896
rect 6814 16836 6818 16892
rect 6818 16836 6874 16892
rect 6874 16836 6878 16892
rect 6814 16832 6878 16836
rect 10322 16892 10386 16896
rect 10322 16836 10326 16892
rect 10326 16836 10382 16892
rect 10382 16836 10386 16892
rect 10322 16832 10386 16836
rect 10402 16892 10466 16896
rect 10402 16836 10406 16892
rect 10406 16836 10462 16892
rect 10462 16836 10466 16892
rect 10402 16832 10466 16836
rect 10482 16892 10546 16896
rect 10482 16836 10486 16892
rect 10486 16836 10542 16892
rect 10542 16836 10546 16892
rect 10482 16832 10546 16836
rect 10562 16892 10626 16896
rect 10562 16836 10566 16892
rect 10566 16836 10622 16892
rect 10622 16836 10626 16892
rect 10562 16832 10626 16836
rect 14070 16892 14134 16896
rect 14070 16836 14074 16892
rect 14074 16836 14130 16892
rect 14130 16836 14134 16892
rect 14070 16832 14134 16836
rect 14150 16892 14214 16896
rect 14150 16836 14154 16892
rect 14154 16836 14210 16892
rect 14210 16836 14214 16892
rect 14150 16832 14214 16836
rect 14230 16892 14294 16896
rect 14230 16836 14234 16892
rect 14234 16836 14290 16892
rect 14290 16836 14294 16892
rect 14230 16832 14294 16836
rect 14310 16892 14374 16896
rect 14310 16836 14314 16892
rect 14314 16836 14370 16892
rect 14370 16836 14374 16892
rect 14310 16832 14374 16836
rect 4292 16628 4356 16692
rect 4700 16348 4764 16352
rect 4700 16292 4704 16348
rect 4704 16292 4760 16348
rect 4760 16292 4764 16348
rect 4700 16288 4764 16292
rect 4780 16348 4844 16352
rect 4780 16292 4784 16348
rect 4784 16292 4840 16348
rect 4840 16292 4844 16348
rect 4780 16288 4844 16292
rect 4860 16348 4924 16352
rect 4860 16292 4864 16348
rect 4864 16292 4920 16348
rect 4920 16292 4924 16348
rect 4860 16288 4924 16292
rect 4940 16348 5004 16352
rect 4940 16292 4944 16348
rect 4944 16292 5000 16348
rect 5000 16292 5004 16348
rect 4940 16288 5004 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 12196 16348 12260 16352
rect 12196 16292 12200 16348
rect 12200 16292 12256 16348
rect 12256 16292 12260 16348
rect 12196 16288 12260 16292
rect 12276 16348 12340 16352
rect 12276 16292 12280 16348
rect 12280 16292 12336 16348
rect 12336 16292 12340 16348
rect 12276 16288 12340 16292
rect 12356 16348 12420 16352
rect 12356 16292 12360 16348
rect 12360 16292 12416 16348
rect 12416 16292 12420 16348
rect 12356 16288 12420 16292
rect 12436 16348 12500 16352
rect 12436 16292 12440 16348
rect 12440 16292 12496 16348
rect 12496 16292 12500 16348
rect 12436 16288 12500 16292
rect 9076 16084 9140 16148
rect 7052 16008 7116 16012
rect 7052 15952 7066 16008
rect 7066 15952 7116 16008
rect 7052 15948 7116 15952
rect 1164 15812 1228 15876
rect 2826 15804 2890 15808
rect 2826 15748 2830 15804
rect 2830 15748 2886 15804
rect 2886 15748 2890 15804
rect 2826 15744 2890 15748
rect 2906 15804 2970 15808
rect 2906 15748 2910 15804
rect 2910 15748 2966 15804
rect 2966 15748 2970 15804
rect 2906 15744 2970 15748
rect 2986 15804 3050 15808
rect 2986 15748 2990 15804
rect 2990 15748 3046 15804
rect 3046 15748 3050 15804
rect 2986 15744 3050 15748
rect 3066 15804 3130 15808
rect 3066 15748 3070 15804
rect 3070 15748 3126 15804
rect 3126 15748 3130 15804
rect 3066 15744 3130 15748
rect 6574 15804 6638 15808
rect 6574 15748 6578 15804
rect 6578 15748 6634 15804
rect 6634 15748 6638 15804
rect 6574 15744 6638 15748
rect 6654 15804 6718 15808
rect 6654 15748 6658 15804
rect 6658 15748 6714 15804
rect 6714 15748 6718 15804
rect 6654 15744 6718 15748
rect 6734 15804 6798 15808
rect 6734 15748 6738 15804
rect 6738 15748 6794 15804
rect 6794 15748 6798 15804
rect 6734 15744 6798 15748
rect 6814 15804 6878 15808
rect 6814 15748 6818 15804
rect 6818 15748 6874 15804
rect 6874 15748 6878 15804
rect 6814 15744 6878 15748
rect 10322 15804 10386 15808
rect 10322 15748 10326 15804
rect 10326 15748 10382 15804
rect 10382 15748 10386 15804
rect 10322 15744 10386 15748
rect 10402 15804 10466 15808
rect 10402 15748 10406 15804
rect 10406 15748 10462 15804
rect 10462 15748 10466 15804
rect 10402 15744 10466 15748
rect 10482 15804 10546 15808
rect 10482 15748 10486 15804
rect 10486 15748 10542 15804
rect 10542 15748 10546 15804
rect 10482 15744 10546 15748
rect 10562 15804 10626 15808
rect 10562 15748 10566 15804
rect 10566 15748 10622 15804
rect 10622 15748 10626 15804
rect 10562 15744 10626 15748
rect 14070 15804 14134 15808
rect 14070 15748 14074 15804
rect 14074 15748 14130 15804
rect 14130 15748 14134 15804
rect 14070 15744 14134 15748
rect 14150 15804 14214 15808
rect 14150 15748 14154 15804
rect 14154 15748 14210 15804
rect 14210 15748 14214 15804
rect 14150 15744 14214 15748
rect 14230 15804 14294 15808
rect 14230 15748 14234 15804
rect 14234 15748 14290 15804
rect 14290 15748 14294 15804
rect 14230 15744 14294 15748
rect 14310 15804 14374 15808
rect 14310 15748 14314 15804
rect 14314 15748 14370 15804
rect 14370 15748 14374 15804
rect 14310 15744 14374 15748
rect 1348 15676 1412 15740
rect 4476 15676 4540 15740
rect 9812 15676 9876 15740
rect 5396 15464 5460 15468
rect 5396 15408 5410 15464
rect 5410 15408 5460 15464
rect 5396 15404 5460 15408
rect 11468 15404 11532 15468
rect 4700 15260 4764 15264
rect 4700 15204 4704 15260
rect 4704 15204 4760 15260
rect 4760 15204 4764 15260
rect 4700 15200 4764 15204
rect 4780 15260 4844 15264
rect 4780 15204 4784 15260
rect 4784 15204 4840 15260
rect 4840 15204 4844 15260
rect 4780 15200 4844 15204
rect 4860 15260 4924 15264
rect 4860 15204 4864 15260
rect 4864 15204 4920 15260
rect 4920 15204 4924 15260
rect 4860 15200 4924 15204
rect 4940 15260 5004 15264
rect 4940 15204 4944 15260
rect 4944 15204 5000 15260
rect 5000 15204 5004 15260
rect 4940 15200 5004 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 12196 15260 12260 15264
rect 12196 15204 12200 15260
rect 12200 15204 12256 15260
rect 12256 15204 12260 15260
rect 12196 15200 12260 15204
rect 12276 15260 12340 15264
rect 12276 15204 12280 15260
rect 12280 15204 12336 15260
rect 12336 15204 12340 15260
rect 12276 15200 12340 15204
rect 12356 15260 12420 15264
rect 12356 15204 12360 15260
rect 12360 15204 12416 15260
rect 12416 15204 12420 15260
rect 12356 15200 12420 15204
rect 12436 15260 12500 15264
rect 12436 15204 12440 15260
rect 12440 15204 12496 15260
rect 12496 15204 12500 15260
rect 12436 15200 12500 15204
rect 7972 14996 8036 15060
rect 13860 14996 13924 15060
rect 5764 14724 5828 14788
rect 9260 14724 9324 14788
rect 2826 14716 2890 14720
rect 2826 14660 2830 14716
rect 2830 14660 2886 14716
rect 2886 14660 2890 14716
rect 2826 14656 2890 14660
rect 2906 14716 2970 14720
rect 2906 14660 2910 14716
rect 2910 14660 2966 14716
rect 2966 14660 2970 14716
rect 2906 14656 2970 14660
rect 2986 14716 3050 14720
rect 2986 14660 2990 14716
rect 2990 14660 3046 14716
rect 3046 14660 3050 14716
rect 2986 14656 3050 14660
rect 3066 14716 3130 14720
rect 3066 14660 3070 14716
rect 3070 14660 3126 14716
rect 3126 14660 3130 14716
rect 3066 14656 3130 14660
rect 6574 14716 6638 14720
rect 6574 14660 6578 14716
rect 6578 14660 6634 14716
rect 6634 14660 6638 14716
rect 6574 14656 6638 14660
rect 6654 14716 6718 14720
rect 6654 14660 6658 14716
rect 6658 14660 6714 14716
rect 6714 14660 6718 14716
rect 6654 14656 6718 14660
rect 6734 14716 6798 14720
rect 6734 14660 6738 14716
rect 6738 14660 6794 14716
rect 6794 14660 6798 14716
rect 6734 14656 6798 14660
rect 6814 14716 6878 14720
rect 6814 14660 6818 14716
rect 6818 14660 6874 14716
rect 6874 14660 6878 14716
rect 6814 14656 6878 14660
rect 10322 14716 10386 14720
rect 10322 14660 10326 14716
rect 10326 14660 10382 14716
rect 10382 14660 10386 14716
rect 10322 14656 10386 14660
rect 10402 14716 10466 14720
rect 10402 14660 10406 14716
rect 10406 14660 10462 14716
rect 10462 14660 10466 14716
rect 10402 14656 10466 14660
rect 10482 14716 10546 14720
rect 10482 14660 10486 14716
rect 10486 14660 10542 14716
rect 10542 14660 10546 14716
rect 10482 14656 10546 14660
rect 10562 14716 10626 14720
rect 10562 14660 10566 14716
rect 10566 14660 10622 14716
rect 10622 14660 10626 14716
rect 10562 14656 10626 14660
rect 14070 14716 14134 14720
rect 14070 14660 14074 14716
rect 14074 14660 14130 14716
rect 14130 14660 14134 14716
rect 14070 14656 14134 14660
rect 14150 14716 14214 14720
rect 14150 14660 14154 14716
rect 14154 14660 14210 14716
rect 14210 14660 14214 14716
rect 14150 14656 14214 14660
rect 14230 14716 14294 14720
rect 14230 14660 14234 14716
rect 14234 14660 14290 14716
rect 14290 14660 14294 14716
rect 14230 14656 14294 14660
rect 14310 14716 14374 14720
rect 14310 14660 14314 14716
rect 14314 14660 14370 14716
rect 14370 14660 14374 14716
rect 14310 14656 14374 14660
rect 980 14588 1044 14652
rect 3372 14648 3436 14652
rect 3372 14592 3386 14648
rect 3386 14592 3436 14648
rect 3372 14588 3436 14592
rect 1716 14452 1780 14516
rect 1532 14180 1596 14244
rect 4108 14316 4172 14380
rect 7604 14180 7668 14244
rect 4700 14172 4764 14176
rect 4700 14116 4704 14172
rect 4704 14116 4760 14172
rect 4760 14116 4764 14172
rect 4700 14112 4764 14116
rect 4780 14172 4844 14176
rect 4780 14116 4784 14172
rect 4784 14116 4840 14172
rect 4840 14116 4844 14172
rect 4780 14112 4844 14116
rect 4860 14172 4924 14176
rect 4860 14116 4864 14172
rect 4864 14116 4920 14172
rect 4920 14116 4924 14172
rect 4860 14112 4924 14116
rect 4940 14172 5004 14176
rect 4940 14116 4944 14172
rect 4944 14116 5000 14172
rect 5000 14116 5004 14172
rect 4940 14112 5004 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 12196 14172 12260 14176
rect 12196 14116 12200 14172
rect 12200 14116 12256 14172
rect 12256 14116 12260 14172
rect 12196 14112 12260 14116
rect 12276 14172 12340 14176
rect 12276 14116 12280 14172
rect 12280 14116 12336 14172
rect 12336 14116 12340 14172
rect 12276 14112 12340 14116
rect 12356 14172 12420 14176
rect 12356 14116 12360 14172
rect 12360 14116 12416 14172
rect 12416 14116 12420 14172
rect 12356 14112 12420 14116
rect 12436 14172 12500 14176
rect 12436 14116 12440 14172
rect 12440 14116 12496 14172
rect 12496 14116 12500 14172
rect 12436 14112 12500 14116
rect 3924 14044 3988 14108
rect 9260 14044 9324 14108
rect 3740 13832 3804 13836
rect 3740 13776 3790 13832
rect 3790 13776 3804 13832
rect 3740 13772 3804 13776
rect 4108 13772 4172 13836
rect 5580 13772 5644 13836
rect 9628 13772 9692 13836
rect 11100 13772 11164 13836
rect 2826 13628 2890 13632
rect 2826 13572 2830 13628
rect 2830 13572 2886 13628
rect 2886 13572 2890 13628
rect 2826 13568 2890 13572
rect 2906 13628 2970 13632
rect 2906 13572 2910 13628
rect 2910 13572 2966 13628
rect 2966 13572 2970 13628
rect 2906 13568 2970 13572
rect 2986 13628 3050 13632
rect 2986 13572 2990 13628
rect 2990 13572 3046 13628
rect 3046 13572 3050 13628
rect 2986 13568 3050 13572
rect 3066 13628 3130 13632
rect 3066 13572 3070 13628
rect 3070 13572 3126 13628
rect 3126 13572 3130 13628
rect 3066 13568 3130 13572
rect 6574 13628 6638 13632
rect 6574 13572 6578 13628
rect 6578 13572 6634 13628
rect 6634 13572 6638 13628
rect 6574 13568 6638 13572
rect 6654 13628 6718 13632
rect 6654 13572 6658 13628
rect 6658 13572 6714 13628
rect 6714 13572 6718 13628
rect 6654 13568 6718 13572
rect 6734 13628 6798 13632
rect 6734 13572 6738 13628
rect 6738 13572 6794 13628
rect 6794 13572 6798 13628
rect 6734 13568 6798 13572
rect 6814 13628 6878 13632
rect 6814 13572 6818 13628
rect 6818 13572 6874 13628
rect 6874 13572 6878 13628
rect 6814 13568 6878 13572
rect 9444 13500 9508 13564
rect 10322 13628 10386 13632
rect 10322 13572 10326 13628
rect 10326 13572 10382 13628
rect 10382 13572 10386 13628
rect 10322 13568 10386 13572
rect 10402 13628 10466 13632
rect 10402 13572 10406 13628
rect 10406 13572 10462 13628
rect 10462 13572 10466 13628
rect 10402 13568 10466 13572
rect 10482 13628 10546 13632
rect 10482 13572 10486 13628
rect 10486 13572 10542 13628
rect 10542 13572 10546 13628
rect 10482 13568 10546 13572
rect 10562 13628 10626 13632
rect 10562 13572 10566 13628
rect 10566 13572 10622 13628
rect 10622 13572 10626 13628
rect 10562 13568 10626 13572
rect 14070 13628 14134 13632
rect 14070 13572 14074 13628
rect 14074 13572 14130 13628
rect 14130 13572 14134 13628
rect 14070 13568 14134 13572
rect 14150 13628 14214 13632
rect 14150 13572 14154 13628
rect 14154 13572 14210 13628
rect 14210 13572 14214 13628
rect 14150 13568 14214 13572
rect 14230 13628 14294 13632
rect 14230 13572 14234 13628
rect 14234 13572 14290 13628
rect 14290 13572 14294 13628
rect 14230 13568 14294 13572
rect 14310 13628 14374 13632
rect 14310 13572 14314 13628
rect 14314 13572 14370 13628
rect 14370 13572 14374 13628
rect 14310 13568 14374 13572
rect 10180 13560 10244 13564
rect 10180 13504 10194 13560
rect 10194 13504 10244 13560
rect 10180 13500 10244 13504
rect 13676 13500 13740 13564
rect 4292 13364 4356 13428
rect 9996 13288 10060 13292
rect 9996 13232 10010 13288
rect 10010 13232 10060 13288
rect 9996 13228 10060 13232
rect 4700 13084 4764 13088
rect 4700 13028 4704 13084
rect 4704 13028 4760 13084
rect 4760 13028 4764 13084
rect 4700 13024 4764 13028
rect 4780 13084 4844 13088
rect 4780 13028 4784 13084
rect 4784 13028 4840 13084
rect 4840 13028 4844 13084
rect 4780 13024 4844 13028
rect 4860 13084 4924 13088
rect 4860 13028 4864 13084
rect 4864 13028 4920 13084
rect 4920 13028 4924 13084
rect 4860 13024 4924 13028
rect 4940 13084 5004 13088
rect 4940 13028 4944 13084
rect 4944 13028 5000 13084
rect 5000 13028 5004 13084
rect 4940 13024 5004 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 12196 13084 12260 13088
rect 12196 13028 12200 13084
rect 12200 13028 12256 13084
rect 12256 13028 12260 13084
rect 12196 13024 12260 13028
rect 12276 13084 12340 13088
rect 12276 13028 12280 13084
rect 12280 13028 12336 13084
rect 12336 13028 12340 13084
rect 12276 13024 12340 13028
rect 12356 13084 12420 13088
rect 12356 13028 12360 13084
rect 12360 13028 12416 13084
rect 12416 13028 12420 13084
rect 12356 13024 12420 13028
rect 12436 13084 12500 13088
rect 12436 13028 12440 13084
rect 12440 13028 12496 13084
rect 12496 13028 12500 13084
rect 12436 13024 12500 13028
rect 5396 12956 5460 13020
rect 7236 12956 7300 13020
rect 9444 12956 9508 13020
rect 12020 12956 12084 13020
rect 5396 12684 5460 12748
rect 2452 12548 2516 12612
rect 5212 12548 5276 12612
rect 11284 12880 11348 12884
rect 11284 12824 11298 12880
rect 11298 12824 11348 12880
rect 11284 12820 11348 12824
rect 12940 12820 13004 12884
rect 8156 12548 8220 12612
rect 2826 12540 2890 12544
rect 2826 12484 2830 12540
rect 2830 12484 2886 12540
rect 2886 12484 2890 12540
rect 2826 12480 2890 12484
rect 2906 12540 2970 12544
rect 2906 12484 2910 12540
rect 2910 12484 2966 12540
rect 2966 12484 2970 12540
rect 2906 12480 2970 12484
rect 2986 12540 3050 12544
rect 2986 12484 2990 12540
rect 2990 12484 3046 12540
rect 3046 12484 3050 12540
rect 2986 12480 3050 12484
rect 3066 12540 3130 12544
rect 3066 12484 3070 12540
rect 3070 12484 3126 12540
rect 3126 12484 3130 12540
rect 3066 12480 3130 12484
rect 6574 12540 6638 12544
rect 6574 12484 6578 12540
rect 6578 12484 6634 12540
rect 6634 12484 6638 12540
rect 6574 12480 6638 12484
rect 6654 12540 6718 12544
rect 6654 12484 6658 12540
rect 6658 12484 6714 12540
rect 6714 12484 6718 12540
rect 6654 12480 6718 12484
rect 6734 12540 6798 12544
rect 6734 12484 6738 12540
rect 6738 12484 6794 12540
rect 6794 12484 6798 12540
rect 6734 12480 6798 12484
rect 6814 12540 6878 12544
rect 6814 12484 6818 12540
rect 6818 12484 6874 12540
rect 6874 12484 6878 12540
rect 6814 12480 6878 12484
rect 3556 12412 3620 12476
rect 10322 12540 10386 12544
rect 10322 12484 10326 12540
rect 10326 12484 10382 12540
rect 10382 12484 10386 12540
rect 10322 12480 10386 12484
rect 10402 12540 10466 12544
rect 10402 12484 10406 12540
rect 10406 12484 10462 12540
rect 10462 12484 10466 12540
rect 10402 12480 10466 12484
rect 10482 12540 10546 12544
rect 10482 12484 10486 12540
rect 10486 12484 10542 12540
rect 10542 12484 10546 12540
rect 10482 12480 10546 12484
rect 10562 12540 10626 12544
rect 10562 12484 10566 12540
rect 10566 12484 10622 12540
rect 10622 12484 10626 12540
rect 10562 12480 10626 12484
rect 14070 12540 14134 12544
rect 14070 12484 14074 12540
rect 14074 12484 14130 12540
rect 14130 12484 14134 12540
rect 14070 12480 14134 12484
rect 14150 12540 14214 12544
rect 14150 12484 14154 12540
rect 14154 12484 14210 12540
rect 14210 12484 14214 12540
rect 14150 12480 14214 12484
rect 14230 12540 14294 12544
rect 14230 12484 14234 12540
rect 14234 12484 14290 12540
rect 14290 12484 14294 12540
rect 14230 12480 14294 12484
rect 14310 12540 14374 12544
rect 14310 12484 14314 12540
rect 14314 12484 14370 12540
rect 14370 12484 14374 12540
rect 14310 12480 14374 12484
rect 10732 12412 10796 12476
rect 13492 12412 13556 12476
rect 5212 12276 5276 12340
rect 7788 12276 7852 12340
rect 8892 12276 8956 12340
rect 9076 12336 9140 12340
rect 9076 12280 9090 12336
rect 9090 12280 9140 12336
rect 9076 12276 9140 12280
rect 9260 12276 9324 12340
rect 13860 12276 13924 12340
rect 796 12004 860 12068
rect 1164 12004 1228 12068
rect 5764 12064 5828 12068
rect 5764 12008 5778 12064
rect 5778 12008 5828 12064
rect 5764 12004 5828 12008
rect 4700 11996 4764 12000
rect 4700 11940 4704 11996
rect 4704 11940 4760 11996
rect 4760 11940 4764 11996
rect 4700 11936 4764 11940
rect 4780 11996 4844 12000
rect 4780 11940 4784 11996
rect 4784 11940 4840 11996
rect 4840 11940 4844 11996
rect 4780 11936 4844 11940
rect 4860 11996 4924 12000
rect 4860 11940 4864 11996
rect 4864 11940 4920 11996
rect 4920 11940 4924 11996
rect 4860 11936 4924 11940
rect 4940 11996 5004 12000
rect 4940 11940 4944 11996
rect 4944 11940 5000 11996
rect 5000 11940 5004 11996
rect 4940 11936 5004 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 1164 11868 1228 11932
rect 2636 11928 2700 11932
rect 2636 11872 2686 11928
rect 2686 11872 2700 11928
rect 2636 11868 2700 11872
rect 7420 11868 7484 11932
rect 9260 11868 9324 11932
rect 11652 12140 11716 12204
rect 9628 12004 9692 12068
rect 11284 12004 11348 12068
rect 12196 11996 12260 12000
rect 12196 11940 12200 11996
rect 12200 11940 12256 11996
rect 12256 11940 12260 11996
rect 12196 11936 12260 11940
rect 12276 11996 12340 12000
rect 12276 11940 12280 11996
rect 12280 11940 12336 11996
rect 12336 11940 12340 11996
rect 12276 11936 12340 11940
rect 12356 11996 12420 12000
rect 12356 11940 12360 11996
rect 12360 11940 12416 11996
rect 12416 11940 12420 11996
rect 12356 11936 12420 11940
rect 12436 11996 12500 12000
rect 12436 11940 12440 11996
rect 12440 11940 12496 11996
rect 12496 11940 12500 11996
rect 12436 11936 12500 11940
rect 7788 11732 7852 11796
rect 9260 11792 9324 11796
rect 9260 11736 9274 11792
rect 9274 11736 9324 11792
rect 9260 11732 9324 11736
rect 9812 11732 9876 11796
rect 3556 11596 3620 11660
rect 7604 11460 7668 11524
rect 2826 11452 2890 11456
rect 2826 11396 2830 11452
rect 2830 11396 2886 11452
rect 2886 11396 2890 11452
rect 2826 11392 2890 11396
rect 2906 11452 2970 11456
rect 2906 11396 2910 11452
rect 2910 11396 2966 11452
rect 2966 11396 2970 11452
rect 2906 11392 2970 11396
rect 2986 11452 3050 11456
rect 2986 11396 2990 11452
rect 2990 11396 3046 11452
rect 3046 11396 3050 11452
rect 2986 11392 3050 11396
rect 3066 11452 3130 11456
rect 3066 11396 3070 11452
rect 3070 11396 3126 11452
rect 3126 11396 3130 11452
rect 3066 11392 3130 11396
rect 6574 11452 6638 11456
rect 6574 11396 6578 11452
rect 6578 11396 6634 11452
rect 6634 11396 6638 11452
rect 6574 11392 6638 11396
rect 6654 11452 6718 11456
rect 6654 11396 6658 11452
rect 6658 11396 6714 11452
rect 6714 11396 6718 11452
rect 6654 11392 6718 11396
rect 6734 11452 6798 11456
rect 6734 11396 6738 11452
rect 6738 11396 6794 11452
rect 6794 11396 6798 11452
rect 6734 11392 6798 11396
rect 6814 11452 6878 11456
rect 6814 11396 6818 11452
rect 6818 11396 6874 11452
rect 6874 11396 6878 11452
rect 6814 11392 6878 11396
rect 4476 11324 4540 11388
rect 6316 11324 6380 11388
rect 9628 11460 9692 11524
rect 10322 11452 10386 11456
rect 10322 11396 10326 11452
rect 10326 11396 10382 11452
rect 10382 11396 10386 11452
rect 10322 11392 10386 11396
rect 10402 11452 10466 11456
rect 10402 11396 10406 11452
rect 10406 11396 10462 11452
rect 10462 11396 10466 11452
rect 10402 11392 10466 11396
rect 10482 11452 10546 11456
rect 10482 11396 10486 11452
rect 10486 11396 10542 11452
rect 10542 11396 10546 11452
rect 10482 11392 10546 11396
rect 10562 11452 10626 11456
rect 10562 11396 10566 11452
rect 10566 11396 10622 11452
rect 10622 11396 10626 11452
rect 10562 11392 10626 11396
rect 9996 11384 10060 11388
rect 9996 11328 10010 11384
rect 10010 11328 10060 11384
rect 9996 11324 10060 11328
rect 7972 11188 8036 11252
rect 9996 11188 10060 11252
rect 13860 11928 13924 11932
rect 13860 11872 13874 11928
rect 13874 11872 13924 11928
rect 13860 11868 13924 11872
rect 12756 11596 12820 11660
rect 11836 11324 11900 11388
rect 13492 11384 13556 11388
rect 13492 11328 13542 11384
rect 13542 11328 13556 11384
rect 13492 11324 13556 11328
rect 11468 11188 11532 11252
rect 14070 11452 14134 11456
rect 14070 11396 14074 11452
rect 14074 11396 14130 11452
rect 14130 11396 14134 11452
rect 14070 11392 14134 11396
rect 14150 11452 14214 11456
rect 14150 11396 14154 11452
rect 14154 11396 14210 11452
rect 14210 11396 14214 11452
rect 14150 11392 14214 11396
rect 14230 11452 14294 11456
rect 14230 11396 14234 11452
rect 14234 11396 14290 11452
rect 14290 11396 14294 11452
rect 14230 11392 14294 11396
rect 14310 11452 14374 11456
rect 14310 11396 14314 11452
rect 14314 11396 14370 11452
rect 14370 11396 14374 11452
rect 14310 11392 14374 11396
rect 14780 11384 14844 11388
rect 14780 11328 14794 11384
rect 14794 11328 14844 11384
rect 14780 11324 14844 11328
rect 1900 11112 1964 11116
rect 1900 11056 1914 11112
rect 1914 11056 1964 11112
rect 1900 11052 1964 11056
rect 10916 11052 10980 11116
rect 12572 11052 12636 11116
rect 4700 10908 4764 10912
rect 4700 10852 4704 10908
rect 4704 10852 4760 10908
rect 4760 10852 4764 10908
rect 4700 10848 4764 10852
rect 4780 10908 4844 10912
rect 4780 10852 4784 10908
rect 4784 10852 4840 10908
rect 4840 10852 4844 10908
rect 4780 10848 4844 10852
rect 4860 10908 4924 10912
rect 4860 10852 4864 10908
rect 4864 10852 4920 10908
rect 4920 10852 4924 10908
rect 4860 10848 4924 10852
rect 4940 10908 5004 10912
rect 4940 10852 4944 10908
rect 4944 10852 5000 10908
rect 5000 10852 5004 10908
rect 4940 10848 5004 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 3372 10780 3436 10844
rect 7420 10780 7484 10844
rect 9444 10780 9508 10844
rect 13860 10916 13924 10980
rect 12196 10908 12260 10912
rect 12196 10852 12200 10908
rect 12200 10852 12256 10908
rect 12256 10852 12260 10908
rect 12196 10848 12260 10852
rect 12276 10908 12340 10912
rect 12276 10852 12280 10908
rect 12280 10852 12336 10908
rect 12336 10852 12340 10908
rect 12276 10848 12340 10852
rect 12356 10908 12420 10912
rect 12356 10852 12360 10908
rect 12360 10852 12416 10908
rect 12416 10852 12420 10908
rect 12356 10848 12420 10852
rect 12436 10908 12500 10912
rect 12436 10852 12440 10908
rect 12440 10852 12496 10908
rect 12496 10852 12500 10908
rect 12436 10848 12500 10852
rect 13124 10780 13188 10844
rect 14596 10780 14660 10844
rect 9076 10508 9140 10572
rect 9996 10508 10060 10572
rect 11652 10508 11716 10572
rect 13676 10644 13740 10708
rect 13492 10508 13556 10572
rect 2826 10364 2890 10368
rect 2826 10308 2830 10364
rect 2830 10308 2886 10364
rect 2886 10308 2890 10364
rect 2826 10304 2890 10308
rect 2906 10364 2970 10368
rect 2906 10308 2910 10364
rect 2910 10308 2966 10364
rect 2966 10308 2970 10364
rect 2906 10304 2970 10308
rect 2986 10364 3050 10368
rect 2986 10308 2990 10364
rect 2990 10308 3046 10364
rect 3046 10308 3050 10364
rect 2986 10304 3050 10308
rect 3066 10364 3130 10368
rect 3066 10308 3070 10364
rect 3070 10308 3126 10364
rect 3126 10308 3130 10364
rect 3066 10304 3130 10308
rect 6574 10364 6638 10368
rect 6574 10308 6578 10364
rect 6578 10308 6634 10364
rect 6634 10308 6638 10364
rect 6574 10304 6638 10308
rect 6654 10364 6718 10368
rect 6654 10308 6658 10364
rect 6658 10308 6714 10364
rect 6714 10308 6718 10364
rect 6654 10304 6718 10308
rect 6734 10364 6798 10368
rect 6734 10308 6738 10364
rect 6738 10308 6794 10364
rect 6794 10308 6798 10364
rect 6734 10304 6798 10308
rect 6814 10364 6878 10368
rect 6814 10308 6818 10364
rect 6818 10308 6874 10364
rect 6874 10308 6878 10364
rect 6814 10304 6878 10308
rect 10322 10364 10386 10368
rect 10322 10308 10326 10364
rect 10326 10308 10382 10364
rect 10382 10308 10386 10364
rect 10322 10304 10386 10308
rect 10402 10364 10466 10368
rect 10402 10308 10406 10364
rect 10406 10308 10462 10364
rect 10462 10308 10466 10364
rect 10402 10304 10466 10308
rect 10482 10364 10546 10368
rect 10482 10308 10486 10364
rect 10486 10308 10542 10364
rect 10542 10308 10546 10364
rect 10482 10304 10546 10308
rect 10562 10364 10626 10368
rect 10562 10308 10566 10364
rect 10566 10308 10622 10364
rect 10622 10308 10626 10364
rect 10562 10304 10626 10308
rect 14070 10364 14134 10368
rect 14070 10308 14074 10364
rect 14074 10308 14130 10364
rect 14130 10308 14134 10364
rect 14070 10304 14134 10308
rect 14150 10364 14214 10368
rect 14150 10308 14154 10364
rect 14154 10308 14210 10364
rect 14210 10308 14214 10364
rect 14150 10304 14214 10308
rect 14230 10364 14294 10368
rect 14230 10308 14234 10364
rect 14234 10308 14290 10364
rect 14290 10308 14294 10364
rect 14230 10304 14294 10308
rect 14310 10364 14374 10368
rect 14310 10308 14314 10364
rect 14314 10308 14370 10364
rect 14370 10308 14374 10364
rect 14310 10304 14374 10308
rect 13860 10236 13924 10300
rect 8892 10100 8956 10164
rect 12756 10100 12820 10164
rect 4108 9828 4172 9892
rect 4476 9828 4540 9892
rect 10180 9828 10244 9892
rect 11100 9888 11164 9892
rect 11100 9832 11150 9888
rect 11150 9832 11164 9888
rect 11100 9828 11164 9832
rect 13492 9828 13556 9892
rect 13860 9828 13924 9892
rect 4700 9820 4764 9824
rect 4700 9764 4704 9820
rect 4704 9764 4760 9820
rect 4760 9764 4764 9820
rect 4700 9760 4764 9764
rect 4780 9820 4844 9824
rect 4780 9764 4784 9820
rect 4784 9764 4840 9820
rect 4840 9764 4844 9820
rect 4780 9760 4844 9764
rect 4860 9820 4924 9824
rect 4860 9764 4864 9820
rect 4864 9764 4920 9820
rect 4920 9764 4924 9820
rect 4860 9760 4924 9764
rect 4940 9820 5004 9824
rect 4940 9764 4944 9820
rect 4944 9764 5000 9820
rect 5000 9764 5004 9820
rect 4940 9760 5004 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 12196 9820 12260 9824
rect 12196 9764 12200 9820
rect 12200 9764 12256 9820
rect 12256 9764 12260 9820
rect 12196 9760 12260 9764
rect 12276 9820 12340 9824
rect 12276 9764 12280 9820
rect 12280 9764 12336 9820
rect 12336 9764 12340 9820
rect 12276 9760 12340 9764
rect 12356 9820 12420 9824
rect 12356 9764 12360 9820
rect 12360 9764 12416 9820
rect 12416 9764 12420 9820
rect 12356 9760 12420 9764
rect 12436 9820 12500 9824
rect 12436 9764 12440 9820
rect 12440 9764 12496 9820
rect 12496 9764 12500 9820
rect 12436 9760 12500 9764
rect 7420 9556 7484 9620
rect 10916 9556 10980 9620
rect 13124 9692 13188 9756
rect 13308 9556 13372 9620
rect 7236 9344 7300 9348
rect 7236 9288 7286 9344
rect 7286 9288 7300 9344
rect 7236 9284 7300 9288
rect 12020 9284 12084 9348
rect 2826 9276 2890 9280
rect 2826 9220 2830 9276
rect 2830 9220 2886 9276
rect 2886 9220 2890 9276
rect 2826 9216 2890 9220
rect 2906 9276 2970 9280
rect 2906 9220 2910 9276
rect 2910 9220 2966 9276
rect 2966 9220 2970 9276
rect 2906 9216 2970 9220
rect 2986 9276 3050 9280
rect 2986 9220 2990 9276
rect 2990 9220 3046 9276
rect 3046 9220 3050 9276
rect 2986 9216 3050 9220
rect 3066 9276 3130 9280
rect 3066 9220 3070 9276
rect 3070 9220 3126 9276
rect 3126 9220 3130 9276
rect 3066 9216 3130 9220
rect 6574 9276 6638 9280
rect 6574 9220 6578 9276
rect 6578 9220 6634 9276
rect 6634 9220 6638 9276
rect 6574 9216 6638 9220
rect 6654 9276 6718 9280
rect 6654 9220 6658 9276
rect 6658 9220 6714 9276
rect 6714 9220 6718 9276
rect 6654 9216 6718 9220
rect 6734 9276 6798 9280
rect 6734 9220 6738 9276
rect 6738 9220 6794 9276
rect 6794 9220 6798 9276
rect 6734 9216 6798 9220
rect 6814 9276 6878 9280
rect 6814 9220 6818 9276
rect 6818 9220 6874 9276
rect 6874 9220 6878 9276
rect 6814 9216 6878 9220
rect 10322 9276 10386 9280
rect 10322 9220 10326 9276
rect 10326 9220 10382 9276
rect 10382 9220 10386 9276
rect 10322 9216 10386 9220
rect 10402 9276 10466 9280
rect 10402 9220 10406 9276
rect 10406 9220 10462 9276
rect 10462 9220 10466 9276
rect 10402 9216 10466 9220
rect 10482 9276 10546 9280
rect 10482 9220 10486 9276
rect 10486 9220 10542 9276
rect 10542 9220 10546 9276
rect 10482 9216 10546 9220
rect 10562 9276 10626 9280
rect 10562 9220 10566 9276
rect 10566 9220 10622 9276
rect 10622 9220 10626 9276
rect 10562 9216 10626 9220
rect 14070 9276 14134 9280
rect 14070 9220 14074 9276
rect 14074 9220 14130 9276
rect 14130 9220 14134 9276
rect 14070 9216 14134 9220
rect 14150 9276 14214 9280
rect 14150 9220 14154 9276
rect 14154 9220 14210 9276
rect 14210 9220 14214 9276
rect 14150 9216 14214 9220
rect 14230 9276 14294 9280
rect 14230 9220 14234 9276
rect 14234 9220 14290 9276
rect 14290 9220 14294 9276
rect 14230 9216 14294 9220
rect 14310 9276 14374 9280
rect 14310 9220 14314 9276
rect 14314 9220 14370 9276
rect 14370 9220 14374 9276
rect 14310 9216 14374 9220
rect 7236 9148 7300 9212
rect 12572 9148 12636 9212
rect 6316 8876 6380 8940
rect 9812 8740 9876 8804
rect 11836 8800 11900 8804
rect 11836 8744 11850 8800
rect 11850 8744 11900 8800
rect 11836 8740 11900 8744
rect 4700 8732 4764 8736
rect 4700 8676 4704 8732
rect 4704 8676 4760 8732
rect 4760 8676 4764 8732
rect 4700 8672 4764 8676
rect 4780 8732 4844 8736
rect 4780 8676 4784 8732
rect 4784 8676 4840 8732
rect 4840 8676 4844 8732
rect 4780 8672 4844 8676
rect 4860 8732 4924 8736
rect 4860 8676 4864 8732
rect 4864 8676 4920 8732
rect 4920 8676 4924 8732
rect 4860 8672 4924 8676
rect 4940 8732 5004 8736
rect 4940 8676 4944 8732
rect 4944 8676 5000 8732
rect 5000 8676 5004 8732
rect 4940 8672 5004 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 12196 8732 12260 8736
rect 12196 8676 12200 8732
rect 12200 8676 12256 8732
rect 12256 8676 12260 8732
rect 12196 8672 12260 8676
rect 12276 8732 12340 8736
rect 12276 8676 12280 8732
rect 12280 8676 12336 8732
rect 12336 8676 12340 8732
rect 12276 8672 12340 8676
rect 12356 8732 12420 8736
rect 12356 8676 12360 8732
rect 12360 8676 12416 8732
rect 12416 8676 12420 8732
rect 12356 8672 12420 8676
rect 12436 8732 12500 8736
rect 12436 8676 12440 8732
rect 12440 8676 12496 8732
rect 12496 8676 12500 8732
rect 12436 8672 12500 8676
rect 12940 8604 13004 8668
rect 5580 8392 5644 8396
rect 5580 8336 5594 8392
rect 5594 8336 5644 8392
rect 5580 8332 5644 8336
rect 6316 8332 6380 8396
rect 11836 8332 11900 8396
rect 13124 8392 13188 8396
rect 13124 8336 13174 8392
rect 13174 8336 13188 8392
rect 13124 8332 13188 8336
rect 13676 8332 13740 8396
rect 3924 8196 3988 8260
rect 2826 8188 2890 8192
rect 2826 8132 2830 8188
rect 2830 8132 2886 8188
rect 2886 8132 2890 8188
rect 2826 8128 2890 8132
rect 2906 8188 2970 8192
rect 2906 8132 2910 8188
rect 2910 8132 2966 8188
rect 2966 8132 2970 8188
rect 2906 8128 2970 8132
rect 2986 8188 3050 8192
rect 2986 8132 2990 8188
rect 2990 8132 3046 8188
rect 3046 8132 3050 8188
rect 2986 8128 3050 8132
rect 3066 8188 3130 8192
rect 3066 8132 3070 8188
rect 3070 8132 3126 8188
rect 3126 8132 3130 8188
rect 3066 8128 3130 8132
rect 3740 8060 3804 8124
rect 5396 8060 5460 8124
rect 7972 8196 8036 8260
rect 11284 8196 11348 8260
rect 12940 8196 13004 8260
rect 6574 8188 6638 8192
rect 6574 8132 6578 8188
rect 6578 8132 6634 8188
rect 6634 8132 6638 8188
rect 6574 8128 6638 8132
rect 6654 8188 6718 8192
rect 6654 8132 6658 8188
rect 6658 8132 6714 8188
rect 6714 8132 6718 8188
rect 6654 8128 6718 8132
rect 6734 8188 6798 8192
rect 6734 8132 6738 8188
rect 6738 8132 6794 8188
rect 6794 8132 6798 8188
rect 6734 8128 6798 8132
rect 6814 8188 6878 8192
rect 6814 8132 6818 8188
rect 6818 8132 6874 8188
rect 6874 8132 6878 8188
rect 6814 8128 6878 8132
rect 10322 8188 10386 8192
rect 10322 8132 10326 8188
rect 10326 8132 10382 8188
rect 10382 8132 10386 8188
rect 10322 8128 10386 8132
rect 10402 8188 10466 8192
rect 10402 8132 10406 8188
rect 10406 8132 10462 8188
rect 10462 8132 10466 8188
rect 10402 8128 10466 8132
rect 10482 8188 10546 8192
rect 10482 8132 10486 8188
rect 10486 8132 10542 8188
rect 10542 8132 10546 8188
rect 10482 8128 10546 8132
rect 10562 8188 10626 8192
rect 10562 8132 10566 8188
rect 10566 8132 10622 8188
rect 10622 8132 10626 8188
rect 10562 8128 10626 8132
rect 8156 8060 8220 8124
rect 9260 8060 9324 8124
rect 12020 8060 12084 8124
rect 12572 8120 12636 8124
rect 14070 8188 14134 8192
rect 14070 8132 14074 8188
rect 14074 8132 14130 8188
rect 14130 8132 14134 8188
rect 14070 8128 14134 8132
rect 14150 8188 14214 8192
rect 14150 8132 14154 8188
rect 14154 8132 14210 8188
rect 14210 8132 14214 8188
rect 14150 8128 14214 8132
rect 14230 8188 14294 8192
rect 14230 8132 14234 8188
rect 14234 8132 14290 8188
rect 14290 8132 14294 8188
rect 14230 8128 14294 8132
rect 14310 8188 14374 8192
rect 14310 8132 14314 8188
rect 14314 8132 14370 8188
rect 14370 8132 14374 8188
rect 14310 8128 14374 8132
rect 12572 8064 12586 8120
rect 12586 8064 12636 8120
rect 12572 8060 12636 8064
rect 14964 8060 15028 8124
rect 15332 8060 15396 8124
rect 1348 7788 1412 7852
rect 5396 7788 5460 7852
rect 3556 7712 3620 7716
rect 3556 7656 3606 7712
rect 3606 7656 3620 7712
rect 3556 7652 3620 7656
rect 9812 7652 9876 7716
rect 4700 7644 4764 7648
rect 4700 7588 4704 7644
rect 4704 7588 4760 7644
rect 4760 7588 4764 7644
rect 4700 7584 4764 7588
rect 4780 7644 4844 7648
rect 4780 7588 4784 7644
rect 4784 7588 4840 7644
rect 4840 7588 4844 7644
rect 4780 7584 4844 7588
rect 4860 7644 4924 7648
rect 4860 7588 4864 7644
rect 4864 7588 4920 7644
rect 4920 7588 4924 7644
rect 4860 7584 4924 7588
rect 4940 7644 5004 7648
rect 4940 7588 4944 7644
rect 4944 7588 5000 7644
rect 5000 7588 5004 7644
rect 4940 7584 5004 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 12196 7644 12260 7648
rect 12196 7588 12200 7644
rect 12200 7588 12256 7644
rect 12256 7588 12260 7644
rect 12196 7584 12260 7588
rect 12276 7644 12340 7648
rect 12276 7588 12280 7644
rect 12280 7588 12336 7644
rect 12336 7588 12340 7644
rect 12276 7584 12340 7588
rect 12356 7644 12420 7648
rect 12356 7588 12360 7644
rect 12360 7588 12416 7644
rect 12416 7588 12420 7644
rect 12356 7584 12420 7588
rect 12436 7644 12500 7648
rect 12436 7588 12440 7644
rect 12440 7588 12496 7644
rect 12496 7588 12500 7644
rect 12436 7584 12500 7588
rect 8892 7516 8956 7580
rect 5948 7380 6012 7444
rect 13308 7516 13372 7580
rect 13676 7576 13740 7580
rect 13676 7520 13726 7576
rect 13726 7520 13740 7576
rect 13676 7516 13740 7520
rect 11468 7244 11532 7308
rect 12572 7244 12636 7308
rect 13124 7244 13188 7308
rect 2826 7100 2890 7104
rect 2826 7044 2830 7100
rect 2830 7044 2886 7100
rect 2886 7044 2890 7100
rect 2826 7040 2890 7044
rect 2906 7100 2970 7104
rect 2906 7044 2910 7100
rect 2910 7044 2966 7100
rect 2966 7044 2970 7100
rect 2906 7040 2970 7044
rect 2986 7100 3050 7104
rect 2986 7044 2990 7100
rect 2990 7044 3046 7100
rect 3046 7044 3050 7100
rect 2986 7040 3050 7044
rect 3066 7100 3130 7104
rect 3066 7044 3070 7100
rect 3070 7044 3126 7100
rect 3126 7044 3130 7100
rect 3066 7040 3130 7044
rect 6574 7100 6638 7104
rect 6574 7044 6578 7100
rect 6578 7044 6634 7100
rect 6634 7044 6638 7100
rect 6574 7040 6638 7044
rect 6654 7100 6718 7104
rect 6654 7044 6658 7100
rect 6658 7044 6714 7100
rect 6714 7044 6718 7100
rect 6654 7040 6718 7044
rect 6734 7100 6798 7104
rect 6734 7044 6738 7100
rect 6738 7044 6794 7100
rect 6794 7044 6798 7100
rect 6734 7040 6798 7044
rect 6814 7100 6878 7104
rect 6814 7044 6818 7100
rect 6818 7044 6874 7100
rect 6874 7044 6878 7100
rect 6814 7040 6878 7044
rect 10322 7100 10386 7104
rect 10322 7044 10326 7100
rect 10326 7044 10382 7100
rect 10382 7044 10386 7100
rect 10322 7040 10386 7044
rect 10402 7100 10466 7104
rect 10402 7044 10406 7100
rect 10406 7044 10462 7100
rect 10462 7044 10466 7100
rect 10402 7040 10466 7044
rect 10482 7100 10546 7104
rect 10482 7044 10486 7100
rect 10486 7044 10542 7100
rect 10542 7044 10546 7100
rect 10482 7040 10546 7044
rect 10562 7100 10626 7104
rect 10562 7044 10566 7100
rect 10566 7044 10622 7100
rect 10622 7044 10626 7100
rect 10562 7040 10626 7044
rect 14070 7100 14134 7104
rect 14070 7044 14074 7100
rect 14074 7044 14130 7100
rect 14130 7044 14134 7100
rect 14070 7040 14134 7044
rect 14150 7100 14214 7104
rect 14150 7044 14154 7100
rect 14154 7044 14210 7100
rect 14210 7044 14214 7100
rect 14150 7040 14214 7044
rect 14230 7100 14294 7104
rect 14230 7044 14234 7100
rect 14234 7044 14290 7100
rect 14290 7044 14294 7100
rect 14230 7040 14294 7044
rect 14310 7100 14374 7104
rect 14310 7044 14314 7100
rect 14314 7044 14370 7100
rect 14370 7044 14374 7100
rect 14310 7040 14374 7044
rect 3740 7032 3804 7036
rect 3740 6976 3790 7032
rect 3790 6976 3804 7032
rect 3740 6972 3804 6976
rect 1716 6896 1780 6900
rect 1716 6840 1766 6896
rect 1766 6840 1780 6896
rect 1716 6836 1780 6840
rect 4476 6896 4540 6900
rect 4476 6840 4490 6896
rect 4490 6840 4540 6896
rect 4476 6836 4540 6840
rect 5764 6836 5828 6900
rect 12020 6836 12084 6900
rect 12756 6972 12820 7036
rect 13492 6972 13556 7036
rect 14964 6836 15028 6900
rect 14964 6760 15028 6764
rect 14964 6704 14978 6760
rect 14978 6704 15028 6760
rect 14964 6700 15028 6704
rect 12756 6564 12820 6628
rect 13860 6564 13924 6628
rect 15516 6564 15580 6628
rect 4700 6556 4764 6560
rect 4700 6500 4704 6556
rect 4704 6500 4760 6556
rect 4760 6500 4764 6556
rect 4700 6496 4764 6500
rect 4780 6556 4844 6560
rect 4780 6500 4784 6556
rect 4784 6500 4840 6556
rect 4840 6500 4844 6556
rect 4780 6496 4844 6500
rect 4860 6556 4924 6560
rect 4860 6500 4864 6556
rect 4864 6500 4920 6556
rect 4920 6500 4924 6556
rect 4860 6496 4924 6500
rect 4940 6556 5004 6560
rect 4940 6500 4944 6556
rect 4944 6500 5000 6556
rect 5000 6500 5004 6556
rect 4940 6496 5004 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 12196 6556 12260 6560
rect 12196 6500 12200 6556
rect 12200 6500 12256 6556
rect 12256 6500 12260 6556
rect 12196 6496 12260 6500
rect 12276 6556 12340 6560
rect 12276 6500 12280 6556
rect 12280 6500 12336 6556
rect 12336 6500 12340 6556
rect 12276 6496 12340 6500
rect 12356 6556 12420 6560
rect 12356 6500 12360 6556
rect 12360 6500 12416 6556
rect 12416 6500 12420 6556
rect 12356 6496 12420 6500
rect 12436 6556 12500 6560
rect 12436 6500 12440 6556
rect 12440 6500 12496 6556
rect 12496 6500 12500 6556
rect 12436 6496 12500 6500
rect 796 6156 860 6220
rect 10916 6428 10980 6492
rect 11100 6488 11164 6492
rect 11100 6432 11150 6488
rect 11150 6432 11164 6488
rect 11100 6428 11164 6432
rect 11284 6428 11348 6492
rect 12756 6428 12820 6492
rect 13860 6428 13924 6492
rect 9996 6292 10060 6356
rect 5580 6020 5644 6084
rect 10916 6020 10980 6084
rect 11100 6080 11164 6084
rect 11100 6024 11114 6080
rect 11114 6024 11164 6080
rect 11100 6020 11164 6024
rect 11284 6020 11348 6084
rect 2826 6012 2890 6016
rect 2826 5956 2830 6012
rect 2830 5956 2886 6012
rect 2886 5956 2890 6012
rect 2826 5952 2890 5956
rect 2906 6012 2970 6016
rect 2906 5956 2910 6012
rect 2910 5956 2966 6012
rect 2966 5956 2970 6012
rect 2906 5952 2970 5956
rect 2986 6012 3050 6016
rect 2986 5956 2990 6012
rect 2990 5956 3046 6012
rect 3046 5956 3050 6012
rect 2986 5952 3050 5956
rect 3066 6012 3130 6016
rect 3066 5956 3070 6012
rect 3070 5956 3126 6012
rect 3126 5956 3130 6012
rect 3066 5952 3130 5956
rect 6574 6012 6638 6016
rect 6574 5956 6578 6012
rect 6578 5956 6634 6012
rect 6634 5956 6638 6012
rect 6574 5952 6638 5956
rect 6654 6012 6718 6016
rect 6654 5956 6658 6012
rect 6658 5956 6714 6012
rect 6714 5956 6718 6012
rect 6654 5952 6718 5956
rect 6734 6012 6798 6016
rect 6734 5956 6738 6012
rect 6738 5956 6794 6012
rect 6794 5956 6798 6012
rect 6734 5952 6798 5956
rect 6814 6012 6878 6016
rect 6814 5956 6818 6012
rect 6818 5956 6874 6012
rect 6874 5956 6878 6012
rect 6814 5952 6878 5956
rect 10322 6012 10386 6016
rect 10322 5956 10326 6012
rect 10326 5956 10382 6012
rect 10382 5956 10386 6012
rect 10322 5952 10386 5956
rect 10402 6012 10466 6016
rect 10402 5956 10406 6012
rect 10406 5956 10462 6012
rect 10462 5956 10466 6012
rect 10402 5952 10466 5956
rect 10482 6012 10546 6016
rect 10482 5956 10486 6012
rect 10486 5956 10542 6012
rect 10542 5956 10546 6012
rect 10482 5952 10546 5956
rect 10562 6012 10626 6016
rect 10562 5956 10566 6012
rect 10566 5956 10622 6012
rect 10622 5956 10626 6012
rect 10562 5952 10626 5956
rect 14070 6012 14134 6016
rect 14070 5956 14074 6012
rect 14074 5956 14130 6012
rect 14130 5956 14134 6012
rect 14070 5952 14134 5956
rect 14150 6012 14214 6016
rect 14150 5956 14154 6012
rect 14154 5956 14210 6012
rect 14210 5956 14214 6012
rect 14150 5952 14214 5956
rect 14230 6012 14294 6016
rect 14230 5956 14234 6012
rect 14234 5956 14290 6012
rect 14290 5956 14294 6012
rect 14230 5952 14294 5956
rect 14310 6012 14374 6016
rect 14310 5956 14314 6012
rect 14314 5956 14370 6012
rect 14370 5956 14374 6012
rect 14310 5952 14374 5956
rect 4476 5884 4540 5948
rect 7788 5884 7852 5948
rect 7972 5884 8036 5948
rect 14780 5884 14844 5948
rect 1348 5748 1412 5812
rect 13308 5808 13372 5812
rect 13308 5752 13358 5808
rect 13358 5752 13372 5808
rect 13308 5748 13372 5752
rect 2268 5672 2332 5676
rect 2268 5616 2318 5672
rect 2318 5616 2332 5672
rect 2268 5612 2332 5616
rect 6132 5612 6196 5676
rect 9628 5612 9692 5676
rect 10180 5612 10244 5676
rect 10732 5476 10796 5540
rect 4700 5468 4764 5472
rect 4700 5412 4704 5468
rect 4704 5412 4760 5468
rect 4760 5412 4764 5468
rect 4700 5408 4764 5412
rect 4780 5468 4844 5472
rect 4780 5412 4784 5468
rect 4784 5412 4840 5468
rect 4840 5412 4844 5468
rect 4780 5408 4844 5412
rect 4860 5468 4924 5472
rect 4860 5412 4864 5468
rect 4864 5412 4920 5468
rect 4920 5412 4924 5468
rect 4860 5408 4924 5412
rect 4940 5468 5004 5472
rect 4940 5412 4944 5468
rect 4944 5412 5000 5468
rect 5000 5412 5004 5468
rect 4940 5408 5004 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 5212 5340 5276 5404
rect 11652 5400 11716 5404
rect 11652 5344 11666 5400
rect 11666 5344 11716 5400
rect 11652 5340 11716 5344
rect 10180 5068 10244 5132
rect 10732 5204 10796 5268
rect 11100 5204 11164 5268
rect 13308 5476 13372 5540
rect 13676 5476 13740 5540
rect 14780 5536 14844 5540
rect 14780 5480 14830 5536
rect 14830 5480 14844 5536
rect 14780 5476 14844 5480
rect 12196 5468 12260 5472
rect 12196 5412 12200 5468
rect 12200 5412 12256 5468
rect 12256 5412 12260 5468
rect 12196 5408 12260 5412
rect 12276 5468 12340 5472
rect 12276 5412 12280 5468
rect 12280 5412 12336 5468
rect 12336 5412 12340 5468
rect 12276 5408 12340 5412
rect 12356 5468 12420 5472
rect 12356 5412 12360 5468
rect 12360 5412 12416 5468
rect 12416 5412 12420 5468
rect 12356 5408 12420 5412
rect 12436 5468 12500 5472
rect 12436 5412 12440 5468
rect 12440 5412 12496 5468
rect 12496 5412 12500 5468
rect 12436 5408 12500 5412
rect 12756 5340 12820 5404
rect 15516 5264 15580 5268
rect 15516 5208 15530 5264
rect 15530 5208 15580 5264
rect 15516 5204 15580 5208
rect 15148 5068 15212 5132
rect 9628 4932 9692 4996
rect 11100 4932 11164 4996
rect 2826 4924 2890 4928
rect 2826 4868 2830 4924
rect 2830 4868 2886 4924
rect 2886 4868 2890 4924
rect 2826 4864 2890 4868
rect 2906 4924 2970 4928
rect 2906 4868 2910 4924
rect 2910 4868 2966 4924
rect 2966 4868 2970 4924
rect 2906 4864 2970 4868
rect 2986 4924 3050 4928
rect 2986 4868 2990 4924
rect 2990 4868 3046 4924
rect 3046 4868 3050 4924
rect 2986 4864 3050 4868
rect 3066 4924 3130 4928
rect 3066 4868 3070 4924
rect 3070 4868 3126 4924
rect 3126 4868 3130 4924
rect 3066 4864 3130 4868
rect 6574 4924 6638 4928
rect 6574 4868 6578 4924
rect 6578 4868 6634 4924
rect 6634 4868 6638 4924
rect 6574 4864 6638 4868
rect 6654 4924 6718 4928
rect 6654 4868 6658 4924
rect 6658 4868 6714 4924
rect 6714 4868 6718 4924
rect 6654 4864 6718 4868
rect 6734 4924 6798 4928
rect 6734 4868 6738 4924
rect 6738 4868 6794 4924
rect 6794 4868 6798 4924
rect 6734 4864 6798 4868
rect 6814 4924 6878 4928
rect 6814 4868 6818 4924
rect 6818 4868 6874 4924
rect 6874 4868 6878 4924
rect 6814 4864 6878 4868
rect 10322 4924 10386 4928
rect 10322 4868 10326 4924
rect 10326 4868 10382 4924
rect 10382 4868 10386 4924
rect 10322 4864 10386 4868
rect 10402 4924 10466 4928
rect 10402 4868 10406 4924
rect 10406 4868 10462 4924
rect 10462 4868 10466 4924
rect 10402 4864 10466 4868
rect 10482 4924 10546 4928
rect 10482 4868 10486 4924
rect 10486 4868 10542 4924
rect 10542 4868 10546 4924
rect 10482 4864 10546 4868
rect 10562 4924 10626 4928
rect 10562 4868 10566 4924
rect 10566 4868 10622 4924
rect 10622 4868 10626 4924
rect 10562 4864 10626 4868
rect 9628 4796 9692 4860
rect 13492 4932 13556 4996
rect 14070 4924 14134 4928
rect 14070 4868 14074 4924
rect 14074 4868 14130 4924
rect 14130 4868 14134 4924
rect 14070 4864 14134 4868
rect 14150 4924 14214 4928
rect 14150 4868 14154 4924
rect 14154 4868 14210 4924
rect 14210 4868 14214 4924
rect 14150 4864 14214 4868
rect 14230 4924 14294 4928
rect 14230 4868 14234 4924
rect 14234 4868 14290 4924
rect 14290 4868 14294 4924
rect 14230 4864 14294 4868
rect 14310 4924 14374 4928
rect 14310 4868 14314 4924
rect 14314 4868 14370 4924
rect 14370 4868 14374 4924
rect 14310 4864 14374 4868
rect 980 4660 1044 4724
rect 10180 4524 10244 4588
rect 11468 4524 11532 4588
rect 3372 4388 3436 4452
rect 12756 4388 12820 4452
rect 4700 4380 4764 4384
rect 4700 4324 4704 4380
rect 4704 4324 4760 4380
rect 4760 4324 4764 4380
rect 4700 4320 4764 4324
rect 4780 4380 4844 4384
rect 4780 4324 4784 4380
rect 4784 4324 4840 4380
rect 4840 4324 4844 4380
rect 4780 4320 4844 4324
rect 4860 4380 4924 4384
rect 4860 4324 4864 4380
rect 4864 4324 4920 4380
rect 4920 4324 4924 4380
rect 4860 4320 4924 4324
rect 4940 4380 5004 4384
rect 4940 4324 4944 4380
rect 4944 4324 5000 4380
rect 5000 4324 5004 4380
rect 4940 4320 5004 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 12196 4380 12260 4384
rect 12196 4324 12200 4380
rect 12200 4324 12256 4380
rect 12256 4324 12260 4380
rect 12196 4320 12260 4324
rect 12276 4380 12340 4384
rect 12276 4324 12280 4380
rect 12280 4324 12336 4380
rect 12336 4324 12340 4380
rect 12276 4320 12340 4324
rect 12356 4380 12420 4384
rect 12356 4324 12360 4380
rect 12360 4324 12416 4380
rect 12416 4324 12420 4380
rect 12356 4320 12420 4324
rect 12436 4380 12500 4384
rect 12436 4324 12440 4380
rect 12440 4324 12496 4380
rect 12496 4324 12500 4380
rect 12436 4320 12500 4324
rect 7604 4252 7668 4316
rect 10916 4116 10980 4180
rect 11468 4116 11532 4180
rect 12572 4116 12636 4180
rect 1532 3980 1596 4044
rect 5396 3980 5460 4044
rect 7052 3980 7116 4044
rect 15332 4252 15396 4316
rect 13308 4116 13372 4180
rect 14964 4040 15028 4044
rect 14964 3984 14978 4040
rect 14978 3984 15028 4040
rect 14964 3980 15028 3984
rect 2826 3836 2890 3840
rect 2826 3780 2830 3836
rect 2830 3780 2886 3836
rect 2886 3780 2890 3836
rect 2826 3776 2890 3780
rect 2906 3836 2970 3840
rect 2906 3780 2910 3836
rect 2910 3780 2966 3836
rect 2966 3780 2970 3836
rect 2906 3776 2970 3780
rect 2986 3836 3050 3840
rect 2986 3780 2990 3836
rect 2990 3780 3046 3836
rect 3046 3780 3050 3836
rect 2986 3776 3050 3780
rect 3066 3836 3130 3840
rect 3066 3780 3070 3836
rect 3070 3780 3126 3836
rect 3126 3780 3130 3836
rect 3066 3776 3130 3780
rect 6574 3836 6638 3840
rect 6574 3780 6578 3836
rect 6578 3780 6634 3836
rect 6634 3780 6638 3836
rect 6574 3776 6638 3780
rect 6654 3836 6718 3840
rect 6654 3780 6658 3836
rect 6658 3780 6714 3836
rect 6714 3780 6718 3836
rect 6654 3776 6718 3780
rect 6734 3836 6798 3840
rect 6734 3780 6738 3836
rect 6738 3780 6794 3836
rect 6794 3780 6798 3836
rect 6734 3776 6798 3780
rect 6814 3836 6878 3840
rect 6814 3780 6818 3836
rect 6818 3780 6874 3836
rect 6874 3780 6878 3836
rect 6814 3776 6878 3780
rect 10322 3836 10386 3840
rect 10322 3780 10326 3836
rect 10326 3780 10382 3836
rect 10382 3780 10386 3836
rect 10322 3776 10386 3780
rect 10402 3836 10466 3840
rect 10402 3780 10406 3836
rect 10406 3780 10462 3836
rect 10462 3780 10466 3836
rect 10402 3776 10466 3780
rect 10482 3836 10546 3840
rect 10482 3780 10486 3836
rect 10486 3780 10542 3836
rect 10542 3780 10546 3836
rect 10482 3776 10546 3780
rect 10562 3836 10626 3840
rect 10562 3780 10566 3836
rect 10566 3780 10622 3836
rect 10622 3780 10626 3836
rect 10562 3776 10626 3780
rect 14070 3836 14134 3840
rect 14070 3780 14074 3836
rect 14074 3780 14130 3836
rect 14130 3780 14134 3836
rect 14070 3776 14134 3780
rect 14150 3836 14214 3840
rect 14150 3780 14154 3836
rect 14154 3780 14210 3836
rect 14210 3780 14214 3836
rect 14150 3776 14214 3780
rect 14230 3836 14294 3840
rect 14230 3780 14234 3836
rect 14234 3780 14290 3836
rect 14290 3780 14294 3836
rect 14230 3776 14294 3780
rect 14310 3836 14374 3840
rect 14310 3780 14314 3836
rect 14314 3780 14370 3836
rect 14370 3780 14374 3836
rect 14310 3776 14374 3780
rect 8156 3708 8220 3772
rect 9996 3708 10060 3772
rect 12020 3708 12084 3772
rect 9260 3572 9324 3636
rect 11468 3436 11532 3500
rect 11652 3436 11716 3500
rect 4700 3292 4764 3296
rect 4700 3236 4704 3292
rect 4704 3236 4760 3292
rect 4760 3236 4764 3292
rect 4700 3232 4764 3236
rect 4780 3292 4844 3296
rect 4780 3236 4784 3292
rect 4784 3236 4840 3292
rect 4840 3236 4844 3292
rect 4780 3232 4844 3236
rect 4860 3292 4924 3296
rect 4860 3236 4864 3292
rect 4864 3236 4920 3292
rect 4920 3236 4924 3292
rect 4860 3232 4924 3236
rect 4940 3292 5004 3296
rect 4940 3236 4944 3292
rect 4944 3236 5000 3292
rect 5000 3236 5004 3292
rect 4940 3232 5004 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 12196 3292 12260 3296
rect 12196 3236 12200 3292
rect 12200 3236 12256 3292
rect 12256 3236 12260 3292
rect 12196 3232 12260 3236
rect 12276 3292 12340 3296
rect 12276 3236 12280 3292
rect 12280 3236 12336 3292
rect 12336 3236 12340 3292
rect 12276 3232 12340 3236
rect 12356 3292 12420 3296
rect 12356 3236 12360 3292
rect 12360 3236 12416 3292
rect 12416 3236 12420 3292
rect 12356 3232 12420 3236
rect 12436 3292 12500 3296
rect 12436 3236 12440 3292
rect 12440 3236 12496 3292
rect 12496 3236 12500 3292
rect 12436 3232 12500 3236
rect 5948 3224 6012 3228
rect 5948 3168 5962 3224
rect 5962 3168 6012 3224
rect 5948 3164 6012 3168
rect 7236 3164 7300 3228
rect 9996 3164 10060 3228
rect 11468 3164 11532 3228
rect 2452 3028 2516 3092
rect 8892 2892 8956 2956
rect 12940 3028 13004 3092
rect 9628 2892 9692 2956
rect 4476 2756 4540 2820
rect 7420 2756 7484 2820
rect 9996 2756 10060 2820
rect 10732 2816 10796 2820
rect 13492 3164 13556 3228
rect 10732 2760 10782 2816
rect 10782 2760 10796 2816
rect 10732 2756 10796 2760
rect 2826 2748 2890 2752
rect 2826 2692 2830 2748
rect 2830 2692 2886 2748
rect 2886 2692 2890 2748
rect 2826 2688 2890 2692
rect 2906 2748 2970 2752
rect 2906 2692 2910 2748
rect 2910 2692 2966 2748
rect 2966 2692 2970 2748
rect 2906 2688 2970 2692
rect 2986 2748 3050 2752
rect 2986 2692 2990 2748
rect 2990 2692 3046 2748
rect 3046 2692 3050 2748
rect 2986 2688 3050 2692
rect 3066 2748 3130 2752
rect 3066 2692 3070 2748
rect 3070 2692 3126 2748
rect 3126 2692 3130 2748
rect 3066 2688 3130 2692
rect 6574 2748 6638 2752
rect 6574 2692 6578 2748
rect 6578 2692 6634 2748
rect 6634 2692 6638 2748
rect 6574 2688 6638 2692
rect 6654 2748 6718 2752
rect 6654 2692 6658 2748
rect 6658 2692 6714 2748
rect 6714 2692 6718 2748
rect 6654 2688 6718 2692
rect 6734 2748 6798 2752
rect 6734 2692 6738 2748
rect 6738 2692 6794 2748
rect 6794 2692 6798 2748
rect 6734 2688 6798 2692
rect 6814 2748 6878 2752
rect 6814 2692 6818 2748
rect 6818 2692 6874 2748
rect 6874 2692 6878 2748
rect 6814 2688 6878 2692
rect 10322 2748 10386 2752
rect 10322 2692 10326 2748
rect 10326 2692 10382 2748
rect 10382 2692 10386 2748
rect 10322 2688 10386 2692
rect 10402 2748 10466 2752
rect 10402 2692 10406 2748
rect 10406 2692 10462 2748
rect 10462 2692 10466 2748
rect 10402 2688 10466 2692
rect 10482 2748 10546 2752
rect 10482 2692 10486 2748
rect 10486 2692 10542 2748
rect 10542 2692 10546 2748
rect 10482 2688 10546 2692
rect 10562 2748 10626 2752
rect 10562 2692 10566 2748
rect 10566 2692 10622 2748
rect 10622 2692 10626 2748
rect 10562 2688 10626 2692
rect 1900 2620 1964 2684
rect 1348 2484 1412 2548
rect 2268 2544 2332 2548
rect 5212 2620 5276 2684
rect 6316 2620 6380 2684
rect 9076 2620 9140 2684
rect 15148 3028 15212 3092
rect 14596 2892 14660 2956
rect 14070 2748 14134 2752
rect 14070 2692 14074 2748
rect 14074 2692 14130 2748
rect 14130 2692 14134 2748
rect 14070 2688 14134 2692
rect 14150 2748 14214 2752
rect 14150 2692 14154 2748
rect 14154 2692 14210 2748
rect 14210 2692 14214 2748
rect 14150 2688 14214 2692
rect 14230 2748 14294 2752
rect 14230 2692 14234 2748
rect 14234 2692 14290 2748
rect 14290 2692 14294 2748
rect 14230 2688 14294 2692
rect 14310 2748 14374 2752
rect 14310 2692 14314 2748
rect 14314 2692 14370 2748
rect 14370 2692 14374 2748
rect 14310 2688 14374 2692
rect 2268 2488 2318 2544
rect 2318 2488 2332 2544
rect 2268 2484 2332 2488
rect 5764 2544 5828 2548
rect 5764 2488 5814 2544
rect 5814 2488 5828 2544
rect 5764 2484 5828 2488
rect 7236 2484 7300 2548
rect 9260 2544 9324 2548
rect 9260 2488 9310 2544
rect 9310 2488 9324 2544
rect 9260 2484 9324 2488
rect 9812 2484 9876 2548
rect 11468 2484 11532 2548
rect 5580 2212 5644 2276
rect 7972 2272 8036 2276
rect 7972 2216 7986 2272
rect 7986 2216 8036 2272
rect 7972 2212 8036 2216
rect 13860 2348 13924 2412
rect 4700 2204 4764 2208
rect 4700 2148 4704 2204
rect 4704 2148 4760 2204
rect 4760 2148 4764 2204
rect 4700 2144 4764 2148
rect 4780 2204 4844 2208
rect 4780 2148 4784 2204
rect 4784 2148 4840 2204
rect 4840 2148 4844 2204
rect 4780 2144 4844 2148
rect 4860 2204 4924 2208
rect 4860 2148 4864 2204
rect 4864 2148 4920 2204
rect 4920 2148 4924 2204
rect 4860 2144 4924 2148
rect 4940 2204 5004 2208
rect 4940 2148 4944 2204
rect 4944 2148 5000 2204
rect 5000 2148 5004 2204
rect 4940 2144 5004 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 12196 2204 12260 2208
rect 12196 2148 12200 2204
rect 12200 2148 12256 2204
rect 12256 2148 12260 2204
rect 12196 2144 12260 2148
rect 12276 2204 12340 2208
rect 12276 2148 12280 2204
rect 12280 2148 12336 2204
rect 12336 2148 12340 2204
rect 12276 2144 12340 2148
rect 12356 2204 12420 2208
rect 12356 2148 12360 2204
rect 12360 2148 12416 2204
rect 12416 2148 12420 2204
rect 12356 2144 12420 2148
rect 12436 2204 12500 2208
rect 12436 2148 12440 2204
rect 12440 2148 12496 2204
rect 12496 2148 12500 2204
rect 12436 2144 12500 2148
rect 10916 2076 10980 2140
rect 7788 1940 7852 2004
rect 11836 1940 11900 2004
rect 11468 1804 11532 1868
rect 7604 1668 7668 1732
rect 12940 1532 13004 1596
rect 13676 1396 13740 1460
rect 1164 1260 1228 1324
rect 14780 1260 14844 1324
rect 3372 1124 3436 1188
rect 7052 852 7116 916
rect 6132 716 6196 780
rect 13308 580 13372 644
rect 12756 172 12820 236
<< metal4 >>
rect 4107 18324 4173 18325
rect 4107 18260 4108 18324
rect 4172 18260 4173 18324
rect 4107 18259 4173 18260
rect 2635 17236 2701 17237
rect 2635 17172 2636 17236
rect 2700 17172 2701 17236
rect 2635 17171 2701 17172
rect 1163 15876 1229 15877
rect 1163 15812 1164 15876
rect 1228 15812 1229 15876
rect 1163 15811 1229 15812
rect 979 14652 1045 14653
rect 979 14588 980 14652
rect 1044 14588 1045 14652
rect 979 14587 1045 14588
rect 795 12068 861 12069
rect 795 12004 796 12068
rect 860 12004 861 12068
rect 795 12003 861 12004
rect 798 6221 858 12003
rect 795 6220 861 6221
rect 795 6156 796 6220
rect 860 6156 861 6220
rect 795 6155 861 6156
rect 982 4725 1042 14587
rect 1166 12069 1226 15811
rect 1347 15740 1413 15741
rect 1347 15676 1348 15740
rect 1412 15676 1413 15740
rect 1347 15675 1413 15676
rect 1163 12068 1229 12069
rect 1163 12004 1164 12068
rect 1228 12004 1229 12068
rect 1163 12003 1229 12004
rect 1163 11932 1229 11933
rect 1163 11868 1164 11932
rect 1228 11868 1229 11932
rect 1163 11867 1229 11868
rect 979 4724 1045 4725
rect 979 4660 980 4724
rect 1044 4660 1045 4724
rect 979 4659 1045 4660
rect 1166 1325 1226 11867
rect 1350 7853 1410 15675
rect 1715 14516 1781 14517
rect 1715 14452 1716 14516
rect 1780 14452 1781 14516
rect 1715 14451 1781 14452
rect 1531 14244 1597 14245
rect 1531 14180 1532 14244
rect 1596 14180 1597 14244
rect 1531 14179 1597 14180
rect 1347 7852 1413 7853
rect 1347 7788 1348 7852
rect 1412 7788 1413 7852
rect 1347 7787 1413 7788
rect 1347 5812 1413 5813
rect 1347 5748 1348 5812
rect 1412 5748 1413 5812
rect 1347 5747 1413 5748
rect 1350 2549 1410 5747
rect 1534 4045 1594 14179
rect 1718 6901 1778 14451
rect 2451 12612 2517 12613
rect 2451 12548 2452 12612
rect 2516 12548 2517 12612
rect 2451 12547 2517 12548
rect 1899 11116 1965 11117
rect 1899 11052 1900 11116
rect 1964 11052 1965 11116
rect 1899 11051 1965 11052
rect 1715 6900 1781 6901
rect 1715 6836 1716 6900
rect 1780 6836 1781 6900
rect 1715 6835 1781 6836
rect 1531 4044 1597 4045
rect 1531 3980 1532 4044
rect 1596 3980 1597 4044
rect 1531 3979 1597 3980
rect 1902 2685 1962 11051
rect 2267 5676 2333 5677
rect 2267 5612 2268 5676
rect 2332 5612 2333 5676
rect 2267 5611 2333 5612
rect 1899 2684 1965 2685
rect 1899 2620 1900 2684
rect 1964 2620 1965 2684
rect 1899 2619 1965 2620
rect 2270 2549 2330 5611
rect 2454 3093 2514 12547
rect 2638 11933 2698 17171
rect 2818 16896 3138 17456
rect 2818 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3138 16896
rect 2818 15808 3138 16832
rect 2818 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3138 15808
rect 2818 14720 3138 15744
rect 2818 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3138 14720
rect 2818 13632 3138 14656
rect 3371 14652 3437 14653
rect 3371 14588 3372 14652
rect 3436 14588 3437 14652
rect 3371 14587 3437 14588
rect 2818 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3138 13632
rect 2818 12544 3138 13568
rect 2818 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3138 12544
rect 2635 11932 2701 11933
rect 2635 11868 2636 11932
rect 2700 11868 2701 11932
rect 2635 11867 2701 11868
rect 2818 11456 3138 12480
rect 2818 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3138 11456
rect 2818 10368 3138 11392
rect 3374 10845 3434 14587
rect 4110 14381 4170 18259
rect 10731 18052 10797 18053
rect 10731 17988 10732 18052
rect 10796 17988 10797 18052
rect 10731 17987 10797 17988
rect 7787 17508 7853 17509
rect 4692 17440 5012 17456
rect 4692 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5012 17440
rect 4291 16692 4357 16693
rect 4291 16628 4292 16692
rect 4356 16628 4357 16692
rect 4291 16627 4357 16628
rect 4107 14380 4173 14381
rect 4107 14316 4108 14380
rect 4172 14316 4173 14380
rect 4107 14315 4173 14316
rect 3923 14108 3989 14109
rect 3923 14044 3924 14108
rect 3988 14044 3989 14108
rect 3923 14043 3989 14044
rect 3739 13836 3805 13837
rect 3739 13772 3740 13836
rect 3804 13772 3805 13836
rect 3739 13771 3805 13772
rect 3555 12476 3621 12477
rect 3555 12412 3556 12476
rect 3620 12412 3621 12476
rect 3555 12411 3621 12412
rect 3558 11661 3618 12411
rect 3555 11660 3621 11661
rect 3555 11596 3556 11660
rect 3620 11596 3621 11660
rect 3555 11595 3621 11596
rect 3371 10844 3437 10845
rect 3371 10780 3372 10844
rect 3436 10780 3437 10844
rect 3371 10779 3437 10780
rect 2818 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3138 10368
rect 2818 9280 3138 10304
rect 2818 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3138 9280
rect 2818 8192 3138 9216
rect 2818 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3138 8192
rect 2818 7104 3138 8128
rect 3558 7717 3618 11595
rect 3742 8125 3802 13771
rect 3926 8261 3986 14043
rect 4107 13836 4173 13837
rect 4107 13772 4108 13836
rect 4172 13772 4173 13836
rect 4107 13771 4173 13772
rect 4110 9893 4170 13771
rect 4294 13429 4354 16627
rect 4692 16352 5012 17376
rect 4692 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5012 16352
rect 4475 15740 4541 15741
rect 4475 15676 4476 15740
rect 4540 15676 4541 15740
rect 4475 15675 4541 15676
rect 4291 13428 4357 13429
rect 4291 13364 4292 13428
rect 4356 13364 4357 13428
rect 4291 13363 4357 13364
rect 4478 11389 4538 15675
rect 4692 15264 5012 16288
rect 6566 16896 6886 17456
rect 7787 17444 7788 17508
rect 7852 17444 7853 17508
rect 7787 17443 7853 17444
rect 6566 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6886 16896
rect 6566 15808 6886 16832
rect 7051 16012 7117 16013
rect 7051 15948 7052 16012
rect 7116 15948 7117 16012
rect 7051 15947 7117 15948
rect 6566 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6886 15808
rect 5395 15468 5461 15469
rect 5395 15404 5396 15468
rect 5460 15404 5461 15468
rect 5395 15403 5461 15404
rect 4692 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5012 15264
rect 4692 14176 5012 15200
rect 4692 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5012 14176
rect 4692 13088 5012 14112
rect 4692 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5012 13088
rect 4692 12000 5012 13024
rect 5398 13021 5458 15403
rect 5763 14788 5829 14789
rect 5763 14724 5764 14788
rect 5828 14724 5829 14788
rect 5763 14723 5829 14724
rect 5579 13836 5645 13837
rect 5579 13772 5580 13836
rect 5644 13772 5645 13836
rect 5579 13771 5645 13772
rect 5395 13020 5461 13021
rect 5395 12956 5396 13020
rect 5460 12956 5461 13020
rect 5395 12955 5461 12956
rect 5395 12748 5461 12749
rect 5395 12684 5396 12748
rect 5460 12684 5461 12748
rect 5395 12683 5461 12684
rect 5211 12612 5277 12613
rect 5211 12548 5212 12612
rect 5276 12548 5277 12612
rect 5211 12547 5277 12548
rect 5214 12341 5274 12547
rect 5211 12340 5277 12341
rect 5211 12276 5212 12340
rect 5276 12276 5277 12340
rect 5211 12275 5277 12276
rect 4692 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5012 12000
rect 4475 11388 4541 11389
rect 4475 11324 4476 11388
rect 4540 11324 4541 11388
rect 4475 11323 4541 11324
rect 4692 10912 5012 11936
rect 4692 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5012 10912
rect 4107 9892 4173 9893
rect 4107 9828 4108 9892
rect 4172 9828 4173 9892
rect 4107 9827 4173 9828
rect 4475 9892 4541 9893
rect 4475 9828 4476 9892
rect 4540 9828 4541 9892
rect 4475 9827 4541 9828
rect 3923 8260 3989 8261
rect 3923 8196 3924 8260
rect 3988 8196 3989 8260
rect 3923 8195 3989 8196
rect 3739 8124 3805 8125
rect 3739 8060 3740 8124
rect 3804 8060 3805 8124
rect 3739 8059 3805 8060
rect 3555 7716 3621 7717
rect 3555 7652 3556 7716
rect 3620 7652 3621 7716
rect 3555 7651 3621 7652
rect 2818 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3138 7104
rect 2818 6016 3138 7040
rect 3742 7037 3802 8059
rect 3739 7036 3805 7037
rect 3739 6972 3740 7036
rect 3804 6972 3805 7036
rect 3739 6971 3805 6972
rect 4478 6901 4538 9827
rect 4692 9824 5012 10848
rect 4692 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5012 9824
rect 4692 8736 5012 9760
rect 4692 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5012 8736
rect 4692 7648 5012 8672
rect 5398 8125 5458 12683
rect 5582 8397 5642 13771
rect 5766 12069 5826 14723
rect 6566 14720 6886 15744
rect 6566 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6886 14720
rect 6566 13632 6886 14656
rect 6566 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6886 13632
rect 6566 12544 6886 13568
rect 6566 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6886 12544
rect 5763 12068 5829 12069
rect 5763 12004 5764 12068
rect 5828 12066 5829 12068
rect 5828 12006 6194 12066
rect 5828 12004 5829 12006
rect 5763 12003 5829 12004
rect 5579 8396 5645 8397
rect 5579 8332 5580 8396
rect 5644 8332 5645 8396
rect 5579 8331 5645 8332
rect 5395 8124 5461 8125
rect 5395 8060 5396 8124
rect 5460 8060 5461 8124
rect 5395 8059 5461 8060
rect 5395 7852 5461 7853
rect 5395 7788 5396 7852
rect 5460 7788 5461 7852
rect 5395 7787 5461 7788
rect 4692 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5012 7648
rect 4475 6900 4541 6901
rect 4475 6836 4476 6900
rect 4540 6836 4541 6900
rect 4475 6835 4541 6836
rect 2818 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3138 6016
rect 2818 4928 3138 5952
rect 4692 6560 5012 7584
rect 4692 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5012 6560
rect 4475 5948 4541 5949
rect 4475 5884 4476 5948
rect 4540 5884 4541 5948
rect 4475 5883 4541 5884
rect 2818 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3138 4928
rect 2818 3840 3138 4864
rect 3371 4452 3437 4453
rect 3371 4388 3372 4452
rect 3436 4388 3437 4452
rect 3371 4387 3437 4388
rect 2818 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3138 3840
rect 2451 3092 2517 3093
rect 2451 3028 2452 3092
rect 2516 3028 2517 3092
rect 2451 3027 2517 3028
rect 2818 2752 3138 3776
rect 2818 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3138 2752
rect 1347 2548 1413 2549
rect 1347 2484 1348 2548
rect 1412 2484 1413 2548
rect 1347 2483 1413 2484
rect 2267 2548 2333 2549
rect 2267 2484 2268 2548
rect 2332 2484 2333 2548
rect 2267 2483 2333 2484
rect 2818 2128 3138 2688
rect 1163 1324 1229 1325
rect 1163 1260 1164 1324
rect 1228 1260 1229 1324
rect 1163 1259 1229 1260
rect 3374 1189 3434 4387
rect 4478 2821 4538 5883
rect 4692 5472 5012 6496
rect 4692 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5012 5472
rect 4692 4384 5012 5408
rect 5211 5404 5277 5405
rect 5211 5340 5212 5404
rect 5276 5340 5277 5404
rect 5211 5339 5277 5340
rect 4692 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5012 4384
rect 4692 3296 5012 4320
rect 4692 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5012 3296
rect 4475 2820 4541 2821
rect 4475 2756 4476 2820
rect 4540 2756 4541 2820
rect 4475 2755 4541 2756
rect 4692 2208 5012 3232
rect 5214 2685 5274 5339
rect 5398 4045 5458 7787
rect 5947 7444 6013 7445
rect 5947 7380 5948 7444
rect 6012 7380 6013 7444
rect 5947 7379 6013 7380
rect 5763 6900 5829 6901
rect 5763 6836 5764 6900
rect 5828 6836 5829 6900
rect 5763 6835 5829 6836
rect 5579 6084 5645 6085
rect 5579 6020 5580 6084
rect 5644 6020 5645 6084
rect 5579 6019 5645 6020
rect 5395 4044 5461 4045
rect 5395 3980 5396 4044
rect 5460 3980 5461 4044
rect 5395 3979 5461 3980
rect 5211 2684 5277 2685
rect 5211 2620 5212 2684
rect 5276 2620 5277 2684
rect 5211 2619 5277 2620
rect 5582 2277 5642 6019
rect 5766 2549 5826 6835
rect 5950 3229 6010 7379
rect 6134 5677 6194 12006
rect 6566 11456 6886 12480
rect 6566 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6886 11456
rect 6315 11388 6381 11389
rect 6315 11324 6316 11388
rect 6380 11324 6381 11388
rect 6315 11323 6381 11324
rect 6318 8941 6378 11323
rect 6566 10368 6886 11392
rect 6566 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6886 10368
rect 6566 9280 6886 10304
rect 6566 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6886 9280
rect 6315 8940 6381 8941
rect 6315 8876 6316 8940
rect 6380 8876 6381 8940
rect 6315 8875 6381 8876
rect 6315 8396 6381 8397
rect 6315 8332 6316 8396
rect 6380 8332 6381 8396
rect 6315 8331 6381 8332
rect 6131 5676 6197 5677
rect 6131 5612 6132 5676
rect 6196 5612 6197 5676
rect 6131 5611 6197 5612
rect 5947 3228 6013 3229
rect 5947 3164 5948 3228
rect 6012 3164 6013 3228
rect 5947 3163 6013 3164
rect 5763 2548 5829 2549
rect 5763 2484 5764 2548
rect 5828 2484 5829 2548
rect 5763 2483 5829 2484
rect 5579 2276 5645 2277
rect 5579 2212 5580 2276
rect 5644 2212 5645 2276
rect 5579 2211 5645 2212
rect 4692 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5012 2208
rect 4692 2128 5012 2144
rect 3371 1188 3437 1189
rect 3371 1124 3372 1188
rect 3436 1124 3437 1188
rect 3371 1123 3437 1124
rect 6134 781 6194 5611
rect 6318 2685 6378 8331
rect 6566 8192 6886 9216
rect 6566 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6886 8192
rect 6566 7104 6886 8128
rect 6566 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6886 7104
rect 6566 6016 6886 7040
rect 6566 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6886 6016
rect 6566 4928 6886 5952
rect 6566 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6886 4928
rect 6566 3840 6886 4864
rect 7054 4045 7114 15947
rect 7603 14244 7669 14245
rect 7603 14180 7604 14244
rect 7668 14180 7669 14244
rect 7603 14179 7669 14180
rect 7235 13020 7301 13021
rect 7235 12956 7236 13020
rect 7300 12956 7301 13020
rect 7235 12955 7301 12956
rect 7238 9349 7298 12955
rect 7419 11932 7485 11933
rect 7419 11868 7420 11932
rect 7484 11868 7485 11932
rect 7419 11867 7485 11868
rect 7422 10845 7482 11867
rect 7606 11525 7666 14179
rect 7790 12341 7850 17443
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 15264 8760 16288
rect 10314 16896 10634 17456
rect 10314 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10634 16896
rect 9075 16148 9141 16149
rect 9075 16084 9076 16148
rect 9140 16084 9141 16148
rect 9075 16083 9141 16084
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 7971 15060 8037 15061
rect 7971 14996 7972 15060
rect 8036 14996 8037 15060
rect 7971 14995 8037 14996
rect 7787 12340 7853 12341
rect 7787 12276 7788 12340
rect 7852 12276 7853 12340
rect 7787 12275 7853 12276
rect 7787 11796 7853 11797
rect 7787 11732 7788 11796
rect 7852 11794 7853 11796
rect 7974 11794 8034 14995
rect 8440 14176 8760 15200
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 9078 13830 9138 16083
rect 10314 15808 10634 16832
rect 10314 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10634 15808
rect 9811 15740 9877 15741
rect 9811 15676 9812 15740
rect 9876 15676 9877 15740
rect 9811 15675 9877 15676
rect 9259 14788 9325 14789
rect 9259 14724 9260 14788
rect 9324 14724 9325 14788
rect 9259 14723 9325 14724
rect 9262 14109 9322 14723
rect 9259 14108 9325 14109
rect 9259 14044 9260 14108
rect 9324 14044 9325 14108
rect 9259 14043 9325 14044
rect 9627 13836 9693 13837
rect 9078 13770 9322 13830
rect 9627 13772 9628 13836
rect 9692 13772 9693 13836
rect 9627 13771 9693 13772
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8155 12612 8221 12613
rect 8155 12548 8156 12612
rect 8220 12548 8221 12612
rect 8155 12547 8221 12548
rect 7852 11734 8034 11794
rect 7852 11732 7853 11734
rect 7787 11731 7853 11732
rect 7603 11524 7669 11525
rect 7603 11460 7604 11524
rect 7668 11460 7669 11524
rect 7603 11459 7669 11460
rect 7419 10844 7485 10845
rect 7419 10780 7420 10844
rect 7484 10780 7485 10844
rect 7419 10779 7485 10780
rect 7419 9620 7485 9621
rect 7419 9556 7420 9620
rect 7484 9556 7485 9620
rect 7419 9555 7485 9556
rect 7235 9348 7301 9349
rect 7235 9284 7236 9348
rect 7300 9284 7301 9348
rect 7235 9283 7301 9284
rect 7235 9212 7301 9213
rect 7235 9148 7236 9212
rect 7300 9148 7301 9212
rect 7235 9147 7301 9148
rect 7051 4044 7117 4045
rect 7051 3980 7052 4044
rect 7116 3980 7117 4044
rect 7051 3979 7117 3980
rect 6566 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6886 3840
rect 6566 2752 6886 3776
rect 6566 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6886 2752
rect 6315 2684 6381 2685
rect 6315 2620 6316 2684
rect 6380 2620 6381 2684
rect 6315 2619 6381 2620
rect 6566 2128 6886 2688
rect 7054 917 7114 3979
rect 7238 3229 7298 9147
rect 7235 3228 7301 3229
rect 7235 3164 7236 3228
rect 7300 3164 7301 3228
rect 7235 3163 7301 3164
rect 7422 2821 7482 9555
rect 7790 6490 7850 11731
rect 7971 11252 8037 11253
rect 7971 11188 7972 11252
rect 8036 11188 8037 11252
rect 7971 11187 8037 11188
rect 7974 8261 8034 11187
rect 7971 8260 8037 8261
rect 7971 8196 7972 8260
rect 8036 8196 8037 8260
rect 7971 8195 8037 8196
rect 8158 8125 8218 12547
rect 8440 12000 8760 13024
rect 9262 12341 9322 13770
rect 9443 13564 9509 13565
rect 9443 13500 9444 13564
rect 9508 13500 9509 13564
rect 9443 13499 9509 13500
rect 9446 13021 9506 13499
rect 9443 13020 9509 13021
rect 9443 12956 9444 13020
rect 9508 12956 9509 13020
rect 9443 12955 9509 12956
rect 8891 12340 8957 12341
rect 8891 12276 8892 12340
rect 8956 12276 8957 12340
rect 8891 12275 8957 12276
rect 9075 12340 9141 12341
rect 9075 12276 9076 12340
rect 9140 12276 9141 12340
rect 9075 12275 9141 12276
rect 9259 12340 9325 12341
rect 9259 12276 9260 12340
rect 9324 12276 9325 12340
rect 9259 12275 9325 12276
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 8894 10165 8954 12275
rect 9078 10573 9138 12275
rect 9630 12069 9690 13771
rect 9627 12068 9693 12069
rect 9627 12004 9628 12068
rect 9692 12004 9693 12068
rect 9627 12003 9693 12004
rect 9259 11932 9325 11933
rect 9259 11868 9260 11932
rect 9324 11930 9325 11932
rect 9324 11870 9690 11930
rect 9324 11868 9325 11870
rect 9259 11867 9325 11868
rect 9259 11796 9325 11797
rect 9259 11732 9260 11796
rect 9324 11732 9325 11796
rect 9259 11731 9325 11732
rect 9075 10572 9141 10573
rect 9075 10508 9076 10572
rect 9140 10508 9141 10572
rect 9075 10507 9141 10508
rect 9262 10298 9322 11731
rect 9630 11525 9690 11870
rect 9814 11797 9874 15675
rect 10314 14720 10634 15744
rect 10314 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10634 14720
rect 10314 13632 10634 14656
rect 10314 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10634 13632
rect 10179 13564 10245 13565
rect 10179 13500 10180 13564
rect 10244 13500 10245 13564
rect 10179 13499 10245 13500
rect 9995 13292 10061 13293
rect 9995 13228 9996 13292
rect 10060 13228 10061 13292
rect 9995 13227 10061 13228
rect 9811 11796 9877 11797
rect 9811 11732 9812 11796
rect 9876 11732 9877 11796
rect 9811 11731 9877 11732
rect 9627 11524 9693 11525
rect 9627 11460 9628 11524
rect 9692 11460 9693 11524
rect 9627 11459 9693 11460
rect 9443 10844 9509 10845
rect 9443 10780 9444 10844
rect 9508 10780 9509 10844
rect 9443 10779 9509 10780
rect 9078 10238 9322 10298
rect 8891 10164 8957 10165
rect 8891 10100 8892 10164
rect 8956 10100 8957 10164
rect 8891 10099 8957 10100
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 8736 8760 9760
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8155 8124 8221 8125
rect 8155 8060 8156 8124
rect 8220 8060 8221 8124
rect 8155 8059 8221 8060
rect 8440 7648 8760 8672
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 6560 8760 7584
rect 8891 7580 8957 7581
rect 8891 7516 8892 7580
rect 8956 7516 8957 7580
rect 8891 7515 8957 7516
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 7790 6430 8218 6490
rect 7787 5948 7853 5949
rect 7787 5884 7788 5948
rect 7852 5884 7853 5948
rect 7787 5883 7853 5884
rect 7971 5948 8037 5949
rect 7971 5884 7972 5948
rect 8036 5884 8037 5948
rect 7971 5883 8037 5884
rect 7603 4316 7669 4317
rect 7603 4252 7604 4316
rect 7668 4252 7669 4316
rect 7603 4251 7669 4252
rect 7419 2820 7485 2821
rect 7419 2790 7420 2820
rect 7238 2756 7420 2790
rect 7484 2756 7485 2820
rect 7238 2755 7485 2756
rect 7238 2730 7482 2755
rect 7238 2549 7298 2730
rect 7235 2548 7301 2549
rect 7235 2484 7236 2548
rect 7300 2484 7301 2548
rect 7235 2483 7301 2484
rect 7606 1733 7666 4251
rect 7790 2005 7850 5883
rect 7974 2277 8034 5883
rect 8158 3773 8218 6430
rect 8440 5472 8760 6496
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8155 3772 8221 3773
rect 8155 3708 8156 3772
rect 8220 3708 8221 3772
rect 8155 3707 8221 3708
rect 8440 3296 8760 4320
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 7971 2276 8037 2277
rect 7971 2212 7972 2276
rect 8036 2212 8037 2276
rect 7971 2211 8037 2212
rect 8440 2208 8760 3232
rect 8894 2957 8954 7515
rect 8891 2956 8957 2957
rect 8891 2892 8892 2956
rect 8956 2892 8957 2956
rect 8891 2891 8957 2892
rect 9078 2685 9138 10238
rect 9259 8124 9325 8125
rect 9259 8060 9260 8124
rect 9324 8060 9325 8124
rect 9259 8059 9325 8060
rect 9262 3637 9322 8059
rect 9259 3636 9325 3637
rect 9259 3572 9260 3636
rect 9324 3572 9325 3636
rect 9259 3571 9325 3572
rect 9446 3362 9506 10779
rect 9814 8805 9874 11731
rect 9998 11389 10058 13227
rect 9995 11388 10061 11389
rect 9995 11324 9996 11388
rect 10060 11324 10061 11388
rect 9995 11323 10061 11324
rect 9995 11252 10061 11253
rect 9995 11188 9996 11252
rect 10060 11188 10061 11252
rect 9995 11187 10061 11188
rect 9998 10573 10058 11187
rect 9995 10572 10061 10573
rect 9995 10508 9996 10572
rect 10060 10508 10061 10572
rect 9995 10507 10061 10508
rect 10182 9893 10242 13499
rect 10314 12544 10634 13568
rect 10314 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10634 12544
rect 10314 11456 10634 12480
rect 10734 12477 10794 17987
rect 12571 17644 12637 17645
rect 12571 17580 12572 17644
rect 12636 17580 12637 17644
rect 12571 17579 12637 17580
rect 12188 17440 12508 17456
rect 12188 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12508 17440
rect 12188 16352 12508 17376
rect 12188 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12508 16352
rect 11467 15468 11533 15469
rect 11467 15404 11468 15468
rect 11532 15404 11533 15468
rect 11467 15403 11533 15404
rect 11099 13836 11165 13837
rect 11099 13772 11100 13836
rect 11164 13772 11165 13836
rect 11099 13771 11165 13772
rect 10731 12476 10797 12477
rect 10731 12412 10732 12476
rect 10796 12412 10797 12476
rect 10731 12411 10797 12412
rect 10314 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10634 11456
rect 10314 10368 10634 11392
rect 10314 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10634 10368
rect 10179 9892 10245 9893
rect 10179 9828 10180 9892
rect 10244 9828 10245 9892
rect 10179 9827 10245 9828
rect 9811 8804 9877 8805
rect 9811 8740 9812 8804
rect 9876 8740 9877 8804
rect 9811 8739 9877 8740
rect 9811 7716 9877 7717
rect 9811 7652 9812 7716
rect 9876 7652 9877 7716
rect 9811 7651 9877 7652
rect 9627 5676 9693 5677
rect 9627 5612 9628 5676
rect 9692 5612 9693 5676
rect 9627 5611 9693 5612
rect 9630 4997 9690 5611
rect 9627 4996 9693 4997
rect 9627 4932 9628 4996
rect 9692 4932 9693 4996
rect 9627 4931 9693 4932
rect 9627 4860 9693 4861
rect 9627 4796 9628 4860
rect 9692 4796 9693 4860
rect 9627 4795 9693 4796
rect 9262 3302 9506 3362
rect 9075 2684 9141 2685
rect 9075 2620 9076 2684
rect 9140 2620 9141 2684
rect 9075 2619 9141 2620
rect 9262 2549 9322 3302
rect 9630 2957 9690 4795
rect 9627 2956 9693 2957
rect 9627 2892 9628 2956
rect 9692 2892 9693 2956
rect 9627 2891 9693 2892
rect 9814 2549 9874 7651
rect 9995 6356 10061 6357
rect 9995 6292 9996 6356
rect 10060 6292 10061 6356
rect 9995 6291 10061 6292
rect 9998 3773 10058 6291
rect 10182 5677 10242 9827
rect 10314 9280 10634 10304
rect 10314 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10634 9280
rect 10314 8192 10634 9216
rect 10314 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10634 8192
rect 10314 7104 10634 8128
rect 10314 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10634 7104
rect 10314 6016 10634 7040
rect 10314 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10634 6016
rect 10179 5676 10245 5677
rect 10179 5612 10180 5676
rect 10244 5612 10245 5676
rect 10179 5611 10245 5612
rect 10179 5132 10245 5133
rect 10179 5068 10180 5132
rect 10244 5068 10245 5132
rect 10179 5067 10245 5068
rect 10182 4589 10242 5067
rect 10314 4928 10634 5952
rect 10734 5541 10794 12411
rect 10915 11116 10981 11117
rect 10915 11052 10916 11116
rect 10980 11052 10981 11116
rect 10915 11051 10981 11052
rect 10918 9621 10978 11051
rect 11102 9893 11162 13771
rect 11283 12884 11349 12885
rect 11283 12820 11284 12884
rect 11348 12820 11349 12884
rect 11283 12819 11349 12820
rect 11286 12069 11346 12819
rect 11283 12068 11349 12069
rect 11283 12004 11284 12068
rect 11348 12004 11349 12068
rect 11283 12003 11349 12004
rect 11099 9892 11165 9893
rect 11099 9828 11100 9892
rect 11164 9828 11165 9892
rect 11099 9827 11165 9828
rect 10915 9620 10981 9621
rect 10915 9556 10916 9620
rect 10980 9556 10981 9620
rect 10915 9555 10981 9556
rect 11286 8261 11346 12003
rect 11470 11253 11530 15403
rect 12188 15264 12508 16288
rect 12188 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12508 15264
rect 12188 14176 12508 15200
rect 12188 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12508 14176
rect 12188 13088 12508 14112
rect 12188 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12508 13088
rect 12019 13020 12085 13021
rect 12019 12956 12020 13020
rect 12084 12956 12085 13020
rect 12019 12955 12085 12956
rect 11651 12204 11717 12205
rect 11651 12140 11652 12204
rect 11716 12140 11717 12204
rect 11651 12139 11717 12140
rect 11467 11252 11533 11253
rect 11467 11188 11468 11252
rect 11532 11188 11533 11252
rect 11467 11187 11533 11188
rect 11654 10573 11714 12139
rect 11835 11388 11901 11389
rect 11835 11324 11836 11388
rect 11900 11324 11901 11388
rect 11835 11323 11901 11324
rect 11651 10572 11717 10573
rect 11651 10508 11652 10572
rect 11716 10508 11717 10572
rect 11651 10507 11717 10508
rect 11283 8260 11349 8261
rect 11283 8196 11284 8260
rect 11348 8196 11349 8260
rect 11283 8195 11349 8196
rect 10918 7382 11530 7442
rect 10918 6493 10978 7382
rect 11470 7309 11530 7382
rect 11467 7308 11533 7309
rect 11467 7244 11468 7308
rect 11532 7244 11533 7308
rect 11467 7243 11533 7244
rect 11102 6702 11530 6762
rect 11102 6493 11162 6702
rect 10915 6492 10981 6493
rect 10915 6428 10916 6492
rect 10980 6428 10981 6492
rect 10915 6427 10981 6428
rect 11099 6492 11165 6493
rect 11099 6428 11100 6492
rect 11164 6428 11165 6492
rect 11099 6427 11165 6428
rect 11283 6492 11349 6493
rect 11283 6428 11284 6492
rect 11348 6428 11349 6492
rect 11283 6427 11349 6428
rect 11286 6085 11346 6427
rect 10915 6084 10981 6085
rect 10915 6020 10916 6084
rect 10980 6020 10981 6084
rect 10915 6019 10981 6020
rect 11099 6084 11165 6085
rect 11099 6020 11100 6084
rect 11164 6020 11165 6084
rect 11099 6019 11165 6020
rect 11283 6084 11349 6085
rect 11283 6020 11284 6084
rect 11348 6020 11349 6084
rect 11283 6019 11349 6020
rect 10731 5540 10797 5541
rect 10731 5476 10732 5540
rect 10796 5476 10797 5540
rect 10731 5475 10797 5476
rect 10731 5268 10797 5269
rect 10731 5204 10732 5268
rect 10796 5204 10797 5268
rect 10731 5203 10797 5204
rect 10314 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10634 4928
rect 10179 4588 10245 4589
rect 10179 4524 10180 4588
rect 10244 4524 10245 4588
rect 10179 4523 10245 4524
rect 10314 3840 10634 4864
rect 10314 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10634 3840
rect 9995 3772 10061 3773
rect 9995 3708 9996 3772
rect 10060 3708 10061 3772
rect 9995 3707 10061 3708
rect 9995 3228 10061 3229
rect 9995 3164 9996 3228
rect 10060 3164 10061 3228
rect 9995 3163 10061 3164
rect 9998 2821 10058 3163
rect 9995 2820 10061 2821
rect 9995 2756 9996 2820
rect 10060 2756 10061 2820
rect 9995 2755 10061 2756
rect 10314 2752 10634 3776
rect 10734 2821 10794 5203
rect 10918 4181 10978 6019
rect 11102 5269 11162 6019
rect 11099 5268 11165 5269
rect 11099 5204 11100 5268
rect 11164 5204 11165 5268
rect 11099 5203 11165 5204
rect 11099 4996 11165 4997
rect 11099 4932 11100 4996
rect 11164 4994 11165 4996
rect 11470 4994 11530 6702
rect 11654 5405 11714 10507
rect 11838 8805 11898 11323
rect 12022 9349 12082 12955
rect 12188 12000 12508 13024
rect 12188 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12508 12000
rect 12188 10912 12508 11936
rect 12574 11117 12634 17579
rect 13307 17236 13373 17237
rect 13307 17172 13308 17236
rect 13372 17172 13373 17236
rect 13307 17171 13373 17172
rect 13123 17100 13189 17101
rect 13123 17036 13124 17100
rect 13188 17036 13189 17100
rect 13123 17035 13189 17036
rect 12939 12884 13005 12885
rect 12939 12820 12940 12884
rect 13004 12820 13005 12884
rect 12939 12819 13005 12820
rect 12755 11660 12821 11661
rect 12755 11596 12756 11660
rect 12820 11596 12821 11660
rect 12755 11595 12821 11596
rect 12571 11116 12637 11117
rect 12571 11052 12572 11116
rect 12636 11052 12637 11116
rect 12571 11051 12637 11052
rect 12188 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12508 10912
rect 12188 9824 12508 10848
rect 12758 10165 12818 11595
rect 12755 10164 12821 10165
rect 12755 10100 12756 10164
rect 12820 10100 12821 10164
rect 12755 10099 12821 10100
rect 12188 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12508 9824
rect 12019 9348 12085 9349
rect 12019 9284 12020 9348
rect 12084 9284 12085 9348
rect 12019 9283 12085 9284
rect 11835 8804 11901 8805
rect 11835 8740 11836 8804
rect 11900 8740 11901 8804
rect 11835 8739 11901 8740
rect 12188 8736 12508 9760
rect 12571 9212 12637 9213
rect 12571 9148 12572 9212
rect 12636 9148 12637 9212
rect 12571 9147 12637 9148
rect 12188 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12508 8736
rect 11835 8396 11901 8397
rect 11835 8332 11836 8396
rect 11900 8332 11901 8396
rect 11835 8331 11901 8332
rect 11651 5404 11717 5405
rect 11651 5340 11652 5404
rect 11716 5340 11717 5404
rect 11651 5339 11717 5340
rect 11164 4934 11530 4994
rect 11164 4932 11165 4934
rect 11099 4931 11165 4932
rect 11467 4588 11533 4589
rect 11467 4524 11468 4588
rect 11532 4524 11533 4588
rect 11467 4523 11533 4524
rect 11470 4181 11530 4523
rect 10915 4180 10981 4181
rect 10915 4116 10916 4180
rect 10980 4116 10981 4180
rect 10915 4115 10981 4116
rect 11467 4180 11533 4181
rect 11467 4116 11468 4180
rect 11532 4116 11533 4180
rect 11467 4115 11533 4116
rect 10731 2820 10797 2821
rect 10731 2756 10732 2820
rect 10796 2756 10797 2820
rect 10731 2755 10797 2756
rect 10314 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10634 2752
rect 9259 2548 9325 2549
rect 9259 2484 9260 2548
rect 9324 2484 9325 2548
rect 9259 2483 9325 2484
rect 9811 2548 9877 2549
rect 9811 2484 9812 2548
rect 9876 2484 9877 2548
rect 9811 2483 9877 2484
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 10314 2128 10634 2688
rect 10918 2141 10978 4115
rect 11654 3501 11714 5339
rect 11467 3500 11533 3501
rect 11467 3436 11468 3500
rect 11532 3436 11533 3500
rect 11467 3435 11533 3436
rect 11651 3500 11717 3501
rect 11651 3436 11652 3500
rect 11716 3436 11717 3500
rect 11651 3435 11717 3436
rect 11470 3229 11530 3435
rect 11467 3228 11533 3229
rect 11467 3164 11468 3228
rect 11532 3164 11533 3228
rect 11467 3163 11533 3164
rect 11467 2548 11533 2549
rect 11467 2484 11468 2548
rect 11532 2484 11533 2548
rect 11467 2483 11533 2484
rect 10915 2140 10981 2141
rect 10915 2076 10916 2140
rect 10980 2076 10981 2140
rect 10915 2075 10981 2076
rect 7787 2004 7853 2005
rect 7787 1940 7788 2004
rect 7852 1940 7853 2004
rect 7787 1939 7853 1940
rect 11470 1869 11530 2483
rect 11838 2005 11898 8331
rect 12019 8124 12085 8125
rect 12019 8060 12020 8124
rect 12084 8060 12085 8124
rect 12019 8059 12085 8060
rect 12022 6901 12082 8059
rect 12188 7648 12508 8672
rect 12574 8125 12634 9147
rect 12942 8669 13002 12819
rect 13126 10845 13186 17035
rect 13123 10844 13189 10845
rect 13123 10780 13124 10844
rect 13188 10780 13189 10844
rect 13123 10779 13189 10780
rect 13123 9756 13189 9757
rect 13123 9692 13124 9756
rect 13188 9692 13189 9756
rect 13123 9691 13189 9692
rect 12939 8668 13005 8669
rect 12939 8604 12940 8668
rect 13004 8604 13005 8668
rect 12939 8603 13005 8604
rect 13126 8397 13186 9691
rect 13310 9621 13370 17171
rect 14062 16896 14382 17456
rect 14062 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14382 16896
rect 14062 15808 14382 16832
rect 14062 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14382 15808
rect 13859 15060 13925 15061
rect 13859 14996 13860 15060
rect 13924 14996 13925 15060
rect 13859 14995 13925 14996
rect 13675 13564 13741 13565
rect 13675 13500 13676 13564
rect 13740 13500 13741 13564
rect 13675 13499 13741 13500
rect 13491 12476 13557 12477
rect 13491 12412 13492 12476
rect 13556 12412 13557 12476
rect 13491 12411 13557 12412
rect 13494 11389 13554 12411
rect 13491 11388 13557 11389
rect 13491 11324 13492 11388
rect 13556 11324 13557 11388
rect 13491 11323 13557 11324
rect 13678 11250 13738 13499
rect 13862 12341 13922 14995
rect 14062 14720 14382 15744
rect 14062 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14382 14720
rect 14062 13632 14382 14656
rect 14062 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14382 13632
rect 14062 12544 14382 13568
rect 14062 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14382 12544
rect 13859 12340 13925 12341
rect 13859 12276 13860 12340
rect 13924 12276 13925 12340
rect 13859 12275 13925 12276
rect 13859 11932 13925 11933
rect 13859 11868 13860 11932
rect 13924 11868 13925 11932
rect 13859 11867 13925 11868
rect 13494 11190 13738 11250
rect 13494 10573 13554 11190
rect 13862 10981 13922 11867
rect 14062 11456 14382 12480
rect 14062 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14382 11456
rect 13859 10980 13925 10981
rect 13859 10916 13860 10980
rect 13924 10916 13925 10980
rect 13859 10915 13925 10916
rect 13675 10708 13741 10709
rect 13675 10644 13676 10708
rect 13740 10644 13741 10708
rect 13675 10643 13741 10644
rect 13491 10572 13557 10573
rect 13491 10508 13492 10572
rect 13556 10508 13557 10572
rect 13491 10507 13557 10508
rect 13491 9892 13557 9893
rect 13491 9828 13492 9892
rect 13556 9828 13557 9892
rect 13491 9827 13557 9828
rect 13307 9620 13373 9621
rect 13307 9556 13308 9620
rect 13372 9556 13373 9620
rect 13307 9555 13373 9556
rect 13123 8396 13189 8397
rect 13123 8332 13124 8396
rect 13188 8332 13189 8396
rect 13123 8331 13189 8332
rect 12939 8260 13005 8261
rect 12939 8196 12940 8260
rect 13004 8196 13005 8260
rect 12939 8195 13005 8196
rect 12571 8124 12637 8125
rect 12571 8060 12572 8124
rect 12636 8060 12637 8124
rect 12571 8059 12637 8060
rect 12188 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12508 7648
rect 12019 6900 12085 6901
rect 12019 6836 12020 6900
rect 12084 6836 12085 6900
rect 12019 6835 12085 6836
rect 12022 3773 12082 6835
rect 12188 6560 12508 7584
rect 12571 7308 12637 7309
rect 12571 7244 12572 7308
rect 12636 7244 12637 7308
rect 12571 7243 12637 7244
rect 12188 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12508 6560
rect 12188 5472 12508 6496
rect 12188 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12508 5472
rect 12188 4384 12508 5408
rect 12188 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12508 4384
rect 12019 3772 12085 3773
rect 12019 3708 12020 3772
rect 12084 3708 12085 3772
rect 12019 3707 12085 3708
rect 12188 3296 12508 4320
rect 12574 4181 12634 7243
rect 12755 7036 12821 7037
rect 12755 6972 12756 7036
rect 12820 6972 12821 7036
rect 12755 6971 12821 6972
rect 12758 6629 12818 6971
rect 12755 6628 12821 6629
rect 12755 6564 12756 6628
rect 12820 6564 12821 6628
rect 12755 6563 12821 6564
rect 12755 6492 12821 6493
rect 12755 6428 12756 6492
rect 12820 6428 12821 6492
rect 12755 6427 12821 6428
rect 12758 5405 12818 6427
rect 12755 5404 12821 5405
rect 12755 5340 12756 5404
rect 12820 5340 12821 5404
rect 12755 5339 12821 5340
rect 12755 4452 12821 4453
rect 12755 4388 12756 4452
rect 12820 4388 12821 4452
rect 12755 4387 12821 4388
rect 12571 4180 12637 4181
rect 12571 4116 12572 4180
rect 12636 4116 12637 4180
rect 12571 4115 12637 4116
rect 12188 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12508 3296
rect 12188 2208 12508 3232
rect 12188 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12508 2208
rect 12188 2128 12508 2144
rect 11835 2004 11901 2005
rect 11835 1940 11836 2004
rect 11900 1940 11901 2004
rect 11835 1939 11901 1940
rect 11467 1868 11533 1869
rect 11467 1804 11468 1868
rect 11532 1804 11533 1868
rect 11467 1803 11533 1804
rect 7603 1732 7669 1733
rect 7603 1668 7604 1732
rect 7668 1668 7669 1732
rect 7603 1667 7669 1668
rect 7051 916 7117 917
rect 7051 852 7052 916
rect 7116 852 7117 916
rect 7051 851 7117 852
rect 6131 780 6197 781
rect 6131 716 6132 780
rect 6196 716 6197 780
rect 6131 715 6197 716
rect 12758 237 12818 4387
rect 12942 3093 13002 8195
rect 13307 7580 13373 7581
rect 13307 7516 13308 7580
rect 13372 7516 13373 7580
rect 13307 7515 13373 7516
rect 13123 7308 13189 7309
rect 13123 7244 13124 7308
rect 13188 7244 13189 7308
rect 13123 7243 13189 7244
rect 12939 3092 13005 3093
rect 12939 3028 12940 3092
rect 13004 3028 13005 3092
rect 12939 3027 13005 3028
rect 13126 2790 13186 7243
rect 13310 5813 13370 7515
rect 13494 7037 13554 9827
rect 13678 8397 13738 10643
rect 14062 10368 14382 11392
rect 14779 11388 14845 11389
rect 14779 11324 14780 11388
rect 14844 11324 14845 11388
rect 14779 11323 14845 11324
rect 14595 10844 14661 10845
rect 14595 10780 14596 10844
rect 14660 10780 14661 10844
rect 14595 10779 14661 10780
rect 14062 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14382 10368
rect 13859 10300 13925 10301
rect 13859 10236 13860 10300
rect 13924 10236 13925 10300
rect 13859 10235 13925 10236
rect 13862 9893 13922 10235
rect 13859 9892 13925 9893
rect 13859 9828 13860 9892
rect 13924 9828 13925 9892
rect 13859 9827 13925 9828
rect 13675 8396 13741 8397
rect 13675 8332 13676 8396
rect 13740 8332 13741 8396
rect 13675 8331 13741 8332
rect 13675 7580 13741 7581
rect 13675 7516 13676 7580
rect 13740 7516 13741 7580
rect 13675 7515 13741 7516
rect 13491 7036 13557 7037
rect 13491 6972 13492 7036
rect 13556 6972 13557 7036
rect 13491 6971 13557 6972
rect 13307 5812 13373 5813
rect 13307 5748 13308 5812
rect 13372 5748 13373 5812
rect 13307 5747 13373 5748
rect 13307 5540 13373 5541
rect 13307 5476 13308 5540
rect 13372 5476 13373 5540
rect 13307 5475 13373 5476
rect 13310 4858 13370 5475
rect 13494 4997 13554 6971
rect 13678 5541 13738 7515
rect 13862 6629 13922 9827
rect 14062 9280 14382 10304
rect 14062 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14382 9280
rect 14062 8192 14382 9216
rect 14062 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14382 8192
rect 14062 7104 14382 8128
rect 14062 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14382 7104
rect 13859 6628 13925 6629
rect 13859 6564 13860 6628
rect 13924 6564 13925 6628
rect 13859 6563 13925 6564
rect 13859 6492 13925 6493
rect 13859 6428 13860 6492
rect 13924 6428 13925 6492
rect 13859 6427 13925 6428
rect 13675 5540 13741 5541
rect 13675 5476 13676 5540
rect 13740 5476 13741 5540
rect 13675 5475 13741 5476
rect 13491 4996 13557 4997
rect 13491 4932 13492 4996
rect 13556 4932 13557 4996
rect 13491 4931 13557 4932
rect 13310 4798 13554 4858
rect 13307 4180 13373 4181
rect 13307 4116 13308 4180
rect 13372 4116 13373 4180
rect 13307 4115 13373 4116
rect 12942 2730 13186 2790
rect 12942 1597 13002 2730
rect 12939 1596 13005 1597
rect 12939 1532 12940 1596
rect 13004 1532 13005 1596
rect 12939 1531 13005 1532
rect 13310 645 13370 4115
rect 13494 3229 13554 4798
rect 13491 3228 13557 3229
rect 13491 3164 13492 3228
rect 13556 3164 13557 3228
rect 13491 3163 13557 3164
rect 13678 1461 13738 5475
rect 13862 2413 13922 6427
rect 14062 6016 14382 7040
rect 14062 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14382 6016
rect 14062 4928 14382 5952
rect 14062 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14382 4928
rect 14062 3840 14382 4864
rect 14062 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14382 3840
rect 14062 2752 14382 3776
rect 14598 2957 14658 10779
rect 14782 5949 14842 11323
rect 14963 8124 15029 8125
rect 14963 8060 14964 8124
rect 15028 8060 15029 8124
rect 14963 8059 15029 8060
rect 15331 8124 15397 8125
rect 15331 8060 15332 8124
rect 15396 8060 15397 8124
rect 15331 8059 15397 8060
rect 14966 6901 15026 8059
rect 14963 6900 15029 6901
rect 14963 6836 14964 6900
rect 15028 6836 15029 6900
rect 14963 6835 15029 6836
rect 14963 6764 15029 6765
rect 14963 6700 14964 6764
rect 15028 6700 15029 6764
rect 14963 6699 15029 6700
rect 14779 5948 14845 5949
rect 14779 5884 14780 5948
rect 14844 5884 14845 5948
rect 14779 5883 14845 5884
rect 14779 5540 14845 5541
rect 14779 5476 14780 5540
rect 14844 5476 14845 5540
rect 14779 5475 14845 5476
rect 14595 2956 14661 2957
rect 14595 2892 14596 2956
rect 14660 2892 14661 2956
rect 14595 2891 14661 2892
rect 14062 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14382 2752
rect 13859 2412 13925 2413
rect 13859 2348 13860 2412
rect 13924 2348 13925 2412
rect 13859 2347 13925 2348
rect 14062 2128 14382 2688
rect 13675 1460 13741 1461
rect 13675 1396 13676 1460
rect 13740 1396 13741 1460
rect 13675 1395 13741 1396
rect 14782 1325 14842 5475
rect 14966 4045 15026 6699
rect 15147 5132 15213 5133
rect 15147 5068 15148 5132
rect 15212 5068 15213 5132
rect 15147 5067 15213 5068
rect 14963 4044 15029 4045
rect 14963 3980 14964 4044
rect 15028 3980 15029 4044
rect 14963 3979 15029 3980
rect 15150 3093 15210 5067
rect 15334 4317 15394 8059
rect 15515 6628 15581 6629
rect 15515 6564 15516 6628
rect 15580 6564 15581 6628
rect 15515 6563 15581 6564
rect 15518 5269 15578 6563
rect 15515 5268 15581 5269
rect 15515 5204 15516 5268
rect 15580 5204 15581 5268
rect 15515 5203 15581 5204
rect 15331 4316 15397 4317
rect 15331 4252 15332 4316
rect 15396 4252 15397 4316
rect 15331 4251 15397 4252
rect 15147 3092 15213 3093
rect 15147 3028 15148 3092
rect 15212 3028 15213 3092
rect 15147 3027 15213 3028
rect 14779 1324 14845 1325
rect 14779 1260 14780 1324
rect 14844 1260 14845 1324
rect 14779 1259 14845 1260
rect 13307 644 13373 645
rect 13307 580 13308 644
rect 13372 580 13373 644
rect 13307 579 13373 580
rect 12755 236 12821 237
rect 12755 172 12756 236
rect 12820 172 12821 236
rect 12755 171 12821 172
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_E_FTB01_A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14628 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_N_FTB01_A
timestamp 1649977179
transform 1 0 5244 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_W_FTB01_A
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1649977179
transform 1 0 15364 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__33__A
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A
timestamp 1649977179
transform -1 0 15180 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1649977179
transform 1 0 15180 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1649977179
transform 1 0 1564 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1649977179
transform -1 0 3680 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform -1 0 1564 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1649977179
transform 1 0 3404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform 1 0 1656 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform 1 0 14628 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform 1 0 1840 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform 1 0 3312 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1649977179
transform -1 0 15732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform 1 0 3956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform 1 0 4508 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform -1 0 3864 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1649977179
transform 1 0 4324 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1649977179
transform -1 0 4876 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1649977179
transform -1 0 5336 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1649977179
transform -1 0 4784 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1649977179
transform 1 0 5704 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1649977179
transform -1 0 5704 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1649977179
transform 1 0 10948 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1649977179
transform -1 0 6440 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1649977179
transform -1 0 9292 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1649977179
transform 1 0 6440 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1649977179
transform -1 0 7912 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform 1 0 8740 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform -1 0 8556 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1649977179
transform -1 0 10304 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform -1 0 10488 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform 1 0 9844 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform -1 0 10120 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_N_FTB01_A
timestamp 1649977179
transform -1 0 7084 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_2_S_FTB01_A
timestamp 1649977179
transform -1 0 14628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_N_FTB01_A
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clk_3_S_FTB01_A
timestamp 1649977179
transform -1 0 14996 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_0_W_in_A
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 2760 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2__D
timestamp 1649977179
transform 1 0 11132 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10856 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 1840 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12420 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 15456 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8372 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 14260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__S
timestamp 1649977179
transform 1 0 12604 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12052 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__S
timestamp 1649977179
transform -1 0 1656 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 9476 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__S
timestamp 1649977179
transform -1 0 9476 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 12788 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 5244 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 15364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 15088 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 2944 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 2760 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 11868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 5612 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 5336 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14720 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 15272 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15456 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 15088 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 15364 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 14720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 14352 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 15272 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14628 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 15640 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14076 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 9016 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 12052 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 8096 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14168 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 15456 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 15732 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 15732 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 1840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 15548 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 15732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 15548 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 15088 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 15732 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5060 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3128 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 10672 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 15180 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 15364 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14812 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4968 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4784 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 3312 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3128 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 15640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 15456 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 6624 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7360 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 7360 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 2208 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 10028 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__S
timestamp 1649977179
transform -1 0 7728 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 15180 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 15364 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__S
timestamp 1649977179
transform -1 0 14444 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11684 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__S
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l3_in_0__A1
timestamp 1649977179
transform -1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14996 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 9752 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 15732 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 14812 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 1656 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10580 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 2944 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 14996 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14628 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 1564 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 2392 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 2576 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10120 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10488 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 14168 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 12420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12788 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12052 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 2576 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 2760 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9476 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 13984 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14444 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11316 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4416 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4692 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 8188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13708 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3128 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12972 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 11684 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12604 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 11500 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13892 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14076 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 10764 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 12420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13708 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_N_FTB01_A
timestamp 1649977179
transform 1 0 15364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_2_S_FTB01_A
timestamp 1649977179
transform -1 0 15732 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_N_FTB01_A
timestamp 1649977179
transform -1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_3_S_FTB01_A
timestamp 1649977179
transform -1 0 15364 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_81
timestamp 1649977179
transform 1 0 8556 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_81
timestamp 1649977179
transform 1 0 8556 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_158
timestamp 1649977179
transform 1 0 15640 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_158
timestamp 1649977179
transform 1 0 15640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_23
timestamp 1649977179
transform 1 0 3220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_158
timestamp 1649977179
transform 1 0 15640 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_35
timestamp 1649977179
transform 1 0 4324 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_158
timestamp 1649977179
transform 1 0 15640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_23
timestamp 1649977179
transform 1 0 3220 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_158
timestamp 1649977179
transform 1 0 15640 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_35
timestamp 1649977179
transform 1 0 4324 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_158
timestamp 1649977179
transform 1 0 15640 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_129 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_147 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_151
timestamp 1649977179
transform 1 0 14996 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_155
timestamp 1649977179
transform 1 0 15364 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_119 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12052 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_131
timestamp 1649977179
transform 1 0 13156 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_143
timestamp 1649977179
transform 1 0 14260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_155
timestamp 1649977179
transform 1 0 15364 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_18
timestamp 1649977179
transform 1 0 2760 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_38
timestamp 1649977179
transform 1 0 4600 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp 1649977179
transform 1 0 9292 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_108
timestamp 1649977179
transform 1 0 11040 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_120
timestamp 1649977179
transform 1 0 12144 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_132 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13248 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_153 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_24
timestamp 1649977179
transform 1 0 3312 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_82
timestamp 1649977179
transform 1 0 8648 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_99
timestamp 1649977179
transform 1 0 10212 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1649977179
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_33
timestamp 1649977179
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_95
timestamp 1649977179
transform 1 0 9844 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_107
timestamp 1649977179
transform 1 0 10948 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_119
timestamp 1649977179
transform 1 0 12052 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_131
timestamp 1649977179
transform 1 0 13156 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_30
timestamp 1649977179
transform 1 0 3864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_76
timestamp 1649977179
transform 1 0 8096 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_85
timestamp 1649977179
transform 1 0 8924 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_97
timestamp 1649977179
transform 1 0 10028 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_109
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_157
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_23
timestamp 1649977179
transform 1 0 3220 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_45
timestamp 1649977179
transform 1 0 5244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_49
timestamp 1649977179
transform 1 0 5612 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_55
timestamp 1649977179
transform 1 0 6164 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_60
timestamp 1649977179
transform 1 0 6624 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_76
timestamp 1649977179
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_30
timestamp 1649977179
transform 1 0 3864 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_38
timestamp 1649977179
transform 1 0 4600 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_47
timestamp 1649977179
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_157
timestamp 1649977179
transform 1 0 15548 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_29
timestamp 1649977179
transform 1 0 3772 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_41
timestamp 1649977179
transform 1 0 4876 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 1649977179
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_85
timestamp 1649977179
transform 1 0 8924 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_97
timestamp 1649977179
transform 1 0 10028 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_141
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_153
timestamp 1649977179
transform 1 0 15180 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 16008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 16008 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 16008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 16008 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 16008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 16008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__buf_4  Test_en_E_FTB01 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13156 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  Test_en_N_FTB01
timestamp 1649977179
transform -1 0 5244 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  Test_en_W_FTB01
timestamp 1649977179
transform -1 0 4324 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _16_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13708 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _17_
timestamp 1649977179
transform -1 0 13984 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1649977179
transform 1 0 13524 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1649977179
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1649977179
transform -1 0 1840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1649977179
transform 1 0 14720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1649977179
transform 1 0 14444 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1649977179
transform -1 0 7360 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1649977179
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1649977179
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1649977179
transform -1 0 5152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1649977179
transform -1 0 8740 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1649977179
transform -1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1649977179
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _32_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15364 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _33_
timestamp 1649977179
transform -1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _34_
timestamp 1649977179
transform -1 0 14720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1649977179
transform -1 0 14996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1649977179
transform -1 0 1840 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1649977179
transform -1 0 14628 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1649977179
transform -1 0 4600 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1649977179
transform 1 0 1472 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1649977179
transform -1 0 3680 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1649977179
transform -1 0 1840 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1649977179
transform -1 0 14352 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1649977179
transform -1 0 1840 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1649977179
transform -1 0 3680 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1649977179
transform -1 0 14444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1649977179
transform -1 0 11316 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1649977179
transform -1 0 11408 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1649977179
transform -1 0 13800 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1649977179
transform -1 0 3680 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1649977179
transform -1 0 13432 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1649977179
transform -1 0 3864 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1649977179
transform -1 0 3680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1649977179
transform -1 0 4324 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1649977179
transform -1 0 4692 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1649977179
transform -1 0 5152 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1649977179
transform -1 0 4600 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1649977179
transform -1 0 5520 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1649977179
transform -1 0 5520 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1649977179
transform -1 0 8832 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1649977179
transform -1 0 6256 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1649977179
transform -1 0 8740 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1649977179
transform -1 0 6808 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1649977179
transform -1 0 7728 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1649977179
transform -1 0 8096 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1649977179
transform -1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1649977179
transform -1 0 9292 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1649977179
transform -1 0 8832 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1649977179
transform -1 0 9476 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1649977179
transform -1 0 9108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1649977179
transform -1 0 9752 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  clk_2_N_FTB01
timestamp 1649977179
transform -1 0 6900 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_2_S_FTB01
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_N_FTB01
timestamp 1649977179
transform -1 0 11316 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  clk_3_S_FTB01
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_right_ipin_0.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk_0_W_in
timestamp 1649977179
transform 1 0 6624 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk_0_W_in
timestamp 1649977179
transform -1 0 4416 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk_0_W_in
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_mem_right_ipin_0.prog_clk
timestamp 1649977179
transform -1 0 3220 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_mem_right_ipin_0.prog_clk
timestamp 1649977179
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_mem_right_ipin_0.prog_clk
timestamp 1649977179
transform -1 0 3220 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_mem_right_ipin_0.prog_clk
timestamp 1649977179
transform -1 0 6348 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_mem_right_ipin_0.prog_clk
timestamp 1649977179
transform 1 0 5244 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_mem_right_ipin_0.prog_clk
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_mem_right_ipin_0.prog_clk
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_mem_right_ipin_0.prog_clk
timestamp 1649977179
transform 1 0 7820 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2760 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10396 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2208 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9292 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6900 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7820 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7820 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 3312 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 2208 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4784 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 1840 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8832 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3680 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 1840 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 1840 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10396 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5428 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7820 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 3312 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8556 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 6256 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 3312 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 4784 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 1840 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7360 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10396 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 3312 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9292 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7820 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 3312 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6992 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6256 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5888 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 2208 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5888 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 6256 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 5244 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 6256 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 3312 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 6992 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 3312 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7360 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 6164 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4784 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 9292 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8832 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 4784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4784 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7636 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10672 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13064 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 10120 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13984 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 8556 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform -1 0 7728 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 9844 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 13156 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13156 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10212 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform -1 0 11408 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 13064 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13156 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform -1 0 13156 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 2760 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11408 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5428 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 13984 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform -1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14904 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 12236 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 13156 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12880 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9292 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8004 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform -1 0 11224 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11868 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 11408 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13156 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13984 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13156 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7176 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform -1 0 13524 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13064 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9752 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10580 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11224 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12052 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 11040 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 10580 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12328 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13984 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8832 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform -1 0 10580 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1932 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4784 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform -1 0 3680 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6256 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2852 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4324 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12880 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2208 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8004 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 9476 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5428 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2484 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9292 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13984 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 4692 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2852 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2208 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12328 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3312 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5520 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10304 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3772 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1649977179
transform -1 0 2484 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1649977179
transform -1 0 8188 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7636 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3128 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6348 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2576 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1649977179
transform -1 0 2208 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1649977179
transform -1 0 8464 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6532 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1649977179
transform 1 0 10396 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7820 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2852 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7176 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1649977179
transform 1 0 10396 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1649977179
transform 1 0 6808 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3956 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2208 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 2208 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1649977179
transform 1 0 11408 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10488 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2576 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12052 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12880 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1649977179
transform -1 0 9476 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11224 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12052 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1649977179
transform -1 0 4784 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7360 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3128 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1649977179
transform -1 0 2484 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1649977179
transform -1 0 14628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1649977179
transform 1 0 15180 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_N_FTB01
timestamp 1649977179
transform -1 0 8832 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_3_S_FTB01
timestamp 1649977179
transform 1 0 14628 0 -1 3264
box -38 -48 590 592
<< labels >>
rlabel metal3 s 16400 16600 17200 16720 6 Test_en_E_in
port 0 nsew signal input
rlabel metal3 s 16400 9936 17200 10056 6 Test_en_E_out
port 1 nsew signal tristate
rlabel metal2 s 2042 19200 2098 20000 6 Test_en_N_out
port 2 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 Test_en_S_in
port 3 nsew signal input
rlabel metal3 s 0 17280 800 17400 6 Test_en_W_in
port 4 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 Test_en_W_out
port 5 nsew signal tristate
rlabel metal4 s 4692 2128 5012 17456 6 VGND
port 6 nsew ground input
rlabel metal4 s 8440 2128 8760 17456 6 VGND
port 6 nsew ground input
rlabel metal4 s 12188 2128 12508 17456 6 VGND
port 6 nsew ground input
rlabel metal4 s 2818 2128 3138 17456 6 VPWR
port 7 nsew power input
rlabel metal4 s 6566 2128 6886 17456 6 VPWR
port 7 nsew power input
rlabel metal4 s 10314 2128 10634 17456 6 VPWR
port 7 nsew power input
rlabel metal4 s 14062 2128 14382 17456 6 VPWR
port 7 nsew power input
rlabel metal3 s 0 416 800 536 6 ccff_head
port 8 nsew signal input
rlabel metal3 s 16400 3272 17200 3392 6 ccff_tail
port 9 nsew signal tristate
rlabel metal2 s 6918 0 6974 800 6 chany_bottom_in[0]
port 10 nsew signal input
rlabel metal2 s 10414 0 10470 800 6 chany_bottom_in[10]
port 11 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 chany_bottom_in[11]
port 12 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[12]
port 13 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[13]
port 14 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[14]
port 15 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 chany_bottom_in[15]
port 16 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 chany_bottom_in[16]
port 17 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 chany_bottom_in[17]
port 18 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 chany_bottom_in[18]
port 19 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 chany_bottom_in[19]
port 20 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[1]
port 21 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[2]
port 22 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 chany_bottom_in[3]
port 23 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_in[4]
port 24 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 chany_bottom_in[5]
port 25 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 chany_bottom_in[6]
port 26 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 chany_bottom_in[7]
port 27 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 chany_bottom_in[8]
port 28 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[9]
port 29 nsew signal input
rlabel metal2 s 110 0 166 800 6 chany_bottom_out[0]
port 30 nsew signal tristate
rlabel metal2 s 3514 0 3570 800 6 chany_bottom_out[10]
port 31 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 chany_bottom_out[11]
port 32 nsew signal tristate
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_out[12]
port 33 nsew signal tristate
rlabel metal2 s 4526 0 4582 800 6 chany_bottom_out[13]
port 34 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 chany_bottom_out[14]
port 35 nsew signal tristate
rlabel metal2 s 5262 0 5318 800 6 chany_bottom_out[15]
port 36 nsew signal tristate
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_out[16]
port 37 nsew signal tristate
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_out[17]
port 38 nsew signal tristate
rlabel metal2 s 6274 0 6330 800 6 chany_bottom_out[18]
port 39 nsew signal tristate
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_out[19]
port 40 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 chany_bottom_out[1]
port 41 nsew signal tristate
rlabel metal2 s 754 0 810 800 6 chany_bottom_out[2]
port 42 nsew signal tristate
rlabel metal2 s 1122 0 1178 800 6 chany_bottom_out[3]
port 43 nsew signal tristate
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_out[4]
port 44 nsew signal tristate
rlabel metal2 s 1766 0 1822 800 6 chany_bottom_out[5]
port 45 nsew signal tristate
rlabel metal2 s 2134 0 2190 800 6 chany_bottom_out[6]
port 46 nsew signal tristate
rlabel metal2 s 2502 0 2558 800 6 chany_bottom_out[7]
port 47 nsew signal tristate
rlabel metal2 s 2778 0 2834 800 6 chany_bottom_out[8]
port 48 nsew signal tristate
rlabel metal2 s 3146 0 3202 800 6 chany_bottom_out[9]
port 49 nsew signal tristate
rlabel metal2 s 9862 19200 9918 20000 6 chany_top_in[0]
port 50 nsew signal input
rlabel metal2 s 13634 19200 13690 20000 6 chany_top_in[10]
port 51 nsew signal input
rlabel metal2 s 14002 19200 14058 20000 6 chany_top_in[11]
port 52 nsew signal input
rlabel metal2 s 14370 19200 14426 20000 6 chany_top_in[12]
port 53 nsew signal input
rlabel metal2 s 14738 19200 14794 20000 6 chany_top_in[13]
port 54 nsew signal input
rlabel metal2 s 15106 19200 15162 20000 6 chany_top_in[14]
port 55 nsew signal input
rlabel metal2 s 15474 19200 15530 20000 6 chany_top_in[15]
port 56 nsew signal input
rlabel metal2 s 15842 19200 15898 20000 6 chany_top_in[16]
port 57 nsew signal input
rlabel metal2 s 16210 19200 16266 20000 6 chany_top_in[17]
port 58 nsew signal input
rlabel metal2 s 16578 19200 16634 20000 6 chany_top_in[18]
port 59 nsew signal input
rlabel metal2 s 16946 19200 17002 20000 6 chany_top_in[19]
port 60 nsew signal input
rlabel metal2 s 10230 19200 10286 20000 6 chany_top_in[1]
port 61 nsew signal input
rlabel metal2 s 10598 19200 10654 20000 6 chany_top_in[2]
port 62 nsew signal input
rlabel metal2 s 10966 19200 11022 20000 6 chany_top_in[3]
port 63 nsew signal input
rlabel metal2 s 11334 19200 11390 20000 6 chany_top_in[4]
port 64 nsew signal input
rlabel metal2 s 11794 19200 11850 20000 6 chany_top_in[5]
port 65 nsew signal input
rlabel metal2 s 12162 19200 12218 20000 6 chany_top_in[6]
port 66 nsew signal input
rlabel metal2 s 12530 19200 12586 20000 6 chany_top_in[7]
port 67 nsew signal input
rlabel metal2 s 12898 19200 12954 20000 6 chany_top_in[8]
port 68 nsew signal input
rlabel metal2 s 13266 19200 13322 20000 6 chany_top_in[9]
port 69 nsew signal input
rlabel metal2 s 2410 19200 2466 20000 6 chany_top_out[0]
port 70 nsew signal tristate
rlabel metal2 s 6182 19200 6238 20000 6 chany_top_out[10]
port 71 nsew signal tristate
rlabel metal2 s 6550 19200 6606 20000 6 chany_top_out[11]
port 72 nsew signal tristate
rlabel metal2 s 6918 19200 6974 20000 6 chany_top_out[12]
port 73 nsew signal tristate
rlabel metal2 s 7286 19200 7342 20000 6 chany_top_out[13]
port 74 nsew signal tristate
rlabel metal2 s 7654 19200 7710 20000 6 chany_top_out[14]
port 75 nsew signal tristate
rlabel metal2 s 8022 19200 8078 20000 6 chany_top_out[15]
port 76 nsew signal tristate
rlabel metal2 s 8390 19200 8446 20000 6 chany_top_out[16]
port 77 nsew signal tristate
rlabel metal2 s 8758 19200 8814 20000 6 chany_top_out[17]
port 78 nsew signal tristate
rlabel metal2 s 9126 19200 9182 20000 6 chany_top_out[18]
port 79 nsew signal tristate
rlabel metal2 s 9494 19200 9550 20000 6 chany_top_out[19]
port 80 nsew signal tristate
rlabel metal2 s 2778 19200 2834 20000 6 chany_top_out[1]
port 81 nsew signal tristate
rlabel metal2 s 3146 19200 3202 20000 6 chany_top_out[2]
port 82 nsew signal tristate
rlabel metal2 s 3514 19200 3570 20000 6 chany_top_out[3]
port 83 nsew signal tristate
rlabel metal2 s 3882 19200 3938 20000 6 chany_top_out[4]
port 84 nsew signal tristate
rlabel metal2 s 4250 19200 4306 20000 6 chany_top_out[5]
port 85 nsew signal tristate
rlabel metal2 s 4618 19200 4674 20000 6 chany_top_out[6]
port 86 nsew signal tristate
rlabel metal2 s 4986 19200 5042 20000 6 chany_top_out[7]
port 87 nsew signal tristate
rlabel metal2 s 5354 19200 5410 20000 6 chany_top_out[8]
port 88 nsew signal tristate
rlabel metal2 s 5722 19200 5778 20000 6 chany_top_out[9]
port 89 nsew signal tristate
rlabel metal2 s 202 19200 258 20000 6 clk_2_N_out
port 90 nsew signal tristate
rlabel metal2 s 14186 0 14242 800 6 clk_2_S_in
port 91 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 clk_2_S_out
port 92 nsew signal tristate
rlabel metal2 s 570 19200 626 20000 6 clk_3_N_out
port 93 nsew signal tristate
rlabel metal2 s 14554 0 14610 800 6 clk_3_S_in
port 94 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 clk_3_S_out
port 95 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 left_grid_pin_16_
port 96 nsew signal tristate
rlabel metal3 s 0 2320 800 2440 6 left_grid_pin_17_
port 97 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 left_grid_pin_18_
port 98 nsew signal tristate
rlabel metal3 s 0 4360 800 4480 6 left_grid_pin_19_
port 99 nsew signal tristate
rlabel metal3 s 0 5312 800 5432 6 left_grid_pin_20_
port 100 nsew signal tristate
rlabel metal3 s 0 6400 800 6520 6 left_grid_pin_21_
port 101 nsew signal tristate
rlabel metal3 s 0 7352 800 7472 6 left_grid_pin_22_
port 102 nsew signal tristate
rlabel metal3 s 0 8304 800 8424 6 left_grid_pin_23_
port 103 nsew signal tristate
rlabel metal3 s 0 9392 800 9512 6 left_grid_pin_24_
port 104 nsew signal tristate
rlabel metal3 s 0 10344 800 10464 6 left_grid_pin_25_
port 105 nsew signal tristate
rlabel metal3 s 0 11296 800 11416 6 left_grid_pin_26_
port 106 nsew signal tristate
rlabel metal3 s 0 12384 800 12504 6 left_grid_pin_27_
port 107 nsew signal tristate
rlabel metal3 s 0 13336 800 13456 6 left_grid_pin_28_
port 108 nsew signal tristate
rlabel metal3 s 0 14288 800 14408 6 left_grid_pin_29_
port 109 nsew signal tristate
rlabel metal3 s 0 15376 800 15496 6 left_grid_pin_30_
port 110 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 left_grid_pin_31_
port 111 nsew signal tristate
rlabel metal2 s 938 19200 994 20000 6 prog_clk_0_N_out
port 112 nsew signal tristate
rlabel metal2 s 16210 0 16266 800 6 prog_clk_0_S_out
port 113 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 prog_clk_0_W_in
port 114 nsew signal input
rlabel metal2 s 1306 19200 1362 20000 6 prog_clk_2_N_out
port 115 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 prog_clk_2_S_in
port 116 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 prog_clk_2_S_out
port 117 nsew signal tristate
rlabel metal2 s 1674 19200 1730 20000 6 prog_clk_3_N_out
port 118 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 prog_clk_3_S_in
port 119 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 prog_clk_3_S_out
port 120 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
