* NGSPICE file created from sb_2__0_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

.subckt sb_2__0_ VGND VPWR ccff_head ccff_tail chanx_left_in[0] chanx_left_in[10]
+ chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14] chanx_left_in[15]
+ chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19] chanx_left_in[1]
+ chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5] chanx_left_in[6]
+ chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0] chanx_left_out[10]
+ chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14] chanx_left_out[15]
+ chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19] chanx_left_out[1]
+ chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5] chanx_left_out[6]
+ chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_top_in[0] chany_top_in[10]
+ chany_top_in[11] chany_top_in[12] chany_top_in[13] chany_top_in[14] chany_top_in[15]
+ chany_top_in[16] chany_top_in[17] chany_top_in[18] chany_top_in[19] chany_top_in[1]
+ chany_top_in[2] chany_top_in[3] chany_top_in[4] chany_top_in[5] chany_top_in[6]
+ chany_top_in[7] chany_top_in[8] chany_top_in[9] chany_top_out[0] chany_top_out[10]
+ chany_top_out[11] chany_top_out[12] chany_top_out[13] chany_top_out[14] chany_top_out[15]
+ chany_top_out[16] chany_top_out[17] chany_top_out[18] chany_top_out[19] chany_top_out[1]
+ chany_top_out[2] chany_top_out[3] chany_top_out[4] chany_top_out[5] chany_top_out[6]
+ chany_top_out[7] chany_top_out[8] chany_top_out[9] left_bottom_grid_pin_11_ left_bottom_grid_pin_13_
+ left_bottom_grid_pin_15_ left_bottom_grid_pin_17_ left_bottom_grid_pin_1_ left_bottom_grid_pin_3_
+ left_bottom_grid_pin_5_ left_bottom_grid_pin_7_ left_bottom_grid_pin_9_ prog_clk_0_N_in
+ top_left_grid_pin_42_ top_left_grid_pin_43_ top_left_grid_pin_44_ top_left_grid_pin_45_
+ top_left_grid_pin_46_ top_left_grid_pin_47_ top_left_grid_pin_48_ top_left_grid_pin_49_
+ top_right_grid_pin_1_
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7__f_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_3_7__f_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3__f_mem_left_track_1.prog_clk/X
+ hold35/X VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A0 input53/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input55_A top_left_grid_pin_46_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_27.mux_l2_in_0__133 VGND VGND VPWR VPWR mux_left_track_27.mux_l2_in_0_/A0
+ mux_left_track_27.mux_l2_in_0__133/LO sky130_fd_sc_hd__conb_1
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input18_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput64 _080_/X VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
Xoutput75 _072_/X VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
Xoutput97 _094_/X VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
Xoutput86 _102_/X VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
XFILLER_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_104 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_31.mux_l2_in_0__102 VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/A0
+ mux_left_track_31.mux_l2_in_0__102/LO sky130_fd_sc_hd__conb_1
XFILLER_24_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input48_A left_bottom_grid_pin_5_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _072_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_31.sky130_fd_sc_hd__buf_4_0_ mux_left_track_31.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _083_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_top_track_10.mux_l2_in_0_ mux_top_track_10.mux_l2_in_0_/A0 mux_top_track_10.mux_l1_in_0_/X
+ hold9/A VGND VGND VPWR VPWR mux_top_track_10.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold36/X VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput98 _095_/X VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
Xoutput65 _081_/X VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
Xoutput76 _073_/X VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
Xoutput87 _103_/X VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
XANTENNA_input30_A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _080_/A sky130_fd_sc_hd__clkbuf_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_19.sky130_fd_sc_hd__buf_4_0_ mux_left_track_19.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_7.mux_l3_in_0_ mux_left_track_7.mux_l2_in_1_/X mux_left_track_7.mux_l2_in_0_/X
+ hold60/A VGND VGND VPWR VPWR mux_left_track_7.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_5.mux_l2_in_1__107 VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/A0
+ mux_left_track_5.mux_l2_in_1__107/LO sky130_fd_sc_hd__conb_1
Xclkbuf_0_mem_left_track_1.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_left_track_1.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1__f_mem_left_track_1.prog_clk/X
+ hold44/X VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_7.mux_l2_in_1_ mux_left_track_7.mux_l2_in_1_/A0 input44/X hold15/A
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_14.mux_l2_in_0__113 VGND VGND VPWR VPWR mux_top_track_14.mux_l2_in_0_/A0
+ mux_top_track_14.mux_l2_in_0__113/LO sky130_fd_sc_hd__conb_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold30/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput99 _096_/X VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput77 _074_/X VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
Xoutput66 _082_/X VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
Xoutput88 _104_/X VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
XANTENNA_input23_A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_10.mux_l1_in_0_ input8/X input52/X hold44/A VGND VGND VPWR VPWR mux_top_track_10.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_2.mux_l1_in_1__A0 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_22.mux_l2_in_0_ mux_top_track_22.mux_l2_in_0_/A0 mux_top_track_22.mux_l1_in_0_/X
+ hold13/A VGND VGND VPWR VPWR mux_top_track_22.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_15.mux_l2_in_0_ mux_left_track_15.mux_l2_in_0_/A0 mux_left_track_15.mux_l1_in_0_/X
+ hold35/A VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l2_in_1__101 VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/A0
+ mux_left_track_3.mux_l2_in_1__101/LO sky130_fd_sc_hd__conb_1
XFILLER_15_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1__f_mem_left_track_1.prog_clk/X
+ hold7/X VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xprog_clk_0_FTB00 prog_clk_0_N_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_7.mux_l2_in_0_ mux_left_track_7.mux_l1_in_1_/X mux_left_track_7.mux_l1_in_0_/X
+ hold15/A VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input53_A top_left_grid_pin_44_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ hold59/A VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_59 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6__f_mem_left_track_1.prog_clk/X
+ hold12/X VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_7.mux_l1_in_1_ input42/X input49/X mux_left_track_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput78 _075_/X VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
Xoutput67 _083_/X VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
Xoutput89 _105_/X VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
XANTENNA_input16_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ mux_top_track_0.mux_l2_in_1_/A0 mux_top_track_0.mux_l1_in_2_/X
+ hold61/A VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_80 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input8_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_1__A1 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_22.sky130_fd_sc_hd__buf_4_0_ mux_top_track_22.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _099_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_1__132 VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/A0
+ mux_left_track_25.mux_l1_in_1__132/LO sky130_fd_sc_hd__conb_1
XFILLER_18_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_0.mux_l1_in_2_ input2/X input59/X mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_14.mux_l1_in_0__A0 input6/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_22.mux_l1_in_0_ input21/X input58/X hold41/A VGND VGND VPWR VPWR mux_top_track_22.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _096_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_23_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_15.mux_l1_in_0_ input49/X input26/X hold23/A VGND VGND VPWR VPWR mux_left_track_15.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input46_A left_bottom_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_27.mux_l2_in_0_ mux_left_track_27.mux_l2_in_0_/A0 mux_left_track_27.mux_l1_in_0_/X
+ hold45/A VGND VGND VPWR VPWR mux_left_track_27.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4__f_mem_left_track_1.prog_clk/X
+ hold6/X VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_13.mux_l2_in_0__126 VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_0_/A0
+ mux_left_track_13.mux_l2_in_0__126/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_7.mux_l1_in_0_ input47/X input30/X mux_left_track_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _088_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_31_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput79 _076_/X VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
Xoutput68 _084_/X VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ hold61/A VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_92 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_22.mux_l1_in_0__A0 input21/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l1_in_1_ input57/X input55/X mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_left_track_1.prog_clk/X
+ hold25/X VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_14.mux_l1_in_0__A1 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_26.mux_l2_in_0__120 VGND VGND VPWR VPWR mux_top_track_26.mux_l2_in_0_/A0
+ mux_top_track_26.mux_l2_in_0__120/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_6.mux_l1_in_0__A0 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input39_A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_3__f_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_3_3__f_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_27.mux_l1_in_0_ input47/X input39/X hold48/A VGND VGND VPWR VPWR mux_left_track_27.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput69 _085_/X VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
XFILLER_16_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_39.mux_l2_in_0_ mux_left_track_39.mux_l2_in_0_/A0 mux_left_track_39.mux_l1_in_0_/X
+ output60/A VGND VGND VPWR VPWR mux_left_track_39.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input21_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_22.mux_l1_in_0__A1 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_15.mux_l1_in_0__A0 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l1_in_0_ input53/X input51/X mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold1/X VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l1_in_0__A1 input52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_099_ _099_/A VGND VGND VPWR VPWR _099_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_left_track_1.prog_clk/X
+ hold48/X VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input51_A top_left_grid_pin_42_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input14_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input6_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_39.mux_l1_in_0_ input44/X input33/X hold24/A VGND VGND VPWR VPWR mux_left_track_39.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 input31/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_098_ _098_/A VGND VGND VPWR VPWR _098_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0__f_mem_left_track_1.prog_clk/X
+ hold26/X VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input44_A left_bottom_grid_pin_15_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_31.mux_l1_in_0__A0 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _070_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0__f_mem_left_track_1.prog_clk/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_21.sky130_fd_sc_hd__buf_4_0_ mux_left_track_21.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_097_ _097_/A VGND VGND VPWR VPWR _097_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_top_track_12.mux_l2_in_0__112 VGND VGND VPWR VPWR mux_top_track_12.mux_l2_in_0_/A0
+ mux_top_track_12.mux_l2_in_0__112/LO sky130_fd_sc_hd__conb_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3__f_mem_left_track_1.prog_clk/X
+ hold47/X VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_15.sky130_fd_sc_hd__buf_4_0_ mux_left_track_15.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _075_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_24.mux_l1_in_1__A1 input20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input37_A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ hold55/A VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_7.mux_l1_in_1__A0 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_left_track_1.prog_clk/X
+ mux_left_track_1.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_1_ mux_left_track_3.mux_l2_in_1_/A0 input44/X mux_left_track_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_096_ _096_/A VGND VGND VPWR VPWR _096_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0__f_mem_left_track_1.prog_clk/X
+ hold15/X VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l2_in_0_/A0 mux_top_track_16.mux_l1_in_0_/X
+ hold5/A VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6__f_mem_left_track_1.prog_clk/X
+ mux_top_track_4.mux_l1_in_2_/S VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_079_ _079_/A VGND VGND VPWR VPWR _079_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_11.mux_l2_in_0_ mux_left_track_11.mux_l2_in_0_/A0 mux_left_track_11.mux_l1_in_0_/X
+ hold14/A VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_37.sky130_fd_sc_hd__buf_4_0_ mux_left_track_37.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _086_/A sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7__f_mem_left_track_1.prog_clk/X
+ hold29/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__dfxtp_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_7.mux_l1_in_1__A1 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__103__A _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_left_track_1.prog_clk/X
+ hold4/X VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5__f_mem_left_track_1.prog_clk/X
+ hold18/X VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ mux_left_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input12_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input4_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.mux_l1_in_1_ input42/X input49/X mux_left_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_095_ _095_/A VGND VGND VPWR VPWR _095_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1__f_mem_left_track_1.prog_clk/X
+ mux_left_track_7.mux_l1_in_1_/S VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_left_track_1.prog_clk/X
+ hold43/X VGND VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_11.mux_l2_in_0__125 VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_0_/A0
+ mux_left_track_11.mux_l2_in_0__125/LO sky130_fd_sc_hd__conb_1
XANTENNA__106__A _106_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_078_ _078_/A VGND VGND VPWR VPWR _078_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_12.sky130_fd_sc_hd__buf_4_0_ mux_top_track_12.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _094_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input42_A left_bottom_grid_pin_11_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_16.mux_l1_in_0_ input5/X input55/X hold12/A VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_left_track_1.prog_clk/X
+ hold28/X VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__dfxtp_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_185 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6__f_mem_left_track_1.prog_clk/X
+ hold14/X VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_11.mux_l1_in_0_ input47/X input28/X hold17/A VGND VGND VPWR VPWR mux_left_track_11.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_23.mux_l2_in_0_ mux_left_track_23.mux_l2_in_0_/A0 mux_left_track_23.mux_l1_in_0_/X
+ hold51/A VGND VGND VPWR VPWR mux_left_track_23.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_55 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_left_track_1.prog_clk/X
+ hold33/X VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_1.mux_l2_in_1__124 VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/A0
+ mux_left_track_1.mux_l2_in_1__124/LO sky130_fd_sc_hd__conb_1
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_3.mux_l1_in_0_ input47/X input32/X mux_left_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_left_track_1.prog_clk/X
+ hold34/X VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_6.mux_l3_in_0_ mux_top_track_6.mux_l2_in_1_/X mux_top_track_6.mux_l2_in_0_/X
+ hold49/A VGND VGND VPWR VPWR mux_top_track_6.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
X_094_ _094_/A VGND VGND VPWR VPWR _094_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1__f_mem_left_track_1.prog_clk/X
+ hold20/X VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_3_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_077_ _077_/A VGND VGND VPWR VPWR _077_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_6.mux_l2_in_1_ mux_top_track_6.mux_l2_in_1_/A0 input10/X hold52/A VGND
+ VGND VPWR VPWR mux_top_track_6.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input35_A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_112 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_29.mux_l1_in_0__A0 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_67 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5__f_mem_left_track_1.prog_clk/X
+ hold38/X VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_23.mux_l2_in_0__131 VGND VGND VPWR VPWR mux_left_track_23.mux_l2_in_0_/A0
+ mux_left_track_23.mux_l2_in_0__131/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_23.mux_l1_in_0_ input44/X input41/X hold56/A VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3__f_mem_left_track_1.prog_clk/X
+ hold57/X VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_093_ _093_/A VGND VGND VPWR VPWR _093_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_35.mux_l2_in_0_ mux_left_track_35.mux_l2_in_0_/A0 mux_left_track_35.mux_l1_in_0_/X
+ hold58/A VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 ccff_head VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_076_ _076_/A VGND VGND VPWR VPWR _076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold42/X VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_37.mux_l1_in_0__A0 input43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l2_in_0_ mux_top_track_6.mux_l1_in_1_/X mux_top_track_6.mux_l1_in_0_/X
+ hold52/A VGND VGND VPWR VPWR mux_top_track_6.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input28_A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_6.mux_l2_in_1__122 VGND VGND VPWR VPWR mux_top_track_6.mux_l2_in_1_/A0
+ mux_top_track_6.mux_l2_in_1__122/LO sky130_fd_sc_hd__conb_1
XFILLER_12_124 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_6.sky130_fd_sc_hd__buf_4_0_ mux_top_track_6.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _091_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_6.mux_l1_in_1_ input58/X input56/X mux_top_track_6.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_6.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_39.mux_l2_in_0__106 VGND VGND VPWR VPWR mux_left_track_39.mux_l2_in_0_/A0
+ mux_left_track_39.mux_l2_in_0__106/LO sky130_fd_sc_hd__conb_1
Xclkbuf_3_4__f_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_3_4__f_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input10_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input2_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_211 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input58_A top_left_grid_pin_49_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_092_ _092_/A VGND VGND VPWR VPWR _092_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 chanx_left_in[0] VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_075_ _075_/A VGND VGND VPWR VPWR _075_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold40/X VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_10.mux_l1_in_0__A1 input52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_35.mux_l1_in_0_ input42/X input35/X hold36/A VGND VGND VPWR VPWR mux_left_track_35.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A0 input54/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input40_A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_6.mux_l1_in_0_ input54/X input52/X mux_top_track_6.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_6.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold37/X VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_0.mux_l1_in_2__A0 input2/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _068_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_091_ _091_/A VGND VGND VPWR VPWR _091_/X sky130_fd_sc_hd__clkbuf_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 chanx_left_in[10] VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_10.mux_l2_in_0__111 VGND VGND VPWR VPWR mux_top_track_10.mux_l2_in_0_/A0
+ mux_top_track_10.mux_l2_in_0__111/LO sky130_fd_sc_hd__conb_1
XFILLER_19_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_074_ _074_/A VGND VGND VPWR VPWR _074_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_11.mux_l1_in_0__A0 input47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4__f_mem_left_track_1.prog_clk/X
+ hold22/X VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput50 left_bottom_grid_pin_9_ VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 input52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input33_A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_11.sky130_fd_sc_hd__buf_4_0_ mux_left_track_11.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _073_/A sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold58/X VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_090_ _090_/A VGND VGND VPWR VPWR _090_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput4 chanx_left_in[11] VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.mux_l1_in_1__123 VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_1_/A0
+ mux_top_track_8.mux_l1_in_1__123/LO sky130_fd_sc_hd__conb_1
X_073_ _073_/A VGND VGND VPWR VPWR _073_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4__f_mem_left_track_1.prog_clk/X
+ hold9/X VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput40 chany_top_in[8] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
Xinput51 top_left_grid_pin_42_ VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input26_A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7__f_mem_left_track_1.prog_clk/X
+ hold32/X VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_12.mux_l2_in_0_ mux_top_track_12.mux_l2_in_0_/A0 mux_top_track_12.mux_l1_in_0_/X
+ hold27/A VGND VGND VPWR VPWR mux_top_track_12.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _084_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_9_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 chanx_left_in[12] VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A0 input57/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_27.sky130_fd_sc_hd__buf_4_0_ mux_left_track_27.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input56_A top_left_grid_pin_47_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_072_ _072_/A VGND VGND VPWR VPWR _072_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput41 chany_top_in[9] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_1
Xinput52 top_left_grid_pin_43_ VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__clkbuf_2
Xinput30 chany_top_in[17] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input19_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_107_ _107_/A VGND VGND VPWR VPWR _107_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_left_track_1.prog_clk/X
+ hold5/X VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_12.mux_l1_in_0_ input7/X input53/X hold22/A VGND VGND VPWR VPWR mux_top_track_12.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xinput6 chanx_left_in[13] VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_4.mux_l1_in_1__A1 input55/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ hold38/A VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_3.mux_l1_in_1__A0 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold56/X VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__dfxtp_1
X_071_ _071_/A VGND VGND VPWR VPWR _071_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input49_A left_bottom_grid_pin_7_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l2_in_0_/A0 mux_left_track_17.mux_l1_in_0_/X
+ hold57/A VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l1_in_1_ mux_top_track_24.mux_l1_in_1_/A0 input20/X mux_top_track_24.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A0 input5/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput20 chanx_left_in[8] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_1
Xinput31 chany_top_in[18] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_1
Xinput42 left_bottom_grid_pin_11_ VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_2
Xinput53 top_left_grid_pin_44_ VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_106_ _106_/A VGND VGND VPWR VPWR _106_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_9.mux_l2_in_0_ mux_left_track_9.mux_l1_in_1_/X mux_left_track_9.mux_l1_in_0_/X
+ hold2/A VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input31_A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ hold43/A VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l1_in_1_ mux_left_track_9.mux_l1_in_1_/A0 input45/X mux_left_track_9.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_21.mux_l2_in_0__130 VGND VGND VPWR VPWR mux_left_track_21.mux_l2_in_0_/A0
+ mux_left_track_21.mux_l2_in_0__130/LO sky130_fd_sc_hd__conb_1
XFILLER_6_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l2_in_1_ mux_top_track_2.mux_l2_in_1_/A0 input12/X mux_top_track_2.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput7 chanx_left_in[14] VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l1_in_1__A1 input49/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold3/X VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__dfxtp_1
X_070_ _070_/A VGND VGND VPWR VPWR _070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _100_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_51 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_0__f_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_3_0__f_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
Xmux_top_track_24.mux_l1_in_0_ input59/X input51/X mux_top_track_24.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A1 input55/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l2_in_1__121 VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/A0
+ mux_top_track_4.mux_l2_in_1__121/LO sky130_fd_sc_hd__conb_1
Xinput32 chany_top_in[19] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_1
Xinput21 chanx_left_in[9] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_1
Xinput43 left_bottom_grid_pin_13_ VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_2
Xinput10 chanx_left_in[17] VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_1
Xinput54 top_left_grid_pin_45_ VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_18.sky130_fd_sc_hd__buf_4_0_ mux_top_track_18.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _097_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_32_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_105_ _105_/A VGND VGND VPWR VPWR _105_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold10/X VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_17.mux_l1_in_0_ input50/X input25/X hold31/A VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_37.mux_l2_in_0__105 VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/A0
+ mux_left_track_37.mux_l2_in_0__105/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_29.mux_l2_in_0_ mux_left_track_29.mux_l2_in_0_/A0 mux_left_track_29.mux_l1_in_0_/X
+ hold40/A VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input24_A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_31.mux_l2_in_0_ mux_left_track_31.mux_l2_in_0_/A0 mux_left_track_31.mux_l1_in_0_/X
+ hold39/A VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l1_in_0_ input46/X input29/X mux_left_track_9.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l2_in_0_ mux_top_track_2.mux_l1_in_1_/X mux_top_track_2.mux_l1_in_0_/X
+ mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _089_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 chanx_left_in[15] VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6__f_mem_left_track_1.prog_clk/X
+ hold61/X VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_24.mux_l1_in_0__A1 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_63 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_2.mux_l1_in_1_ input58/X input56/X hold21/A VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input54_A top_left_grid_pin_45_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput55 top_left_grid_pin_46_ VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput44 left_bottom_grid_pin_15_ VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput11 chanx_left_in[18] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_1
Xinput33 chany_top_in[1] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
Xinput22 chany_top_in[0] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_24.mux_l1_in_1__119 VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/A0
+ mux_top_track_24.mux_l1_in_1__119/LO sky130_fd_sc_hd__conb_1
XFILLER_20_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0__f_mem_left_track_1.prog_clk/X
+ hold45/X VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_104_ _104_/A VGND VGND VPWR VPWR _104_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_7.mux_l1_in_0__A0 input47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input17_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input9_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_29.mux_l1_in_0_ input48/X input38/X hold10/A VGND VGND VPWR VPWR mux_left_track_29.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_31.mux_l1_in_0_ input49/X input37/X hold42/A VGND VGND VPWR VPWR mux_left_track_31.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 chanx_left_in[16] VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0__f_mem_left_track_1.prog_clk/X
+ mux_left_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4__f_mem_left_track_1.prog_clk/X
+ mux_top_track_0.mux_l1_in_2_/S VGND VGND VPWR VPWR hold61/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5__f_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_3_5__f_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_25_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_2.mux_l1_in_0_ input54/X input52/X hold21/A VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input47_A left_bottom_grid_pin_3_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput45 left_bottom_grid_pin_17_ VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput12 chanx_left_in[19] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_1
Xinput23 chany_top_in[10] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_1
Xinput34 chany_top_in[2] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_1
Xinput56 top_left_grid_pin_47_ VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_103_ _103_/A VGND VGND VPWR VPWR _103_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_7.mux_l1_in_0__A1 input30/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4__f_mem_left_track_1.prog_clk/X
+ hold52/X VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__dfxtp_1
XFILLER_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 input43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_left_track_1.prog_clk/X
+ mux_left_track_3.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5__f_mem_left_track_1.prog_clk/X
+ input1/X VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output60_A output60/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput100 _097_/X VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
Xinput13 chanx_left_in[1] VGND VGND VPWR VPWR _107_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput35 chany_top_in[3] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
Xinput57 top_left_grid_pin_48_ VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput46 left_bottom_grid_pin_1_ VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput24 chany_top_in[11] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_102_ _102_/A VGND VGND VPWR VPWR _102_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6__f_mem_left_track_1.prog_clk/X
+ mux_top_track_6.mux_l1_in_1_/S VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_22_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7__f_mem_left_track_1.prog_clk/X
+ hold41/X VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input22_A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_left_track_1.prog_clk/X
+ hold23/X VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__dfxtp_1
XFILLER_30_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0__f_mem_left_track_1.prog_clk/X
+ hold53/X VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_19.mux_l2_in_0__129 VGND VGND VPWR VPWR mux_left_track_19.mux_l2_in_0_/A0
+ mux_left_track_19.mux_l2_in_0__129/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_7.sky130_fd_sc_hd__buf_4_0_ mux_left_track_7.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _071_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__107__A _107_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput14 chanx_left_in[2] VGND VGND VPWR VPWR _106_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput25 chany_top_in[12] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
Xinput36 chany_top_in[4] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__clkbuf_1
Xinput58 top_left_grid_pin_49_ VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput47 left_bottom_grid_pin_3_ VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__dlymetal6s2s_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1__f_mem_left_track_1.prog_clk/X
+ mux_left_track_9.mux_l1_in_1_/S VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_101_ _101_/A VGND VGND VPWR VPWR _101_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input52_A top_left_grid_pin_43_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6__f_mem_left_track_1.prog_clk/X
+ hold11/X VGND VGND VPWR VPWR mux_top_track_6.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_8_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_87 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_23.sky130_fd_sc_hd__buf_4_0_ mux_left_track_23.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _079_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_33_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_left_track_1.prog_clk/X
+ hold46/X VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _076_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input15_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input7_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ hold20/A VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3__f_mem_left_track_1.prog_clk/X
+ hold19/X VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__dfxtp_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l2_in_1_/A0 mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput59 top_right_grid_pin_1_ VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput15 chanx_left_in[3] VGND VGND VPWR VPWR _105_/A sky130_fd_sc_hd__clkbuf_1
Xinput48 left_bottom_grid_pin_5_ VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_2
Xinput37 chany_top_in[5] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
Xinput26 chany_top_in[13] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1__f_mem_left_track_1.prog_clk/X
+ hold60/X VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_11_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_100_ _100_/A VGND VGND VPWR VPWR _100_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input45_A left_bottom_grid_pin_17_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_2_ input45/X input43/X mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_99 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_18.mux_l2_in_0_ mux_top_track_18.mux_l2_in_0_/A0 mux_top_track_18.mux_l1_in_0_/X
+ hold28/A VGND VGND VPWR VPWR mux_top_track_18.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_top_track_20.mux_l2_in_0_ mux_top_track_20.mux_l2_in_0_/A0 mux_top_track_20.mux_l1_in_0_/X
+ hold46/A VGND VGND VPWR VPWR mux_top_track_20.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_13.mux_l2_in_0_ mux_left_track_13.mux_l2_in_0_/A0 mux_left_track_13.mux_l1_in_0_/X
+ hold19/A VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_39.sky130_fd_sc_hd__buf_4_0_ mux_left_track_39.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _087_/A sky130_fd_sc_hd__clkbuf_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput16 chanx_left_in[4] VGND VGND VPWR VPWR _104_/A sky130_fd_sc_hd__clkbuf_1
Xinput49 left_bottom_grid_pin_7_ VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_2
Xinput38 chany_top_in[6] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_1
Xinput27 chany_top_in[14] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input38_A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_1_ input50/X input48/X mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_35.mux_l2_in_0__104 VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/A0
+ mux_left_track_35.mux_l2_in_0__104/LO sky130_fd_sc_hd__conb_1
XFILLER_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1__A0 input57/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_20.sky130_fd_sc_hd__buf_4_0_ mux_top_track_20.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _098_/A sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold50/X VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__dfxtp_1
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_14.sky130_fd_sc_hd__buf_4_0_ mux_top_track_14.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _095_/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_18.mux_l1_in_0_ input4/X input56/X hold32/A VGND VGND VPWR VPWR mux_top_track_18.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input20_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_20.mux_l1_in_0_ input3/X input57/X hold29/A VGND VGND VPWR VPWR mux_top_track_20.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_13.mux_l1_in_0_ input48/X input27/X hold4/A VGND VGND VPWR VPWR mux_left_track_13.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_32_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ hold26/A VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput17 chanx_left_in[5] VGND VGND VPWR VPWR _103_/A sky130_fd_sc_hd__clkbuf_1
Xinput39 chany_top_in[7] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__clkbuf_1
Xinput28 chany_top_in[15] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l1_in_0_ input46/X input31/X mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_1_ mux_left_track_25.mux_l1_in_1_/A0 input45/X hold16/A
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_089_ _089_/A VGND VGND VPWR VPWR _089_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_0.mux_l1_in_1__A1 input55/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold39/X VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input50_A left_bottom_grid_pin_9_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_1__f_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_3_1__f_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_30_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input13_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_18.mux_l2_in_0__115 VGND VGND VPWR VPWR mux_top_track_18.mux_l2_in_0_/A0
+ mux_top_track_18.mux_l2_in_0__115/LO sky130_fd_sc_hd__conb_1
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold24/X VGND VGND VPWR VPWR output60/A sky130_fd_sc_hd__dfxtp_1
XFILLER_2_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input5_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 chanx_left_in[6] VGND VGND VPWR VPWR _102_/A sky130_fd_sc_hd__clkbuf_1
Xinput29 chany_top_in[16] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_0_ input46/X input40/X hold16/A VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_088_ _088_/A VGND VGND VPWR VPWR _088_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_37.mux_l2_in_0_ mux_left_track_37.mux_l2_in_0_/A0 mux_left_track_37.mux_l1_in_0_/X
+ hold54/A VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_left_track_1.prog_clk/X
+ hold8/X VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input43_A left_bottom_grid_pin_13_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_30_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_20.mux_l1_in_0__A0 input3/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_8.mux_l2_in_0_ mux_top_track_8.mux_l1_in_1_/X mux_top_track_8.mux_l1_in_0_/X
+ hold7/A VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_12.mux_l1_in_0__A1 input53/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_left_track_1.prog_clk/X
+ hold54/X VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 input53/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_1_ mux_top_track_8.mux_l1_in_1_/A0 input9/X mux_top_track_8.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _092_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_32_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 chanx_left_in[7] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_087_ _087_/A VGND VGND VPWR VPWR _087_/X sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4__f_mem_left_track_1.prog_clk/X
+ hold27/X VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dfxtp_1
XFILLER_16_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input36_A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xclkbuf_3_6__f_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_3_6__f_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XANTENNA_mux_top_track_20.mux_l1_in_0__A1 input57/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_22.mux_l2_in_0__118 VGND VGND VPWR VPWR mux_top_track_22.mux_l2_in_0_/A0
+ mux_top_track_22.mux_l2_in_0__118/LO sky130_fd_sc_hd__conb_1
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_13.mux_l1_in_0__A0 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_37.mux_l1_in_0_ input43/X input34/X hold37/A VGND VGND VPWR VPWR mux_left_track_37.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_17.mux_l2_in_0__128 VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/A0
+ mux_left_track_17.mux_l2_in_0__128/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_3.mux_l1_in_0__A0 input47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__077__A _077_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_0_ input59/X input51/X mux_top_track_8.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_086_ _086_/A VGND VGND VPWR VPWR _086_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_2.mux_l2_in_1__A1 input12/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _069_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_21.mux_l1_in_0__A0 input43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_15_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input29_A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_069_ _069_/A VGND VGND VPWR VPWR _069_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_71 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 input32/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input11_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput90 _106_/X VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
XFILLER_23_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input3_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_2__A1 input43/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_13.sky130_fd_sc_hd__buf_4_0_ mux_left_track_13.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _074_/A sky130_fd_sc_hd__clkbuf_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input59_A top_right_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_left_track_1.prog_clk/X
+ hold16/X VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__dfxtp_1
X_085_ _085_/A VGND VGND VPWR VPWR _085_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ hold53/A VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_068_ _068_/A VGND VGND VPWR VPWR _068_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_6.mux_l1_in_1__A0 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_29.mux_l2_in_0__134 VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/A0
+ mux_left_track_29.mux_l2_in_0__134/LO sky130_fd_sc_hd__conb_1
XFILLER_28_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input41_A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_1_ mux_left_track_1.mux_l2_in_1_/A0 mux_left_track_1.mux_l1_in_2_/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_2_ input45/X input43/X mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xoutput80 _077_/X VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
Xoutput91 _107_/X VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
XFILLER_23_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_14.mux_l2_in_0_ mux_top_track_14.mux_l2_in_0_/A0 mux_top_track_14.mux_l1_in_0_/X
+ hold6/A VGND VGND VPWR VPWR mux_top_track_14.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_35.sky130_fd_sc_hd__buf_4_0_ mux_left_track_35.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _085_/A sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1__f_mem_left_track_1.prog_clk/X
+ hold51/X VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dfxtp_1
X_084_ _084_/A VGND VGND VPWR VPWR _084_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.mux_l2_in_0__103 VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/A0
+ mux_left_track_33.mux_l2_in_0__103/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_39.mux_l2_in_0__S output60/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_6.mux_l1_in_1__A1 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_29.sky130_fd_sc_hd__buf_4_0_ mux_left_track_29.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _082_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input34_A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_18.mux_l1_in_0__A0 input4/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_1.mux_l1_in_1_ input50/X input48/X mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput70 _086_/X VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
Xoutput92 _089_/X VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
Xoutput81 _088_/X VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
XFILLER_31_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_2.mux_l2_in_1__116 VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/A0
+ mux_top_track_2.mux_l2_in_1__116/LO sky130_fd_sc_hd__conb_1
XFILLER_9_100 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_10.sky130_fd_sc_hd__buf_4_0_ mux_top_track_10.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _093_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_083_ _083_/A VGND VGND VPWR VPWR _083_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7__f_mem_left_track_1.prog_clk/X
+ mux_top_track_2.mux_l2_in_1_/S VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_14.mux_l1_in_0_ input6/X input54/X hold8/A VGND VGND VPWR VPWR mux_top_track_14.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_7.mux_l2_in_1__108 VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/A0
+ mux_left_track_7.mux_l2_in_1__108/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_26.mux_l2_in_0_ mux_top_track_26.mux_l2_in_0_/A0 mux_top_track_26.mux_l1_in_0_/X
+ hold18/A VGND VGND VPWR VPWR mux_top_track_26.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A1 input48/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_26.mux_l1_in_0__A0 input19/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_19.mux_l2_in_0_ mux_left_track_19.mux_l2_in_0_/A0 mux_left_track_19.mux_l1_in_0_/X
+ hold1/A VGND VGND VPWR VPWR mux_left_track_19.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input27_A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_21.mux_l2_in_0_ mux_left_track_21.mux_l2_in_0_/A0 mux_left_track_21.mux_l1_in_0_/X
+ hold3/A VGND VGND VPWR VPWR mux_left_track_21.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_16.mux_l2_in_0__114 VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/A0
+ mux_top_track_16.mux_l2_in_0__114/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_18.mux_l1_in_0__A1 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_0_ input46/X input22/X mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xoutput82 _098_/X VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
Xoutput93 _090_/X VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
Xoutput71 _087_/X VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
Xoutput60 output60/A VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_2
XFILLER_31_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ hold11/A VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1__110 VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/A0
+ mux_top_track_0.mux_l2_in_1__110/LO sky130_fd_sc_hd__conb_1
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input1_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1__f_mem_left_track_1.prog_clk/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_082_ _082_/A VGND VGND VPWR VPWR _082_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input57_A top_left_grid_pin_48_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7__f_mem_left_track_1.prog_clk/X
+ hold21/X VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_1_ mux_top_track_4.mux_l2_in_1_/A0 mux_top_track_4.mux_l1_in_2_/X
+ hold47/A VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_26.mux_l1_in_0__A1 input52/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_2_ input11/X input59/X mux_top_track_4.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_26.sky130_fd_sc_hd__buf_4_0_ mux_top_track_26.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _101_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_19.mux_l1_in_0__A0 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_26.mux_l1_in_0_ input19/X input52/X hold33/A VGND VGND VPWR VPWR mux_top_track_26.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1__f_mem_left_track_1.prog_clk/X
+ hold17/X VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dfxtp_1
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_19.mux_l1_in_0_ input42/X input24/X hold34/A VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_1_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput94 _091_/X VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
Xoutput83 _099_/X VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
XANTENNA__102__A _102_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput61 _068_/X VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
Xoutput72 _069_/X VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
Xmux_left_track_21.mux_l1_in_0_ input43/X input23/X hold25/A VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_16_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l2_in_0_/A0 mux_left_track_33.mux_l1_in_0_/X
+ hold30/A VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2__f_mem_left_track_1.prog_clk clkbuf_0_mem_left_track_1.prog_clk/X VGND
+ VGND VPWR VPWR clkbuf_3_2__f_mem_left_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_left_track_1.prog_clk/X
+ mux_left_track_5.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_081_ _081_/A VGND VGND VPWR VPWR _081_/X sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6__f_mem_left_track_1.prog_clk/X
+ hold59/X VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ hold47/A VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _090_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_2_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_27.mux_l1_in_0__A0 input47/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_20.mux_l2_in_0__117 VGND VGND VPWR VPWR mux_top_track_20.mux_l2_in_0_/A0
+ mux_top_track_20.mux_l2_in_0__117/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_4.mux_l1_in_1_ input57/X input55/X mux_top_track_4.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4__f_mem_left_track_1.prog_clk/X
+ mux_top_track_8.mux_l1_in_1_/S VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0__f_mem_left_track_1.prog_clk/X
+ hold2/X VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input32_A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold61 hold61/A VGND VGND VPWR VPWR hold61/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_15.mux_l2_in_0__127 VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_0_/A0
+ mux_left_track_15.mux_l2_in_0__127/LO sky130_fd_sc_hd__conb_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_left_track_1.prog_clk/X
+ mux_top_track_24.mux_l1_in_1_/S VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__dfxtp_1
XFILLER_25_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput84 _100_/X VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
Xoutput95 _092_/X VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
Xoutput62 _078_/X VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
Xoutput73 _070_/X VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
XFILLER_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_9.mux_l1_in_1__109 VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_1_/A0
+ mux_left_track_9.mux_l1_in_1__109/LO sky130_fd_sc_hd__conb_1
XFILLER_3_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_left_track_1.prog_clk/X
+ hold31/X VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0__f_mem_left_track_1.prog_clk/X
+ hold55/X VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_35.mux_l1_in_0__A0 input42/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_080_ _080_/A VGND VGND VPWR VPWR _080_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_33.mux_l1_in_0_ input50/X input36/X hold50/A VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l1_in_0_ input53/X input51/X mux_top_track_4.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4__f_mem_left_track_1.prog_clk/X
+ hold49/X VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input25_A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5__f_mem_left_track_1.prog_clk/X
+ hold13/X VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_25_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput85 _101_/X VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
Xoutput96 _093_/X VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
Xoutput63 _079_/X VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
Xoutput74 _071_/X VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
XFILLER_16_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

