magic
tech sky130A
magscale 1 2
timestamp 1650625003
<< viali >>
rect 4537 20553 4571 20587
rect 11161 20553 11195 20587
rect 13001 20553 13035 20587
rect 13645 20553 13679 20587
rect 15577 20553 15611 20587
rect 16773 20553 16807 20587
rect 17325 20553 17359 20587
rect 19349 20553 19383 20587
rect 20545 20553 20579 20587
rect 21097 20553 21131 20587
rect 1685 20485 1719 20519
rect 9045 20485 9079 20519
rect 2329 20417 2363 20451
rect 2789 20417 2823 20451
rect 3249 20417 3283 20451
rect 3893 20417 3927 20451
rect 4353 20417 4387 20451
rect 5457 20417 5491 20451
rect 5825 20417 5859 20451
rect 6561 20417 6595 20451
rect 7021 20417 7055 20451
rect 7481 20417 7515 20451
rect 7941 20417 7975 20451
rect 9321 20417 9355 20451
rect 9873 20417 9907 20451
rect 10425 20417 10459 20451
rect 10977 20417 11011 20451
rect 11529 20417 11563 20451
rect 12633 20417 12667 20451
rect 13185 20417 13219 20451
rect 13461 20417 13495 20451
rect 14841 20417 14875 20451
rect 15761 20417 15795 20451
rect 16313 20417 16347 20451
rect 16957 20417 16991 20451
rect 17509 20417 17543 20451
rect 18061 20417 18095 20451
rect 18613 20417 18647 20451
rect 19533 20417 19567 20451
rect 20085 20417 20119 20451
rect 20361 20417 20395 20451
rect 20913 20417 20947 20451
rect 1869 20349 1903 20383
rect 14657 20349 14691 20383
rect 14749 20349 14783 20383
rect 6745 20281 6779 20315
rect 10609 20281 10643 20315
rect 15209 20281 15243 20315
rect 18429 20281 18463 20315
rect 2513 20213 2547 20247
rect 2973 20213 3007 20247
rect 3433 20213 3467 20247
rect 4077 20213 4111 20247
rect 4813 20213 4847 20247
rect 6009 20213 6043 20247
rect 7205 20213 7239 20247
rect 7665 20213 7699 20247
rect 8585 20213 8619 20247
rect 9505 20213 9539 20247
rect 10057 20213 10091 20247
rect 11713 20213 11747 20247
rect 11989 20213 12023 20247
rect 14197 20213 14231 20247
rect 16129 20213 16163 20247
rect 17877 20213 17911 20247
rect 19901 20213 19935 20247
rect 1685 20009 1719 20043
rect 2789 20009 2823 20043
rect 10333 20009 10367 20043
rect 11989 20009 12023 20043
rect 12449 20009 12483 20043
rect 14197 20009 14231 20043
rect 19349 20009 19383 20043
rect 19901 20009 19935 20043
rect 8033 19941 8067 19975
rect 16129 19941 16163 19975
rect 4169 19873 4203 19907
rect 4261 19873 4295 19907
rect 9045 19873 9079 19907
rect 16865 19873 16899 19907
rect 16957 19873 16991 19907
rect 1501 19805 1535 19839
rect 1961 19805 1995 19839
rect 2605 19805 2639 19839
rect 3249 19805 3283 19839
rect 4997 19805 5031 19839
rect 6653 19805 6687 19839
rect 10609 19805 10643 19839
rect 12265 19805 12299 19839
rect 13093 19805 13127 19839
rect 14381 19805 14415 19839
rect 14749 19805 14783 19839
rect 18889 19805 18923 19839
rect 19533 19805 19567 19839
rect 20085 19805 20119 19839
rect 20545 19805 20579 19839
rect 21097 19805 21131 19839
rect 5264 19737 5298 19771
rect 6920 19737 6954 19771
rect 8585 19737 8619 19771
rect 9321 19737 9355 19771
rect 10876 19737 10910 19771
rect 15016 19737 15050 19771
rect 16773 19737 16807 19771
rect 17417 19737 17451 19771
rect 18061 19737 18095 19771
rect 2145 19669 2179 19703
rect 3433 19669 3467 19703
rect 4353 19669 4387 19703
rect 4721 19669 4755 19703
rect 6377 19669 6411 19703
rect 9229 19669 9263 19703
rect 9689 19669 9723 19703
rect 13737 19669 13771 19703
rect 16405 19669 16439 19703
rect 20729 19669 20763 19703
rect 21281 19669 21315 19703
rect 1777 19465 1811 19499
rect 3157 19465 3191 19499
rect 7021 19465 7055 19499
rect 8585 19465 8619 19499
rect 9045 19465 9079 19499
rect 9597 19465 9631 19499
rect 13093 19465 13127 19499
rect 16129 19465 16163 19499
rect 20085 19465 20119 19499
rect 20729 19465 20763 19499
rect 2789 19397 2823 19431
rect 2053 19329 2087 19363
rect 3433 19329 3467 19363
rect 3700 19329 3734 19363
rect 5457 19329 5491 19363
rect 6377 19329 6411 19363
rect 7297 19329 7331 19363
rect 8677 19329 8711 19363
rect 9689 19329 9723 19363
rect 10333 19329 10367 19363
rect 11713 19329 11747 19363
rect 11980 19329 12014 19363
rect 13369 19329 13403 19363
rect 13636 19329 13670 19363
rect 15025 19329 15059 19363
rect 15945 19329 15979 19363
rect 17325 19329 17359 19363
rect 17601 19329 17635 19363
rect 18613 19329 18647 19363
rect 18889 19329 18923 19363
rect 19717 19329 19751 19363
rect 20269 19329 20303 19363
rect 20545 19329 20579 19363
rect 21097 19329 21131 19363
rect 5549 19261 5583 19295
rect 5641 19261 5675 19295
rect 8401 19261 8435 19295
rect 9505 19261 9539 19295
rect 15669 19261 15703 19295
rect 4813 19193 4847 19227
rect 10977 19193 11011 19227
rect 14749 19193 14783 19227
rect 18429 19193 18463 19227
rect 19073 19193 19107 19227
rect 19533 19193 19567 19227
rect 2237 19125 2271 19159
rect 5089 19125 5123 19159
rect 7481 19125 7515 19159
rect 8033 19125 8067 19159
rect 10057 19125 10091 19159
rect 16681 19125 16715 19159
rect 17785 19125 17819 19159
rect 21281 19125 21315 19159
rect 1777 18921 1811 18955
rect 3801 18921 3835 18955
rect 5273 18921 5307 18955
rect 5733 18921 5767 18955
rect 6193 18921 6227 18955
rect 7389 18921 7423 18955
rect 7849 18921 7883 18955
rect 8125 18921 8159 18955
rect 8585 18921 8619 18955
rect 13737 18921 13771 18955
rect 15393 18921 15427 18955
rect 18705 18921 18739 18955
rect 20177 18921 20211 18955
rect 20637 18921 20671 18955
rect 6653 18853 6687 18887
rect 7113 18853 7147 18887
rect 19533 18853 19567 18887
rect 4997 18785 5031 18819
rect 11989 18785 12023 18819
rect 13093 18785 13127 18819
rect 15669 18785 15703 18819
rect 2053 18717 2087 18751
rect 4445 18717 4479 18751
rect 6929 18717 6963 18751
rect 9505 18717 9539 18751
rect 15209 18717 15243 18751
rect 15936 18717 15970 18751
rect 17325 18717 17359 18751
rect 18245 18717 18279 18751
rect 18889 18717 18923 18751
rect 19717 18717 19751 18751
rect 19993 18717 20027 18751
rect 20821 18717 20855 18751
rect 21097 18717 21131 18751
rect 2320 18649 2354 18683
rect 9772 18649 9806 18683
rect 12081 18649 12115 18683
rect 12173 18649 12207 18683
rect 13369 18649 13403 18683
rect 14105 18649 14139 18683
rect 3433 18581 3467 18615
rect 9229 18581 9263 18615
rect 10885 18581 10919 18615
rect 11161 18581 11195 18615
rect 12541 18581 12575 18615
rect 13277 18581 13311 18615
rect 14565 18581 14599 18615
rect 17049 18581 17083 18615
rect 17969 18581 18003 18615
rect 18429 18581 18463 18615
rect 21281 18581 21315 18615
rect 2053 18377 2087 18411
rect 2697 18377 2731 18411
rect 3157 18377 3191 18411
rect 4261 18377 4295 18411
rect 7205 18377 7239 18411
rect 9505 18377 9539 18411
rect 10701 18377 10735 18411
rect 10793 18377 10827 18411
rect 12173 18377 12207 18411
rect 18337 18377 18371 18411
rect 19625 18377 19659 18411
rect 20729 18377 20763 18411
rect 3433 18309 3467 18343
rect 17224 18309 17258 18343
rect 1685 18241 1719 18275
rect 4813 18241 4847 18275
rect 6837 18241 6871 18275
rect 7481 18241 7515 18275
rect 8125 18241 8159 18275
rect 8392 18241 8426 18275
rect 10057 18241 10091 18275
rect 11529 18241 11563 18275
rect 16129 18241 16163 18275
rect 18981 18241 19015 18275
rect 19993 18241 20027 18275
rect 20545 18241 20579 18275
rect 21097 18241 21131 18275
rect 6561 18173 6595 18207
rect 6745 18173 6779 18207
rect 10609 18173 10643 18207
rect 16957 18173 16991 18207
rect 19073 18173 19107 18207
rect 19165 18173 19199 18207
rect 11161 18105 11195 18139
rect 18613 18105 18647 18139
rect 20177 18105 20211 18139
rect 21281 18105 21315 18139
rect 1501 18037 1535 18071
rect 4997 18037 5031 18071
rect 12725 18037 12759 18071
rect 15301 18037 15335 18071
rect 16313 18037 16347 18071
rect 2329 17833 2363 17867
rect 7113 17833 7147 17867
rect 10333 17833 10367 17867
rect 17509 17833 17543 17867
rect 19441 17833 19475 17867
rect 2605 17765 2639 17799
rect 17969 17765 18003 17799
rect 18889 17765 18923 17799
rect 6285 17697 6319 17731
rect 7573 17697 7607 17731
rect 7757 17697 7791 17731
rect 11621 17697 11655 17731
rect 11805 17697 11839 17731
rect 16957 17697 16991 17731
rect 1685 17629 1719 17663
rect 17049 17629 17083 17663
rect 17785 17629 17819 17663
rect 18245 17629 18279 17663
rect 18705 17629 18739 17663
rect 19257 17629 19291 17663
rect 19717 17629 19751 17663
rect 20545 17629 20579 17663
rect 21097 17629 21131 17663
rect 6040 17561 6074 17595
rect 11897 17561 11931 17595
rect 3157 17493 3191 17527
rect 4905 17493 4939 17527
rect 7481 17493 7515 17527
rect 8217 17493 8251 17527
rect 12265 17493 12299 17527
rect 12633 17493 12667 17527
rect 14749 17493 14783 17527
rect 16497 17493 16531 17527
rect 17141 17493 17175 17527
rect 18429 17493 18463 17527
rect 19901 17493 19935 17527
rect 20729 17493 20763 17527
rect 21281 17493 21315 17527
rect 3709 17289 3743 17323
rect 4997 17289 5031 17323
rect 14657 17289 14691 17323
rect 15209 17289 15243 17323
rect 17785 17289 17819 17323
rect 18981 17289 19015 17323
rect 19625 17289 19659 17323
rect 20085 17289 20119 17323
rect 3617 17221 3651 17255
rect 4353 17221 4387 17255
rect 12633 17221 12667 17255
rect 14197 17221 14231 17255
rect 2717 17153 2751 17187
rect 5641 17153 5675 17187
rect 9229 17153 9263 17187
rect 12725 17153 12759 17187
rect 13369 17153 13403 17187
rect 14289 17153 14323 17187
rect 15301 17153 15335 17187
rect 15945 17153 15979 17187
rect 16681 17153 16715 17187
rect 18705 17153 18739 17187
rect 19165 17153 19199 17187
rect 19441 17153 19475 17187
rect 19901 17153 19935 17187
rect 20545 17153 20579 17187
rect 21097 17153 21131 17187
rect 2973 17085 3007 17119
rect 3893 17085 3927 17119
rect 10149 17085 10183 17119
rect 12449 17085 12483 17119
rect 14013 17085 14047 17119
rect 15117 17085 15151 17119
rect 20361 17017 20395 17051
rect 1593 16949 1627 16983
rect 3249 16949 3283 16983
rect 8677 16949 8711 16983
rect 9873 16949 9907 16983
rect 13093 16949 13127 16983
rect 15669 16949 15703 16983
rect 17325 16949 17359 16983
rect 18061 16949 18095 16983
rect 21281 16949 21315 16983
rect 20821 16745 20855 16779
rect 15485 16677 15519 16711
rect 17233 16677 17267 16711
rect 2789 16609 2823 16643
rect 2973 16609 3007 16643
rect 4537 16609 4571 16643
rect 7941 16609 7975 16643
rect 8125 16609 8159 16643
rect 9229 16609 9263 16643
rect 10701 16609 10735 16643
rect 12357 16609 12391 16643
rect 14105 16609 14139 16643
rect 16681 16609 16715 16643
rect 18153 16609 18187 16643
rect 18245 16609 18279 16643
rect 3065 16541 3099 16575
rect 3801 16541 3835 16575
rect 4804 16541 4838 16575
rect 6193 16541 6227 16575
rect 8217 16541 8251 16575
rect 10149 16541 10183 16575
rect 16773 16541 16807 16575
rect 19901 16541 19935 16575
rect 20177 16541 20211 16575
rect 20637 16541 20671 16575
rect 21097 16541 21131 16575
rect 9505 16473 9539 16507
rect 10968 16473 11002 16507
rect 12624 16473 12658 16507
rect 14372 16473 14406 16507
rect 18337 16473 18371 16507
rect 19257 16473 19291 16507
rect 3433 16405 3467 16439
rect 3985 16405 4019 16439
rect 5917 16405 5951 16439
rect 6837 16405 6871 16439
rect 8585 16405 8619 16439
rect 9413 16405 9447 16439
rect 9873 16405 9907 16439
rect 10333 16405 10367 16439
rect 12081 16405 12115 16439
rect 13737 16405 13771 16439
rect 16865 16405 16899 16439
rect 17509 16405 17543 16439
rect 18705 16405 18739 16439
rect 19717 16405 19751 16439
rect 20361 16405 20395 16439
rect 21281 16405 21315 16439
rect 9229 16201 9263 16235
rect 12725 16201 12759 16235
rect 14381 16201 14415 16235
rect 16313 16201 16347 16235
rect 18061 16201 18095 16235
rect 19441 16201 19475 16235
rect 20085 16201 20119 16235
rect 20637 16201 20671 16235
rect 8094 16133 8128 16167
rect 16948 16133 16982 16167
rect 1777 16065 1811 16099
rect 2044 16065 2078 16099
rect 4077 16065 4111 16099
rect 6929 16065 6963 16099
rect 9781 16065 9815 16099
rect 10037 16065 10071 16099
rect 12081 16065 12115 16099
rect 13737 16065 13771 16099
rect 14933 16065 14967 16099
rect 15200 16065 15234 16099
rect 16681 16065 16715 16099
rect 19625 16065 19659 16099
rect 19901 16065 19935 16099
rect 20821 16065 20855 16099
rect 21097 16065 21131 16099
rect 3433 15997 3467 16031
rect 6745 15997 6779 16031
rect 6837 15997 6871 16031
rect 7849 15997 7883 16031
rect 3157 15929 3191 15963
rect 11161 15929 11195 15963
rect 7297 15861 7331 15895
rect 21281 15861 21315 15895
rect 2237 15657 2271 15691
rect 5733 15657 5767 15691
rect 8401 15657 8435 15691
rect 11161 15657 11195 15691
rect 16129 15657 16163 15691
rect 20361 15657 20395 15691
rect 19901 15589 19935 15623
rect 20821 15589 20855 15623
rect 3893 15521 3927 15555
rect 7297 15521 7331 15555
rect 17509 15521 17543 15555
rect 2881 15453 2915 15487
rect 7757 15453 7791 15487
rect 11805 15453 11839 15487
rect 15485 15453 15519 15487
rect 17776 15453 17810 15487
rect 19717 15453 19751 15487
rect 20177 15453 20211 15487
rect 20637 15453 20671 15487
rect 21097 15453 21131 15487
rect 4169 15385 4203 15419
rect 4813 15385 4847 15419
rect 7021 15385 7055 15419
rect 4077 15317 4111 15351
rect 4537 15317 4571 15351
rect 18889 15317 18923 15351
rect 21281 15317 21315 15351
rect 2145 15113 2179 15147
rect 4169 15113 4203 15147
rect 7757 15113 7791 15147
rect 20269 15113 20303 15147
rect 20821 15113 20855 15147
rect 4629 15045 4663 15079
rect 3258 14977 3292 15011
rect 3525 14977 3559 15011
rect 4537 14977 4571 15011
rect 6644 14977 6678 15011
rect 8677 14977 8711 15011
rect 9413 14977 9447 15011
rect 12817 14977 12851 15011
rect 14841 14977 14875 15011
rect 20085 14977 20119 15011
rect 20637 14977 20671 15011
rect 21097 14977 21131 15011
rect 4721 14909 4755 14943
rect 6377 14909 6411 14943
rect 12541 14909 12575 14943
rect 12725 14909 12759 14943
rect 15669 14909 15703 14943
rect 9597 14841 9631 14875
rect 5273 14773 5307 14807
rect 8033 14773 8067 14807
rect 13185 14773 13219 14807
rect 14197 14773 14231 14807
rect 21281 14773 21315 14807
rect 3801 14569 3835 14603
rect 7021 14569 7055 14603
rect 9689 14569 9723 14603
rect 15485 14569 15519 14603
rect 20269 14569 20303 14603
rect 20821 14569 20855 14603
rect 6745 14501 6779 14535
rect 8125 14501 8159 14535
rect 7573 14433 7607 14467
rect 9045 14433 9079 14467
rect 11437 14433 11471 14467
rect 12081 14433 12115 14467
rect 16313 14433 16347 14467
rect 4445 14365 4479 14399
rect 5365 14365 5399 14399
rect 7389 14365 7423 14399
rect 7481 14365 7515 14399
rect 14105 14365 14139 14399
rect 16129 14365 16163 14399
rect 20085 14365 20119 14399
rect 20637 14365 20671 14399
rect 21097 14365 21131 14399
rect 5632 14297 5666 14331
rect 9229 14297 9263 14331
rect 11192 14297 11226 14331
rect 12326 14297 12360 14331
rect 14372 14297 14406 14331
rect 9321 14229 9355 14263
rect 10057 14229 10091 14263
rect 13461 14229 13495 14263
rect 15761 14229 15795 14263
rect 16221 14229 16255 14263
rect 16865 14229 16899 14263
rect 21281 14229 21315 14263
rect 3709 14025 3743 14059
rect 6745 14025 6779 14059
rect 9045 14025 9079 14059
rect 9781 14025 9815 14059
rect 13093 14025 13127 14059
rect 15117 14025 15151 14059
rect 15485 14025 15519 14059
rect 16037 14025 16071 14059
rect 19717 14025 19751 14059
rect 4844 13957 4878 13991
rect 10241 13957 10275 13991
rect 15025 13957 15059 13991
rect 17592 13957 17626 13991
rect 19349 13957 19383 13991
rect 5089 13889 5123 13923
rect 7389 13889 7423 13923
rect 7932 13889 7966 13923
rect 10149 13889 10183 13923
rect 10793 13889 10827 13923
rect 12725 13889 12759 13923
rect 13369 13889 13403 13923
rect 15853 13889 15887 13923
rect 17325 13889 17359 13923
rect 19257 13889 19291 13923
rect 20637 13889 20671 13923
rect 21097 13889 21131 13923
rect 7665 13821 7699 13855
rect 10333 13821 10367 13855
rect 11621 13821 11655 13855
rect 12541 13821 12575 13855
rect 12633 13821 12667 13855
rect 13829 13821 13863 13855
rect 14933 13821 14967 13855
rect 19073 13821 19107 13855
rect 19993 13821 20027 13855
rect 18705 13685 18739 13719
rect 20821 13685 20855 13719
rect 21281 13685 21315 13719
rect 5917 13481 5951 13515
rect 9689 13481 9723 13515
rect 13093 13481 13127 13515
rect 18521 13481 18555 13515
rect 19257 13481 19291 13515
rect 20545 13481 20579 13515
rect 20821 13481 20855 13515
rect 17417 13413 17451 13447
rect 9045 13345 9079 13379
rect 9229 13345 9263 13379
rect 10333 13345 10367 13379
rect 12541 13345 12575 13379
rect 17969 13345 18003 13379
rect 19809 13345 19843 13379
rect 7297 13277 7331 13311
rect 12081 13277 12115 13311
rect 19625 13277 19659 13311
rect 20361 13277 20395 13311
rect 21005 13277 21039 13311
rect 7030 13209 7064 13243
rect 12633 13209 12667 13243
rect 18153 13209 18187 13243
rect 18797 13209 18831 13243
rect 19717 13209 19751 13243
rect 21281 13209 21315 13243
rect 9321 13141 9355 13175
rect 9965 13141 9999 13175
rect 12725 13141 12759 13175
rect 13369 13141 13403 13175
rect 18061 13141 18095 13175
rect 6377 12937 6411 12971
rect 12081 12937 12115 12971
rect 19625 12937 19659 12971
rect 20545 12937 20579 12971
rect 20821 12937 20855 12971
rect 21373 12937 21407 12971
rect 13001 12869 13035 12903
rect 14749 12869 14783 12903
rect 17693 12869 17727 12903
rect 7021 12801 7055 12835
rect 11621 12801 11655 12835
rect 12725 12801 12759 12835
rect 17049 12801 17083 12835
rect 19165 12801 19199 12835
rect 19441 12801 19475 12835
rect 19901 12801 19935 12835
rect 20361 12801 20395 12835
rect 21005 12801 21039 12835
rect 17141 12733 17175 12767
rect 17233 12733 17267 12767
rect 11805 12665 11839 12699
rect 20085 12665 20119 12699
rect 16681 12597 16715 12631
rect 18429 12597 18463 12631
rect 9045 12393 9079 12427
rect 12909 12393 12943 12427
rect 14289 12393 14323 12427
rect 17049 12393 17083 12427
rect 17325 12393 17359 12427
rect 20545 12393 20579 12427
rect 21005 12393 21039 12427
rect 7941 12257 7975 12291
rect 8125 12257 8159 12291
rect 16405 12257 16439 12291
rect 17877 12257 17911 12291
rect 9413 12189 9447 12223
rect 9669 12189 9703 12223
rect 11529 12189 11563 12223
rect 14105 12189 14139 12223
rect 16037 12189 16071 12223
rect 16589 12189 16623 12223
rect 16681 12189 16715 12223
rect 19901 12189 19935 12223
rect 20361 12189 20395 12223
rect 20821 12189 20855 12223
rect 8217 12121 8251 12155
rect 11774 12121 11808 12155
rect 15792 12121 15826 12155
rect 17785 12121 17819 12155
rect 8585 12053 8619 12087
rect 10793 12053 10827 12087
rect 11069 12053 11103 12087
rect 14657 12053 14691 12087
rect 17693 12053 17727 12087
rect 18337 12053 18371 12087
rect 18889 12053 18923 12087
rect 19625 12053 19659 12087
rect 20085 12053 20119 12087
rect 21373 12053 21407 12087
rect 8677 11849 8711 11883
rect 8769 11849 8803 11883
rect 9413 11849 9447 11883
rect 9781 11849 9815 11883
rect 11161 11849 11195 11883
rect 11529 11849 11563 11883
rect 16957 11849 16991 11883
rect 17049 11849 17083 11883
rect 17693 11849 17727 11883
rect 18061 11849 18095 11883
rect 18153 11849 18187 11883
rect 18705 11849 18739 11883
rect 19073 11849 19107 11883
rect 19717 11849 19751 11883
rect 20361 11849 20395 11883
rect 20821 11849 20855 11883
rect 9873 11781 9907 11815
rect 14320 11781 14354 11815
rect 14841 11781 14875 11815
rect 10517 11713 10551 11747
rect 11897 11713 11931 11747
rect 15485 11713 15519 11747
rect 19165 11713 19199 11747
rect 19901 11713 19935 11747
rect 20545 11713 20579 11747
rect 21005 11713 21039 11747
rect 8585 11645 8619 11679
rect 9965 11645 9999 11679
rect 11989 11645 12023 11679
rect 12081 11645 12115 11679
rect 14565 11645 14599 11679
rect 16773 11645 16807 11679
rect 18245 11645 18279 11679
rect 19257 11645 19291 11679
rect 9137 11577 9171 11611
rect 17417 11577 17451 11611
rect 13185 11509 13219 11543
rect 21281 11509 21315 11543
rect 10333 11305 10367 11339
rect 11345 11305 11379 11339
rect 12633 11305 12667 11339
rect 19441 11305 19475 11339
rect 20545 11305 20579 11339
rect 20821 11305 20855 11339
rect 12357 11237 12391 11271
rect 13737 11237 13771 11271
rect 14841 11237 14875 11271
rect 20085 11237 20119 11271
rect 10701 11169 10735 11203
rect 13185 11169 13219 11203
rect 14289 11169 14323 11203
rect 14381 11169 14415 11203
rect 8953 11101 8987 11135
rect 9209 11101 9243 11135
rect 10885 11101 10919 11135
rect 13277 11101 13311 11135
rect 19257 11101 19291 11135
rect 19901 11101 19935 11135
rect 20361 11101 20395 11135
rect 21005 11101 21039 11135
rect 10977 11033 11011 11067
rect 11621 11033 11655 11067
rect 13369 11033 13403 11067
rect 14473 11033 14507 11067
rect 15209 11033 15243 11067
rect 21373 11033 21407 11067
rect 10241 10761 10275 10795
rect 11529 10761 11563 10795
rect 11897 10761 11931 10795
rect 12541 10761 12575 10795
rect 15025 10761 15059 10795
rect 15485 10761 15519 10795
rect 16681 10761 16715 10795
rect 19349 10761 19383 10795
rect 20913 10761 20947 10795
rect 21189 10761 21223 10795
rect 9597 10693 9631 10727
rect 13001 10693 13035 10727
rect 17794 10693 17828 10727
rect 11989 10625 12023 10659
rect 15393 10625 15427 10659
rect 18613 10625 18647 10659
rect 18889 10625 18923 10659
rect 19717 10625 19751 10659
rect 20361 10625 20395 10659
rect 21373 10625 21407 10659
rect 12081 10557 12115 10591
rect 15577 10557 15611 10591
rect 18061 10557 18095 10591
rect 19809 10557 19843 10591
rect 19993 10557 20027 10591
rect 8309 10421 8343 10455
rect 14289 10421 14323 10455
rect 19073 10421 19107 10455
rect 10149 10217 10183 10251
rect 15761 10217 15795 10251
rect 17141 10217 17175 10251
rect 19533 10217 19567 10251
rect 11529 10081 11563 10115
rect 16313 10081 16347 10115
rect 20085 10081 20119 10115
rect 13185 10013 13219 10047
rect 14105 10013 14139 10047
rect 18521 10013 18555 10047
rect 19901 10013 19935 10047
rect 20545 10013 20579 10047
rect 11284 9945 11318 9979
rect 12940 9945 12974 9979
rect 14350 9945 14384 9979
rect 18276 9945 18310 9979
rect 21189 9945 21223 9979
rect 11805 9877 11839 9911
rect 15485 9877 15519 9911
rect 16129 9877 16163 9911
rect 16221 9877 16255 9911
rect 16865 9877 16899 9911
rect 18797 9877 18831 9911
rect 19993 9877 20027 9911
rect 11897 9673 11931 9707
rect 15485 9673 15519 9707
rect 20177 9673 20211 9707
rect 21373 9673 21407 9707
rect 14105 9605 14139 9639
rect 14841 9605 14875 9639
rect 12541 9537 12575 9571
rect 16221 9537 16255 9571
rect 19064 9537 19098 9571
rect 21005 9537 21039 9571
rect 13829 9469 13863 9503
rect 14013 9469 14047 9503
rect 18797 9469 18831 9503
rect 14473 9401 14507 9435
rect 16037 9401 16071 9435
rect 20821 9401 20855 9435
rect 20545 9333 20579 9367
rect 11805 9129 11839 9163
rect 13461 9129 13495 9163
rect 16313 9129 16347 9163
rect 19625 9129 19659 9163
rect 21005 9129 21039 9163
rect 11621 8925 11655 8959
rect 13277 8925 13311 8959
rect 16497 8925 16531 8959
rect 20269 8925 20303 8959
rect 20545 8925 20579 8959
rect 21189 8925 21223 8959
rect 14841 8789 14875 8823
rect 17417 8789 17451 8823
rect 20729 8789 20763 8823
rect 11161 8585 11195 8619
rect 13461 8585 13495 8619
rect 19625 8585 19659 8619
rect 20085 8585 20119 8619
rect 20821 8585 20855 8619
rect 21373 8585 21407 8619
rect 9413 8449 9447 8483
rect 10977 8449 11011 8483
rect 11529 8449 11563 8483
rect 13645 8449 13679 8483
rect 15485 8449 15519 8483
rect 17141 8449 17175 8483
rect 18512 8449 18546 8483
rect 19901 8449 19935 8483
rect 20545 8449 20579 8483
rect 21005 8449 21039 8483
rect 12449 8381 12483 8415
rect 14473 8381 14507 8415
rect 18245 8381 18279 8415
rect 20361 8313 20395 8347
rect 10057 8245 10091 8279
rect 12173 8245 12207 8279
rect 16129 8245 16163 8279
rect 17785 8245 17819 8279
rect 19901 8041 19935 8075
rect 20821 7973 20855 8007
rect 21373 7905 21407 7939
rect 9781 7837 9815 7871
rect 10048 7837 10082 7871
rect 11713 7837 11747 7871
rect 14105 7837 14139 7871
rect 15761 7837 15795 7871
rect 17417 7837 17451 7871
rect 19257 7837 19291 7871
rect 20177 7837 20211 7871
rect 21005 7837 21039 7871
rect 11980 7769 12014 7803
rect 14350 7769 14384 7803
rect 16028 7769 16062 7803
rect 17684 7769 17718 7803
rect 11161 7701 11195 7735
rect 13093 7701 13127 7735
rect 15485 7701 15519 7735
rect 17141 7701 17175 7735
rect 18797 7701 18831 7735
rect 20361 7701 20395 7735
rect 9413 7497 9447 7531
rect 11529 7497 11563 7531
rect 11897 7497 11931 7531
rect 13737 7497 13771 7531
rect 14013 7497 14047 7531
rect 14381 7497 14415 7531
rect 15485 7497 15519 7531
rect 16957 7497 16991 7531
rect 17325 7497 17359 7531
rect 17417 7497 17451 7531
rect 17969 7497 18003 7531
rect 18337 7497 18371 7531
rect 20085 7497 20119 7531
rect 21189 7497 21223 7531
rect 20913 7429 20947 7463
rect 8033 7361 8067 7395
rect 8300 7361 8334 7395
rect 13093 7361 13127 7395
rect 15393 7361 15427 7395
rect 19625 7361 19659 7395
rect 19901 7361 19935 7395
rect 20545 7361 20579 7395
rect 21373 7361 21407 7395
rect 11989 7293 12023 7327
rect 12081 7293 12115 7327
rect 14473 7293 14507 7327
rect 14657 7293 14691 7327
rect 15577 7293 15611 7327
rect 17601 7293 17635 7327
rect 18429 7293 18463 7327
rect 18521 7293 18555 7327
rect 15025 7225 15059 7259
rect 20361 7157 20395 7191
rect 11897 6953 11931 6987
rect 21373 6953 21407 6987
rect 20361 6885 20395 6919
rect 11253 6817 11287 6851
rect 14841 6749 14875 6783
rect 17785 6749 17819 6783
rect 20545 6749 20579 6783
rect 21005 6749 21039 6783
rect 10793 6613 10827 6647
rect 11437 6613 11471 6647
rect 11529 6613 11563 6647
rect 20821 6613 20855 6647
rect 1593 6409 1627 6443
rect 20453 6409 20487 6443
rect 21189 6409 21223 6443
rect 1409 6273 1443 6307
rect 1869 6273 1903 6307
rect 19993 6273 20027 6307
rect 20269 6273 20303 6307
rect 20913 6273 20947 6307
rect 21373 6273 21407 6307
rect 19625 6205 19659 6239
rect 20729 6137 20763 6171
rect 20821 5797 20855 5831
rect 20085 5661 20119 5695
rect 20361 5661 20395 5695
rect 21005 5593 21039 5627
rect 20545 5525 20579 5559
rect 20729 5321 20763 5355
rect 21189 5321 21223 5355
rect 20453 5253 20487 5287
rect 20913 5185 20947 5219
rect 21373 5185 21407 5219
rect 20269 4777 20303 4811
rect 20913 4777 20947 4811
rect 21189 4777 21223 4811
rect 20453 4573 20487 4607
rect 20729 4573 20763 4607
rect 21373 4573 21407 4607
rect 19993 4505 20027 4539
rect 20545 4233 20579 4267
rect 21189 4233 21223 4267
rect 21281 4165 21315 4199
rect 19901 4097 19935 4131
rect 20269 4097 20303 4131
rect 19993 3621 20027 3655
rect 20821 3553 20855 3587
rect 19349 3485 19383 3519
rect 20545 3485 20579 3519
rect 19717 3417 19751 3451
rect 20177 3417 20211 3451
rect 20085 3145 20119 3179
rect 18981 3077 19015 3111
rect 20729 3077 20763 3111
rect 19349 3009 19383 3043
rect 20177 3009 20211 3043
rect 21281 3009 21315 3043
rect 18613 2941 18647 2975
rect 20545 2873 20579 2907
rect 19625 2805 19659 2839
rect 21189 2805 21223 2839
rect 19993 2533 20027 2567
rect 18521 2465 18555 2499
rect 20821 2465 20855 2499
rect 19441 2397 19475 2431
rect 20545 2397 20579 2431
rect 19625 2329 19659 2363
rect 20177 2329 20211 2363
rect 18889 2261 18923 2295
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21896 20698
rect 1104 20624 21896 20646
rect 3234 20544 3240 20596
rect 3292 20584 3298 20596
rect 4430 20584 4436 20596
rect 3292 20556 4436 20584
rect 3292 20544 3298 20556
rect 4430 20544 4436 20556
rect 4488 20544 4494 20596
rect 4525 20587 4583 20593
rect 4525 20553 4537 20587
rect 4571 20584 4583 20587
rect 11149 20587 11207 20593
rect 4571 20556 11100 20584
rect 4571 20553 4583 20556
rect 4525 20547 4583 20553
rect 290 20476 296 20528
rect 348 20516 354 20528
rect 1673 20519 1731 20525
rect 1673 20516 1685 20519
rect 348 20488 1685 20516
rect 348 20476 354 20488
rect 1673 20485 1685 20488
rect 1719 20516 1731 20519
rect 2406 20516 2412 20528
rect 1719 20488 2412 20516
rect 1719 20485 1731 20488
rect 1673 20479 1731 20485
rect 2406 20476 2412 20488
rect 2464 20476 2470 20528
rect 3142 20516 3148 20528
rect 2792 20488 3148 20516
rect 2317 20451 2375 20457
rect 2317 20417 2329 20451
rect 2363 20448 2375 20451
rect 2682 20448 2688 20460
rect 2363 20420 2688 20448
rect 2363 20417 2375 20420
rect 2317 20411 2375 20417
rect 2682 20408 2688 20420
rect 2740 20408 2746 20460
rect 2792 20457 2820 20488
rect 3142 20476 3148 20488
rect 3200 20516 3206 20528
rect 4062 20516 4068 20528
rect 3200 20488 4068 20516
rect 3200 20476 3206 20488
rect 4062 20476 4068 20488
rect 4120 20476 4126 20528
rect 5718 20516 5724 20528
rect 4356 20488 5724 20516
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20417 2835 20451
rect 3234 20448 3240 20460
rect 3195 20420 3240 20448
rect 2777 20411 2835 20417
rect 3234 20408 3240 20420
rect 3292 20408 3298 20460
rect 4356 20457 4384 20488
rect 5718 20476 5724 20488
rect 5776 20476 5782 20528
rect 8110 20516 8116 20528
rect 7024 20488 8116 20516
rect 3881 20451 3939 20457
rect 3881 20417 3893 20451
rect 3927 20417 3939 20451
rect 3881 20411 3939 20417
rect 4341 20451 4399 20457
rect 4341 20417 4353 20451
rect 4387 20417 4399 20451
rect 4341 20411 4399 20417
rect 1857 20383 1915 20389
rect 1857 20349 1869 20383
rect 1903 20380 1915 20383
rect 3786 20380 3792 20392
rect 1903 20352 3792 20380
rect 1903 20349 1915 20352
rect 1857 20343 1915 20349
rect 3786 20340 3792 20352
rect 3844 20340 3850 20392
rect 3896 20380 3924 20411
rect 5350 20408 5356 20460
rect 5408 20448 5414 20460
rect 5445 20451 5503 20457
rect 5445 20448 5457 20451
rect 5408 20420 5457 20448
rect 5408 20408 5414 20420
rect 5445 20417 5457 20420
rect 5491 20417 5503 20451
rect 5445 20411 5503 20417
rect 5813 20451 5871 20457
rect 5813 20417 5825 20451
rect 5859 20417 5871 20451
rect 5813 20411 5871 20417
rect 4246 20380 4252 20392
rect 3896 20352 4252 20380
rect 4246 20340 4252 20352
rect 4304 20380 4310 20392
rect 5258 20380 5264 20392
rect 4304 20352 5264 20380
rect 4304 20340 4310 20352
rect 5258 20340 5264 20352
rect 5316 20340 5322 20392
rect 5828 20380 5856 20411
rect 6454 20408 6460 20460
rect 6512 20448 6518 20460
rect 7024 20457 7052 20488
rect 8110 20476 8116 20488
rect 8168 20476 8174 20528
rect 9033 20519 9091 20525
rect 9033 20485 9045 20519
rect 9079 20516 9091 20519
rect 9079 20488 10916 20516
rect 9079 20485 9091 20488
rect 9033 20479 9091 20485
rect 10888 20460 10916 20488
rect 6549 20451 6607 20457
rect 6549 20448 6561 20451
rect 6512 20420 6561 20448
rect 6512 20408 6518 20420
rect 6549 20417 6561 20420
rect 6595 20417 6607 20451
rect 6549 20411 6607 20417
rect 7009 20451 7067 20457
rect 7009 20417 7021 20451
rect 7055 20417 7067 20451
rect 7009 20411 7067 20417
rect 7469 20451 7527 20457
rect 7469 20417 7481 20451
rect 7515 20417 7527 20451
rect 7926 20448 7932 20460
rect 7887 20420 7932 20448
rect 7469 20411 7527 20417
rect 6822 20380 6828 20392
rect 5828 20352 6828 20380
rect 6822 20340 6828 20352
rect 6880 20340 6886 20392
rect 7484 20380 7512 20411
rect 7926 20408 7932 20420
rect 7984 20408 7990 20460
rect 9214 20408 9220 20460
rect 9272 20448 9278 20460
rect 9309 20451 9367 20457
rect 9309 20448 9321 20451
rect 9272 20420 9321 20448
rect 9272 20408 9278 20420
rect 9309 20417 9321 20420
rect 9355 20417 9367 20451
rect 9309 20411 9367 20417
rect 9766 20408 9772 20460
rect 9824 20448 9830 20460
rect 9861 20451 9919 20457
rect 9861 20448 9873 20451
rect 9824 20420 9873 20448
rect 9824 20408 9830 20420
rect 9861 20417 9873 20420
rect 9907 20417 9919 20451
rect 9861 20411 9919 20417
rect 10318 20408 10324 20460
rect 10376 20448 10382 20460
rect 10413 20451 10471 20457
rect 10413 20448 10425 20451
rect 10376 20420 10425 20448
rect 10376 20408 10382 20420
rect 10413 20417 10425 20420
rect 10459 20417 10471 20451
rect 10413 20411 10471 20417
rect 10870 20408 10876 20460
rect 10928 20448 10934 20460
rect 10965 20451 11023 20457
rect 10965 20448 10977 20451
rect 10928 20420 10977 20448
rect 10928 20408 10934 20420
rect 10965 20417 10977 20420
rect 11011 20417 11023 20451
rect 10965 20411 11023 20417
rect 7834 20380 7840 20392
rect 7484 20352 7840 20380
rect 7834 20340 7840 20352
rect 7892 20380 7898 20392
rect 8202 20380 8208 20392
rect 7892 20352 8208 20380
rect 7892 20340 7898 20352
rect 8202 20340 8208 20352
rect 8260 20340 8266 20392
rect 11072 20380 11100 20556
rect 11149 20553 11161 20587
rect 11195 20553 11207 20587
rect 11149 20547 11207 20553
rect 11164 20516 11192 20547
rect 12618 20544 12624 20596
rect 12676 20584 12682 20596
rect 12989 20587 13047 20593
rect 12989 20584 13001 20587
rect 12676 20556 13001 20584
rect 12676 20544 12682 20556
rect 12989 20553 13001 20556
rect 13035 20553 13047 20587
rect 12989 20547 13047 20553
rect 13170 20544 13176 20596
rect 13228 20584 13234 20596
rect 13633 20587 13691 20593
rect 13633 20584 13645 20587
rect 13228 20556 13645 20584
rect 13228 20544 13234 20556
rect 13633 20553 13645 20556
rect 13679 20553 13691 20587
rect 13633 20547 13691 20553
rect 14274 20544 14280 20596
rect 14332 20584 14338 20596
rect 15565 20587 15623 20593
rect 15565 20584 15577 20587
rect 14332 20556 15577 20584
rect 14332 20544 14338 20556
rect 15565 20553 15577 20556
rect 15611 20553 15623 20587
rect 15565 20547 15623 20553
rect 15746 20544 15752 20596
rect 15804 20584 15810 20596
rect 16761 20587 16819 20593
rect 16761 20584 16773 20587
rect 15804 20556 16773 20584
rect 15804 20544 15810 20556
rect 16761 20553 16773 20556
rect 16807 20553 16819 20587
rect 16761 20547 16819 20553
rect 17313 20587 17371 20593
rect 17313 20553 17325 20587
rect 17359 20553 17371 20587
rect 17313 20547 17371 20553
rect 12894 20516 12900 20528
rect 11164 20488 12900 20516
rect 12894 20476 12900 20488
rect 12952 20476 12958 20528
rect 13814 20516 13820 20528
rect 13188 20488 13820 20516
rect 11238 20408 11244 20460
rect 11296 20448 11302 20460
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 11296 20420 11529 20448
rect 11296 20408 11302 20420
rect 11517 20417 11529 20420
rect 11563 20417 11575 20451
rect 11517 20411 11575 20417
rect 12066 20408 12072 20460
rect 12124 20448 12130 20460
rect 13188 20457 13216 20488
rect 13814 20476 13820 20488
rect 13872 20476 13878 20528
rect 16022 20476 16028 20528
rect 16080 20516 16086 20528
rect 17328 20516 17356 20547
rect 17678 20544 17684 20596
rect 17736 20584 17742 20596
rect 19337 20587 19395 20593
rect 19337 20584 19349 20587
rect 17736 20556 19349 20584
rect 17736 20544 17742 20556
rect 19337 20553 19349 20556
rect 19383 20553 19395 20587
rect 19337 20547 19395 20553
rect 19886 20544 19892 20596
rect 19944 20584 19950 20596
rect 20533 20587 20591 20593
rect 20533 20584 20545 20587
rect 19944 20556 20545 20584
rect 19944 20544 19950 20556
rect 20533 20553 20545 20556
rect 20579 20553 20591 20587
rect 20533 20547 20591 20553
rect 20714 20544 20720 20596
rect 20772 20584 20778 20596
rect 21085 20587 21143 20593
rect 21085 20584 21097 20587
rect 20772 20556 21097 20584
rect 20772 20544 20778 20556
rect 21085 20553 21097 20556
rect 21131 20553 21143 20587
rect 21085 20547 21143 20553
rect 16080 20488 17356 20516
rect 16080 20476 16086 20488
rect 12621 20451 12679 20457
rect 12621 20448 12633 20451
rect 12124 20420 12633 20448
rect 12124 20408 12130 20420
rect 12621 20417 12633 20420
rect 12667 20417 12679 20451
rect 12621 20411 12679 20417
rect 13173 20451 13231 20457
rect 13173 20417 13185 20451
rect 13219 20417 13231 20451
rect 13446 20448 13452 20460
rect 13407 20420 13452 20448
rect 13173 20411 13231 20417
rect 13446 20408 13452 20420
rect 13504 20408 13510 20460
rect 14829 20451 14887 20457
rect 14829 20417 14841 20451
rect 14875 20448 14887 20451
rect 14918 20448 14924 20460
rect 14875 20420 14924 20448
rect 14875 20417 14887 20420
rect 14829 20411 14887 20417
rect 14918 20408 14924 20420
rect 14976 20408 14982 20460
rect 15749 20451 15807 20457
rect 15749 20417 15761 20451
rect 15795 20448 15807 20451
rect 15930 20448 15936 20460
rect 15795 20420 15936 20448
rect 15795 20417 15807 20420
rect 15749 20411 15807 20417
rect 15930 20408 15936 20420
rect 15988 20408 15994 20460
rect 16298 20448 16304 20460
rect 16259 20420 16304 20448
rect 16298 20408 16304 20420
rect 16356 20408 16362 20460
rect 16945 20451 17003 20457
rect 16945 20417 16957 20451
rect 16991 20417 17003 20451
rect 17494 20448 17500 20460
rect 17455 20420 17500 20448
rect 16945 20411 17003 20417
rect 14274 20380 14280 20392
rect 11072 20352 14280 20380
rect 14274 20340 14280 20352
rect 14332 20340 14338 20392
rect 14642 20380 14648 20392
rect 14603 20352 14648 20380
rect 14642 20340 14648 20352
rect 14700 20340 14706 20392
rect 14737 20383 14795 20389
rect 14737 20349 14749 20383
rect 14783 20349 14795 20383
rect 16960 20380 16988 20411
rect 17494 20408 17500 20420
rect 17552 20408 17558 20460
rect 18049 20451 18107 20457
rect 18049 20417 18061 20451
rect 18095 20417 18107 20451
rect 18598 20448 18604 20460
rect 18559 20420 18604 20448
rect 18049 20411 18107 20417
rect 17586 20380 17592 20392
rect 16960 20352 17592 20380
rect 14737 20343 14795 20349
rect 1670 20272 1676 20324
rect 1728 20312 1734 20324
rect 6733 20315 6791 20321
rect 1728 20284 6132 20312
rect 1728 20272 1734 20284
rect 2498 20244 2504 20256
rect 2459 20216 2504 20244
rect 2498 20204 2504 20216
rect 2556 20204 2562 20256
rect 2958 20244 2964 20256
rect 2919 20216 2964 20244
rect 2958 20204 2964 20216
rect 3016 20204 3022 20256
rect 3326 20204 3332 20256
rect 3384 20244 3390 20256
rect 3421 20247 3479 20253
rect 3421 20244 3433 20247
rect 3384 20216 3433 20244
rect 3384 20204 3390 20216
rect 3421 20213 3433 20216
rect 3467 20213 3479 20247
rect 4062 20244 4068 20256
rect 4023 20216 4068 20244
rect 3421 20207 3479 20213
rect 4062 20204 4068 20216
rect 4120 20204 4126 20256
rect 4798 20244 4804 20256
rect 4759 20216 4804 20244
rect 4798 20204 4804 20216
rect 4856 20204 4862 20256
rect 5994 20244 6000 20256
rect 5955 20216 6000 20244
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 6104 20244 6132 20284
rect 6733 20281 6745 20315
rect 6779 20312 6791 20315
rect 10597 20315 10655 20321
rect 6779 20284 8248 20312
rect 6779 20281 6791 20284
rect 6733 20275 6791 20281
rect 8220 20256 8248 20284
rect 10597 20281 10609 20315
rect 10643 20312 10655 20315
rect 14752 20312 14780 20343
rect 17586 20340 17592 20352
rect 17644 20340 17650 20392
rect 18064 20380 18092 20411
rect 18598 20408 18604 20420
rect 18656 20408 18662 20460
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20417 19579 20451
rect 19521 20411 19579 20417
rect 20073 20451 20131 20457
rect 20073 20417 20085 20451
rect 20119 20417 20131 20451
rect 20073 20411 20131 20417
rect 18506 20380 18512 20392
rect 18064 20352 18512 20380
rect 18506 20340 18512 20352
rect 18564 20340 18570 20392
rect 10643 20284 14780 20312
rect 15197 20315 15255 20321
rect 10643 20281 10655 20284
rect 10597 20275 10655 20281
rect 15197 20281 15209 20315
rect 15243 20312 15255 20315
rect 16850 20312 16856 20324
rect 15243 20284 16856 20312
rect 15243 20281 15255 20284
rect 15197 20275 15255 20281
rect 16850 20272 16856 20284
rect 16908 20272 16914 20324
rect 17034 20272 17040 20324
rect 17092 20312 17098 20324
rect 18417 20315 18475 20321
rect 18417 20312 18429 20315
rect 17092 20284 18429 20312
rect 17092 20272 17098 20284
rect 18417 20281 18429 20284
rect 18463 20281 18475 20315
rect 19536 20312 19564 20411
rect 20088 20380 20116 20411
rect 20254 20408 20260 20460
rect 20312 20448 20318 20460
rect 20349 20451 20407 20457
rect 20349 20448 20361 20451
rect 20312 20420 20361 20448
rect 20312 20408 20318 20420
rect 20349 20417 20361 20420
rect 20395 20417 20407 20451
rect 20349 20411 20407 20417
rect 20901 20451 20959 20457
rect 20901 20417 20913 20451
rect 20947 20448 20959 20451
rect 21634 20448 21640 20460
rect 20947 20420 21640 20448
rect 20947 20417 20959 20420
rect 20901 20411 20959 20417
rect 21634 20408 21640 20420
rect 21692 20408 21698 20460
rect 21726 20380 21732 20392
rect 20088 20352 21732 20380
rect 21726 20340 21732 20352
rect 21784 20340 21790 20392
rect 21818 20312 21824 20324
rect 19536 20284 21824 20312
rect 18417 20275 18475 20281
rect 21818 20272 21824 20284
rect 21876 20272 21882 20324
rect 6822 20244 6828 20256
rect 6104 20216 6828 20244
rect 6822 20204 6828 20216
rect 6880 20204 6886 20256
rect 7193 20247 7251 20253
rect 7193 20213 7205 20247
rect 7239 20244 7251 20247
rect 7374 20244 7380 20256
rect 7239 20216 7380 20244
rect 7239 20213 7251 20216
rect 7193 20207 7251 20213
rect 7374 20204 7380 20216
rect 7432 20204 7438 20256
rect 7650 20244 7656 20256
rect 7611 20216 7656 20244
rect 7650 20204 7656 20216
rect 7708 20204 7714 20256
rect 8202 20204 8208 20256
rect 8260 20204 8266 20256
rect 8386 20204 8392 20256
rect 8444 20244 8450 20256
rect 8573 20247 8631 20253
rect 8573 20244 8585 20247
rect 8444 20216 8585 20244
rect 8444 20204 8450 20216
rect 8573 20213 8585 20216
rect 8619 20213 8631 20247
rect 8573 20207 8631 20213
rect 9493 20247 9551 20253
rect 9493 20213 9505 20247
rect 9539 20244 9551 20247
rect 9674 20244 9680 20256
rect 9539 20216 9680 20244
rect 9539 20213 9551 20216
rect 9493 20207 9551 20213
rect 9674 20204 9680 20216
rect 9732 20204 9738 20256
rect 10045 20247 10103 20253
rect 10045 20213 10057 20247
rect 10091 20244 10103 20247
rect 11054 20244 11060 20256
rect 10091 20216 11060 20244
rect 10091 20213 10103 20216
rect 10045 20207 10103 20213
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 11698 20244 11704 20256
rect 11659 20216 11704 20244
rect 11698 20204 11704 20216
rect 11756 20204 11762 20256
rect 11974 20244 11980 20256
rect 11935 20216 11980 20244
rect 11974 20204 11980 20216
rect 12032 20204 12038 20256
rect 13814 20204 13820 20256
rect 13872 20244 13878 20256
rect 14185 20247 14243 20253
rect 14185 20244 14197 20247
rect 13872 20216 14197 20244
rect 13872 20204 13878 20216
rect 14185 20213 14197 20216
rect 14231 20244 14243 20247
rect 14734 20244 14740 20256
rect 14231 20216 14740 20244
rect 14231 20213 14243 20216
rect 14185 20207 14243 20213
rect 14734 20204 14740 20216
rect 14792 20204 14798 20256
rect 14826 20204 14832 20256
rect 14884 20244 14890 20256
rect 16117 20247 16175 20253
rect 16117 20244 16129 20247
rect 14884 20216 16129 20244
rect 14884 20204 14890 20216
rect 16117 20213 16129 20216
rect 16163 20213 16175 20247
rect 16117 20207 16175 20213
rect 16574 20204 16580 20256
rect 16632 20244 16638 20256
rect 17865 20247 17923 20253
rect 17865 20244 17877 20247
rect 16632 20216 17877 20244
rect 16632 20204 16638 20216
rect 17865 20213 17877 20216
rect 17911 20213 17923 20247
rect 17865 20207 17923 20213
rect 18230 20204 18236 20256
rect 18288 20244 18294 20256
rect 19889 20247 19947 20253
rect 19889 20244 19901 20247
rect 18288 20216 19901 20244
rect 18288 20204 18294 20216
rect 19889 20213 19901 20216
rect 19935 20213 19947 20247
rect 19889 20207 19947 20213
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 1670 20040 1676 20052
rect 1631 20012 1676 20040
rect 1670 20000 1676 20012
rect 1728 20000 1734 20052
rect 2777 20043 2835 20049
rect 2777 20009 2789 20043
rect 2823 20040 2835 20043
rect 2823 20012 6684 20040
rect 2823 20009 2835 20012
rect 2777 20003 2835 20009
rect 2958 19932 2964 19984
rect 3016 19972 3022 19984
rect 3016 19944 4292 19972
rect 3016 19932 3022 19944
rect 1394 19864 1400 19916
rect 1452 19904 1458 19916
rect 1452 19876 1992 19904
rect 1452 19864 1458 19876
rect 1486 19836 1492 19848
rect 1447 19808 1492 19836
rect 1486 19796 1492 19808
rect 1544 19796 1550 19848
rect 1964 19845 1992 19876
rect 3326 19864 3332 19916
rect 3384 19904 3390 19916
rect 4154 19904 4160 19916
rect 3384 19876 4016 19904
rect 4115 19876 4160 19904
rect 3384 19864 3390 19876
rect 1949 19839 2007 19845
rect 1949 19805 1961 19839
rect 1995 19836 2007 19839
rect 2038 19836 2044 19848
rect 1995 19808 2044 19836
rect 1995 19805 2007 19808
rect 1949 19799 2007 19805
rect 2038 19796 2044 19808
rect 2096 19796 2102 19848
rect 2590 19836 2596 19848
rect 2551 19808 2596 19836
rect 2590 19796 2596 19808
rect 2648 19796 2654 19848
rect 3237 19839 3295 19845
rect 3237 19805 3249 19839
rect 3283 19836 3295 19839
rect 3418 19836 3424 19848
rect 3283 19808 3424 19836
rect 3283 19805 3295 19808
rect 3237 19799 3295 19805
rect 3418 19796 3424 19808
rect 3476 19796 3482 19848
rect 3988 19768 4016 19876
rect 4154 19864 4160 19876
rect 4212 19864 4218 19916
rect 4264 19913 4292 19944
rect 4249 19907 4307 19913
rect 4249 19873 4261 19907
rect 4295 19873 4307 19907
rect 6656 19904 6684 20012
rect 6822 20000 6828 20052
rect 6880 20040 6886 20052
rect 7742 20040 7748 20052
rect 6880 20012 7748 20040
rect 6880 20000 6886 20012
rect 7742 20000 7748 20012
rect 7800 20000 7806 20052
rect 10321 20043 10379 20049
rect 10321 20009 10333 20043
rect 10367 20040 10379 20043
rect 11238 20040 11244 20052
rect 10367 20012 11244 20040
rect 10367 20009 10379 20012
rect 10321 20003 10379 20009
rect 11238 20000 11244 20012
rect 11296 20000 11302 20052
rect 11977 20043 12035 20049
rect 11977 20009 11989 20043
rect 12023 20040 12035 20043
rect 12066 20040 12072 20052
rect 12023 20012 12072 20040
rect 12023 20009 12035 20012
rect 11977 20003 12035 20009
rect 12066 20000 12072 20012
rect 12124 20000 12130 20052
rect 12434 20000 12440 20052
rect 12492 20040 12498 20052
rect 12492 20012 12537 20040
rect 12492 20000 12498 20012
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 14185 20043 14243 20049
rect 14185 20040 14197 20043
rect 13872 20012 14197 20040
rect 13872 20000 13878 20012
rect 14185 20009 14197 20012
rect 14231 20009 14243 20043
rect 14185 20003 14243 20009
rect 18782 20000 18788 20052
rect 18840 20040 18846 20052
rect 19337 20043 19395 20049
rect 19337 20040 19349 20043
rect 18840 20012 19349 20040
rect 18840 20000 18846 20012
rect 19337 20009 19349 20012
rect 19383 20009 19395 20043
rect 19337 20003 19395 20009
rect 19518 20000 19524 20052
rect 19576 20040 19582 20052
rect 19889 20043 19947 20049
rect 19889 20040 19901 20043
rect 19576 20012 19901 20040
rect 19576 20000 19582 20012
rect 19889 20009 19901 20012
rect 19935 20009 19947 20043
rect 19889 20003 19947 20009
rect 7926 19932 7932 19984
rect 7984 19972 7990 19984
rect 8021 19975 8079 19981
rect 8021 19972 8033 19975
rect 7984 19944 8033 19972
rect 7984 19932 7990 19944
rect 8021 19941 8033 19944
rect 8067 19941 8079 19975
rect 8021 19935 8079 19941
rect 16117 19975 16175 19981
rect 16117 19941 16129 19975
rect 16163 19972 16175 19975
rect 16163 19944 16988 19972
rect 16163 19941 16175 19944
rect 16117 19935 16175 19941
rect 8036 19904 8064 19935
rect 9033 19907 9091 19913
rect 9033 19904 9045 19907
rect 6656 19876 6776 19904
rect 8036 19876 9045 19904
rect 4249 19867 4307 19873
rect 4985 19839 5043 19845
rect 4985 19805 4997 19839
rect 5031 19836 5043 19839
rect 6638 19836 6644 19848
rect 5031 19808 6644 19836
rect 5031 19805 5043 19808
rect 4985 19799 5043 19805
rect 6638 19796 6644 19808
rect 6696 19796 6702 19848
rect 6748 19836 6776 19876
rect 9033 19873 9045 19876
rect 9079 19873 9091 19907
rect 9033 19867 9091 19873
rect 12894 19864 12900 19916
rect 12952 19904 12958 19916
rect 16850 19904 16856 19916
rect 12952 19876 14872 19904
rect 16811 19876 16856 19904
rect 12952 19864 12958 19876
rect 9122 19836 9128 19848
rect 6748 19808 9128 19836
rect 9122 19796 9128 19808
rect 9180 19796 9186 19848
rect 10594 19836 10600 19848
rect 10555 19808 10600 19836
rect 10594 19796 10600 19808
rect 10652 19796 10658 19848
rect 12250 19836 12256 19848
rect 12211 19808 12256 19836
rect 12250 19796 12256 19808
rect 12308 19796 12314 19848
rect 13078 19836 13084 19848
rect 13039 19808 13084 19836
rect 13078 19796 13084 19808
rect 13136 19796 13142 19848
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19836 14427 19839
rect 14550 19836 14556 19848
rect 14415 19808 14556 19836
rect 14415 19805 14427 19808
rect 14369 19799 14427 19805
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 14734 19836 14740 19848
rect 14695 19808 14740 19836
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 14844 19836 14872 19876
rect 16850 19864 16856 19876
rect 16908 19864 16914 19916
rect 16960 19913 16988 19944
rect 16945 19907 17003 19913
rect 16945 19873 16957 19907
rect 16991 19904 17003 19907
rect 17310 19904 17316 19916
rect 16991 19876 17316 19904
rect 16991 19873 17003 19876
rect 16945 19867 17003 19873
rect 17310 19864 17316 19876
rect 17368 19864 17374 19916
rect 21910 19904 21916 19916
rect 20088 19876 21916 19904
rect 16390 19836 16396 19848
rect 14844 19808 16396 19836
rect 16390 19796 16396 19808
rect 16448 19796 16454 19848
rect 18874 19836 18880 19848
rect 18835 19808 18880 19836
rect 18874 19796 18880 19808
rect 18932 19796 18938 19848
rect 19521 19839 19579 19845
rect 19521 19805 19533 19839
rect 19567 19836 19579 19839
rect 19886 19836 19892 19848
rect 19567 19808 19892 19836
rect 19567 19805 19579 19808
rect 19521 19799 19579 19805
rect 19886 19796 19892 19808
rect 19944 19796 19950 19848
rect 20088 19845 20116 19876
rect 21910 19864 21916 19876
rect 21968 19864 21974 19916
rect 20073 19839 20131 19845
rect 20073 19805 20085 19839
rect 20119 19805 20131 19839
rect 20073 19799 20131 19805
rect 20346 19796 20352 19848
rect 20404 19836 20410 19848
rect 20533 19839 20591 19845
rect 20533 19836 20545 19839
rect 20404 19808 20545 19836
rect 20404 19796 20410 19808
rect 20533 19805 20545 19808
rect 20579 19805 20591 19839
rect 21082 19836 21088 19848
rect 21043 19808 21088 19836
rect 20533 19799 20591 19805
rect 21082 19796 21088 19808
rect 21140 19796 21146 19848
rect 5258 19777 5264 19780
rect 3988 19740 5212 19768
rect 2130 19700 2136 19712
rect 2091 19672 2136 19700
rect 2130 19660 2136 19672
rect 2188 19660 2194 19712
rect 3326 19660 3332 19712
rect 3384 19700 3390 19712
rect 3421 19703 3479 19709
rect 3421 19700 3433 19703
rect 3384 19672 3433 19700
rect 3384 19660 3390 19672
rect 3421 19669 3433 19672
rect 3467 19669 3479 19703
rect 4338 19700 4344 19712
rect 4299 19672 4344 19700
rect 3421 19663 3479 19669
rect 4338 19660 4344 19672
rect 4396 19660 4402 19712
rect 4706 19700 4712 19712
rect 4667 19672 4712 19700
rect 4706 19660 4712 19672
rect 4764 19660 4770 19712
rect 5184 19700 5212 19740
rect 5252 19731 5264 19777
rect 5316 19768 5322 19780
rect 5316 19740 5352 19768
rect 5258 19728 5264 19731
rect 5316 19728 5322 19740
rect 6454 19728 6460 19780
rect 6512 19768 6518 19780
rect 6730 19768 6736 19780
rect 6512 19740 6736 19768
rect 6512 19728 6518 19740
rect 6730 19728 6736 19740
rect 6788 19728 6794 19780
rect 6908 19771 6966 19777
rect 6908 19737 6920 19771
rect 6954 19768 6966 19771
rect 7006 19768 7012 19780
rect 6954 19740 7012 19768
rect 6954 19737 6966 19740
rect 6908 19731 6966 19737
rect 7006 19728 7012 19740
rect 7064 19728 7070 19780
rect 8573 19771 8631 19777
rect 8573 19737 8585 19771
rect 8619 19768 8631 19771
rect 9309 19771 9367 19777
rect 9309 19768 9321 19771
rect 8619 19740 9321 19768
rect 8619 19737 8631 19740
rect 8573 19731 8631 19737
rect 9309 19737 9321 19740
rect 9355 19737 9367 19771
rect 9309 19731 9367 19737
rect 10864 19771 10922 19777
rect 10864 19737 10876 19771
rect 10910 19768 10922 19771
rect 12158 19768 12164 19780
rect 10910 19740 12164 19768
rect 10910 19737 10922 19740
rect 10864 19731 10922 19737
rect 12158 19728 12164 19740
rect 12216 19728 12222 19780
rect 15004 19771 15062 19777
rect 15004 19737 15016 19771
rect 15050 19768 15062 19771
rect 15562 19768 15568 19780
rect 15050 19740 15568 19768
rect 15050 19737 15062 19740
rect 15004 19731 15062 19737
rect 15562 19728 15568 19740
rect 15620 19728 15626 19780
rect 16761 19771 16819 19777
rect 16761 19737 16773 19771
rect 16807 19768 16819 19771
rect 17405 19771 17463 19777
rect 17405 19768 17417 19771
rect 16807 19740 17417 19768
rect 16807 19737 16819 19740
rect 16761 19731 16819 19737
rect 17405 19737 17417 19740
rect 17451 19737 17463 19771
rect 18046 19768 18052 19780
rect 18007 19740 18052 19768
rect 17405 19731 17463 19737
rect 18046 19728 18052 19740
rect 18104 19728 18110 19780
rect 18414 19728 18420 19780
rect 18472 19768 18478 19780
rect 22646 19768 22652 19780
rect 18472 19740 22652 19768
rect 18472 19728 18478 19740
rect 22646 19728 22652 19740
rect 22704 19728 22710 19780
rect 5810 19700 5816 19712
rect 5184 19672 5816 19700
rect 5810 19660 5816 19672
rect 5868 19660 5874 19712
rect 6365 19703 6423 19709
rect 6365 19669 6377 19703
rect 6411 19700 6423 19703
rect 6546 19700 6552 19712
rect 6411 19672 6552 19700
rect 6411 19669 6423 19672
rect 6365 19663 6423 19669
rect 6546 19660 6552 19672
rect 6604 19660 6610 19712
rect 9030 19660 9036 19712
rect 9088 19700 9094 19712
rect 9217 19703 9275 19709
rect 9217 19700 9229 19703
rect 9088 19672 9229 19700
rect 9088 19660 9094 19672
rect 9217 19669 9229 19672
rect 9263 19669 9275 19703
rect 9217 19663 9275 19669
rect 9677 19703 9735 19709
rect 9677 19669 9689 19703
rect 9723 19700 9735 19703
rect 10962 19700 10968 19712
rect 9723 19672 10968 19700
rect 9723 19669 9735 19672
rect 9677 19663 9735 19669
rect 10962 19660 10968 19672
rect 11020 19660 11026 19712
rect 13630 19660 13636 19712
rect 13688 19700 13694 19712
rect 13725 19703 13783 19709
rect 13725 19700 13737 19703
rect 13688 19672 13737 19700
rect 13688 19660 13694 19672
rect 13725 19669 13737 19672
rect 13771 19669 13783 19703
rect 13725 19663 13783 19669
rect 15194 19660 15200 19712
rect 15252 19700 15258 19712
rect 16393 19703 16451 19709
rect 16393 19700 16405 19703
rect 15252 19672 16405 19700
rect 15252 19660 15258 19672
rect 16393 19669 16405 19672
rect 16439 19669 16451 19703
rect 20714 19700 20720 19712
rect 20675 19672 20720 19700
rect 16393 19663 16451 19669
rect 20714 19660 20720 19672
rect 20772 19660 20778 19712
rect 21266 19700 21272 19712
rect 21227 19672 21272 19700
rect 21266 19660 21272 19672
rect 21324 19660 21330 19712
rect 1104 19610 21896 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21896 19610
rect 1104 19536 21896 19558
rect 1765 19499 1823 19505
rect 1765 19465 1777 19499
rect 1811 19496 1823 19499
rect 2590 19496 2596 19508
rect 1811 19468 2596 19496
rect 1811 19465 1823 19468
rect 1765 19459 1823 19465
rect 2590 19456 2596 19468
rect 2648 19456 2654 19508
rect 3145 19499 3203 19505
rect 3145 19465 3157 19499
rect 3191 19496 3203 19499
rect 3418 19496 3424 19508
rect 3191 19468 3424 19496
rect 3191 19465 3203 19468
rect 3145 19459 3203 19465
rect 3418 19456 3424 19468
rect 3476 19456 3482 19508
rect 7006 19496 7012 19508
rect 6967 19468 7012 19496
rect 7006 19456 7012 19468
rect 7064 19456 7070 19508
rect 7558 19496 7564 19508
rect 7116 19468 7564 19496
rect 2777 19431 2835 19437
rect 2777 19397 2789 19431
rect 2823 19428 2835 19431
rect 3234 19428 3240 19440
rect 2823 19400 3240 19428
rect 2823 19397 2835 19400
rect 2777 19391 2835 19397
rect 3234 19388 3240 19400
rect 3292 19388 3298 19440
rect 6730 19388 6736 19440
rect 6788 19428 6794 19440
rect 7116 19428 7144 19468
rect 7558 19456 7564 19468
rect 7616 19456 7622 19508
rect 7650 19456 7656 19508
rect 7708 19496 7714 19508
rect 8573 19499 8631 19505
rect 8573 19496 8585 19499
rect 7708 19468 8585 19496
rect 7708 19456 7714 19468
rect 8573 19465 8585 19468
rect 8619 19465 8631 19499
rect 9030 19496 9036 19508
rect 8991 19468 9036 19496
rect 8573 19459 8631 19465
rect 9030 19456 9036 19468
rect 9088 19456 9094 19508
rect 9585 19499 9643 19505
rect 9585 19465 9597 19499
rect 9631 19496 9643 19499
rect 9674 19496 9680 19508
rect 9631 19468 9680 19496
rect 9631 19465 9643 19468
rect 9585 19459 9643 19465
rect 9674 19456 9680 19468
rect 9732 19456 9738 19508
rect 13078 19496 13084 19508
rect 13039 19468 13084 19496
rect 13078 19456 13084 19468
rect 13136 19456 13142 19508
rect 13814 19456 13820 19508
rect 13872 19496 13878 19508
rect 16117 19499 16175 19505
rect 13872 19468 15884 19496
rect 13872 19456 13878 19468
rect 14734 19428 14740 19440
rect 6788 19400 7144 19428
rect 7208 19400 8432 19428
rect 6788 19388 6794 19400
rect 1946 19320 1952 19372
rect 2004 19360 2010 19372
rect 2041 19363 2099 19369
rect 2041 19360 2053 19363
rect 2004 19332 2053 19360
rect 2004 19320 2010 19332
rect 2041 19329 2053 19332
rect 2087 19329 2099 19363
rect 3418 19360 3424 19372
rect 3379 19332 3424 19360
rect 2041 19323 2099 19329
rect 3418 19320 3424 19332
rect 3476 19320 3482 19372
rect 3688 19363 3746 19369
rect 3688 19329 3700 19363
rect 3734 19360 3746 19363
rect 3970 19360 3976 19372
rect 3734 19332 3976 19360
rect 3734 19329 3746 19332
rect 3688 19323 3746 19329
rect 3970 19320 3976 19332
rect 4028 19320 4034 19372
rect 5442 19360 5448 19372
rect 5403 19332 5448 19360
rect 5442 19320 5448 19332
rect 5500 19320 5506 19372
rect 6365 19363 6423 19369
rect 6365 19329 6377 19363
rect 6411 19360 6423 19363
rect 6546 19360 6552 19372
rect 6411 19332 6552 19360
rect 6411 19329 6423 19332
rect 6365 19323 6423 19329
rect 6546 19320 6552 19332
rect 6604 19360 6610 19372
rect 7208 19360 7236 19400
rect 6604 19332 7236 19360
rect 6604 19320 6610 19332
rect 7282 19320 7288 19372
rect 7340 19360 7346 19372
rect 7340 19332 7385 19360
rect 7340 19320 7346 19332
rect 4706 19252 4712 19304
rect 4764 19292 4770 19304
rect 8404 19301 8432 19400
rect 11716 19400 12434 19428
rect 8665 19363 8723 19369
rect 8665 19329 8677 19363
rect 8711 19360 8723 19363
rect 9306 19360 9312 19372
rect 8711 19332 9312 19360
rect 8711 19329 8723 19332
rect 8665 19323 8723 19329
rect 9306 19320 9312 19332
rect 9364 19320 9370 19372
rect 9677 19363 9735 19369
rect 9677 19329 9689 19363
rect 9723 19360 9735 19363
rect 9950 19360 9956 19372
rect 9723 19332 9956 19360
rect 9723 19329 9735 19332
rect 9677 19323 9735 19329
rect 9950 19320 9956 19332
rect 10008 19320 10014 19372
rect 11716 19369 11744 19400
rect 11974 19369 11980 19372
rect 10321 19363 10379 19369
rect 10321 19329 10333 19363
rect 10367 19329 10379 19363
rect 10321 19323 10379 19329
rect 11701 19363 11759 19369
rect 11701 19329 11713 19363
rect 11747 19329 11759 19363
rect 11968 19360 11980 19369
rect 11935 19332 11980 19360
rect 11701 19323 11759 19329
rect 11968 19323 11980 19332
rect 5537 19295 5595 19301
rect 5537 19292 5549 19295
rect 4764 19264 5549 19292
rect 4764 19252 4770 19264
rect 5537 19261 5549 19264
rect 5583 19261 5595 19295
rect 5537 19255 5595 19261
rect 5629 19295 5687 19301
rect 5629 19261 5641 19295
rect 5675 19261 5687 19295
rect 5629 19255 5687 19261
rect 8389 19295 8447 19301
rect 8389 19261 8401 19295
rect 8435 19261 8447 19295
rect 8389 19255 8447 19261
rect 9493 19295 9551 19301
rect 9493 19261 9505 19295
rect 9539 19292 9551 19295
rect 10336 19292 10364 19323
rect 11974 19320 11980 19323
rect 12032 19320 12038 19372
rect 12406 19360 12434 19400
rect 13372 19400 14740 19428
rect 13372 19369 13400 19400
rect 14734 19388 14740 19400
rect 14792 19428 14798 19440
rect 15654 19428 15660 19440
rect 14792 19400 15660 19428
rect 14792 19388 14798 19400
rect 15654 19388 15660 19400
rect 15712 19388 15718 19440
rect 13630 19369 13636 19372
rect 13357 19363 13415 19369
rect 13357 19360 13369 19363
rect 12406 19332 13369 19360
rect 13357 19329 13369 19332
rect 13403 19329 13415 19363
rect 13624 19360 13636 19369
rect 13591 19332 13636 19360
rect 13357 19323 13415 19329
rect 13624 19323 13636 19332
rect 13630 19320 13636 19323
rect 13688 19320 13694 19372
rect 14642 19320 14648 19372
rect 14700 19360 14706 19372
rect 15013 19363 15071 19369
rect 15013 19360 15025 19363
rect 14700 19332 15025 19360
rect 14700 19320 14706 19332
rect 9539 19264 10364 19292
rect 9539 19261 9551 19264
rect 9493 19255 9551 19261
rect 4801 19227 4859 19233
rect 4801 19193 4813 19227
rect 4847 19224 4859 19227
rect 5350 19224 5356 19236
rect 4847 19196 5356 19224
rect 4847 19193 4859 19196
rect 4801 19187 4859 19193
rect 5350 19184 5356 19196
rect 5408 19224 5414 19236
rect 5644 19224 5672 19255
rect 5408 19196 5672 19224
rect 9508 19224 9536 19255
rect 9674 19224 9680 19236
rect 9508 19196 9680 19224
rect 5408 19184 5414 19196
rect 9674 19184 9680 19196
rect 9732 19184 9738 19236
rect 9766 19184 9772 19236
rect 9824 19224 9830 19236
rect 14752 19233 14780 19332
rect 15013 19329 15025 19332
rect 15059 19329 15071 19363
rect 15013 19323 15071 19329
rect 15562 19320 15568 19372
rect 15620 19360 15626 19372
rect 15620 19332 15700 19360
rect 15620 19320 15626 19332
rect 15672 19301 15700 19332
rect 15657 19295 15715 19301
rect 15657 19261 15669 19295
rect 15703 19261 15715 19295
rect 15856 19292 15884 19468
rect 16117 19465 16129 19499
rect 16163 19496 16175 19499
rect 19978 19496 19984 19508
rect 16163 19468 19984 19496
rect 16163 19465 16175 19468
rect 16117 19459 16175 19465
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 20070 19456 20076 19508
rect 20128 19496 20134 19508
rect 20717 19499 20775 19505
rect 20128 19468 20173 19496
rect 20128 19456 20134 19468
rect 20717 19465 20729 19499
rect 20763 19496 20775 19499
rect 20990 19496 20996 19508
rect 20763 19468 20996 19496
rect 20763 19465 20775 19468
rect 20717 19459 20775 19465
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 18690 19428 18696 19440
rect 15948 19400 18696 19428
rect 15948 19369 15976 19400
rect 18690 19388 18696 19400
rect 18748 19388 18754 19440
rect 19610 19428 19616 19440
rect 19536 19400 19616 19428
rect 15933 19363 15991 19369
rect 15933 19329 15945 19363
rect 15979 19329 15991 19363
rect 17310 19360 17316 19372
rect 15933 19323 15991 19329
rect 16040 19332 17172 19360
rect 17271 19332 17316 19360
rect 16040 19292 16068 19332
rect 15856 19264 16068 19292
rect 17144 19292 17172 19332
rect 17310 19320 17316 19332
rect 17368 19320 17374 19372
rect 17589 19363 17647 19369
rect 17589 19360 17601 19363
rect 17420 19332 17601 19360
rect 17420 19292 17448 19332
rect 17589 19329 17601 19332
rect 17635 19329 17647 19363
rect 17589 19323 17647 19329
rect 18414 19320 18420 19372
rect 18472 19320 18478 19372
rect 18598 19360 18604 19372
rect 18559 19332 18604 19360
rect 18598 19320 18604 19332
rect 18656 19320 18662 19372
rect 18877 19363 18935 19369
rect 18877 19329 18889 19363
rect 18923 19360 18935 19363
rect 18966 19360 18972 19372
rect 18923 19332 18972 19360
rect 18923 19329 18935 19332
rect 18877 19323 18935 19329
rect 18966 19320 18972 19332
rect 19024 19320 19030 19372
rect 19058 19320 19064 19372
rect 19116 19320 19122 19372
rect 17144 19264 17448 19292
rect 15657 19255 15715 19261
rect 18432 19233 18460 19320
rect 19076 19233 19104 19320
rect 19536 19233 19564 19400
rect 19610 19388 19616 19400
rect 19668 19388 19674 19440
rect 19702 19360 19708 19372
rect 19663 19332 19708 19360
rect 19702 19320 19708 19332
rect 19760 19320 19766 19372
rect 20162 19320 20168 19372
rect 20220 19360 20226 19372
rect 20257 19363 20315 19369
rect 20257 19360 20269 19363
rect 20220 19332 20269 19360
rect 20220 19320 20226 19332
rect 20257 19329 20269 19332
rect 20303 19329 20315 19363
rect 20257 19323 20315 19329
rect 20438 19320 20444 19372
rect 20496 19360 20502 19372
rect 20533 19363 20591 19369
rect 20533 19360 20545 19363
rect 20496 19332 20545 19360
rect 20496 19320 20502 19332
rect 20533 19329 20545 19332
rect 20579 19329 20591 19363
rect 20533 19323 20591 19329
rect 20898 19320 20904 19372
rect 20956 19360 20962 19372
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 20956 19332 21097 19360
rect 20956 19320 20962 19332
rect 21085 19329 21097 19332
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 10965 19227 11023 19233
rect 10965 19224 10977 19227
rect 9824 19196 10977 19224
rect 9824 19184 9830 19196
rect 10965 19193 10977 19196
rect 11011 19193 11023 19227
rect 10965 19187 11023 19193
rect 14737 19227 14795 19233
rect 14737 19193 14749 19227
rect 14783 19193 14795 19227
rect 14737 19187 14795 19193
rect 18417 19227 18475 19233
rect 18417 19193 18429 19227
rect 18463 19193 18475 19227
rect 18417 19187 18475 19193
rect 19061 19227 19119 19233
rect 19061 19193 19073 19227
rect 19107 19193 19119 19227
rect 19061 19187 19119 19193
rect 19521 19227 19579 19233
rect 19521 19193 19533 19227
rect 19567 19193 19579 19227
rect 19521 19187 19579 19193
rect 2222 19156 2228 19168
rect 2183 19128 2228 19156
rect 2222 19116 2228 19128
rect 2280 19116 2286 19168
rect 5074 19156 5080 19168
rect 5035 19128 5080 19156
rect 5074 19116 5080 19128
rect 5132 19116 5138 19168
rect 7469 19159 7527 19165
rect 7469 19125 7481 19159
rect 7515 19156 7527 19159
rect 7558 19156 7564 19168
rect 7515 19128 7564 19156
rect 7515 19125 7527 19128
rect 7469 19119 7527 19125
rect 7558 19116 7564 19128
rect 7616 19116 7622 19168
rect 8021 19159 8079 19165
rect 8021 19125 8033 19159
rect 8067 19156 8079 19159
rect 9858 19156 9864 19168
rect 8067 19128 9864 19156
rect 8067 19125 8079 19128
rect 8021 19119 8079 19125
rect 9858 19116 9864 19128
rect 9916 19116 9922 19168
rect 10042 19156 10048 19168
rect 10003 19128 10048 19156
rect 10042 19116 10048 19128
rect 10100 19116 10106 19168
rect 16666 19156 16672 19168
rect 16627 19128 16672 19156
rect 16666 19116 16672 19128
rect 16724 19116 16730 19168
rect 17773 19159 17831 19165
rect 17773 19125 17785 19159
rect 17819 19156 17831 19159
rect 17862 19156 17868 19168
rect 17819 19128 17868 19156
rect 17819 19125 17831 19128
rect 17773 19119 17831 19125
rect 17862 19116 17868 19128
rect 17920 19116 17926 19168
rect 21269 19159 21327 19165
rect 21269 19125 21281 19159
rect 21315 19156 21327 19159
rect 21358 19156 21364 19168
rect 21315 19128 21364 19156
rect 21315 19125 21327 19128
rect 21269 19119 21327 19125
rect 21358 19116 21364 19128
rect 21416 19116 21422 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1765 18955 1823 18961
rect 1765 18921 1777 18955
rect 1811 18952 1823 18955
rect 1946 18952 1952 18964
rect 1811 18924 1952 18952
rect 1811 18921 1823 18924
rect 1765 18915 1823 18921
rect 1946 18912 1952 18924
rect 2004 18912 2010 18964
rect 3789 18955 3847 18961
rect 3789 18921 3801 18955
rect 3835 18952 3847 18955
rect 3970 18952 3976 18964
rect 3835 18924 3976 18952
rect 3835 18921 3847 18924
rect 3789 18915 3847 18921
rect 3970 18912 3976 18924
rect 4028 18912 4034 18964
rect 4338 18912 4344 18964
rect 4396 18952 4402 18964
rect 5261 18955 5319 18961
rect 5261 18952 5273 18955
rect 4396 18924 5273 18952
rect 4396 18912 4402 18924
rect 5261 18921 5273 18924
rect 5307 18921 5319 18955
rect 5718 18952 5724 18964
rect 5679 18924 5724 18952
rect 5261 18915 5319 18921
rect 5276 18884 5304 18915
rect 5718 18912 5724 18924
rect 5776 18912 5782 18964
rect 6181 18955 6239 18961
rect 6181 18921 6193 18955
rect 6227 18952 6239 18955
rect 6914 18952 6920 18964
rect 6227 18924 6920 18952
rect 6227 18921 6239 18924
rect 6181 18915 6239 18921
rect 6914 18912 6920 18924
rect 6972 18912 6978 18964
rect 7282 18912 7288 18964
rect 7340 18952 7346 18964
rect 7377 18955 7435 18961
rect 7377 18952 7389 18955
rect 7340 18924 7389 18952
rect 7340 18912 7346 18924
rect 7377 18921 7389 18924
rect 7423 18921 7435 18955
rect 7834 18952 7840 18964
rect 7795 18924 7840 18952
rect 7377 18915 7435 18921
rect 7834 18912 7840 18924
rect 7892 18912 7898 18964
rect 8110 18952 8116 18964
rect 8071 18924 8116 18952
rect 8110 18912 8116 18924
rect 8168 18912 8174 18964
rect 8573 18955 8631 18961
rect 8573 18921 8585 18955
rect 8619 18952 8631 18955
rect 9214 18952 9220 18964
rect 8619 18924 9220 18952
rect 8619 18921 8631 18924
rect 8573 18915 8631 18921
rect 9214 18912 9220 18924
rect 9272 18912 9278 18964
rect 13725 18955 13783 18961
rect 13725 18921 13737 18955
rect 13771 18952 13783 18955
rect 13814 18952 13820 18964
rect 13771 18924 13820 18952
rect 13771 18921 13783 18924
rect 13725 18915 13783 18921
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 15381 18955 15439 18961
rect 15381 18921 15393 18955
rect 15427 18952 15439 18955
rect 17770 18952 17776 18964
rect 15427 18924 17776 18952
rect 15427 18921 15439 18924
rect 15381 18915 15439 18921
rect 17770 18912 17776 18924
rect 17828 18912 17834 18964
rect 18690 18952 18696 18964
rect 18651 18924 18696 18952
rect 18690 18912 18696 18924
rect 18748 18912 18754 18964
rect 20165 18955 20223 18961
rect 20165 18921 20177 18955
rect 20211 18952 20223 18955
rect 20530 18952 20536 18964
rect 20211 18924 20536 18952
rect 20211 18921 20223 18924
rect 20165 18915 20223 18921
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 20625 18955 20683 18961
rect 20625 18921 20637 18955
rect 20671 18952 20683 18955
rect 21542 18952 21548 18964
rect 20671 18924 21548 18952
rect 20671 18921 20683 18924
rect 20625 18915 20683 18921
rect 21542 18912 21548 18924
rect 21600 18912 21606 18964
rect 6641 18887 6699 18893
rect 5276 18856 5580 18884
rect 4985 18819 5043 18825
rect 4985 18785 4997 18819
rect 5031 18816 5043 18819
rect 5442 18816 5448 18828
rect 5031 18788 5448 18816
rect 5031 18785 5043 18788
rect 4985 18779 5043 18785
rect 5442 18776 5448 18788
rect 5500 18776 5506 18828
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18748 2099 18751
rect 3418 18748 3424 18760
rect 2087 18720 3424 18748
rect 2087 18717 2099 18720
rect 2041 18711 2099 18717
rect 3418 18708 3424 18720
rect 3476 18708 3482 18760
rect 4433 18751 4491 18757
rect 4433 18717 4445 18751
rect 4479 18717 4491 18751
rect 4433 18711 4491 18717
rect 2314 18689 2320 18692
rect 2308 18643 2320 18689
rect 2372 18680 2378 18692
rect 4154 18680 4160 18692
rect 2372 18652 2408 18680
rect 3436 18652 4160 18680
rect 2314 18640 2320 18643
rect 2372 18640 2378 18652
rect 3436 18621 3464 18652
rect 4154 18640 4160 18652
rect 4212 18680 4218 18692
rect 4448 18680 4476 18711
rect 4212 18652 4476 18680
rect 5552 18680 5580 18856
rect 6641 18853 6653 18887
rect 6687 18884 6699 18887
rect 6730 18884 6736 18896
rect 6687 18856 6736 18884
rect 6687 18853 6699 18856
rect 6641 18847 6699 18853
rect 6730 18844 6736 18856
rect 6788 18844 6794 18896
rect 7101 18887 7159 18893
rect 7101 18853 7113 18887
rect 7147 18884 7159 18887
rect 7190 18884 7196 18896
rect 7147 18856 7196 18884
rect 7147 18853 7159 18856
rect 7101 18847 7159 18853
rect 7190 18844 7196 18856
rect 7248 18844 7254 18896
rect 6822 18776 6828 18828
rect 6880 18816 6886 18828
rect 7300 18816 7328 18912
rect 19521 18887 19579 18893
rect 19521 18853 19533 18887
rect 19567 18884 19579 18887
rect 22094 18884 22100 18896
rect 19567 18856 22100 18884
rect 19567 18853 19579 18856
rect 19521 18847 19579 18853
rect 22094 18844 22100 18856
rect 22152 18844 22158 18896
rect 6880 18788 7328 18816
rect 11977 18819 12035 18825
rect 6880 18776 6886 18788
rect 11977 18785 11989 18819
rect 12023 18816 12035 18819
rect 12066 18816 12072 18828
rect 12023 18788 12072 18816
rect 12023 18785 12035 18788
rect 11977 18779 12035 18785
rect 12066 18776 12072 18788
rect 12124 18776 12130 18828
rect 13078 18816 13084 18828
rect 13039 18788 13084 18816
rect 13078 18776 13084 18788
rect 13136 18776 13142 18828
rect 15654 18816 15660 18828
rect 15615 18788 15660 18816
rect 15654 18776 15660 18788
rect 15712 18776 15718 18828
rect 6917 18751 6975 18757
rect 6917 18717 6929 18751
rect 6963 18748 6975 18751
rect 7190 18748 7196 18760
rect 6963 18720 7196 18748
rect 6963 18717 6975 18720
rect 6917 18711 6975 18717
rect 7190 18708 7196 18720
rect 7248 18708 7254 18760
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18748 9551 18751
rect 10594 18748 10600 18760
rect 9539 18720 10600 18748
rect 9539 18717 9551 18720
rect 9493 18711 9551 18717
rect 9876 18692 9904 18720
rect 10594 18708 10600 18720
rect 10652 18708 10658 18760
rect 15194 18748 15200 18760
rect 15155 18720 15200 18748
rect 15194 18708 15200 18720
rect 15252 18708 15258 18760
rect 15924 18751 15982 18757
rect 15924 18717 15936 18751
rect 15970 18748 15982 18751
rect 16666 18748 16672 18760
rect 15970 18720 16672 18748
rect 15970 18717 15982 18720
rect 15924 18711 15982 18717
rect 16666 18708 16672 18720
rect 16724 18708 16730 18760
rect 17313 18751 17371 18757
rect 17313 18748 17325 18751
rect 17052 18720 17325 18748
rect 9766 18689 9772 18692
rect 9760 18680 9772 18689
rect 5552 18652 6914 18680
rect 9727 18652 9772 18680
rect 4212 18640 4218 18652
rect 3421 18615 3479 18621
rect 3421 18581 3433 18615
rect 3467 18581 3479 18615
rect 6886 18612 6914 18652
rect 9760 18643 9772 18652
rect 9766 18640 9772 18643
rect 9824 18640 9830 18692
rect 9858 18640 9864 18692
rect 9916 18640 9922 18692
rect 11054 18640 11060 18692
rect 11112 18680 11118 18692
rect 12069 18683 12127 18689
rect 12069 18680 12081 18683
rect 11112 18652 12081 18680
rect 11112 18640 11118 18652
rect 12069 18649 12081 18652
rect 12115 18649 12127 18683
rect 12069 18643 12127 18649
rect 12161 18683 12219 18689
rect 12161 18649 12173 18683
rect 12207 18680 12219 18683
rect 12802 18680 12808 18692
rect 12207 18652 12808 18680
rect 12207 18649 12219 18652
rect 12161 18643 12219 18649
rect 12802 18640 12808 18652
rect 12860 18640 12866 18692
rect 13357 18683 13415 18689
rect 13357 18649 13369 18683
rect 13403 18680 13415 18683
rect 14093 18683 14151 18689
rect 14093 18680 14105 18683
rect 13403 18652 14105 18680
rect 13403 18649 13415 18652
rect 13357 18643 13415 18649
rect 14093 18649 14105 18652
rect 14139 18649 14151 18683
rect 14093 18643 14151 18649
rect 9217 18615 9275 18621
rect 9217 18612 9229 18615
rect 6886 18584 9229 18612
rect 3421 18575 3479 18581
rect 9217 18581 9229 18584
rect 9263 18612 9275 18615
rect 9306 18612 9312 18624
rect 9263 18584 9312 18612
rect 9263 18581 9275 18584
rect 9217 18575 9275 18581
rect 9306 18572 9312 18584
rect 9364 18572 9370 18624
rect 10870 18612 10876 18624
rect 10831 18584 10876 18612
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 11146 18612 11152 18624
rect 11107 18584 11152 18612
rect 11146 18572 11152 18584
rect 11204 18572 11210 18624
rect 12529 18615 12587 18621
rect 12529 18581 12541 18615
rect 12575 18612 12587 18615
rect 13265 18615 13323 18621
rect 13265 18612 13277 18615
rect 12575 18584 13277 18612
rect 12575 18581 12587 18584
rect 12529 18575 12587 18581
rect 13265 18581 13277 18584
rect 13311 18581 13323 18615
rect 14550 18612 14556 18624
rect 14511 18584 14556 18612
rect 13265 18575 13323 18581
rect 14550 18572 14556 18584
rect 14608 18572 14614 18624
rect 16942 18572 16948 18624
rect 17000 18612 17006 18624
rect 17052 18621 17080 18720
rect 17313 18717 17325 18720
rect 17359 18717 17371 18751
rect 17313 18711 17371 18717
rect 17402 18708 17408 18760
rect 17460 18748 17466 18760
rect 18233 18751 18291 18757
rect 18233 18748 18245 18751
rect 17460 18720 18245 18748
rect 17460 18708 17466 18720
rect 18233 18717 18245 18720
rect 18279 18717 18291 18751
rect 18233 18711 18291 18717
rect 18322 18708 18328 18760
rect 18380 18748 18386 18760
rect 18877 18751 18935 18757
rect 18877 18748 18889 18751
rect 18380 18720 18889 18748
rect 18380 18708 18386 18720
rect 18877 18717 18889 18720
rect 18923 18717 18935 18751
rect 18877 18711 18935 18717
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18717 19763 18751
rect 19978 18748 19984 18760
rect 19939 18720 19984 18748
rect 19705 18711 19763 18717
rect 19720 18680 19748 18711
rect 19978 18708 19984 18720
rect 20036 18708 20042 18760
rect 20806 18748 20812 18760
rect 20767 18720 20812 18748
rect 20806 18708 20812 18720
rect 20864 18708 20870 18760
rect 21085 18751 21143 18757
rect 21085 18717 21097 18751
rect 21131 18748 21143 18751
rect 21174 18748 21180 18760
rect 21131 18720 21180 18748
rect 21131 18717 21143 18720
rect 21085 18711 21143 18717
rect 21174 18708 21180 18720
rect 21232 18708 21238 18760
rect 21542 18680 21548 18692
rect 19720 18652 21548 18680
rect 21542 18640 21548 18652
rect 21600 18640 21606 18692
rect 17037 18615 17095 18621
rect 17037 18612 17049 18615
rect 17000 18584 17049 18612
rect 17000 18572 17006 18584
rect 17037 18581 17049 18584
rect 17083 18581 17095 18615
rect 17954 18612 17960 18624
rect 17915 18584 17960 18612
rect 17037 18575 17095 18581
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 18414 18612 18420 18624
rect 18375 18584 18420 18612
rect 18414 18572 18420 18584
rect 18472 18572 18478 18624
rect 21266 18612 21272 18624
rect 21227 18584 21272 18612
rect 21266 18572 21272 18584
rect 21324 18572 21330 18624
rect 1104 18522 21896 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21896 18522
rect 1104 18448 21896 18470
rect 2038 18408 2044 18420
rect 1999 18380 2044 18408
rect 2038 18368 2044 18380
rect 2096 18368 2102 18420
rect 2682 18408 2688 18420
rect 2643 18380 2688 18408
rect 2682 18368 2688 18380
rect 2740 18368 2746 18420
rect 3142 18408 3148 18420
rect 3103 18380 3148 18408
rect 3142 18368 3148 18380
rect 3200 18368 3206 18420
rect 4246 18408 4252 18420
rect 4207 18380 4252 18408
rect 4246 18368 4252 18380
rect 4304 18368 4310 18420
rect 7190 18408 7196 18420
rect 7151 18380 7196 18408
rect 7190 18368 7196 18380
rect 7248 18368 7254 18420
rect 9493 18411 9551 18417
rect 9493 18377 9505 18411
rect 9539 18408 9551 18411
rect 9674 18408 9680 18420
rect 9539 18380 9680 18408
rect 9539 18377 9551 18380
rect 9493 18371 9551 18377
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 10042 18368 10048 18420
rect 10100 18408 10106 18420
rect 10689 18411 10747 18417
rect 10689 18408 10701 18411
rect 10100 18380 10701 18408
rect 10100 18368 10106 18380
rect 10689 18377 10701 18380
rect 10735 18377 10747 18411
rect 10689 18371 10747 18377
rect 10781 18411 10839 18417
rect 10781 18377 10793 18411
rect 10827 18408 10839 18411
rect 11146 18408 11152 18420
rect 10827 18380 11152 18408
rect 10827 18377 10839 18380
rect 10781 18371 10839 18377
rect 11146 18368 11152 18380
rect 11204 18368 11210 18420
rect 12158 18408 12164 18420
rect 12119 18380 12164 18408
rect 12158 18368 12164 18380
rect 12216 18368 12222 18420
rect 17402 18408 17408 18420
rect 12406 18380 17408 18408
rect 2406 18300 2412 18352
rect 2464 18340 2470 18352
rect 3421 18343 3479 18349
rect 3421 18340 3433 18343
rect 2464 18312 3433 18340
rect 2464 18300 2470 18312
rect 3421 18309 3433 18312
rect 3467 18309 3479 18343
rect 9858 18340 9864 18352
rect 3421 18303 3479 18309
rect 8128 18312 9864 18340
rect 1670 18272 1676 18284
rect 1631 18244 1676 18272
rect 1670 18232 1676 18244
rect 1728 18232 1734 18284
rect 4801 18275 4859 18281
rect 4801 18241 4813 18275
rect 4847 18272 4859 18275
rect 5074 18272 5080 18284
rect 4847 18244 5080 18272
rect 4847 18241 4859 18244
rect 4801 18235 4859 18241
rect 5074 18232 5080 18244
rect 5132 18232 5138 18284
rect 8128 18281 8156 18312
rect 9858 18300 9864 18312
rect 9916 18300 9922 18352
rect 8386 18281 8392 18284
rect 6825 18275 6883 18281
rect 6825 18241 6837 18275
rect 6871 18272 6883 18275
rect 7469 18275 7527 18281
rect 7469 18272 7481 18275
rect 6871 18244 7481 18272
rect 6871 18241 6883 18244
rect 6825 18235 6883 18241
rect 7469 18241 7481 18244
rect 7515 18241 7527 18275
rect 7469 18235 7527 18241
rect 8113 18275 8171 18281
rect 8113 18241 8125 18275
rect 8159 18241 8171 18275
rect 8380 18272 8392 18281
rect 8347 18244 8392 18272
rect 8113 18235 8171 18241
rect 8380 18235 8392 18244
rect 6546 18204 6552 18216
rect 6507 18176 6552 18204
rect 6546 18164 6552 18176
rect 6604 18164 6610 18216
rect 6733 18207 6791 18213
rect 6733 18173 6745 18207
rect 6779 18204 6791 18207
rect 7098 18204 7104 18216
rect 6779 18176 7104 18204
rect 6779 18173 6791 18176
rect 6733 18167 6791 18173
rect 7098 18164 7104 18176
rect 7156 18164 7162 18216
rect 6638 18096 6644 18148
rect 6696 18136 6702 18148
rect 8128 18136 8156 18235
rect 8386 18232 8392 18235
rect 8444 18232 8450 18284
rect 9950 18232 9956 18284
rect 10008 18272 10014 18284
rect 10045 18275 10103 18281
rect 10045 18272 10057 18275
rect 10008 18244 10057 18272
rect 10008 18232 10014 18244
rect 10045 18241 10057 18244
rect 10091 18241 10103 18275
rect 10045 18235 10103 18241
rect 11517 18275 11575 18281
rect 11517 18241 11529 18275
rect 11563 18241 11575 18275
rect 11517 18235 11575 18241
rect 10597 18207 10655 18213
rect 10597 18173 10609 18207
rect 10643 18204 10655 18207
rect 10870 18204 10876 18216
rect 10643 18176 10876 18204
rect 10643 18173 10655 18176
rect 10597 18167 10655 18173
rect 10870 18164 10876 18176
rect 10928 18204 10934 18216
rect 11532 18204 11560 18235
rect 10928 18176 11560 18204
rect 10928 18164 10934 18176
rect 6696 18108 8156 18136
rect 11149 18139 11207 18145
rect 6696 18096 6702 18108
rect 11149 18105 11161 18139
rect 11195 18136 11207 18139
rect 12406 18136 12434 18380
rect 17402 18368 17408 18380
rect 17460 18368 17466 18420
rect 18322 18408 18328 18420
rect 18283 18380 18328 18408
rect 18322 18368 18328 18380
rect 18380 18368 18386 18420
rect 18874 18368 18880 18420
rect 18932 18408 18938 18420
rect 19613 18411 19671 18417
rect 19613 18408 19625 18411
rect 18932 18380 19625 18408
rect 18932 18368 18938 18380
rect 19613 18377 19625 18380
rect 19659 18377 19671 18411
rect 19613 18371 19671 18377
rect 20717 18411 20775 18417
rect 20717 18377 20729 18411
rect 20763 18408 20775 18411
rect 21450 18408 21456 18420
rect 20763 18380 21456 18408
rect 20763 18377 20775 18380
rect 20717 18371 20775 18377
rect 21450 18368 21456 18380
rect 21508 18368 21514 18420
rect 17212 18343 17270 18349
rect 17212 18309 17224 18343
rect 17258 18340 17270 18343
rect 17954 18340 17960 18352
rect 17258 18312 17960 18340
rect 17258 18309 17270 18312
rect 17212 18303 17270 18309
rect 17954 18300 17960 18312
rect 18012 18300 18018 18352
rect 18340 18340 18368 18368
rect 18340 18312 19196 18340
rect 16117 18275 16175 18281
rect 16117 18241 16129 18275
rect 16163 18272 16175 18275
rect 16163 18244 18644 18272
rect 16163 18241 16175 18244
rect 16117 18235 16175 18241
rect 15654 18164 15660 18216
rect 15712 18204 15718 18216
rect 16945 18207 17003 18213
rect 16945 18204 16957 18207
rect 15712 18176 16957 18204
rect 15712 18164 15718 18176
rect 16945 18173 16957 18176
rect 16991 18173 17003 18207
rect 16945 18167 17003 18173
rect 18616 18145 18644 18244
rect 18690 18232 18696 18284
rect 18748 18272 18754 18284
rect 18969 18275 19027 18281
rect 18969 18272 18981 18275
rect 18748 18244 18981 18272
rect 18748 18232 18754 18244
rect 18969 18241 18981 18244
rect 19015 18241 19027 18275
rect 18969 18235 19027 18241
rect 19058 18204 19064 18216
rect 19019 18176 19064 18204
rect 19058 18164 19064 18176
rect 19116 18164 19122 18216
rect 19168 18213 19196 18312
rect 19978 18272 19984 18284
rect 19939 18244 19984 18272
rect 19978 18232 19984 18244
rect 20036 18232 20042 18284
rect 20533 18275 20591 18281
rect 20533 18241 20545 18275
rect 20579 18241 20591 18275
rect 20533 18235 20591 18241
rect 19153 18207 19211 18213
rect 19153 18173 19165 18207
rect 19199 18173 19211 18207
rect 19153 18167 19211 18173
rect 11195 18108 12434 18136
rect 18601 18139 18659 18145
rect 11195 18105 11207 18108
rect 11149 18099 11207 18105
rect 18601 18105 18613 18139
rect 18647 18105 18659 18139
rect 18601 18099 18659 18105
rect 18782 18096 18788 18148
rect 18840 18136 18846 18148
rect 20165 18139 20223 18145
rect 20165 18136 20177 18139
rect 18840 18108 20177 18136
rect 18840 18096 18846 18108
rect 20165 18105 20177 18108
rect 20211 18105 20223 18139
rect 20165 18099 20223 18105
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 4985 18071 5043 18077
rect 4985 18037 4997 18071
rect 5031 18068 5043 18071
rect 5442 18068 5448 18080
rect 5031 18040 5448 18068
rect 5031 18037 5043 18040
rect 4985 18031 5043 18037
rect 5442 18028 5448 18040
rect 5500 18028 5506 18080
rect 12713 18071 12771 18077
rect 12713 18037 12725 18071
rect 12759 18068 12771 18071
rect 12802 18068 12808 18080
rect 12759 18040 12808 18068
rect 12759 18037 12771 18040
rect 12713 18031 12771 18037
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 14734 18028 14740 18080
rect 14792 18068 14798 18080
rect 14918 18068 14924 18080
rect 14792 18040 14924 18068
rect 14792 18028 14798 18040
rect 14918 18028 14924 18040
rect 14976 18068 14982 18080
rect 15289 18071 15347 18077
rect 15289 18068 15301 18071
rect 14976 18040 15301 18068
rect 14976 18028 14982 18040
rect 15289 18037 15301 18040
rect 15335 18037 15347 18071
rect 15289 18031 15347 18037
rect 16301 18071 16359 18077
rect 16301 18037 16313 18071
rect 16347 18068 16359 18071
rect 17678 18068 17684 18080
rect 16347 18040 17684 18068
rect 16347 18037 16359 18040
rect 16301 18031 16359 18037
rect 17678 18028 17684 18040
rect 17736 18028 17742 18080
rect 18874 18028 18880 18080
rect 18932 18068 18938 18080
rect 20548 18068 20576 18235
rect 20990 18232 20996 18284
rect 21048 18272 21054 18284
rect 21085 18275 21143 18281
rect 21085 18272 21097 18275
rect 21048 18244 21097 18272
rect 21048 18232 21054 18244
rect 21085 18241 21097 18244
rect 21131 18241 21143 18275
rect 21085 18235 21143 18241
rect 20622 18096 20628 18148
rect 20680 18136 20686 18148
rect 21269 18139 21327 18145
rect 21269 18136 21281 18139
rect 20680 18108 21281 18136
rect 20680 18096 20686 18108
rect 21269 18105 21281 18108
rect 21315 18105 21327 18139
rect 21269 18099 21327 18105
rect 18932 18040 20576 18068
rect 18932 18028 18938 18040
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 2314 17864 2320 17876
rect 2275 17836 2320 17864
rect 2314 17824 2320 17836
rect 2372 17824 2378 17876
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 7098 17864 7104 17876
rect 4120 17836 6914 17864
rect 7059 17836 7104 17864
rect 4120 17824 4126 17836
rect 1578 17756 1584 17808
rect 1636 17796 1642 17808
rect 2593 17799 2651 17805
rect 2593 17796 2605 17799
rect 1636 17768 2605 17796
rect 1636 17756 1642 17768
rect 2593 17765 2605 17768
rect 2639 17765 2651 17799
rect 6886 17796 6914 17836
rect 7098 17824 7104 17836
rect 7156 17824 7162 17876
rect 10318 17864 10324 17876
rect 10279 17836 10324 17864
rect 10318 17824 10324 17836
rect 10376 17824 10382 17876
rect 17497 17867 17555 17873
rect 17497 17833 17509 17867
rect 17543 17864 17555 17867
rect 19058 17864 19064 17876
rect 17543 17836 19064 17864
rect 17543 17833 17555 17836
rect 17497 17827 17555 17833
rect 19058 17824 19064 17836
rect 19116 17824 19122 17876
rect 19429 17867 19487 17873
rect 19429 17833 19441 17867
rect 19475 17864 19487 17867
rect 19978 17864 19984 17876
rect 19475 17836 19984 17864
rect 19475 17833 19487 17836
rect 19429 17827 19487 17833
rect 19978 17824 19984 17836
rect 20036 17824 20042 17876
rect 17957 17799 18015 17805
rect 6886 17768 11836 17796
rect 2593 17759 2651 17765
rect 6273 17731 6331 17737
rect 6273 17697 6285 17731
rect 6319 17728 6331 17731
rect 6638 17728 6644 17740
rect 6319 17700 6644 17728
rect 6319 17697 6331 17700
rect 6273 17691 6331 17697
rect 1578 17620 1584 17672
rect 1636 17660 1642 17672
rect 1673 17663 1731 17669
rect 1673 17660 1685 17663
rect 1636 17632 1685 17660
rect 1636 17620 1642 17632
rect 1673 17629 1685 17632
rect 1719 17629 1731 17663
rect 1673 17623 1731 17629
rect 5718 17620 5724 17672
rect 5776 17660 5782 17672
rect 6288 17660 6316 17691
rect 6638 17688 6644 17700
rect 6696 17688 6702 17740
rect 7374 17688 7380 17740
rect 7432 17728 7438 17740
rect 7561 17731 7619 17737
rect 7561 17728 7573 17731
rect 7432 17700 7573 17728
rect 7432 17688 7438 17700
rect 7561 17697 7573 17700
rect 7607 17697 7619 17731
rect 7742 17728 7748 17740
rect 7703 17700 7748 17728
rect 7561 17691 7619 17697
rect 7742 17688 7748 17700
rect 7800 17688 7806 17740
rect 11238 17688 11244 17740
rect 11296 17728 11302 17740
rect 11808 17737 11836 17768
rect 17957 17765 17969 17799
rect 18003 17796 18015 17799
rect 18782 17796 18788 17808
rect 18003 17768 18788 17796
rect 18003 17765 18015 17768
rect 17957 17759 18015 17765
rect 18782 17756 18788 17768
rect 18840 17756 18846 17808
rect 18877 17799 18935 17805
rect 18877 17765 18889 17799
rect 18923 17796 18935 17799
rect 18923 17768 21128 17796
rect 18923 17765 18935 17768
rect 18877 17759 18935 17765
rect 11609 17731 11667 17737
rect 11609 17728 11621 17731
rect 11296 17700 11621 17728
rect 11296 17688 11302 17700
rect 11609 17697 11621 17700
rect 11655 17697 11667 17731
rect 11609 17691 11667 17697
rect 11793 17731 11851 17737
rect 11793 17697 11805 17731
rect 11839 17697 11851 17731
rect 16942 17728 16948 17740
rect 16903 17700 16948 17728
rect 11793 17691 11851 17697
rect 16942 17688 16948 17700
rect 17000 17688 17006 17740
rect 17678 17688 17684 17740
rect 17736 17728 17742 17740
rect 17736 17700 18828 17728
rect 17736 17688 17742 17700
rect 5776 17632 6316 17660
rect 5776 17620 5782 17632
rect 16390 17620 16396 17672
rect 16448 17660 16454 17672
rect 17037 17663 17095 17669
rect 17037 17660 17049 17663
rect 16448 17632 17049 17660
rect 16448 17620 16454 17632
rect 17037 17629 17049 17632
rect 17083 17629 17095 17663
rect 17770 17660 17776 17672
rect 17731 17632 17776 17660
rect 17037 17623 17095 17629
rect 17770 17620 17776 17632
rect 17828 17620 17834 17672
rect 18233 17663 18291 17669
rect 18233 17629 18245 17663
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 18693 17663 18751 17669
rect 18693 17629 18705 17663
rect 18739 17629 18751 17663
rect 18800 17660 18828 17700
rect 19245 17663 19303 17669
rect 19245 17660 19257 17663
rect 18800 17632 19257 17660
rect 18693 17623 18751 17629
rect 19245 17629 19257 17632
rect 19291 17629 19303 17663
rect 19245 17623 19303 17629
rect 6028 17595 6086 17601
rect 6028 17561 6040 17595
rect 6074 17592 6086 17595
rect 8018 17592 8024 17604
rect 6074 17564 8024 17592
rect 6074 17561 6086 17564
rect 6028 17555 6086 17561
rect 8018 17552 8024 17564
rect 8076 17552 8082 17604
rect 11885 17595 11943 17601
rect 11885 17561 11897 17595
rect 11931 17592 11943 17595
rect 18248 17592 18276 17623
rect 18708 17592 18736 17623
rect 19610 17620 19616 17672
rect 19668 17660 19674 17672
rect 19705 17663 19763 17669
rect 19705 17660 19717 17663
rect 19668 17632 19717 17660
rect 19668 17620 19674 17632
rect 19705 17629 19717 17632
rect 19751 17629 19763 17663
rect 19705 17623 19763 17629
rect 20070 17620 20076 17672
rect 20128 17660 20134 17672
rect 21100 17669 21128 17768
rect 20533 17663 20591 17669
rect 20533 17660 20545 17663
rect 20128 17632 20545 17660
rect 20128 17620 20134 17632
rect 20533 17629 20545 17632
rect 20579 17629 20591 17663
rect 20533 17623 20591 17629
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 18782 17592 18788 17604
rect 11931 17564 12664 17592
rect 18248 17564 18552 17592
rect 18708 17564 18788 17592
rect 11931 17561 11943 17564
rect 11885 17555 11943 17561
rect 3142 17524 3148 17536
rect 3103 17496 3148 17524
rect 3142 17484 3148 17496
rect 3200 17484 3206 17536
rect 4893 17527 4951 17533
rect 4893 17493 4905 17527
rect 4939 17524 4951 17527
rect 5626 17524 5632 17536
rect 4939 17496 5632 17524
rect 4939 17493 4951 17496
rect 4893 17487 4951 17493
rect 5626 17484 5632 17496
rect 5684 17484 5690 17536
rect 7466 17524 7472 17536
rect 7379 17496 7472 17524
rect 7466 17484 7472 17496
rect 7524 17524 7530 17536
rect 8205 17527 8263 17533
rect 8205 17524 8217 17527
rect 7524 17496 8217 17524
rect 7524 17484 7530 17496
rect 8205 17493 8217 17496
rect 8251 17524 8263 17527
rect 10042 17524 10048 17536
rect 8251 17496 10048 17524
rect 8251 17493 8263 17496
rect 8205 17487 8263 17493
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 12253 17527 12311 17533
rect 12253 17493 12265 17527
rect 12299 17524 12311 17527
rect 12434 17524 12440 17536
rect 12299 17496 12440 17524
rect 12299 17493 12311 17496
rect 12253 17487 12311 17493
rect 12434 17484 12440 17496
rect 12492 17484 12498 17536
rect 12636 17533 12664 17564
rect 12621 17527 12679 17533
rect 12621 17493 12633 17527
rect 12667 17524 12679 17527
rect 12802 17524 12808 17536
rect 12667 17496 12808 17524
rect 12667 17493 12679 17496
rect 12621 17487 12679 17493
rect 12802 17484 12808 17496
rect 12860 17484 12866 17536
rect 14734 17524 14740 17536
rect 14695 17496 14740 17524
rect 14734 17484 14740 17496
rect 14792 17484 14798 17536
rect 16485 17527 16543 17533
rect 16485 17493 16497 17527
rect 16531 17524 16543 17527
rect 16942 17524 16948 17536
rect 16531 17496 16948 17524
rect 16531 17493 16543 17496
rect 16485 17487 16543 17493
rect 16942 17484 16948 17496
rect 17000 17524 17006 17536
rect 17129 17527 17187 17533
rect 17129 17524 17141 17527
rect 17000 17496 17141 17524
rect 17000 17484 17006 17496
rect 17129 17493 17141 17496
rect 17175 17493 17187 17527
rect 17129 17487 17187 17493
rect 18322 17484 18328 17536
rect 18380 17524 18386 17536
rect 18417 17527 18475 17533
rect 18417 17524 18429 17527
rect 18380 17496 18429 17524
rect 18380 17484 18386 17496
rect 18417 17493 18429 17496
rect 18463 17493 18475 17527
rect 18524 17524 18552 17564
rect 18782 17552 18788 17564
rect 18840 17552 18846 17604
rect 20898 17592 20904 17604
rect 19904 17564 20904 17592
rect 19794 17524 19800 17536
rect 18524 17496 19800 17524
rect 18417 17487 18475 17493
rect 19794 17484 19800 17496
rect 19852 17484 19858 17536
rect 19904 17533 19932 17564
rect 20898 17552 20904 17564
rect 20956 17552 20962 17604
rect 19889 17527 19947 17533
rect 19889 17493 19901 17527
rect 19935 17493 19947 17527
rect 20714 17524 20720 17536
rect 20675 17496 20720 17524
rect 19889 17487 19947 17493
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 21266 17524 21272 17536
rect 21227 17496 21272 17524
rect 21266 17484 21272 17496
rect 21324 17484 21330 17536
rect 1104 17434 21896 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21896 17434
rect 1104 17360 21896 17382
rect 3326 17280 3332 17332
rect 3384 17320 3390 17332
rect 3697 17323 3755 17329
rect 3697 17320 3709 17323
rect 3384 17292 3709 17320
rect 3384 17280 3390 17292
rect 3697 17289 3709 17292
rect 3743 17289 3755 17323
rect 3697 17283 3755 17289
rect 4985 17323 5043 17329
rect 4985 17289 4997 17323
rect 5031 17320 5043 17323
rect 5258 17320 5264 17332
rect 5031 17292 5264 17320
rect 5031 17289 5043 17292
rect 4985 17283 5043 17289
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 5442 17280 5448 17332
rect 5500 17320 5506 17332
rect 14090 17320 14096 17332
rect 5500 17292 14096 17320
rect 5500 17280 5506 17292
rect 14090 17280 14096 17292
rect 14148 17280 14154 17332
rect 14645 17323 14703 17329
rect 14645 17289 14657 17323
rect 14691 17320 14703 17323
rect 15197 17323 15255 17329
rect 15197 17320 15209 17323
rect 14691 17292 15209 17320
rect 14691 17289 14703 17292
rect 14645 17283 14703 17289
rect 15197 17289 15209 17292
rect 15243 17289 15255 17323
rect 15197 17283 15255 17289
rect 17773 17323 17831 17329
rect 17773 17289 17785 17323
rect 17819 17320 17831 17323
rect 18690 17320 18696 17332
rect 17819 17292 18696 17320
rect 17819 17289 17831 17292
rect 17773 17283 17831 17289
rect 18690 17280 18696 17292
rect 18748 17280 18754 17332
rect 18966 17320 18972 17332
rect 18927 17292 18972 17320
rect 18966 17280 18972 17292
rect 19024 17280 19030 17332
rect 19610 17320 19616 17332
rect 19571 17292 19616 17320
rect 19610 17280 19616 17292
rect 19668 17280 19674 17332
rect 20070 17320 20076 17332
rect 20031 17292 20076 17320
rect 20070 17280 20076 17292
rect 20128 17280 20134 17332
rect 3605 17255 3663 17261
rect 3605 17221 3617 17255
rect 3651 17252 3663 17255
rect 4341 17255 4399 17261
rect 4341 17252 4353 17255
rect 3651 17224 4353 17252
rect 3651 17221 3663 17224
rect 3605 17215 3663 17221
rect 4341 17221 4353 17224
rect 4387 17252 4399 17255
rect 7466 17252 7472 17264
rect 4387 17224 7472 17252
rect 4387 17221 4399 17224
rect 4341 17215 4399 17221
rect 7466 17212 7472 17224
rect 7524 17212 7530 17264
rect 12434 17212 12440 17264
rect 12492 17252 12498 17264
rect 12621 17255 12679 17261
rect 12621 17252 12633 17255
rect 12492 17224 12633 17252
rect 12492 17212 12498 17224
rect 12621 17221 12633 17224
rect 12667 17221 12679 17255
rect 14182 17252 14188 17264
rect 14143 17224 14188 17252
rect 12621 17215 12679 17221
rect 14182 17212 14188 17224
rect 14240 17212 14246 17264
rect 17862 17212 17868 17264
rect 17920 17252 17926 17264
rect 17920 17224 19196 17252
rect 17920 17212 17926 17224
rect 2705 17187 2763 17193
rect 2705 17153 2717 17187
rect 2751 17184 2763 17187
rect 3326 17184 3332 17196
rect 2751 17156 3332 17184
rect 2751 17153 2763 17156
rect 2705 17147 2763 17153
rect 3326 17144 3332 17156
rect 3384 17144 3390 17196
rect 5626 17184 5632 17196
rect 5539 17156 5632 17184
rect 5626 17144 5632 17156
rect 5684 17184 5690 17196
rect 6546 17184 6552 17196
rect 5684 17156 6552 17184
rect 5684 17144 5690 17156
rect 6546 17144 6552 17156
rect 6604 17144 6610 17196
rect 7282 17144 7288 17196
rect 7340 17184 7346 17196
rect 7834 17184 7840 17196
rect 7340 17156 7840 17184
rect 7340 17144 7346 17156
rect 7834 17144 7840 17156
rect 7892 17144 7898 17196
rect 9214 17184 9220 17196
rect 9175 17156 9220 17184
rect 9214 17144 9220 17156
rect 9272 17144 9278 17196
rect 12713 17187 12771 17193
rect 12713 17153 12725 17187
rect 12759 17184 12771 17187
rect 13357 17187 13415 17193
rect 13357 17184 13369 17187
rect 12759 17156 13369 17184
rect 12759 17153 12771 17156
rect 12713 17147 12771 17153
rect 13357 17153 13369 17156
rect 13403 17153 13415 17187
rect 13357 17147 13415 17153
rect 14277 17187 14335 17193
rect 14277 17153 14289 17187
rect 14323 17184 14335 17187
rect 14458 17184 14464 17196
rect 14323 17156 14464 17184
rect 14323 17153 14335 17156
rect 14277 17147 14335 17153
rect 14458 17144 14464 17156
rect 14516 17184 14522 17196
rect 14734 17184 14740 17196
rect 14516 17156 14740 17184
rect 14516 17144 14522 17156
rect 14734 17144 14740 17156
rect 14792 17144 14798 17196
rect 15289 17187 15347 17193
rect 15289 17153 15301 17187
rect 15335 17184 15347 17187
rect 15933 17187 15991 17193
rect 15933 17184 15945 17187
rect 15335 17156 15945 17184
rect 15335 17153 15347 17156
rect 15289 17147 15347 17153
rect 15933 17153 15945 17156
rect 15979 17153 15991 17187
rect 16666 17184 16672 17196
rect 16627 17156 16672 17184
rect 15933 17147 15991 17153
rect 16666 17144 16672 17156
rect 16724 17144 16730 17196
rect 18138 17144 18144 17196
rect 18196 17184 18202 17196
rect 19168 17193 19196 17224
rect 19812 17224 20576 17252
rect 18693 17187 18751 17193
rect 18693 17184 18705 17187
rect 18196 17156 18705 17184
rect 18196 17144 18202 17156
rect 18693 17153 18705 17156
rect 18739 17153 18751 17187
rect 18693 17147 18751 17153
rect 19153 17187 19211 17193
rect 19153 17153 19165 17187
rect 19199 17153 19211 17187
rect 19153 17147 19211 17153
rect 19429 17187 19487 17193
rect 19429 17153 19441 17187
rect 19475 17184 19487 17187
rect 19518 17184 19524 17196
rect 19475 17156 19524 17184
rect 19475 17153 19487 17156
rect 19429 17147 19487 17153
rect 19518 17144 19524 17156
rect 19576 17144 19582 17196
rect 2961 17119 3019 17125
rect 2961 17085 2973 17119
rect 3007 17116 3019 17119
rect 3418 17116 3424 17128
rect 3007 17088 3424 17116
rect 3007 17085 3019 17088
rect 2961 17079 3019 17085
rect 3418 17076 3424 17088
rect 3476 17076 3482 17128
rect 3878 17116 3884 17128
rect 3839 17088 3884 17116
rect 3878 17076 3884 17088
rect 3936 17076 3942 17128
rect 9766 17076 9772 17128
rect 9824 17116 9830 17128
rect 10137 17119 10195 17125
rect 10137 17116 10149 17119
rect 9824 17088 10149 17116
rect 9824 17076 9830 17088
rect 10137 17085 10149 17088
rect 10183 17085 10195 17119
rect 10137 17079 10195 17085
rect 12434 17076 12440 17128
rect 12492 17116 12498 17128
rect 12492 17088 12537 17116
rect 12492 17076 12498 17088
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 14001 17119 14059 17125
rect 14001 17116 14013 17119
rect 13872 17088 14013 17116
rect 13872 17076 13878 17088
rect 14001 17085 14013 17088
rect 14047 17085 14059 17119
rect 14001 17079 14059 17085
rect 15105 17119 15163 17125
rect 15105 17085 15117 17119
rect 15151 17116 15163 17119
rect 15470 17116 15476 17128
rect 15151 17088 15476 17116
rect 15151 17085 15163 17088
rect 15105 17079 15163 17085
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 19812 17116 19840 17224
rect 20548 17193 20576 17224
rect 19889 17187 19947 17193
rect 19889 17153 19901 17187
rect 19935 17184 19947 17187
rect 20533 17187 20591 17193
rect 19935 17156 20392 17184
rect 19935 17153 19947 17156
rect 19889 17147 19947 17153
rect 15580 17088 19840 17116
rect 7558 17008 7564 17060
rect 7616 17048 7622 17060
rect 15378 17048 15384 17060
rect 7616 17020 15384 17048
rect 7616 17008 7622 17020
rect 15378 17008 15384 17020
rect 15436 17008 15442 17060
rect 1578 16980 1584 16992
rect 1539 16952 1584 16980
rect 1578 16940 1584 16952
rect 1636 16940 1642 16992
rect 2958 16940 2964 16992
rect 3016 16980 3022 16992
rect 3237 16983 3295 16989
rect 3237 16980 3249 16983
rect 3016 16952 3249 16980
rect 3016 16940 3022 16952
rect 3237 16949 3249 16952
rect 3283 16949 3295 16983
rect 8662 16980 8668 16992
rect 8623 16952 8668 16980
rect 3237 16943 3295 16949
rect 8662 16940 8668 16952
rect 8720 16940 8726 16992
rect 9858 16980 9864 16992
rect 9819 16952 9864 16980
rect 9858 16940 9864 16952
rect 9916 16940 9922 16992
rect 13081 16983 13139 16989
rect 13081 16949 13093 16983
rect 13127 16980 13139 16983
rect 15580 16980 15608 17088
rect 19610 17048 19616 17060
rect 17144 17020 19616 17048
rect 13127 16952 15608 16980
rect 15657 16983 15715 16989
rect 13127 16949 13139 16952
rect 13081 16943 13139 16949
rect 15657 16949 15669 16983
rect 15703 16980 15715 16983
rect 17144 16980 17172 17020
rect 19610 17008 19616 17020
rect 19668 17008 19674 17060
rect 20364 17057 20392 17156
rect 20533 17153 20545 17187
rect 20579 17153 20591 17187
rect 21082 17184 21088 17196
rect 21043 17156 21088 17184
rect 20533 17147 20591 17153
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 20349 17051 20407 17057
rect 20349 17017 20361 17051
rect 20395 17017 20407 17051
rect 20349 17011 20407 17017
rect 17310 16980 17316 16992
rect 15703 16952 17172 16980
rect 17271 16952 17316 16980
rect 15703 16949 15715 16952
rect 15657 16943 15715 16949
rect 17310 16940 17316 16952
rect 17368 16940 17374 16992
rect 17770 16940 17776 16992
rect 17828 16980 17834 16992
rect 18049 16983 18107 16989
rect 18049 16980 18061 16983
rect 17828 16952 18061 16980
rect 17828 16940 17834 16952
rect 18049 16949 18061 16952
rect 18095 16949 18107 16983
rect 18049 16943 18107 16949
rect 18322 16940 18328 16992
rect 18380 16980 18386 16992
rect 21174 16980 21180 16992
rect 18380 16952 21180 16980
rect 18380 16940 18386 16952
rect 21174 16940 21180 16952
rect 21232 16940 21238 16992
rect 21269 16983 21327 16989
rect 21269 16949 21281 16983
rect 21315 16980 21327 16983
rect 21358 16980 21364 16992
rect 21315 16952 21364 16980
rect 21315 16949 21327 16952
rect 21269 16943 21327 16949
rect 21358 16940 21364 16952
rect 21416 16940 21422 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 5718 16776 5724 16788
rect 4540 16748 5724 16776
rect 1578 16600 1584 16652
rect 1636 16640 1642 16652
rect 2777 16643 2835 16649
rect 2777 16640 2789 16643
rect 1636 16612 2789 16640
rect 1636 16600 1642 16612
rect 2777 16609 2789 16612
rect 2823 16609 2835 16643
rect 2958 16640 2964 16652
rect 2919 16612 2964 16640
rect 2777 16603 2835 16609
rect 2958 16600 2964 16612
rect 3016 16600 3022 16652
rect 3418 16600 3424 16652
rect 3476 16640 3482 16652
rect 4540 16649 4568 16748
rect 5718 16736 5724 16748
rect 5776 16736 5782 16788
rect 14826 16776 14832 16788
rect 12360 16748 14832 16776
rect 5810 16668 5816 16720
rect 5868 16708 5874 16720
rect 5868 16680 8156 16708
rect 5868 16668 5874 16680
rect 8128 16649 8156 16680
rect 4525 16643 4583 16649
rect 4525 16640 4537 16643
rect 3476 16612 4537 16640
rect 3476 16600 3482 16612
rect 4525 16609 4537 16612
rect 4571 16609 4583 16643
rect 4525 16603 4583 16609
rect 7929 16643 7987 16649
rect 7929 16609 7941 16643
rect 7975 16609 7987 16643
rect 7929 16603 7987 16609
rect 8113 16643 8171 16649
rect 8113 16609 8125 16643
rect 8159 16609 8171 16643
rect 9214 16640 9220 16652
rect 9175 16612 9220 16640
rect 8113 16603 8171 16609
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16572 3111 16575
rect 3142 16572 3148 16584
rect 3099 16544 3148 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 3142 16532 3148 16544
rect 3200 16532 3206 16584
rect 4798 16581 4804 16584
rect 3789 16575 3847 16581
rect 3789 16541 3801 16575
rect 3835 16541 3847 16575
rect 3789 16535 3847 16541
rect 4792 16535 4804 16581
rect 4856 16572 4862 16584
rect 6181 16575 6239 16581
rect 6181 16572 6193 16575
rect 4856 16544 4892 16572
rect 5920 16544 6193 16572
rect 3421 16439 3479 16445
rect 3421 16405 3433 16439
rect 3467 16436 3479 16439
rect 3804 16436 3832 16535
rect 4798 16532 4804 16535
rect 4856 16532 4862 16544
rect 3467 16408 3832 16436
rect 3973 16439 4031 16445
rect 3467 16405 3479 16408
rect 3421 16399 3479 16405
rect 3973 16405 3985 16439
rect 4019 16436 4031 16439
rect 4062 16436 4068 16448
rect 4019 16408 4068 16436
rect 4019 16405 4031 16408
rect 3973 16399 4031 16405
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 5920 16445 5948 16544
rect 6181 16541 6193 16544
rect 6227 16572 6239 16575
rect 7944 16572 7972 16603
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 9950 16640 9956 16652
rect 9646 16612 9956 16640
rect 6227 16544 7972 16572
rect 8205 16575 8263 16581
rect 6227 16541 6239 16544
rect 6181 16535 6239 16541
rect 8205 16541 8217 16575
rect 8251 16572 8263 16575
rect 8662 16572 8668 16584
rect 8251 16544 8668 16572
rect 8251 16541 8263 16544
rect 8205 16535 8263 16541
rect 8662 16532 8668 16544
rect 8720 16572 8726 16584
rect 9646 16572 9674 16612
rect 9950 16600 9956 16612
rect 10008 16640 10014 16652
rect 10226 16640 10232 16652
rect 10008 16612 10232 16640
rect 10008 16600 10014 16612
rect 10226 16600 10232 16612
rect 10284 16600 10290 16652
rect 10594 16600 10600 16652
rect 10652 16640 10658 16652
rect 12360 16649 12388 16748
rect 14108 16649 14136 16748
rect 14826 16736 14832 16748
rect 14884 16776 14890 16788
rect 15654 16776 15660 16788
rect 14884 16748 15660 16776
rect 14884 16736 14890 16748
rect 15654 16736 15660 16748
rect 15712 16776 15718 16788
rect 16390 16776 16396 16788
rect 15712 16748 16396 16776
rect 15712 16736 15718 16748
rect 16390 16736 16396 16748
rect 16448 16736 16454 16788
rect 20809 16779 20867 16785
rect 20809 16745 20821 16779
rect 20855 16776 20867 16779
rect 21082 16776 21088 16788
rect 20855 16748 21088 16776
rect 20855 16745 20867 16748
rect 20809 16739 20867 16745
rect 21082 16736 21088 16748
rect 21140 16736 21146 16788
rect 15470 16708 15476 16720
rect 15431 16680 15476 16708
rect 15470 16668 15476 16680
rect 15528 16668 15534 16720
rect 17221 16711 17279 16717
rect 17221 16677 17233 16711
rect 17267 16708 17279 16711
rect 17267 16680 18276 16708
rect 17267 16677 17279 16680
rect 17221 16671 17279 16677
rect 10689 16643 10747 16649
rect 10689 16640 10701 16643
rect 10652 16612 10701 16640
rect 10652 16600 10658 16612
rect 10689 16609 10701 16612
rect 10735 16609 10747 16643
rect 10689 16603 10747 16609
rect 12345 16643 12403 16649
rect 12345 16609 12357 16643
rect 12391 16609 12403 16643
rect 12345 16603 12403 16609
rect 14093 16643 14151 16649
rect 14093 16609 14105 16643
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 15378 16600 15384 16652
rect 15436 16640 15442 16652
rect 16666 16640 16672 16652
rect 15436 16612 16528 16640
rect 16579 16612 16672 16640
rect 15436 16600 15442 16612
rect 8720 16544 9674 16572
rect 10137 16575 10195 16581
rect 8720 16532 8726 16544
rect 10137 16541 10149 16575
rect 10183 16541 10195 16575
rect 16500 16572 16528 16612
rect 16666 16600 16672 16612
rect 16724 16640 16730 16652
rect 17034 16640 17040 16652
rect 16724 16612 17040 16640
rect 16724 16600 16730 16612
rect 17034 16600 17040 16612
rect 17092 16600 17098 16652
rect 18138 16640 18144 16652
rect 18099 16612 18144 16640
rect 18138 16600 18144 16612
rect 18196 16600 18202 16652
rect 18248 16649 18276 16680
rect 18233 16643 18291 16649
rect 18233 16609 18245 16643
rect 18279 16609 18291 16643
rect 18233 16603 18291 16609
rect 16761 16575 16819 16581
rect 16761 16572 16773 16575
rect 16500 16544 16773 16572
rect 10137 16535 10195 16541
rect 16761 16541 16773 16544
rect 16807 16541 16819 16575
rect 16761 16535 16819 16541
rect 9493 16507 9551 16513
rect 9493 16473 9505 16507
rect 9539 16504 9551 16507
rect 9766 16504 9772 16516
rect 9539 16476 9772 16504
rect 9539 16473 9551 16476
rect 9493 16467 9551 16473
rect 9766 16464 9772 16476
rect 9824 16464 9830 16516
rect 5905 16439 5963 16445
rect 5905 16405 5917 16439
rect 5951 16405 5963 16439
rect 6822 16436 6828 16448
rect 6783 16408 6828 16436
rect 5905 16399 5963 16405
rect 6822 16396 6828 16408
rect 6880 16396 6886 16448
rect 8573 16439 8631 16445
rect 8573 16405 8585 16439
rect 8619 16436 8631 16439
rect 9401 16439 9459 16445
rect 9401 16436 9413 16439
rect 8619 16408 9413 16436
rect 8619 16405 8631 16408
rect 8573 16399 8631 16405
rect 9401 16405 9413 16408
rect 9447 16405 9459 16439
rect 9401 16399 9459 16405
rect 9861 16439 9919 16445
rect 9861 16405 9873 16439
rect 9907 16436 9919 16439
rect 10152 16436 10180 16535
rect 18414 16532 18420 16584
rect 18472 16572 18478 16584
rect 19889 16575 19947 16581
rect 19889 16572 19901 16575
rect 18472 16544 19901 16572
rect 18472 16532 18478 16544
rect 19889 16541 19901 16544
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 20070 16532 20076 16584
rect 20128 16572 20134 16584
rect 20165 16575 20223 16581
rect 20165 16572 20177 16575
rect 20128 16544 20177 16572
rect 20128 16532 20134 16544
rect 20165 16541 20177 16544
rect 20211 16541 20223 16575
rect 20165 16535 20223 16541
rect 20625 16575 20683 16581
rect 20625 16541 20637 16575
rect 20671 16541 20683 16575
rect 21082 16572 21088 16584
rect 21043 16544 21088 16572
rect 20625 16535 20683 16541
rect 10956 16507 11014 16513
rect 10956 16473 10968 16507
rect 11002 16504 11014 16507
rect 11146 16504 11152 16516
rect 11002 16476 11152 16504
rect 11002 16473 11014 16476
rect 10956 16467 11014 16473
rect 11146 16464 11152 16476
rect 11204 16464 11210 16516
rect 12612 16507 12670 16513
rect 12612 16473 12624 16507
rect 12658 16504 12670 16507
rect 12710 16504 12716 16516
rect 12658 16476 12716 16504
rect 12658 16473 12670 16476
rect 12612 16467 12670 16473
rect 12710 16464 12716 16476
rect 12768 16464 12774 16516
rect 14366 16513 14372 16516
rect 14360 16467 14372 16513
rect 14424 16504 14430 16516
rect 18325 16507 18383 16513
rect 14424 16476 14460 16504
rect 14366 16464 14372 16467
rect 14424 16464 14430 16476
rect 18325 16473 18337 16507
rect 18371 16504 18383 16507
rect 19245 16507 19303 16513
rect 19245 16504 19257 16507
rect 18371 16476 19257 16504
rect 18371 16473 18383 16476
rect 18325 16467 18383 16473
rect 19245 16473 19257 16476
rect 19291 16473 19303 16507
rect 19245 16467 19303 16473
rect 19334 16464 19340 16516
rect 19392 16504 19398 16516
rect 20640 16504 20668 16535
rect 21082 16532 21088 16544
rect 21140 16532 21146 16584
rect 19392 16476 20668 16504
rect 19392 16464 19398 16476
rect 9907 16408 10180 16436
rect 10321 16439 10379 16445
rect 9907 16405 9919 16408
rect 9861 16399 9919 16405
rect 10321 16405 10333 16439
rect 10367 16436 10379 16439
rect 10410 16436 10416 16448
rect 10367 16408 10416 16436
rect 10367 16405 10379 16408
rect 10321 16399 10379 16405
rect 10410 16396 10416 16408
rect 10468 16396 10474 16448
rect 12069 16439 12127 16445
rect 12069 16405 12081 16439
rect 12115 16436 12127 16439
rect 12434 16436 12440 16448
rect 12115 16408 12440 16436
rect 12115 16405 12127 16408
rect 12069 16399 12127 16405
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 13725 16439 13783 16445
rect 13725 16405 13737 16439
rect 13771 16436 13783 16439
rect 13814 16436 13820 16448
rect 13771 16408 13820 16436
rect 13771 16405 13783 16408
rect 13725 16399 13783 16405
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 16853 16439 16911 16445
rect 16853 16405 16865 16439
rect 16899 16436 16911 16439
rect 16942 16436 16948 16448
rect 16899 16408 16948 16436
rect 16899 16405 16911 16408
rect 16853 16399 16911 16405
rect 16942 16396 16948 16408
rect 17000 16436 17006 16448
rect 17497 16439 17555 16445
rect 17497 16436 17509 16439
rect 17000 16408 17509 16436
rect 17000 16396 17006 16408
rect 17497 16405 17509 16408
rect 17543 16405 17555 16439
rect 17497 16399 17555 16405
rect 18693 16439 18751 16445
rect 18693 16405 18705 16439
rect 18739 16436 18751 16439
rect 19518 16436 19524 16448
rect 18739 16408 19524 16436
rect 18739 16405 18751 16408
rect 18693 16399 18751 16405
rect 19518 16396 19524 16408
rect 19576 16396 19582 16448
rect 19702 16436 19708 16448
rect 19663 16408 19708 16436
rect 19702 16396 19708 16408
rect 19760 16396 19766 16448
rect 20346 16436 20352 16448
rect 20307 16408 20352 16436
rect 20346 16396 20352 16408
rect 20404 16396 20410 16448
rect 21266 16436 21272 16448
rect 21227 16408 21272 16436
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 21450 16396 21456 16448
rect 21508 16436 21514 16448
rect 21726 16436 21732 16448
rect 21508 16408 21732 16436
rect 21508 16396 21514 16408
rect 21726 16396 21732 16408
rect 21784 16396 21790 16448
rect 1104 16346 21896 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21896 16346
rect 1104 16272 21896 16294
rect 4062 16192 4068 16244
rect 4120 16232 4126 16244
rect 9214 16232 9220 16244
rect 4120 16204 9076 16232
rect 9175 16204 9220 16232
rect 4120 16192 4126 16204
rect 3418 16164 3424 16176
rect 1780 16136 3424 16164
rect 1780 16105 1808 16136
rect 3418 16124 3424 16136
rect 3476 16124 3482 16176
rect 6822 16124 6828 16176
rect 6880 16164 6886 16176
rect 8082 16167 8140 16173
rect 8082 16164 8094 16167
rect 6880 16136 8094 16164
rect 6880 16124 6886 16136
rect 8082 16133 8094 16136
rect 8128 16133 8140 16167
rect 9048 16164 9076 16204
rect 9214 16192 9220 16204
rect 9272 16192 9278 16244
rect 12710 16232 12716 16244
rect 9416 16204 12434 16232
rect 12671 16204 12716 16232
rect 9416 16164 9444 16204
rect 10594 16164 10600 16176
rect 9048 16136 9444 16164
rect 9784 16136 10600 16164
rect 8082 16127 8140 16133
rect 2038 16105 2044 16108
rect 1765 16099 1823 16105
rect 1765 16065 1777 16099
rect 1811 16065 1823 16099
rect 1765 16059 1823 16065
rect 2032 16059 2044 16105
rect 2096 16096 2102 16108
rect 4065 16099 4123 16105
rect 2096 16068 2132 16096
rect 2038 16056 2044 16059
rect 2096 16056 2102 16068
rect 4065 16065 4077 16099
rect 4111 16065 4123 16099
rect 4065 16059 4123 16065
rect 3326 15988 3332 16040
rect 3384 16028 3390 16040
rect 3421 16031 3479 16037
rect 3421 16028 3433 16031
rect 3384 16000 3433 16028
rect 3384 15988 3390 16000
rect 3421 15997 3433 16000
rect 3467 15997 3479 16031
rect 3421 15991 3479 15997
rect 3145 15963 3203 15969
rect 3145 15929 3157 15963
rect 3191 15960 3203 15963
rect 3878 15960 3884 15972
rect 3191 15932 3884 15960
rect 3191 15929 3203 15932
rect 3145 15923 3203 15929
rect 3878 15920 3884 15932
rect 3936 15960 3942 15972
rect 4080 15960 4108 16059
rect 6914 16056 6920 16108
rect 6972 16096 6978 16108
rect 9784 16105 9812 16136
rect 10594 16124 10600 16136
rect 10652 16124 10658 16176
rect 12406 16164 12434 16204
rect 12710 16192 12716 16204
rect 12768 16192 12774 16244
rect 14366 16232 14372 16244
rect 14327 16204 14372 16232
rect 14366 16192 14372 16204
rect 14424 16192 14430 16244
rect 16301 16235 16359 16241
rect 16301 16201 16313 16235
rect 16347 16232 16359 16235
rect 17034 16232 17040 16244
rect 16347 16204 17040 16232
rect 16347 16201 16359 16204
rect 16301 16195 16359 16201
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 18049 16235 18107 16241
rect 18049 16201 18061 16235
rect 18095 16232 18107 16235
rect 18138 16232 18144 16244
rect 18095 16204 18144 16232
rect 18095 16201 18107 16204
rect 18049 16195 18107 16201
rect 18138 16192 18144 16204
rect 18196 16192 18202 16244
rect 19429 16235 19487 16241
rect 19429 16201 19441 16235
rect 19475 16232 19487 16235
rect 19794 16232 19800 16244
rect 19475 16204 19800 16232
rect 19475 16201 19487 16204
rect 19429 16195 19487 16201
rect 19794 16192 19800 16204
rect 19852 16192 19858 16244
rect 20070 16232 20076 16244
rect 20031 16204 20076 16232
rect 20070 16192 20076 16204
rect 20128 16192 20134 16244
rect 20162 16192 20168 16244
rect 20220 16232 20226 16244
rect 20625 16235 20683 16241
rect 20625 16232 20637 16235
rect 20220 16204 20637 16232
rect 20220 16192 20226 16204
rect 20625 16201 20637 16204
rect 20671 16201 20683 16235
rect 20625 16195 20683 16201
rect 20714 16192 20720 16244
rect 20772 16232 20778 16244
rect 20898 16232 20904 16244
rect 20772 16204 20904 16232
rect 20772 16192 20778 16204
rect 20898 16192 20904 16204
rect 20956 16192 20962 16244
rect 16936 16167 16994 16173
rect 12406 16136 16804 16164
rect 9769 16099 9827 16105
rect 6972 16068 7017 16096
rect 6972 16056 6978 16068
rect 9769 16065 9781 16099
rect 9815 16065 9827 16099
rect 9769 16059 9827 16065
rect 9858 16056 9864 16108
rect 9916 16096 9922 16108
rect 10025 16099 10083 16105
rect 10025 16096 10037 16099
rect 9916 16068 10037 16096
rect 9916 16056 9922 16068
rect 10025 16065 10037 16068
rect 10071 16065 10083 16099
rect 10025 16059 10083 16065
rect 12069 16099 12127 16105
rect 12069 16065 12081 16099
rect 12115 16096 12127 16099
rect 12434 16096 12440 16108
rect 12115 16068 12440 16096
rect 12115 16065 12127 16068
rect 12069 16059 12127 16065
rect 12434 16056 12440 16068
rect 12492 16056 12498 16108
rect 13725 16099 13783 16105
rect 13725 16065 13737 16099
rect 13771 16096 13783 16099
rect 13814 16096 13820 16108
rect 13771 16068 13820 16096
rect 13771 16065 13783 16068
rect 13725 16059 13783 16065
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 14826 16056 14832 16108
rect 14884 16096 14890 16108
rect 14921 16099 14979 16105
rect 14921 16096 14933 16099
rect 14884 16068 14933 16096
rect 14884 16056 14890 16068
rect 14921 16065 14933 16068
rect 14967 16065 14979 16099
rect 14921 16059 14979 16065
rect 15188 16099 15246 16105
rect 15188 16065 15200 16099
rect 15234 16096 15246 16099
rect 16114 16096 16120 16108
rect 15234 16068 16120 16096
rect 15234 16065 15246 16068
rect 15188 16059 15246 16065
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 16574 16056 16580 16108
rect 16632 16096 16638 16108
rect 16669 16099 16727 16105
rect 16669 16096 16681 16099
rect 16632 16068 16681 16096
rect 16632 16056 16638 16068
rect 16669 16065 16681 16068
rect 16715 16065 16727 16099
rect 16776 16096 16804 16136
rect 16936 16133 16948 16167
rect 16982 16164 16994 16167
rect 17310 16164 17316 16176
rect 16982 16136 17316 16164
rect 16982 16133 16994 16136
rect 16936 16127 16994 16133
rect 17310 16124 17316 16136
rect 17368 16124 17374 16176
rect 19334 16096 19340 16108
rect 16776 16068 19340 16096
rect 16669 16059 16727 16065
rect 19334 16056 19340 16068
rect 19392 16056 19398 16108
rect 19610 16096 19616 16108
rect 19571 16068 19616 16096
rect 19610 16056 19616 16068
rect 19668 16056 19674 16108
rect 19889 16099 19947 16105
rect 19889 16065 19901 16099
rect 19935 16065 19947 16099
rect 19889 16059 19947 16065
rect 6733 16031 6791 16037
rect 6733 15997 6745 16031
rect 6779 15997 6791 16031
rect 6733 15991 6791 15997
rect 6825 16031 6883 16037
rect 6825 15997 6837 16031
rect 6871 16028 6883 16031
rect 7006 16028 7012 16040
rect 6871 16000 7012 16028
rect 6871 15997 6883 16000
rect 6825 15991 6883 15997
rect 3936 15932 4108 15960
rect 6748 15960 6776 15991
rect 7006 15988 7012 16000
rect 7064 15988 7070 16040
rect 7282 15988 7288 16040
rect 7340 16028 7346 16040
rect 7837 16031 7895 16037
rect 7837 16028 7849 16031
rect 7340 16000 7849 16028
rect 7340 15988 7346 16000
rect 7837 15997 7849 16000
rect 7883 15997 7895 16031
rect 7837 15991 7895 15997
rect 7098 15960 7104 15972
rect 6748 15932 7104 15960
rect 3936 15920 3942 15932
rect 7098 15920 7104 15932
rect 7156 15920 7162 15972
rect 11149 15963 11207 15969
rect 11149 15929 11161 15963
rect 11195 15960 11207 15963
rect 11238 15960 11244 15972
rect 11195 15932 11244 15960
rect 11195 15929 11207 15932
rect 11149 15923 11207 15929
rect 11238 15920 11244 15932
rect 11296 15920 11302 15972
rect 19904 15960 19932 16059
rect 19978 16056 19984 16108
rect 20036 16096 20042 16108
rect 20809 16099 20867 16105
rect 20809 16096 20821 16099
rect 20036 16068 20821 16096
rect 20036 16056 20042 16068
rect 20809 16065 20821 16068
rect 20855 16065 20867 16099
rect 20809 16059 20867 16065
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 20956 16068 21097 16096
rect 20956 16056 20962 16068
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 17604 15932 19932 15960
rect 7285 15895 7343 15901
rect 7285 15861 7297 15895
rect 7331 15892 7343 15895
rect 17604 15892 17632 15932
rect 7331 15864 17632 15892
rect 21269 15895 21327 15901
rect 7331 15861 7343 15864
rect 7285 15855 7343 15861
rect 21269 15861 21281 15895
rect 21315 15892 21327 15895
rect 21358 15892 21364 15904
rect 21315 15864 21364 15892
rect 21315 15861 21327 15864
rect 21269 15855 21327 15861
rect 21358 15852 21364 15864
rect 21416 15852 21422 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 2038 15648 2044 15700
rect 2096 15688 2102 15700
rect 2225 15691 2283 15697
rect 2225 15688 2237 15691
rect 2096 15660 2237 15688
rect 2096 15648 2102 15660
rect 2225 15657 2237 15660
rect 2271 15657 2283 15691
rect 5718 15688 5724 15700
rect 5679 15660 5724 15688
rect 2225 15651 2283 15657
rect 5718 15648 5724 15660
rect 5776 15648 5782 15700
rect 8110 15648 8116 15700
rect 8168 15688 8174 15700
rect 8389 15691 8447 15697
rect 8389 15688 8401 15691
rect 8168 15660 8401 15688
rect 8168 15648 8174 15660
rect 8389 15657 8401 15660
rect 8435 15657 8447 15691
rect 11146 15688 11152 15700
rect 11107 15660 11152 15688
rect 8389 15651 8447 15657
rect 11146 15648 11152 15660
rect 11204 15648 11210 15700
rect 16114 15688 16120 15700
rect 16075 15660 16120 15688
rect 16114 15648 16120 15660
rect 16172 15648 16178 15700
rect 19978 15688 19984 15700
rect 16592 15660 19984 15688
rect 7926 15580 7932 15632
rect 7984 15620 7990 15632
rect 16592 15620 16620 15660
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 20349 15691 20407 15697
rect 20349 15657 20361 15691
rect 20395 15688 20407 15691
rect 21082 15688 21088 15700
rect 20395 15660 21088 15688
rect 20395 15657 20407 15660
rect 20349 15651 20407 15657
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 7984 15592 16620 15620
rect 19889 15623 19947 15629
rect 7984 15580 7990 15592
rect 19889 15589 19901 15623
rect 19935 15620 19947 15623
rect 20714 15620 20720 15632
rect 19935 15592 20720 15620
rect 19935 15589 19947 15592
rect 19889 15583 19947 15589
rect 20714 15580 20720 15592
rect 20772 15580 20778 15632
rect 20809 15623 20867 15629
rect 20809 15589 20821 15623
rect 20855 15620 20867 15623
rect 20990 15620 20996 15632
rect 20855 15592 20996 15620
rect 20855 15589 20867 15592
rect 20809 15583 20867 15589
rect 20990 15580 20996 15592
rect 21048 15580 21054 15632
rect 3881 15555 3939 15561
rect 3881 15521 3893 15555
rect 3927 15521 3939 15555
rect 3881 15515 3939 15521
rect 2866 15484 2872 15496
rect 2827 15456 2872 15484
rect 2866 15444 2872 15456
rect 2924 15484 2930 15496
rect 3896 15484 3924 15515
rect 6914 15512 6920 15564
rect 6972 15552 6978 15564
rect 7285 15555 7343 15561
rect 7285 15552 7297 15555
rect 6972 15524 7297 15552
rect 6972 15512 6978 15524
rect 7285 15521 7297 15524
rect 7331 15521 7343 15555
rect 7285 15515 7343 15521
rect 16574 15512 16580 15564
rect 16632 15552 16638 15564
rect 17310 15552 17316 15564
rect 16632 15524 17316 15552
rect 16632 15512 16638 15524
rect 17310 15512 17316 15524
rect 17368 15552 17374 15564
rect 17497 15555 17555 15561
rect 17497 15552 17509 15555
rect 17368 15524 17509 15552
rect 17368 15512 17374 15524
rect 17497 15521 17509 15524
rect 17543 15521 17555 15555
rect 17497 15515 17555 15521
rect 7742 15484 7748 15496
rect 2924 15456 3924 15484
rect 7703 15456 7748 15484
rect 2924 15444 2930 15456
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 11238 15444 11244 15496
rect 11296 15484 11302 15496
rect 11793 15487 11851 15493
rect 11793 15484 11805 15487
rect 11296 15456 11805 15484
rect 11296 15444 11302 15456
rect 11793 15453 11805 15456
rect 11839 15453 11851 15487
rect 15470 15484 15476 15496
rect 15431 15456 15476 15484
rect 11793 15447 11851 15453
rect 15470 15444 15476 15456
rect 15528 15444 15534 15496
rect 17770 15493 17776 15496
rect 17764 15484 17776 15493
rect 17731 15456 17776 15484
rect 17764 15447 17776 15456
rect 17770 15444 17776 15447
rect 17828 15444 17834 15496
rect 19705 15487 19763 15493
rect 19705 15453 19717 15487
rect 19751 15453 19763 15487
rect 20162 15484 20168 15496
rect 20123 15456 20168 15484
rect 19705 15447 19763 15453
rect 4157 15419 4215 15425
rect 4157 15385 4169 15419
rect 4203 15416 4215 15419
rect 4801 15419 4859 15425
rect 4801 15416 4813 15419
rect 4203 15388 4813 15416
rect 4203 15385 4215 15388
rect 4157 15379 4215 15385
rect 4801 15385 4813 15388
rect 4847 15385 4859 15419
rect 4801 15379 4859 15385
rect 7009 15419 7067 15425
rect 7009 15385 7021 15419
rect 7055 15416 7067 15419
rect 10318 15416 10324 15428
rect 7055 15388 10324 15416
rect 7055 15385 7067 15388
rect 7009 15379 7067 15385
rect 10318 15376 10324 15388
rect 10376 15376 10382 15428
rect 10410 15376 10416 15428
rect 10468 15416 10474 15428
rect 19720 15416 19748 15447
rect 20162 15444 20168 15456
rect 20220 15444 20226 15496
rect 20622 15484 20628 15496
rect 20583 15456 20628 15484
rect 20622 15444 20628 15456
rect 20680 15444 20686 15496
rect 21082 15484 21088 15496
rect 21043 15456 21088 15484
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 10468 15388 19748 15416
rect 10468 15376 10474 15388
rect 4065 15351 4123 15357
rect 4065 15317 4077 15351
rect 4111 15348 4123 15351
rect 4246 15348 4252 15360
rect 4111 15320 4252 15348
rect 4111 15317 4123 15320
rect 4065 15311 4123 15317
rect 4246 15308 4252 15320
rect 4304 15308 4310 15360
rect 4525 15351 4583 15357
rect 4525 15317 4537 15351
rect 4571 15348 4583 15351
rect 5442 15348 5448 15360
rect 4571 15320 5448 15348
rect 4571 15317 4583 15320
rect 4525 15311 4583 15317
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 18874 15348 18880 15360
rect 18835 15320 18880 15348
rect 18874 15308 18880 15320
rect 18932 15308 18938 15360
rect 21266 15348 21272 15360
rect 21227 15320 21272 15348
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 1104 15258 21896 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21896 15258
rect 1104 15184 21896 15206
rect 2133 15147 2191 15153
rect 2133 15113 2145 15147
rect 2179 15144 2191 15147
rect 2866 15144 2872 15156
rect 2179 15116 2872 15144
rect 2179 15113 2191 15116
rect 2133 15107 2191 15113
rect 2866 15104 2872 15116
rect 2924 15104 2930 15156
rect 4157 15147 4215 15153
rect 4157 15113 4169 15147
rect 4203 15144 4215 15147
rect 4246 15144 4252 15156
rect 4203 15116 4252 15144
rect 4203 15113 4215 15116
rect 4157 15107 4215 15113
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 7742 15144 7748 15156
rect 7703 15116 7748 15144
rect 7742 15104 7748 15116
rect 7800 15104 7806 15156
rect 20162 15104 20168 15156
rect 20220 15144 20226 15156
rect 20257 15147 20315 15153
rect 20257 15144 20269 15147
rect 20220 15116 20269 15144
rect 20220 15104 20226 15116
rect 20257 15113 20269 15116
rect 20303 15113 20315 15147
rect 20257 15107 20315 15113
rect 20809 15147 20867 15153
rect 20809 15113 20821 15147
rect 20855 15144 20867 15147
rect 20898 15144 20904 15156
rect 20855 15116 20904 15144
rect 20855 15113 20867 15116
rect 20809 15107 20867 15113
rect 20898 15104 20904 15116
rect 20956 15104 20962 15156
rect 2498 15036 2504 15088
rect 2556 15076 2562 15088
rect 4617 15079 4675 15085
rect 4617 15076 4629 15079
rect 2556 15048 4629 15076
rect 2556 15036 2562 15048
rect 4617 15045 4629 15048
rect 4663 15045 4675 15079
rect 4617 15039 4675 15045
rect 5442 15036 5448 15088
rect 5500 15076 5506 15088
rect 5500 15048 20116 15076
rect 5500 15036 5506 15048
rect 3234 15008 3240 15020
rect 3292 15017 3298 15020
rect 3204 14980 3240 15008
rect 3234 14968 3240 14980
rect 3292 14971 3304 15017
rect 3292 14968 3298 14971
rect 3418 14968 3424 15020
rect 3476 15008 3482 15020
rect 6638 15017 6644 15020
rect 3513 15011 3571 15017
rect 3513 15008 3525 15011
rect 3476 14980 3525 15008
rect 3476 14968 3482 14980
rect 3513 14977 3525 14980
rect 3559 14977 3571 15011
rect 3513 14971 3571 14977
rect 4525 15011 4583 15017
rect 4525 14977 4537 15011
rect 4571 15008 4583 15011
rect 4571 14980 5304 15008
rect 4571 14977 4583 14980
rect 4525 14971 4583 14977
rect 4709 14943 4767 14949
rect 4709 14909 4721 14943
rect 4755 14909 4767 14943
rect 4709 14903 4767 14909
rect 4430 14832 4436 14884
rect 4488 14872 4494 14884
rect 4724 14872 4752 14903
rect 4488 14844 4752 14872
rect 4488 14832 4494 14844
rect 5276 14816 5304 14980
rect 6632 14971 6644 15017
rect 6696 15008 6702 15020
rect 8662 15008 8668 15020
rect 6696 14980 6732 15008
rect 8623 14980 8668 15008
rect 6638 14968 6644 14971
rect 6696 14968 6702 14980
rect 8662 14968 8668 14980
rect 8720 14968 8726 15020
rect 9401 15011 9459 15017
rect 9401 14977 9413 15011
rect 9447 15008 9459 15011
rect 9674 15008 9680 15020
rect 9447 14980 9680 15008
rect 9447 14977 9459 14980
rect 9401 14971 9459 14977
rect 9674 14968 9680 14980
rect 9732 14968 9738 15020
rect 12805 15011 12863 15017
rect 12805 14977 12817 15011
rect 12851 15008 12863 15011
rect 13078 15008 13084 15020
rect 12851 14980 13084 15008
rect 12851 14977 12863 14980
rect 12805 14971 12863 14977
rect 13078 14968 13084 14980
rect 13136 14968 13142 15020
rect 14829 15011 14887 15017
rect 14829 14977 14841 15011
rect 14875 15008 14887 15011
rect 15102 15008 15108 15020
rect 14875 14980 15108 15008
rect 14875 14977 14887 14980
rect 14829 14971 14887 14977
rect 15102 14968 15108 14980
rect 15160 14968 15166 15020
rect 20088 15017 20116 15048
rect 20346 15036 20352 15088
rect 20404 15076 20410 15088
rect 20404 15048 21128 15076
rect 20404 15036 20410 15048
rect 21100 15017 21128 15048
rect 20073 15011 20131 15017
rect 20073 14977 20085 15011
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20625 15011 20683 15017
rect 20625 14977 20637 15011
rect 20671 14977 20683 15011
rect 20625 14971 20683 14977
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 14977 21143 15011
rect 21085 14971 21143 14977
rect 6365 14943 6423 14949
rect 6365 14909 6377 14943
rect 6411 14909 6423 14943
rect 12526 14940 12532 14952
rect 12487 14912 12532 14940
rect 6365 14903 6423 14909
rect 5258 14804 5264 14816
rect 5219 14776 5264 14804
rect 5258 14764 5264 14776
rect 5316 14764 5322 14816
rect 6380 14804 6408 14903
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 12710 14940 12716 14952
rect 12671 14912 12716 14940
rect 12710 14900 12716 14912
rect 12768 14900 12774 14952
rect 15657 14943 15715 14949
rect 15657 14909 15669 14943
rect 15703 14940 15715 14943
rect 16114 14940 16120 14952
rect 15703 14912 16120 14940
rect 15703 14909 15715 14912
rect 15657 14903 15715 14909
rect 16114 14900 16120 14912
rect 16172 14900 16178 14952
rect 9585 14875 9643 14881
rect 9585 14841 9597 14875
rect 9631 14872 9643 14875
rect 20640 14872 20668 14971
rect 9631 14844 20668 14872
rect 9631 14841 9643 14844
rect 9585 14835 9643 14841
rect 7282 14804 7288 14816
rect 6380 14776 7288 14804
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 7466 14764 7472 14816
rect 7524 14804 7530 14816
rect 8021 14807 8079 14813
rect 8021 14804 8033 14807
rect 7524 14776 8033 14804
rect 7524 14764 7530 14776
rect 8021 14773 8033 14776
rect 8067 14773 8079 14807
rect 13170 14804 13176 14816
rect 13131 14776 13176 14804
rect 8021 14767 8079 14773
rect 13170 14764 13176 14776
rect 13228 14764 13234 14816
rect 13262 14764 13268 14816
rect 13320 14804 13326 14816
rect 14185 14807 14243 14813
rect 14185 14804 14197 14807
rect 13320 14776 14197 14804
rect 13320 14764 13326 14776
rect 14185 14773 14197 14776
rect 14231 14773 14243 14807
rect 21266 14804 21272 14816
rect 21227 14776 21272 14804
rect 14185 14767 14243 14773
rect 21266 14764 21272 14776
rect 21324 14764 21330 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 3234 14560 3240 14612
rect 3292 14600 3298 14612
rect 3789 14603 3847 14609
rect 3789 14600 3801 14603
rect 3292 14572 3801 14600
rect 3292 14560 3298 14572
rect 3789 14569 3801 14572
rect 3835 14569 3847 14603
rect 7006 14600 7012 14612
rect 6967 14572 7012 14600
rect 3789 14563 3847 14569
rect 7006 14560 7012 14572
rect 7064 14560 7070 14612
rect 9674 14600 9680 14612
rect 9635 14572 9680 14600
rect 9674 14560 9680 14572
rect 9732 14560 9738 14612
rect 12434 14600 12440 14612
rect 10520 14572 12440 14600
rect 6733 14535 6791 14541
rect 6733 14501 6745 14535
rect 6779 14532 6791 14535
rect 7098 14532 7104 14544
rect 6779 14504 7104 14532
rect 6779 14501 6791 14504
rect 6733 14495 6791 14501
rect 7098 14492 7104 14504
rect 7156 14492 7162 14544
rect 8113 14535 8171 14541
rect 8113 14532 8125 14535
rect 7392 14504 8125 14532
rect 4430 14396 4436 14408
rect 4391 14368 4436 14396
rect 4430 14356 4436 14368
rect 4488 14356 4494 14408
rect 5074 14356 5080 14408
rect 5132 14396 5138 14408
rect 5353 14399 5411 14405
rect 5353 14396 5365 14399
rect 5132 14368 5365 14396
rect 5132 14356 5138 14368
rect 5353 14365 5365 14368
rect 5399 14396 5411 14399
rect 7282 14396 7288 14408
rect 5399 14368 7288 14396
rect 5399 14365 5411 14368
rect 5353 14359 5411 14365
rect 7282 14356 7288 14368
rect 7340 14356 7346 14408
rect 7392 14405 7420 14504
rect 8113 14501 8125 14504
rect 8159 14532 8171 14535
rect 10520 14532 10548 14572
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 15102 14560 15108 14612
rect 15160 14600 15166 14612
rect 15473 14603 15531 14609
rect 15473 14600 15485 14603
rect 15160 14572 15485 14600
rect 15160 14560 15166 14572
rect 15473 14569 15485 14572
rect 15519 14569 15531 14603
rect 15473 14563 15531 14569
rect 20257 14603 20315 14609
rect 20257 14569 20269 14603
rect 20303 14600 20315 14603
rect 20622 14600 20628 14612
rect 20303 14572 20628 14600
rect 20303 14569 20315 14572
rect 20257 14563 20315 14569
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 20809 14603 20867 14609
rect 20809 14569 20821 14603
rect 20855 14600 20867 14603
rect 21082 14600 21088 14612
rect 20855 14572 21088 14600
rect 20855 14569 20867 14572
rect 20809 14563 20867 14569
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 8159 14504 10548 14532
rect 8159 14501 8171 14504
rect 8113 14495 8171 14501
rect 7558 14464 7564 14476
rect 7519 14436 7564 14464
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 8662 14424 8668 14476
rect 8720 14464 8726 14476
rect 9033 14467 9091 14473
rect 9033 14464 9045 14467
rect 8720 14436 9045 14464
rect 8720 14424 8726 14436
rect 9033 14433 9045 14436
rect 9079 14433 9091 14467
rect 9033 14427 9091 14433
rect 11425 14467 11483 14473
rect 11425 14433 11437 14467
rect 11471 14464 11483 14467
rect 12069 14467 12127 14473
rect 12069 14464 12081 14467
rect 11471 14436 12081 14464
rect 11471 14433 11483 14436
rect 11425 14427 11483 14433
rect 12069 14433 12081 14436
rect 12115 14433 12127 14467
rect 16301 14467 16359 14473
rect 16301 14464 16313 14467
rect 12069 14427 12127 14433
rect 15120 14436 16313 14464
rect 7377 14399 7435 14405
rect 7377 14365 7389 14399
rect 7423 14365 7435 14399
rect 7377 14359 7435 14365
rect 7469 14399 7527 14405
rect 7469 14365 7481 14399
rect 7515 14396 7527 14399
rect 8202 14396 8208 14408
rect 7515 14368 8208 14396
rect 7515 14365 7527 14368
rect 7469 14359 7527 14365
rect 5620 14331 5678 14337
rect 5620 14297 5632 14331
rect 5666 14328 5678 14331
rect 5994 14328 6000 14340
rect 5666 14300 6000 14328
rect 5666 14297 5678 14300
rect 5620 14291 5678 14297
rect 5994 14288 6000 14300
rect 6052 14288 6058 14340
rect 5258 14220 5264 14272
rect 5316 14260 5322 14272
rect 7392 14260 7420 14359
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 12084 14396 12112 14427
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 12084 14368 14105 14396
rect 14093 14365 14105 14368
rect 14139 14396 14151 14399
rect 14826 14396 14832 14408
rect 14139 14368 14832 14396
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 14826 14356 14832 14368
rect 14884 14356 14890 14408
rect 15120 14396 15148 14436
rect 16301 14433 16313 14436
rect 16347 14433 16359 14467
rect 16301 14427 16359 14433
rect 16114 14396 16120 14408
rect 14936 14368 15148 14396
rect 16075 14368 16120 14396
rect 9217 14331 9275 14337
rect 9217 14297 9229 14331
rect 9263 14328 9275 14331
rect 9674 14328 9680 14340
rect 9263 14300 9680 14328
rect 9263 14297 9275 14300
rect 9217 14291 9275 14297
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 11180 14331 11238 14337
rect 11180 14297 11192 14331
rect 11226 14328 11238 14331
rect 11226 14300 12020 14328
rect 11226 14297 11238 14300
rect 11180 14291 11238 14297
rect 5316 14232 7420 14260
rect 9309 14263 9367 14269
rect 5316 14220 5322 14232
rect 9309 14229 9321 14263
rect 9355 14260 9367 14263
rect 9766 14260 9772 14272
rect 9355 14232 9772 14260
rect 9355 14229 9367 14232
rect 9309 14223 9367 14229
rect 9766 14220 9772 14232
rect 9824 14220 9830 14272
rect 10042 14260 10048 14272
rect 10003 14232 10048 14260
rect 10042 14220 10048 14232
rect 10100 14220 10106 14272
rect 11992 14260 12020 14300
rect 12066 14288 12072 14340
rect 12124 14328 12130 14340
rect 12314 14331 12372 14337
rect 12314 14328 12326 14331
rect 12124 14300 12326 14328
rect 12124 14288 12130 14300
rect 12314 14297 12326 14300
rect 12360 14297 12372 14331
rect 12314 14291 12372 14297
rect 12526 14288 12532 14340
rect 12584 14328 12590 14340
rect 14360 14331 14418 14337
rect 14360 14328 14372 14331
rect 12584 14300 14372 14328
rect 12584 14288 12590 14300
rect 13262 14260 13268 14272
rect 11992 14232 13268 14260
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 13464 14269 13492 14300
rect 14360 14297 14372 14300
rect 14406 14328 14418 14331
rect 14936 14328 14964 14368
rect 16114 14356 16120 14368
rect 16172 14356 16178 14408
rect 19702 14356 19708 14408
rect 19760 14396 19766 14408
rect 20073 14399 20131 14405
rect 20073 14396 20085 14399
rect 19760 14368 20085 14396
rect 19760 14356 19766 14368
rect 20073 14365 20085 14368
rect 20119 14365 20131 14399
rect 20625 14399 20683 14405
rect 20625 14396 20637 14399
rect 20073 14359 20131 14365
rect 20180 14368 20637 14396
rect 14406 14300 14964 14328
rect 14406 14297 14418 14300
rect 14360 14291 14418 14297
rect 15102 14288 15108 14340
rect 15160 14328 15166 14340
rect 15160 14300 15792 14328
rect 15160 14288 15166 14300
rect 15764 14269 15792 14300
rect 16022 14288 16028 14340
rect 16080 14328 16086 14340
rect 20180 14328 20208 14368
rect 20625 14365 20637 14368
rect 20671 14365 20683 14399
rect 20625 14359 20683 14365
rect 21085 14399 21143 14405
rect 21085 14365 21097 14399
rect 21131 14365 21143 14399
rect 21085 14359 21143 14365
rect 16080 14300 20208 14328
rect 16080 14288 16086 14300
rect 20530 14288 20536 14340
rect 20588 14328 20594 14340
rect 21100 14328 21128 14359
rect 20588 14300 21128 14328
rect 20588 14288 20594 14300
rect 13449 14263 13507 14269
rect 13449 14229 13461 14263
rect 13495 14229 13507 14263
rect 13449 14223 13507 14229
rect 15749 14263 15807 14269
rect 15749 14229 15761 14263
rect 15795 14229 15807 14263
rect 15749 14223 15807 14229
rect 16209 14263 16267 14269
rect 16209 14229 16221 14263
rect 16255 14260 16267 14263
rect 16853 14263 16911 14269
rect 16853 14260 16865 14263
rect 16255 14232 16865 14260
rect 16255 14229 16267 14232
rect 16209 14223 16267 14229
rect 16853 14229 16865 14232
rect 16899 14260 16911 14263
rect 17034 14260 17040 14272
rect 16899 14232 17040 14260
rect 16899 14229 16911 14232
rect 16853 14223 16911 14229
rect 17034 14220 17040 14232
rect 17092 14220 17098 14272
rect 21266 14260 21272 14272
rect 21227 14232 21272 14260
rect 21266 14220 21272 14232
rect 21324 14220 21330 14272
rect 1104 14170 21896 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21896 14170
rect 1104 14096 21896 14118
rect 3697 14059 3755 14065
rect 3697 14025 3709 14059
rect 3743 14056 3755 14059
rect 4430 14056 4436 14068
rect 3743 14028 4436 14056
rect 3743 14025 3755 14028
rect 3697 14019 3755 14025
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 6638 14016 6644 14068
rect 6696 14056 6702 14068
rect 6733 14059 6791 14065
rect 6733 14056 6745 14059
rect 6696 14028 6745 14056
rect 6696 14016 6702 14028
rect 6733 14025 6745 14028
rect 6779 14025 6791 14059
rect 6733 14019 6791 14025
rect 8662 14016 8668 14068
rect 8720 14056 8726 14068
rect 9033 14059 9091 14065
rect 9033 14056 9045 14059
rect 8720 14028 9045 14056
rect 8720 14016 8726 14028
rect 9033 14025 9045 14028
rect 9079 14025 9091 14059
rect 9766 14056 9772 14068
rect 9727 14028 9772 14056
rect 9033 14019 9091 14025
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 13078 14056 13084 14068
rect 10152 14028 12664 14056
rect 13039 14028 13084 14056
rect 4832 13991 4890 13997
rect 4832 13957 4844 13991
rect 4878 13988 4890 13991
rect 7466 13988 7472 14000
rect 4878 13960 7472 13988
rect 4878 13957 4890 13960
rect 4832 13951 4890 13957
rect 7466 13948 7472 13960
rect 7524 13948 7530 14000
rect 9306 13948 9312 14000
rect 9364 13988 9370 14000
rect 10152 13988 10180 14028
rect 9364 13960 10180 13988
rect 10229 13991 10287 13997
rect 9364 13948 9370 13960
rect 10229 13957 10241 13991
rect 10275 13988 10287 13991
rect 10275 13960 11652 13988
rect 10275 13957 10287 13960
rect 10229 13951 10287 13957
rect 5074 13920 5080 13932
rect 5035 13892 5080 13920
rect 5074 13880 5080 13892
rect 5132 13880 5138 13932
rect 7098 13880 7104 13932
rect 7156 13920 7162 13932
rect 7377 13923 7435 13929
rect 7377 13920 7389 13923
rect 7156 13892 7389 13920
rect 7156 13880 7162 13892
rect 7377 13889 7389 13892
rect 7423 13889 7435 13923
rect 7377 13883 7435 13889
rect 7920 13923 7978 13929
rect 7920 13889 7932 13923
rect 7966 13920 7978 13923
rect 8662 13920 8668 13932
rect 7966 13892 8668 13920
rect 7966 13889 7978 13892
rect 7920 13883 7978 13889
rect 8662 13880 8668 13892
rect 8720 13920 8726 13932
rect 10042 13920 10048 13932
rect 8720 13892 10048 13920
rect 8720 13880 8726 13892
rect 10042 13880 10048 13892
rect 10100 13880 10106 13932
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13920 10195 13923
rect 10781 13923 10839 13929
rect 10781 13920 10793 13923
rect 10183 13892 10793 13920
rect 10183 13889 10195 13892
rect 10137 13883 10195 13889
rect 10781 13889 10793 13892
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 7282 13812 7288 13864
rect 7340 13852 7346 13864
rect 7653 13855 7711 13861
rect 7653 13852 7665 13855
rect 7340 13824 7665 13852
rect 7340 13812 7346 13824
rect 7653 13821 7665 13824
rect 7699 13821 7711 13855
rect 7653 13815 7711 13821
rect 10060 13784 10088 13880
rect 11624 13861 11652 13960
rect 10321 13855 10379 13861
rect 10321 13821 10333 13855
rect 10367 13821 10379 13855
rect 10321 13815 10379 13821
rect 11609 13855 11667 13861
rect 11609 13821 11621 13855
rect 11655 13852 11667 13855
rect 12342 13852 12348 13864
rect 11655 13824 12348 13852
rect 11655 13821 11667 13824
rect 11609 13815 11667 13821
rect 10336 13784 10364 13815
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 12636 13861 12664 14028
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 15102 14056 15108 14068
rect 15063 14028 15108 14056
rect 15102 14016 15108 14028
rect 15160 14016 15166 14068
rect 15473 14059 15531 14065
rect 15473 14025 15485 14059
rect 15519 14025 15531 14059
rect 16022 14056 16028 14068
rect 15983 14028 16028 14056
rect 15473 14019 15531 14025
rect 13170 13948 13176 14000
rect 13228 13988 13234 14000
rect 15013 13991 15071 13997
rect 15013 13988 15025 13991
rect 13228 13960 15025 13988
rect 13228 13948 13234 13960
rect 15013 13957 15025 13960
rect 15059 13957 15071 13991
rect 15013 13951 15071 13957
rect 12713 13923 12771 13929
rect 12713 13889 12725 13923
rect 12759 13920 12771 13923
rect 12802 13920 12808 13932
rect 12759 13892 12808 13920
rect 12759 13889 12771 13892
rect 12713 13883 12771 13889
rect 12802 13880 12808 13892
rect 12860 13920 12866 13932
rect 13354 13920 13360 13932
rect 12860 13892 13360 13920
rect 12860 13880 12866 13892
rect 13354 13880 13360 13892
rect 13412 13880 13418 13932
rect 15488 13920 15516 14019
rect 16022 14016 16028 14028
rect 16080 14016 16086 14068
rect 19702 14056 19708 14068
rect 19663 14028 19708 14056
rect 19702 14016 19708 14028
rect 19760 14016 19766 14068
rect 17580 13991 17638 13997
rect 17580 13957 17592 13991
rect 17626 13988 17638 13991
rect 17954 13988 17960 14000
rect 17626 13960 17960 13988
rect 17626 13957 17638 13960
rect 17580 13951 17638 13957
rect 17954 13948 17960 13960
rect 18012 13988 18018 14000
rect 18874 13988 18880 14000
rect 18012 13960 18880 13988
rect 18012 13948 18018 13960
rect 18874 13948 18880 13960
rect 18932 13948 18938 14000
rect 19058 13948 19064 14000
rect 19116 13988 19122 14000
rect 19337 13991 19395 13997
rect 19337 13988 19349 13991
rect 19116 13960 19349 13988
rect 19116 13948 19122 13960
rect 19337 13957 19349 13960
rect 19383 13957 19395 13991
rect 19337 13951 19395 13957
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 15488 13892 15853 13920
rect 15841 13889 15853 13892
rect 15887 13889 15899 13923
rect 17310 13920 17316 13932
rect 17271 13892 17316 13920
rect 15841 13883 15899 13889
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 18506 13880 18512 13932
rect 18564 13920 18570 13932
rect 19245 13923 19303 13929
rect 19245 13920 19257 13923
rect 18564 13892 19257 13920
rect 18564 13880 18570 13892
rect 19245 13889 19257 13892
rect 19291 13889 19303 13923
rect 20622 13920 20628 13932
rect 20583 13892 20628 13920
rect 19245 13883 19303 13889
rect 20622 13880 20628 13892
rect 20680 13880 20686 13932
rect 21082 13920 21088 13932
rect 21043 13892 21088 13920
rect 21082 13880 21088 13892
rect 21140 13880 21146 13932
rect 12529 13855 12587 13861
rect 12529 13821 12541 13855
rect 12575 13821 12587 13855
rect 12529 13815 12587 13821
rect 12621 13855 12679 13861
rect 12621 13821 12633 13855
rect 12667 13852 12679 13855
rect 13817 13855 13875 13861
rect 13817 13852 13829 13855
rect 12667 13824 13829 13852
rect 12667 13821 12679 13824
rect 12621 13815 12679 13821
rect 13817 13821 13829 13824
rect 13863 13852 13875 13855
rect 14366 13852 14372 13864
rect 13863 13824 14372 13852
rect 13863 13821 13875 13824
rect 13817 13815 13875 13821
rect 10060 13756 10364 13784
rect 12544 13784 12572 13815
rect 14366 13812 14372 13824
rect 14424 13812 14430 13864
rect 14918 13852 14924 13864
rect 14879 13824 14924 13852
rect 14918 13812 14924 13824
rect 14976 13812 14982 13864
rect 19061 13855 19119 13861
rect 19061 13852 19073 13855
rect 18708 13824 19073 13852
rect 12894 13784 12900 13796
rect 12544 13756 12900 13784
rect 12894 13744 12900 13756
rect 12952 13744 12958 13796
rect 13280 13756 16804 13784
rect 5902 13676 5908 13728
rect 5960 13716 5966 13728
rect 11606 13716 11612 13728
rect 5960 13688 11612 13716
rect 5960 13676 5966 13688
rect 11606 13676 11612 13688
rect 11664 13676 11670 13728
rect 11790 13676 11796 13728
rect 11848 13716 11854 13728
rect 13280 13716 13308 13756
rect 11848 13688 13308 13716
rect 16776 13716 16804 13756
rect 18708 13725 18736 13824
rect 19061 13821 19073 13824
rect 19107 13821 19119 13855
rect 19978 13852 19984 13864
rect 19939 13824 19984 13852
rect 19061 13815 19119 13821
rect 19978 13812 19984 13824
rect 20036 13812 20042 13864
rect 18693 13719 18751 13725
rect 18693 13716 18705 13719
rect 16776 13688 18705 13716
rect 11848 13676 11854 13688
rect 18693 13685 18705 13688
rect 18739 13685 18751 13719
rect 18693 13679 18751 13685
rect 20809 13719 20867 13725
rect 20809 13685 20821 13719
rect 20855 13716 20867 13719
rect 20990 13716 20996 13728
rect 20855 13688 20996 13716
rect 20855 13685 20867 13688
rect 20809 13679 20867 13685
rect 20990 13676 20996 13688
rect 21048 13676 21054 13728
rect 21266 13716 21272 13728
rect 21227 13688 21272 13716
rect 21266 13676 21272 13688
rect 21324 13676 21330 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 5905 13515 5963 13521
rect 5905 13481 5917 13515
rect 5951 13512 5963 13515
rect 7006 13512 7012 13524
rect 5951 13484 7012 13512
rect 5951 13481 5963 13484
rect 5905 13475 5963 13481
rect 7006 13472 7012 13484
rect 7064 13512 7070 13524
rect 7558 13512 7564 13524
rect 7064 13484 7564 13512
rect 7064 13472 7070 13484
rect 7558 13472 7564 13484
rect 7616 13472 7622 13524
rect 9674 13512 9680 13524
rect 9635 13484 9680 13512
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 12710 13472 12716 13524
rect 12768 13512 12774 13524
rect 13081 13515 13139 13521
rect 13081 13512 13093 13515
rect 12768 13484 13093 13512
rect 12768 13472 12774 13484
rect 13081 13481 13093 13484
rect 13127 13481 13139 13515
rect 18506 13512 18512 13524
rect 18467 13484 18512 13512
rect 13081 13475 13139 13481
rect 18506 13472 18512 13484
rect 18564 13472 18570 13524
rect 19058 13472 19064 13524
rect 19116 13512 19122 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 19116 13484 19257 13512
rect 19116 13472 19122 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 19245 13475 19303 13481
rect 20346 13472 20352 13524
rect 20404 13512 20410 13524
rect 20533 13515 20591 13521
rect 20533 13512 20545 13515
rect 20404 13484 20545 13512
rect 20404 13472 20410 13484
rect 20533 13481 20545 13484
rect 20579 13481 20591 13515
rect 20533 13475 20591 13481
rect 20809 13515 20867 13521
rect 20809 13481 20821 13515
rect 20855 13512 20867 13515
rect 21542 13512 21548 13524
rect 20855 13484 21548 13512
rect 20855 13481 20867 13484
rect 20809 13475 20867 13481
rect 21542 13472 21548 13484
rect 21600 13472 21606 13524
rect 8588 13416 10456 13444
rect 2222 13268 2228 13320
rect 2280 13308 2286 13320
rect 7282 13308 7288 13320
rect 2280 13280 7144 13308
rect 7243 13280 7288 13308
rect 2280 13268 2286 13280
rect 7018 13243 7076 13249
rect 7018 13209 7030 13243
rect 7064 13209 7076 13243
rect 7116 13240 7144 13280
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 8588 13240 8616 13416
rect 8662 13336 8668 13388
rect 8720 13376 8726 13388
rect 9033 13379 9091 13385
rect 9033 13376 9045 13379
rect 8720 13348 9045 13376
rect 8720 13336 8726 13348
rect 9033 13345 9045 13348
rect 9079 13345 9091 13379
rect 9033 13339 9091 13345
rect 9122 13336 9128 13388
rect 9180 13376 9186 13388
rect 9217 13379 9275 13385
rect 9217 13376 9229 13379
rect 9180 13348 9229 13376
rect 9180 13336 9186 13348
rect 9217 13345 9229 13348
rect 9263 13345 9275 13379
rect 10318 13376 10324 13388
rect 10279 13348 10324 13376
rect 9217 13339 9275 13345
rect 10318 13336 10324 13348
rect 10376 13336 10382 13388
rect 10428 13376 10456 13416
rect 11606 13404 11612 13456
rect 11664 13444 11670 13456
rect 17402 13444 17408 13456
rect 11664 13416 17408 13444
rect 11664 13404 11670 13416
rect 17402 13404 17408 13416
rect 17460 13404 17466 13456
rect 12529 13379 12587 13385
rect 10428 13348 11928 13376
rect 11790 13308 11796 13320
rect 7116 13212 8616 13240
rect 9048 13280 11796 13308
rect 7018 13203 7076 13209
rect 7024 13172 7052 13203
rect 9048 13172 9076 13280
rect 11790 13268 11796 13280
rect 11848 13268 11854 13320
rect 11900 13240 11928 13348
rect 12529 13345 12541 13379
rect 12575 13376 12587 13379
rect 12894 13376 12900 13388
rect 12575 13348 12900 13376
rect 12575 13345 12587 13348
rect 12529 13339 12587 13345
rect 12894 13336 12900 13348
rect 12952 13336 12958 13388
rect 17954 13376 17960 13388
rect 17915 13348 17960 13376
rect 17954 13336 17960 13348
rect 18012 13376 18018 13388
rect 19797 13379 19855 13385
rect 19797 13376 19809 13379
rect 18012 13348 19809 13376
rect 18012 13336 18018 13348
rect 19797 13345 19809 13348
rect 19843 13345 19855 13379
rect 19797 13339 19855 13345
rect 12069 13311 12127 13317
rect 12069 13277 12081 13311
rect 12115 13308 12127 13311
rect 18046 13308 18052 13320
rect 12115 13280 15240 13308
rect 12115 13277 12127 13280
rect 12069 13271 12127 13277
rect 12621 13243 12679 13249
rect 12621 13240 12633 13243
rect 11900 13212 12633 13240
rect 12621 13209 12633 13212
rect 12667 13209 12679 13243
rect 15212 13240 15240 13280
rect 17604 13280 18052 13308
rect 17604 13240 17632 13280
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 19613 13311 19671 13317
rect 19613 13277 19625 13311
rect 19659 13308 19671 13311
rect 19978 13308 19984 13320
rect 19659 13280 19984 13308
rect 19659 13277 19671 13280
rect 19613 13271 19671 13277
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 20070 13268 20076 13320
rect 20128 13308 20134 13320
rect 20349 13311 20407 13317
rect 20349 13308 20361 13311
rect 20128 13280 20361 13308
rect 20128 13268 20134 13280
rect 20349 13277 20361 13280
rect 20395 13277 20407 13311
rect 20990 13308 20996 13320
rect 20951 13280 20996 13308
rect 20349 13271 20407 13277
rect 20990 13268 20996 13280
rect 21048 13268 21054 13320
rect 15212 13212 17632 13240
rect 12621 13203 12679 13209
rect 17678 13200 17684 13252
rect 17736 13240 17742 13252
rect 18141 13243 18199 13249
rect 18141 13240 18153 13243
rect 17736 13212 18153 13240
rect 17736 13200 17742 13212
rect 18141 13209 18153 13212
rect 18187 13240 18199 13243
rect 18785 13243 18843 13249
rect 18785 13240 18797 13243
rect 18187 13212 18797 13240
rect 18187 13209 18199 13212
rect 18141 13203 18199 13209
rect 18785 13209 18797 13212
rect 18831 13209 18843 13243
rect 18785 13203 18843 13209
rect 19705 13243 19763 13249
rect 19705 13209 19717 13243
rect 19751 13240 19763 13243
rect 21174 13240 21180 13252
rect 19751 13212 21180 13240
rect 19751 13209 19763 13212
rect 19705 13203 19763 13209
rect 21174 13200 21180 13212
rect 21232 13240 21238 13252
rect 21269 13243 21327 13249
rect 21269 13240 21281 13243
rect 21232 13212 21281 13240
rect 21232 13200 21238 13212
rect 21269 13209 21281 13212
rect 21315 13209 21327 13243
rect 21269 13203 21327 13209
rect 7024 13144 9076 13172
rect 9309 13175 9367 13181
rect 9309 13141 9321 13175
rect 9355 13172 9367 13175
rect 9582 13172 9588 13184
rect 9355 13144 9588 13172
rect 9355 13141 9367 13144
rect 9309 13135 9367 13141
rect 9582 13132 9588 13144
rect 9640 13172 9646 13184
rect 9953 13175 10011 13181
rect 9953 13172 9965 13175
rect 9640 13144 9965 13172
rect 9640 13132 9646 13144
rect 9953 13141 9965 13144
rect 9999 13141 10011 13175
rect 9953 13135 10011 13141
rect 12434 13132 12440 13184
rect 12492 13172 12498 13184
rect 12713 13175 12771 13181
rect 12713 13172 12725 13175
rect 12492 13144 12725 13172
rect 12492 13132 12498 13144
rect 12713 13141 12725 13144
rect 12759 13172 12771 13175
rect 13357 13175 13415 13181
rect 13357 13172 13369 13175
rect 12759 13144 13369 13172
rect 12759 13141 12771 13144
rect 12713 13135 12771 13141
rect 13357 13141 13369 13144
rect 13403 13172 13415 13175
rect 13538 13172 13544 13184
rect 13403 13144 13544 13172
rect 13403 13141 13415 13144
rect 13357 13135 13415 13141
rect 13538 13132 13544 13144
rect 13596 13132 13602 13184
rect 17402 13132 17408 13184
rect 17460 13172 17466 13184
rect 18049 13175 18107 13181
rect 18049 13172 18061 13175
rect 17460 13144 18061 13172
rect 17460 13132 17466 13144
rect 18049 13141 18061 13144
rect 18095 13141 18107 13175
rect 18049 13135 18107 13141
rect 1104 13082 21896 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21896 13082
rect 1104 13008 21896 13030
rect 5994 12928 6000 12980
rect 6052 12968 6058 12980
rect 6365 12971 6423 12977
rect 6365 12968 6377 12971
rect 6052 12940 6377 12968
rect 6052 12928 6058 12940
rect 6365 12937 6377 12940
rect 6411 12937 6423 12971
rect 12066 12968 12072 12980
rect 12027 12940 12072 12968
rect 6365 12931 6423 12937
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 19613 12971 19671 12977
rect 19613 12937 19625 12971
rect 19659 12937 19671 12971
rect 20530 12968 20536 12980
rect 20491 12940 20536 12968
rect 19613 12931 19671 12937
rect 10318 12860 10324 12912
rect 10376 12900 10382 12912
rect 12989 12903 13047 12909
rect 12989 12900 13001 12903
rect 10376 12872 13001 12900
rect 10376 12860 10382 12872
rect 12989 12869 13001 12872
rect 13035 12869 13047 12903
rect 12989 12863 13047 12869
rect 14737 12903 14795 12909
rect 14737 12869 14749 12903
rect 14783 12900 14795 12903
rect 14826 12900 14832 12912
rect 14783 12872 14832 12900
rect 14783 12869 14795 12872
rect 14737 12863 14795 12869
rect 14826 12860 14832 12872
rect 14884 12860 14890 12912
rect 16574 12860 16580 12912
rect 16632 12900 16638 12912
rect 17678 12900 17684 12912
rect 16632 12872 17684 12900
rect 16632 12860 16638 12872
rect 17678 12860 17684 12872
rect 17736 12860 17742 12912
rect 19628 12900 19656 12931
rect 20530 12928 20536 12940
rect 20588 12928 20594 12980
rect 20806 12968 20812 12980
rect 20767 12940 20812 12968
rect 20806 12928 20812 12940
rect 20864 12928 20870 12980
rect 21358 12968 21364 12980
rect 21319 12940 21364 12968
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 19628 12872 21036 12900
rect 7006 12832 7012 12844
rect 6967 12804 7012 12832
rect 7006 12792 7012 12804
rect 7064 12792 7070 12844
rect 11609 12835 11667 12841
rect 11609 12801 11621 12835
rect 11655 12832 11667 12835
rect 11790 12832 11796 12844
rect 11655 12804 11796 12832
rect 11655 12801 11667 12804
rect 11609 12795 11667 12801
rect 11790 12792 11796 12804
rect 11848 12792 11854 12844
rect 12713 12835 12771 12841
rect 12713 12801 12725 12835
rect 12759 12832 12771 12835
rect 12894 12832 12900 12844
rect 12759 12804 12900 12832
rect 12759 12801 12771 12804
rect 12713 12795 12771 12801
rect 12894 12792 12900 12804
rect 12952 12792 12958 12844
rect 17037 12835 17095 12841
rect 17037 12801 17049 12835
rect 17083 12832 17095 12835
rect 17310 12832 17316 12844
rect 17083 12804 17316 12832
rect 17083 12801 17095 12804
rect 17037 12795 17095 12801
rect 17310 12792 17316 12804
rect 17368 12792 17374 12844
rect 19153 12835 19211 12841
rect 19153 12801 19165 12835
rect 19199 12832 19211 12835
rect 19242 12832 19248 12844
rect 19199 12804 19248 12832
rect 19199 12801 19211 12804
rect 19153 12795 19211 12801
rect 19242 12792 19248 12804
rect 19300 12832 19306 12844
rect 19429 12835 19487 12841
rect 19429 12832 19441 12835
rect 19300 12804 19441 12832
rect 19300 12792 19306 12804
rect 19429 12801 19441 12804
rect 19475 12801 19487 12835
rect 19429 12795 19487 12801
rect 19518 12792 19524 12844
rect 19576 12832 19582 12844
rect 21008 12841 21036 12872
rect 19889 12835 19947 12841
rect 19889 12832 19901 12835
rect 19576 12804 19901 12832
rect 19576 12792 19582 12804
rect 19889 12801 19901 12804
rect 19935 12801 19947 12835
rect 19889 12795 19947 12801
rect 20349 12835 20407 12841
rect 20349 12801 20361 12835
rect 20395 12801 20407 12835
rect 20349 12795 20407 12801
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12801 21051 12835
rect 20993 12795 21051 12801
rect 17126 12764 17132 12776
rect 17087 12736 17132 12764
rect 17126 12724 17132 12736
rect 17184 12724 17190 12776
rect 17218 12724 17224 12776
rect 17276 12764 17282 12776
rect 17276 12736 17321 12764
rect 17276 12724 17282 12736
rect 18414 12724 18420 12776
rect 18472 12764 18478 12776
rect 20364 12764 20392 12795
rect 18472 12736 20392 12764
rect 18472 12724 18478 12736
rect 11793 12699 11851 12705
rect 11793 12665 11805 12699
rect 11839 12696 11851 12699
rect 19978 12696 19984 12708
rect 11839 12668 19984 12696
rect 11839 12665 11851 12668
rect 11793 12659 11851 12665
rect 19978 12656 19984 12668
rect 20036 12656 20042 12708
rect 20073 12699 20131 12705
rect 20073 12665 20085 12699
rect 20119 12696 20131 12699
rect 20714 12696 20720 12708
rect 20119 12668 20720 12696
rect 20119 12665 20131 12668
rect 20073 12659 20131 12665
rect 20714 12656 20720 12668
rect 20772 12656 20778 12708
rect 9582 12588 9588 12640
rect 9640 12628 9646 12640
rect 16574 12628 16580 12640
rect 9640 12600 16580 12628
rect 9640 12588 9646 12600
rect 16574 12588 16580 12600
rect 16632 12588 16638 12640
rect 16669 12631 16727 12637
rect 16669 12597 16681 12631
rect 16715 12628 16727 12631
rect 16942 12628 16948 12640
rect 16715 12600 16948 12628
rect 16715 12597 16727 12600
rect 16669 12591 16727 12597
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 18417 12631 18475 12637
rect 18417 12597 18429 12631
rect 18463 12628 18475 12631
rect 18598 12628 18604 12640
rect 18463 12600 18604 12628
rect 18463 12597 18475 12600
rect 18417 12591 18475 12597
rect 18598 12588 18604 12600
rect 18656 12588 18662 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 8294 12384 8300 12436
rect 8352 12424 8358 12436
rect 9033 12427 9091 12433
rect 9033 12424 9045 12427
rect 8352 12396 9045 12424
rect 8352 12384 8358 12396
rect 9033 12393 9045 12396
rect 9079 12424 9091 12427
rect 9582 12424 9588 12436
rect 9079 12396 9588 12424
rect 9079 12393 9091 12396
rect 9033 12387 9091 12393
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 12894 12424 12900 12436
rect 10100 12396 12572 12424
rect 12855 12396 12900 12424
rect 10100 12384 10106 12396
rect 7926 12288 7932 12300
rect 7887 12260 7932 12288
rect 7926 12248 7932 12260
rect 7984 12248 7990 12300
rect 8018 12248 8024 12300
rect 8076 12288 8082 12300
rect 8113 12291 8171 12297
rect 8113 12288 8125 12291
rect 8076 12260 8125 12288
rect 8076 12248 8082 12260
rect 8113 12257 8125 12260
rect 8159 12257 8171 12291
rect 8113 12251 8171 12257
rect 7282 12180 7288 12232
rect 7340 12220 7346 12232
rect 8386 12220 8392 12232
rect 7340 12192 8392 12220
rect 7340 12180 7346 12192
rect 8386 12180 8392 12192
rect 8444 12220 8450 12232
rect 9401 12223 9459 12229
rect 9401 12220 9413 12223
rect 8444 12192 9413 12220
rect 8444 12180 8450 12192
rect 9401 12189 9413 12192
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 9490 12180 9496 12232
rect 9548 12220 9554 12232
rect 9657 12223 9715 12229
rect 9657 12220 9669 12223
rect 9548 12192 9669 12220
rect 9548 12180 9554 12192
rect 9657 12189 9669 12192
rect 9703 12189 9715 12223
rect 9657 12183 9715 12189
rect 11517 12223 11575 12229
rect 11517 12189 11529 12223
rect 11563 12220 11575 12223
rect 11606 12220 11612 12232
rect 11563 12192 11612 12220
rect 11563 12189 11575 12192
rect 11517 12183 11575 12189
rect 11606 12180 11612 12192
rect 11664 12180 11670 12232
rect 8205 12155 8263 12161
rect 8205 12121 8217 12155
rect 8251 12152 8263 12155
rect 8294 12152 8300 12164
rect 8251 12124 8300 12152
rect 8251 12121 8263 12124
rect 8205 12115 8263 12121
rect 8294 12112 8300 12124
rect 8352 12112 8358 12164
rect 11146 12112 11152 12164
rect 11204 12152 11210 12164
rect 11762 12155 11820 12161
rect 11762 12152 11774 12155
rect 11204 12124 11774 12152
rect 11204 12112 11210 12124
rect 11762 12121 11774 12124
rect 11808 12121 11820 12155
rect 12544 12152 12572 12396
rect 12894 12384 12900 12396
rect 12952 12384 12958 12436
rect 14277 12427 14335 12433
rect 14277 12393 14289 12427
rect 14323 12424 14335 12427
rect 17037 12427 17095 12433
rect 14323 12396 16344 12424
rect 14323 12393 14335 12396
rect 14277 12387 14335 12393
rect 16316 12356 16344 12396
rect 17037 12393 17049 12427
rect 17083 12424 17095 12427
rect 17126 12424 17132 12436
rect 17083 12396 17132 12424
rect 17083 12393 17095 12396
rect 17037 12387 17095 12393
rect 17126 12384 17132 12396
rect 17184 12384 17190 12436
rect 17310 12424 17316 12436
rect 17271 12396 17316 12424
rect 17310 12384 17316 12396
rect 17368 12384 17374 12436
rect 20438 12384 20444 12436
rect 20496 12424 20502 12436
rect 20533 12427 20591 12433
rect 20533 12424 20545 12427
rect 20496 12396 20545 12424
rect 20496 12384 20502 12396
rect 20533 12393 20545 12396
rect 20579 12393 20591 12427
rect 20533 12387 20591 12393
rect 20993 12427 21051 12433
rect 20993 12393 21005 12427
rect 21039 12424 21051 12427
rect 21082 12424 21088 12436
rect 21039 12396 21088 12424
rect 21039 12393 21051 12396
rect 20993 12387 21051 12393
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 18414 12356 18420 12368
rect 16316 12328 18420 12356
rect 18414 12316 18420 12328
rect 18472 12316 18478 12368
rect 16393 12291 16451 12297
rect 16393 12257 16405 12291
rect 16439 12288 16451 12291
rect 17770 12288 17776 12300
rect 16439 12260 17776 12288
rect 16439 12257 16451 12260
rect 16393 12251 16451 12257
rect 17770 12248 17776 12260
rect 17828 12288 17834 12300
rect 17865 12291 17923 12297
rect 17865 12288 17877 12291
rect 17828 12260 17877 12288
rect 17828 12248 17834 12260
rect 17865 12257 17877 12260
rect 17911 12257 17923 12291
rect 17865 12251 17923 12257
rect 19904 12260 21404 12288
rect 14093 12223 14151 12229
rect 14093 12189 14105 12223
rect 14139 12220 14151 12223
rect 15010 12220 15016 12232
rect 14139 12192 15016 12220
rect 14139 12189 14151 12192
rect 14093 12183 14151 12189
rect 15010 12180 15016 12192
rect 15068 12180 15074 12232
rect 16022 12220 16028 12232
rect 15983 12192 16028 12220
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 16574 12220 16580 12232
rect 16535 12192 16580 12220
rect 16574 12180 16580 12192
rect 16632 12180 16638 12232
rect 16669 12223 16727 12229
rect 16669 12189 16681 12223
rect 16715 12220 16727 12223
rect 17678 12220 17684 12232
rect 16715 12192 17684 12220
rect 16715 12189 16727 12192
rect 16669 12183 16727 12189
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 17954 12180 17960 12232
rect 18012 12220 18018 12232
rect 18598 12220 18604 12232
rect 18012 12192 18604 12220
rect 18012 12180 18018 12192
rect 18598 12180 18604 12192
rect 18656 12180 18662 12232
rect 19904 12229 19932 12260
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12189 19947 12223
rect 20349 12223 20407 12229
rect 20349 12220 20361 12223
rect 19889 12183 19947 12189
rect 20088 12192 20361 12220
rect 15780 12155 15838 12161
rect 11762 12115 11820 12121
rect 11900 12124 12434 12152
rect 12544 12124 15608 12152
rect 8573 12087 8631 12093
rect 8573 12053 8585 12087
rect 8619 12084 8631 12087
rect 8662 12084 8668 12096
rect 8619 12056 8668 12084
rect 8619 12053 8631 12056
rect 8573 12047 8631 12053
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 10778 12084 10784 12096
rect 10739 12056 10784 12084
rect 10778 12044 10784 12056
rect 10836 12044 10842 12096
rect 10870 12044 10876 12096
rect 10928 12084 10934 12096
rect 11057 12087 11115 12093
rect 11057 12084 11069 12087
rect 10928 12056 11069 12084
rect 10928 12044 10934 12056
rect 11057 12053 11069 12056
rect 11103 12084 11115 12087
rect 11900 12084 11928 12124
rect 11103 12056 11928 12084
rect 12406 12084 12434 12124
rect 14550 12084 14556 12096
rect 12406 12056 14556 12084
rect 11103 12053 11115 12056
rect 11057 12047 11115 12053
rect 14550 12044 14556 12056
rect 14608 12044 14614 12096
rect 14645 12087 14703 12093
rect 14645 12053 14657 12087
rect 14691 12084 14703 12087
rect 15470 12084 15476 12096
rect 14691 12056 15476 12084
rect 14691 12053 14703 12056
rect 14645 12047 14703 12053
rect 15470 12044 15476 12056
rect 15528 12044 15534 12096
rect 15580 12084 15608 12124
rect 15780 12121 15792 12155
rect 15826 12152 15838 12155
rect 17126 12152 17132 12164
rect 15826 12124 17132 12152
rect 15826 12121 15838 12124
rect 15780 12115 15838 12121
rect 17126 12112 17132 12124
rect 17184 12112 17190 12164
rect 17773 12155 17831 12161
rect 17773 12152 17785 12155
rect 17236 12124 17785 12152
rect 17236 12084 17264 12124
rect 17773 12121 17785 12124
rect 17819 12152 17831 12155
rect 17819 12124 18920 12152
rect 17819 12121 17831 12124
rect 17773 12115 17831 12121
rect 15580 12056 17264 12084
rect 17681 12087 17739 12093
rect 17681 12053 17693 12087
rect 17727 12084 17739 12087
rect 17954 12084 17960 12096
rect 17727 12056 17960 12084
rect 17727 12053 17739 12056
rect 17681 12047 17739 12053
rect 17954 12044 17960 12056
rect 18012 12044 18018 12096
rect 18046 12044 18052 12096
rect 18104 12084 18110 12096
rect 18892 12093 18920 12124
rect 18325 12087 18383 12093
rect 18325 12084 18337 12087
rect 18104 12056 18337 12084
rect 18104 12044 18110 12056
rect 18325 12053 18337 12056
rect 18371 12053 18383 12087
rect 18325 12047 18383 12053
rect 18877 12087 18935 12093
rect 18877 12053 18889 12087
rect 18923 12084 18935 12087
rect 19058 12084 19064 12096
rect 18923 12056 19064 12084
rect 18923 12053 18935 12056
rect 18877 12047 18935 12053
rect 19058 12044 19064 12056
rect 19116 12044 19122 12096
rect 19334 12044 19340 12096
rect 19392 12084 19398 12096
rect 19613 12087 19671 12093
rect 19613 12084 19625 12087
rect 19392 12056 19625 12084
rect 19392 12044 19398 12056
rect 19613 12053 19625 12056
rect 19659 12084 19671 12087
rect 19702 12084 19708 12096
rect 19659 12056 19708 12084
rect 19659 12053 19671 12056
rect 19613 12047 19671 12053
rect 19702 12044 19708 12056
rect 19760 12044 19766 12096
rect 20088 12093 20116 12192
rect 20349 12189 20361 12192
rect 20395 12189 20407 12223
rect 20349 12183 20407 12189
rect 20714 12180 20720 12232
rect 20772 12220 20778 12232
rect 20809 12223 20867 12229
rect 20809 12220 20821 12223
rect 20772 12192 20821 12220
rect 20772 12180 20778 12192
rect 20809 12189 20821 12192
rect 20855 12189 20867 12223
rect 20809 12183 20867 12189
rect 21376 12096 21404 12260
rect 20073 12087 20131 12093
rect 20073 12053 20085 12087
rect 20119 12053 20131 12087
rect 21358 12084 21364 12096
rect 21319 12056 21364 12084
rect 20073 12047 20131 12053
rect 21358 12044 21364 12056
rect 21416 12044 21422 12096
rect 1104 11994 21896 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21896 11994
rect 1104 11920 21896 11942
rect 8662 11880 8668 11892
rect 8623 11852 8668 11880
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 8757 11883 8815 11889
rect 8757 11849 8769 11883
rect 8803 11880 8815 11883
rect 9401 11883 9459 11889
rect 9401 11880 9413 11883
rect 8803 11852 9413 11880
rect 8803 11849 8815 11852
rect 8757 11843 8815 11849
rect 9401 11849 9413 11852
rect 9447 11849 9459 11883
rect 9401 11843 9459 11849
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 10226 11880 10232 11892
rect 9815 11852 10232 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 10226 11840 10232 11852
rect 10284 11880 10290 11892
rect 10870 11880 10876 11892
rect 10284 11852 10876 11880
rect 10284 11840 10290 11852
rect 10870 11840 10876 11852
rect 10928 11840 10934 11892
rect 11146 11880 11152 11892
rect 11107 11852 11152 11880
rect 11146 11840 11152 11852
rect 11204 11840 11210 11892
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 11790 11880 11796 11892
rect 11563 11852 11796 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 11790 11840 11796 11852
rect 11848 11840 11854 11892
rect 12342 11840 12348 11892
rect 12400 11880 12406 11892
rect 12400 11852 14228 11880
rect 12400 11840 12406 11852
rect 9861 11815 9919 11821
rect 9861 11781 9873 11815
rect 9907 11812 9919 11815
rect 9950 11812 9956 11824
rect 9907 11784 9956 11812
rect 9907 11781 9919 11784
rect 9861 11775 9919 11781
rect 9950 11772 9956 11784
rect 10008 11772 10014 11824
rect 10778 11812 10784 11824
rect 10520 11784 10784 11812
rect 2130 11704 2136 11756
rect 2188 11744 2194 11756
rect 10520 11753 10548 11784
rect 10778 11772 10784 11784
rect 10836 11812 10842 11824
rect 10836 11784 12112 11812
rect 10836 11772 10842 11784
rect 10505 11747 10563 11753
rect 2188 11716 10456 11744
rect 2188 11704 2194 11716
rect 8573 11679 8631 11685
rect 8573 11645 8585 11679
rect 8619 11676 8631 11679
rect 9490 11676 9496 11688
rect 8619 11648 9496 11676
rect 8619 11645 8631 11648
rect 8573 11639 8631 11645
rect 9490 11636 9496 11648
rect 9548 11636 9554 11688
rect 9950 11636 9956 11688
rect 10008 11676 10014 11688
rect 10428 11676 10456 11716
rect 10505 11713 10517 11747
rect 10551 11713 10563 11747
rect 10505 11707 10563 11713
rect 11330 11704 11336 11756
rect 11388 11744 11394 11756
rect 11885 11747 11943 11753
rect 11885 11744 11897 11747
rect 11388 11716 11897 11744
rect 11388 11704 11394 11716
rect 11885 11713 11897 11716
rect 11931 11713 11943 11747
rect 11885 11707 11943 11713
rect 11790 11676 11796 11688
rect 10008 11648 10053 11676
rect 10428 11648 11796 11676
rect 10008 11636 10014 11648
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 12084 11685 12112 11784
rect 14200 11744 14228 11852
rect 14550 11840 14556 11892
rect 14608 11880 14614 11892
rect 16942 11880 16948 11892
rect 14608 11852 14964 11880
rect 16903 11852 16948 11880
rect 14608 11840 14614 11852
rect 14308 11815 14366 11821
rect 14308 11781 14320 11815
rect 14354 11812 14366 11815
rect 14829 11815 14887 11821
rect 14829 11812 14841 11815
rect 14354 11784 14841 11812
rect 14354 11781 14366 11784
rect 14308 11775 14366 11781
rect 14829 11781 14841 11784
rect 14875 11781 14887 11815
rect 14936 11812 14964 11852
rect 16942 11840 16948 11852
rect 17000 11840 17006 11892
rect 17037 11883 17095 11889
rect 17037 11849 17049 11883
rect 17083 11880 17095 11883
rect 17681 11883 17739 11889
rect 17681 11880 17693 11883
rect 17083 11852 17693 11880
rect 17083 11849 17095 11852
rect 17037 11843 17095 11849
rect 17681 11849 17693 11852
rect 17727 11849 17739 11883
rect 18046 11880 18052 11892
rect 18007 11852 18052 11880
rect 17681 11843 17739 11849
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 18141 11883 18199 11889
rect 18141 11849 18153 11883
rect 18187 11880 18199 11883
rect 18693 11883 18751 11889
rect 18693 11880 18705 11883
rect 18187 11852 18705 11880
rect 18187 11849 18199 11852
rect 18141 11843 18199 11849
rect 18693 11849 18705 11852
rect 18739 11849 18751 11883
rect 18693 11843 18751 11849
rect 19061 11883 19119 11889
rect 19061 11849 19073 11883
rect 19107 11880 19119 11883
rect 19705 11883 19763 11889
rect 19107 11852 19380 11880
rect 19107 11849 19119 11852
rect 19061 11843 19119 11849
rect 14936 11784 16896 11812
rect 14829 11775 14887 11781
rect 15286 11744 15292 11756
rect 14200 11716 15292 11744
rect 15286 11704 15292 11716
rect 15344 11704 15350 11756
rect 15470 11744 15476 11756
rect 15431 11716 15476 11744
rect 15470 11704 15476 11716
rect 15528 11744 15534 11756
rect 16868 11744 16896 11784
rect 17770 11772 17776 11824
rect 17828 11812 17834 11824
rect 19352 11812 19380 11852
rect 19705 11849 19717 11883
rect 19751 11880 19763 11883
rect 19886 11880 19892 11892
rect 19751 11852 19892 11880
rect 19751 11849 19763 11852
rect 19705 11843 19763 11849
rect 19886 11840 19892 11852
rect 19944 11840 19950 11892
rect 20254 11840 20260 11892
rect 20312 11880 20318 11892
rect 20349 11883 20407 11889
rect 20349 11880 20361 11883
rect 20312 11852 20361 11880
rect 20312 11840 20318 11852
rect 20349 11849 20361 11852
rect 20395 11849 20407 11883
rect 20349 11843 20407 11849
rect 20809 11883 20867 11889
rect 20809 11849 20821 11883
rect 20855 11880 20867 11883
rect 21634 11880 21640 11892
rect 20855 11852 21640 11880
rect 20855 11849 20867 11852
rect 20809 11843 20867 11849
rect 21634 11840 21640 11852
rect 21692 11840 21698 11892
rect 21174 11812 21180 11824
rect 17828 11784 19288 11812
rect 19352 11784 21180 11812
rect 17828 11772 17834 11784
rect 17954 11744 17960 11756
rect 15528 11716 16804 11744
rect 16868 11716 17960 11744
rect 15528 11704 15534 11716
rect 11977 11679 12035 11685
rect 11977 11645 11989 11679
rect 12023 11645 12035 11679
rect 11977 11639 12035 11645
rect 12069 11679 12127 11685
rect 12069 11645 12081 11679
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 14553 11679 14611 11685
rect 14553 11645 14565 11679
rect 14599 11676 14611 11679
rect 16022 11676 16028 11688
rect 14599 11648 16028 11676
rect 14599 11645 14611 11648
rect 14553 11639 14611 11645
rect 9125 11611 9183 11617
rect 9125 11577 9137 11611
rect 9171 11608 9183 11611
rect 11992 11608 12020 11639
rect 9171 11580 12020 11608
rect 9171 11577 9183 11580
rect 9125 11571 9183 11577
rect 13170 11540 13176 11552
rect 13131 11512 13176 11540
rect 13170 11500 13176 11512
rect 13228 11500 13234 11552
rect 14274 11500 14280 11552
rect 14332 11540 14338 11552
rect 14568 11540 14596 11639
rect 16022 11636 16028 11648
rect 16080 11636 16086 11688
rect 16776 11685 16804 11716
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 19150 11744 19156 11756
rect 19111 11716 19156 11744
rect 19150 11704 19156 11716
rect 19208 11704 19214 11756
rect 16761 11679 16819 11685
rect 16761 11645 16773 11679
rect 16807 11645 16819 11679
rect 16761 11639 16819 11645
rect 17126 11636 17132 11688
rect 17184 11676 17190 11688
rect 19260 11685 19288 11784
rect 18233 11679 18291 11685
rect 18233 11676 18245 11679
rect 17184 11648 18245 11676
rect 17184 11636 17190 11648
rect 18233 11645 18245 11648
rect 18279 11645 18291 11679
rect 18233 11639 18291 11645
rect 19245 11679 19303 11685
rect 19245 11645 19257 11679
rect 19291 11645 19303 11679
rect 19245 11639 19303 11645
rect 17405 11611 17463 11617
rect 17405 11577 17417 11611
rect 17451 11608 17463 11611
rect 19518 11608 19524 11620
rect 17451 11580 19524 11608
rect 17451 11577 17463 11580
rect 17405 11571 17463 11577
rect 19518 11568 19524 11580
rect 19576 11568 19582 11620
rect 14332 11512 14596 11540
rect 14332 11500 14338 11512
rect 15286 11500 15292 11552
rect 15344 11540 15350 11552
rect 19628 11540 19656 11784
rect 21174 11772 21180 11784
rect 21232 11772 21238 11824
rect 19886 11744 19892 11756
rect 19847 11716 19892 11744
rect 19886 11704 19892 11716
rect 19944 11704 19950 11756
rect 20530 11744 20536 11756
rect 20491 11716 20536 11744
rect 20530 11704 20536 11716
rect 20588 11704 20594 11756
rect 20990 11744 20996 11756
rect 20951 11716 20996 11744
rect 20990 11704 20996 11716
rect 21048 11704 21054 11756
rect 15344 11512 19656 11540
rect 15344 11500 15350 11512
rect 21174 11500 21180 11552
rect 21232 11540 21238 11552
rect 21269 11543 21327 11549
rect 21269 11540 21281 11543
rect 21232 11512 21281 11540
rect 21232 11500 21238 11512
rect 21269 11509 21281 11512
rect 21315 11509 21327 11543
rect 21269 11503 21327 11509
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 9582 11296 9588 11348
rect 9640 11336 9646 11348
rect 10321 11339 10379 11345
rect 10321 11336 10333 11339
rect 9640 11308 10333 11336
rect 9640 11296 9646 11308
rect 10321 11305 10333 11308
rect 10367 11305 10379 11339
rect 11330 11336 11336 11348
rect 11291 11308 11336 11336
rect 10321 11299 10379 11305
rect 7926 11160 7932 11212
rect 7984 11200 7990 11212
rect 10336 11200 10364 11299
rect 11330 11296 11336 11308
rect 11388 11296 11394 11348
rect 11790 11296 11796 11348
rect 11848 11336 11854 11348
rect 12621 11339 12679 11345
rect 12621 11336 12633 11339
rect 11848 11308 12633 11336
rect 11848 11296 11854 11308
rect 10689 11203 10747 11209
rect 10689 11200 10701 11203
rect 7984 11172 9076 11200
rect 10336 11172 10701 11200
rect 7984 11160 7990 11172
rect 8386 11092 8392 11144
rect 8444 11132 8450 11144
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 8444 11104 8953 11132
rect 8444 11092 8450 11104
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 9048 11132 9076 11172
rect 10689 11169 10701 11172
rect 10735 11169 10747 11203
rect 10689 11163 10747 11169
rect 9197 11135 9255 11141
rect 9197 11132 9209 11135
rect 9048 11104 9209 11132
rect 8941 11095 8999 11101
rect 9197 11101 9209 11104
rect 9243 11132 9255 11135
rect 9950 11132 9956 11144
rect 9243 11104 9956 11132
rect 9243 11101 9255 11104
rect 9197 11095 9255 11101
rect 9950 11092 9956 11104
rect 10008 11092 10014 11144
rect 10873 11135 10931 11141
rect 10873 11101 10885 11135
rect 10919 11132 10931 11135
rect 11238 11132 11244 11144
rect 10919 11104 11244 11132
rect 10919 11101 10931 11104
rect 10873 11095 10931 11101
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 11900 11132 11928 11308
rect 12621 11305 12633 11308
rect 12667 11305 12679 11339
rect 14458 11336 14464 11348
rect 12621 11299 12679 11305
rect 13648 11308 14464 11336
rect 11974 11228 11980 11280
rect 12032 11268 12038 11280
rect 12345 11271 12403 11277
rect 12345 11268 12357 11271
rect 12032 11240 12357 11268
rect 12032 11228 12038 11240
rect 12345 11237 12357 11240
rect 12391 11268 12403 11271
rect 13648 11268 13676 11308
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 19429 11339 19487 11345
rect 19429 11305 19441 11339
rect 19475 11336 19487 11339
rect 19886 11336 19892 11348
rect 19475 11308 19892 11336
rect 19475 11305 19487 11308
rect 19429 11299 19487 11305
rect 19886 11296 19892 11308
rect 19944 11296 19950 11348
rect 20530 11336 20536 11348
rect 20491 11308 20536 11336
rect 20530 11296 20536 11308
rect 20588 11296 20594 11348
rect 20809 11339 20867 11345
rect 20809 11305 20821 11339
rect 20855 11336 20867 11339
rect 21910 11336 21916 11348
rect 20855 11308 21916 11336
rect 20855 11305 20867 11308
rect 20809 11299 20867 11305
rect 21910 11296 21916 11308
rect 21968 11296 21974 11348
rect 12391 11240 13676 11268
rect 13725 11271 13783 11277
rect 12391 11237 12403 11240
rect 12345 11231 12403 11237
rect 13725 11237 13737 11271
rect 13771 11268 13783 11271
rect 14829 11271 14887 11277
rect 13771 11240 14412 11268
rect 13771 11237 13783 11240
rect 13725 11231 13783 11237
rect 13170 11200 13176 11212
rect 13131 11172 13176 11200
rect 13170 11160 13176 11172
rect 13228 11200 13234 11212
rect 13814 11200 13820 11212
rect 13228 11172 13820 11200
rect 13228 11160 13234 11172
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 14384 11209 14412 11240
rect 14829 11237 14841 11271
rect 14875 11268 14887 11271
rect 15470 11268 15476 11280
rect 14875 11240 15476 11268
rect 14875 11237 14887 11240
rect 14829 11231 14887 11237
rect 15470 11228 15476 11240
rect 15528 11228 15534 11280
rect 20073 11271 20131 11277
rect 20073 11237 20085 11271
rect 20119 11237 20131 11271
rect 20073 11231 20131 11237
rect 14277 11203 14335 11209
rect 14277 11169 14289 11203
rect 14323 11169 14335 11203
rect 14277 11163 14335 11169
rect 14369 11203 14427 11209
rect 14369 11169 14381 11203
rect 14415 11169 14427 11203
rect 14369 11163 14427 11169
rect 13265 11135 13323 11141
rect 13265 11132 13277 11135
rect 11900 11104 13277 11132
rect 13265 11101 13277 11104
rect 13311 11101 13323 11135
rect 14292 11132 14320 11163
rect 14458 11160 14464 11212
rect 14516 11200 14522 11212
rect 19702 11200 19708 11212
rect 14516 11172 19708 11200
rect 14516 11160 14522 11172
rect 19702 11160 19708 11172
rect 19760 11160 19766 11212
rect 20088 11200 20116 11231
rect 20088 11172 21036 11200
rect 14550 11132 14556 11144
rect 14292 11104 14556 11132
rect 13265 11095 13323 11101
rect 14550 11092 14556 11104
rect 14608 11092 14614 11144
rect 19242 11132 19248 11144
rect 19203 11104 19248 11132
rect 19242 11092 19248 11104
rect 19300 11092 19306 11144
rect 19889 11135 19947 11141
rect 19889 11101 19901 11135
rect 19935 11101 19947 11135
rect 19889 11095 19947 11101
rect 20349 11135 20407 11141
rect 20349 11101 20361 11135
rect 20395 11132 20407 11135
rect 20898 11132 20904 11144
rect 20395 11104 20904 11132
rect 20395 11101 20407 11104
rect 20349 11095 20407 11101
rect 10965 11067 11023 11073
rect 10965 11033 10977 11067
rect 11011 11064 11023 11067
rect 11609 11067 11667 11073
rect 11609 11064 11621 11067
rect 11011 11036 11621 11064
rect 11011 11033 11023 11036
rect 10965 11027 11023 11033
rect 11609 11033 11621 11036
rect 11655 11033 11667 11067
rect 11609 11027 11667 11033
rect 13357 11067 13415 11073
rect 13357 11033 13369 11067
rect 13403 11064 13415 11067
rect 13538 11064 13544 11076
rect 13403 11036 13544 11064
rect 13403 11033 13415 11036
rect 13357 11027 13415 11033
rect 13538 11024 13544 11036
rect 13596 11064 13602 11076
rect 14458 11064 14464 11076
rect 13596 11036 14320 11064
rect 14419 11036 14464 11064
rect 13596 11024 13602 11036
rect 14292 10996 14320 11036
rect 14458 11024 14464 11036
rect 14516 11024 14522 11076
rect 15194 11064 15200 11076
rect 14568 11036 15200 11064
rect 14568 10996 14596 11036
rect 15194 11024 15200 11036
rect 15252 11024 15258 11076
rect 17034 11024 17040 11076
rect 17092 11064 17098 11076
rect 17678 11064 17684 11076
rect 17092 11036 17684 11064
rect 17092 11024 17098 11036
rect 17678 11024 17684 11036
rect 17736 11024 17742 11076
rect 19904 11064 19932 11095
rect 20898 11092 20904 11104
rect 20956 11092 20962 11144
rect 21008 11141 21036 11172
rect 20993 11135 21051 11141
rect 20993 11101 21005 11135
rect 21039 11101 21051 11135
rect 20993 11095 21051 11101
rect 21358 11064 21364 11076
rect 19904 11036 21364 11064
rect 21358 11024 21364 11036
rect 21416 11024 21422 11076
rect 14292 10968 14596 10996
rect 1104 10906 21896 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21896 10906
rect 1104 10832 21896 10854
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10229 10795 10287 10801
rect 10229 10792 10241 10795
rect 10100 10764 10241 10792
rect 10100 10752 10106 10764
rect 10229 10761 10241 10764
rect 10275 10761 10287 10795
rect 10229 10755 10287 10761
rect 11238 10752 11244 10804
rect 11296 10792 11302 10804
rect 11517 10795 11575 10801
rect 11517 10792 11529 10795
rect 11296 10764 11529 10792
rect 11296 10752 11302 10764
rect 11517 10761 11529 10764
rect 11563 10761 11575 10795
rect 11517 10755 11575 10761
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 12342 10792 12348 10804
rect 11931 10764 12348 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 12342 10752 12348 10764
rect 12400 10792 12406 10804
rect 12529 10795 12587 10801
rect 12529 10792 12541 10795
rect 12400 10764 12541 10792
rect 12400 10752 12406 10764
rect 12529 10761 12541 10764
rect 12575 10761 12587 10795
rect 15010 10792 15016 10804
rect 14971 10764 15016 10792
rect 12529 10755 12587 10761
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 15470 10792 15476 10804
rect 15431 10764 15476 10792
rect 15470 10752 15476 10764
rect 15528 10752 15534 10804
rect 16669 10795 16727 10801
rect 16669 10761 16681 10795
rect 16715 10792 16727 10795
rect 17126 10792 17132 10804
rect 16715 10764 17132 10792
rect 16715 10761 16727 10764
rect 16669 10755 16727 10761
rect 17126 10752 17132 10764
rect 17184 10752 17190 10804
rect 19242 10752 19248 10804
rect 19300 10792 19306 10804
rect 19337 10795 19395 10801
rect 19337 10792 19349 10795
rect 19300 10764 19349 10792
rect 19300 10752 19306 10764
rect 19337 10761 19349 10764
rect 19383 10761 19395 10795
rect 20898 10792 20904 10804
rect 20859 10764 20904 10792
rect 19337 10755 19395 10761
rect 20898 10752 20904 10764
rect 20956 10752 20962 10804
rect 20990 10752 20996 10804
rect 21048 10792 21054 10804
rect 21177 10795 21235 10801
rect 21177 10792 21189 10795
rect 21048 10764 21189 10792
rect 21048 10752 21054 10764
rect 21177 10761 21189 10764
rect 21223 10761 21235 10795
rect 21177 10755 21235 10761
rect 9585 10727 9643 10733
rect 9585 10693 9597 10727
rect 9631 10724 9643 10727
rect 10318 10724 10324 10736
rect 9631 10696 10324 10724
rect 9631 10693 9643 10696
rect 9585 10687 9643 10693
rect 10318 10684 10324 10696
rect 10376 10724 10382 10736
rect 12989 10727 13047 10733
rect 12989 10724 13001 10727
rect 10376 10696 13001 10724
rect 10376 10684 10382 10696
rect 12989 10693 13001 10696
rect 13035 10693 13047 10727
rect 12989 10687 13047 10693
rect 17770 10684 17776 10736
rect 17828 10733 17834 10736
rect 17828 10724 17840 10733
rect 17828 10696 17873 10724
rect 17828 10687 17840 10696
rect 17828 10684 17834 10687
rect 11974 10656 11980 10668
rect 11935 10628 11980 10656
rect 11974 10616 11980 10628
rect 12032 10616 12038 10668
rect 15381 10659 15439 10665
rect 15381 10625 15393 10659
rect 15427 10656 15439 10659
rect 15746 10656 15752 10668
rect 15427 10628 15752 10656
rect 15427 10625 15439 10628
rect 15381 10619 15439 10625
rect 15746 10616 15752 10628
rect 15804 10616 15810 10668
rect 18601 10659 18659 10665
rect 18601 10625 18613 10659
rect 18647 10656 18659 10659
rect 18874 10656 18880 10668
rect 18647 10628 18880 10656
rect 18647 10625 18659 10628
rect 18601 10619 18659 10625
rect 18874 10616 18880 10628
rect 18932 10616 18938 10668
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10656 19763 10659
rect 20349 10659 20407 10665
rect 20349 10656 20361 10659
rect 19751 10628 20361 10656
rect 19751 10625 19763 10628
rect 19705 10619 19763 10625
rect 20349 10625 20361 10628
rect 20395 10625 20407 10659
rect 20349 10619 20407 10625
rect 21361 10659 21419 10665
rect 21361 10625 21373 10659
rect 21407 10656 21419 10659
rect 21450 10656 21456 10668
rect 21407 10628 21456 10656
rect 21407 10625 21419 10628
rect 21361 10619 21419 10625
rect 21450 10616 21456 10628
rect 21508 10616 21514 10668
rect 12069 10591 12127 10597
rect 12069 10557 12081 10591
rect 12115 10557 12127 10591
rect 12069 10551 12127 10557
rect 9950 10480 9956 10532
rect 10008 10520 10014 10532
rect 12084 10520 12112 10551
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 15565 10591 15623 10597
rect 15565 10588 15577 10591
rect 12584 10560 15577 10588
rect 12584 10548 12590 10560
rect 15565 10557 15577 10560
rect 15611 10557 15623 10591
rect 15565 10551 15623 10557
rect 18049 10591 18107 10597
rect 18049 10557 18061 10591
rect 18095 10588 18107 10591
rect 18506 10588 18512 10600
rect 18095 10560 18512 10588
rect 18095 10557 18107 10560
rect 18049 10551 18107 10557
rect 18506 10548 18512 10560
rect 18564 10548 18570 10600
rect 19518 10548 19524 10600
rect 19576 10588 19582 10600
rect 19797 10591 19855 10597
rect 19797 10588 19809 10591
rect 19576 10560 19809 10588
rect 19576 10548 19582 10560
rect 19797 10557 19809 10560
rect 19843 10557 19855 10591
rect 19978 10588 19984 10600
rect 19939 10560 19984 10588
rect 19797 10551 19855 10557
rect 19978 10548 19984 10560
rect 20036 10548 20042 10600
rect 10008 10492 12112 10520
rect 10008 10480 10014 10492
rect 8297 10455 8355 10461
rect 8297 10421 8309 10455
rect 8343 10452 8355 10455
rect 8386 10452 8392 10464
rect 8343 10424 8392 10452
rect 8343 10421 8355 10424
rect 8297 10415 8355 10421
rect 8386 10412 8392 10424
rect 8444 10412 8450 10464
rect 14274 10452 14280 10464
rect 14235 10424 14280 10452
rect 14274 10412 14280 10424
rect 14332 10412 14338 10464
rect 19061 10455 19119 10461
rect 19061 10421 19073 10455
rect 19107 10452 19119 10455
rect 19886 10452 19892 10464
rect 19107 10424 19892 10452
rect 19107 10421 19119 10424
rect 19061 10415 19119 10421
rect 19886 10412 19892 10424
rect 19944 10412 19950 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 9950 10208 9956 10260
rect 10008 10248 10014 10260
rect 10137 10251 10195 10257
rect 10137 10248 10149 10251
rect 10008 10220 10149 10248
rect 10008 10208 10014 10220
rect 10137 10217 10149 10220
rect 10183 10217 10195 10251
rect 14274 10248 14280 10260
rect 10137 10211 10195 10217
rect 14108 10220 14280 10248
rect 11517 10115 11575 10121
rect 11517 10081 11529 10115
rect 11563 10112 11575 10115
rect 11698 10112 11704 10124
rect 11563 10084 11704 10112
rect 11563 10081 11575 10084
rect 11517 10075 11575 10081
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 11716 10044 11744 10072
rect 12434 10044 12440 10056
rect 11716 10016 12440 10044
rect 12434 10004 12440 10016
rect 12492 10044 12498 10056
rect 14108 10053 14136 10220
rect 14274 10208 14280 10220
rect 14332 10208 14338 10260
rect 15746 10248 15752 10260
rect 15707 10220 15752 10248
rect 15746 10208 15752 10220
rect 15804 10208 15810 10260
rect 17129 10251 17187 10257
rect 17129 10217 17141 10251
rect 17175 10248 17187 10251
rect 17770 10248 17776 10260
rect 17175 10220 17776 10248
rect 17175 10217 17187 10220
rect 17129 10211 17187 10217
rect 17770 10208 17776 10220
rect 17828 10208 17834 10260
rect 19518 10248 19524 10260
rect 19479 10220 19524 10248
rect 19518 10208 19524 10220
rect 19576 10208 19582 10260
rect 16301 10115 16359 10121
rect 16301 10112 16313 10115
rect 15488 10084 16313 10112
rect 13173 10047 13231 10053
rect 13173 10044 13185 10047
rect 12492 10016 13185 10044
rect 12492 10004 12498 10016
rect 13173 10013 13185 10016
rect 13219 10044 13231 10047
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 13219 10016 14105 10044
rect 13219 10013 13231 10016
rect 13173 10007 13231 10013
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 11272 9979 11330 9985
rect 11272 9945 11284 9979
rect 11318 9976 11330 9979
rect 11882 9976 11888 9988
rect 11318 9948 11888 9976
rect 11318 9945 11330 9948
rect 11272 9939 11330 9945
rect 11882 9936 11888 9948
rect 11940 9936 11946 9988
rect 12928 9979 12986 9985
rect 12928 9945 12940 9979
rect 12974 9976 12986 9979
rect 12974 9948 13768 9976
rect 12974 9945 12986 9948
rect 12928 9939 12986 9945
rect 11793 9911 11851 9917
rect 11793 9877 11805 9911
rect 11839 9908 11851 9911
rect 12526 9908 12532 9920
rect 11839 9880 12532 9908
rect 11839 9877 11851 9880
rect 11793 9871 11851 9877
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 13740 9908 13768 9948
rect 13814 9936 13820 9988
rect 13872 9976 13878 9988
rect 14338 9979 14396 9985
rect 14338 9976 14350 9979
rect 13872 9948 14350 9976
rect 13872 9936 13878 9948
rect 14338 9945 14350 9948
rect 14384 9945 14396 9979
rect 14338 9939 14396 9945
rect 14550 9908 14556 9920
rect 13740 9880 14556 9908
rect 14550 9868 14556 9880
rect 14608 9908 14614 9920
rect 15488 9917 15516 10084
rect 16301 10081 16313 10084
rect 16347 10081 16359 10115
rect 20070 10112 20076 10124
rect 20031 10084 20076 10112
rect 16301 10075 16359 10081
rect 20070 10072 20076 10084
rect 20128 10072 20134 10124
rect 18506 10044 18512 10056
rect 18467 10016 18512 10044
rect 18506 10004 18512 10016
rect 18564 10004 18570 10056
rect 19886 10044 19892 10056
rect 19847 10016 19892 10044
rect 19886 10004 19892 10016
rect 19944 10004 19950 10056
rect 19978 10004 19984 10056
rect 20036 10044 20042 10056
rect 20533 10047 20591 10053
rect 20533 10044 20545 10047
rect 20036 10016 20545 10044
rect 20036 10004 20042 10016
rect 20533 10013 20545 10016
rect 20579 10013 20591 10047
rect 20533 10007 20591 10013
rect 18264 9979 18322 9985
rect 18264 9945 18276 9979
rect 18310 9976 18322 9979
rect 21177 9979 21235 9985
rect 21177 9976 21189 9979
rect 18310 9948 21189 9976
rect 18310 9945 18322 9948
rect 18264 9939 18322 9945
rect 21177 9945 21189 9948
rect 21223 9945 21235 9979
rect 21177 9939 21235 9945
rect 15473 9911 15531 9917
rect 15473 9908 15485 9911
rect 14608 9880 15485 9908
rect 14608 9868 14614 9880
rect 15473 9877 15485 9880
rect 15519 9877 15531 9911
rect 16114 9908 16120 9920
rect 16075 9880 16120 9908
rect 15473 9871 15531 9877
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 16209 9911 16267 9917
rect 16209 9877 16221 9911
rect 16255 9908 16267 9911
rect 16853 9911 16911 9917
rect 16853 9908 16865 9911
rect 16255 9880 16865 9908
rect 16255 9877 16267 9880
rect 16209 9871 16267 9877
rect 16853 9877 16865 9880
rect 16899 9908 16911 9911
rect 16942 9908 16948 9920
rect 16899 9880 16948 9908
rect 16899 9877 16911 9880
rect 16853 9871 16911 9877
rect 16942 9868 16948 9880
rect 17000 9908 17006 9920
rect 17218 9908 17224 9920
rect 17000 9880 17224 9908
rect 17000 9868 17006 9880
rect 17218 9868 17224 9880
rect 17276 9868 17282 9920
rect 18046 9868 18052 9920
rect 18104 9908 18110 9920
rect 18785 9911 18843 9917
rect 18785 9908 18797 9911
rect 18104 9880 18797 9908
rect 18104 9868 18110 9880
rect 18785 9877 18797 9880
rect 18831 9908 18843 9911
rect 19981 9911 20039 9917
rect 19981 9908 19993 9911
rect 18831 9880 19993 9908
rect 18831 9877 18843 9880
rect 18785 9871 18843 9877
rect 19981 9877 19993 9880
rect 20027 9877 20039 9911
rect 19981 9871 20039 9877
rect 1104 9818 21896 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21896 9818
rect 1104 9744 21896 9766
rect 11882 9704 11888 9716
rect 11843 9676 11888 9704
rect 11882 9664 11888 9676
rect 11940 9664 11946 9716
rect 15473 9707 15531 9713
rect 15473 9673 15485 9707
rect 15519 9704 15531 9707
rect 16114 9704 16120 9716
rect 15519 9676 16120 9704
rect 15519 9673 15531 9676
rect 15473 9667 15531 9673
rect 16114 9664 16120 9676
rect 16172 9664 16178 9716
rect 19978 9664 19984 9716
rect 20036 9704 20042 9716
rect 20165 9707 20223 9713
rect 20165 9704 20177 9707
rect 20036 9676 20177 9704
rect 20036 9664 20042 9676
rect 20165 9673 20177 9676
rect 20211 9673 20223 9707
rect 20165 9667 20223 9673
rect 21361 9707 21419 9713
rect 21361 9673 21373 9707
rect 21407 9704 21419 9707
rect 21450 9704 21456 9716
rect 21407 9676 21456 9704
rect 21407 9673 21419 9676
rect 21361 9667 21419 9673
rect 21450 9664 21456 9676
rect 21508 9664 21514 9716
rect 13354 9596 13360 9648
rect 13412 9636 13418 9648
rect 14093 9639 14151 9645
rect 14093 9636 14105 9639
rect 13412 9608 14105 9636
rect 13412 9596 13418 9608
rect 14093 9605 14105 9608
rect 14139 9636 14151 9639
rect 14829 9639 14887 9645
rect 14829 9636 14841 9639
rect 14139 9608 14841 9636
rect 14139 9605 14151 9608
rect 14093 9599 14151 9605
rect 14829 9605 14841 9608
rect 14875 9636 14887 9639
rect 20898 9636 20904 9648
rect 14875 9608 20904 9636
rect 14875 9605 14887 9608
rect 14829 9599 14887 9605
rect 20898 9596 20904 9608
rect 20956 9596 20962 9648
rect 12526 9568 12532 9580
rect 12487 9540 12532 9568
rect 12526 9528 12532 9540
rect 12584 9528 12590 9580
rect 16209 9571 16267 9577
rect 16209 9537 16221 9571
rect 16255 9568 16267 9571
rect 16298 9568 16304 9580
rect 16255 9540 16304 9568
rect 16255 9537 16267 9540
rect 16209 9531 16267 9537
rect 16298 9528 16304 9540
rect 16356 9528 16362 9580
rect 19052 9571 19110 9577
rect 19052 9537 19064 9571
rect 19098 9568 19110 9571
rect 19610 9568 19616 9580
rect 19098 9540 19616 9568
rect 19098 9537 19110 9540
rect 19052 9531 19110 9537
rect 19610 9528 19616 9540
rect 19668 9528 19674 9580
rect 20990 9568 20996 9580
rect 20951 9540 20996 9568
rect 20990 9528 20996 9540
rect 21048 9528 21054 9580
rect 13814 9500 13820 9512
rect 13775 9472 13820 9500
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 14001 9503 14059 9509
rect 14001 9469 14013 9503
rect 14047 9500 14059 9503
rect 14366 9500 14372 9512
rect 14047 9472 14372 9500
rect 14047 9469 14059 9472
rect 14001 9463 14059 9469
rect 14366 9460 14372 9472
rect 14424 9500 14430 9512
rect 14826 9500 14832 9512
rect 14424 9472 14832 9500
rect 14424 9460 14430 9472
rect 14826 9460 14832 9472
rect 14884 9460 14890 9512
rect 18230 9460 18236 9512
rect 18288 9500 18294 9512
rect 18506 9500 18512 9512
rect 18288 9472 18512 9500
rect 18288 9460 18294 9472
rect 18506 9460 18512 9472
rect 18564 9500 18570 9512
rect 18785 9503 18843 9509
rect 18785 9500 18797 9503
rect 18564 9472 18797 9500
rect 18564 9460 18570 9472
rect 18785 9469 18797 9472
rect 18831 9469 18843 9503
rect 18785 9463 18843 9469
rect 14458 9432 14464 9444
rect 14419 9404 14464 9432
rect 14458 9392 14464 9404
rect 14516 9392 14522 9444
rect 15930 9392 15936 9444
rect 15988 9432 15994 9444
rect 16025 9435 16083 9441
rect 16025 9432 16037 9435
rect 15988 9404 16037 9432
rect 15988 9392 15994 9404
rect 16025 9401 16037 9404
rect 16071 9401 16083 9435
rect 16025 9395 16083 9401
rect 20809 9435 20867 9441
rect 20809 9401 20821 9435
rect 20855 9432 20867 9435
rect 21266 9432 21272 9444
rect 20855 9404 21272 9432
rect 20855 9401 20867 9404
rect 20809 9395 20867 9401
rect 21266 9392 21272 9404
rect 21324 9392 21330 9444
rect 20530 9364 20536 9376
rect 20491 9336 20536 9364
rect 20530 9324 20536 9336
rect 20588 9324 20594 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 11793 9163 11851 9169
rect 11793 9129 11805 9163
rect 11839 9160 11851 9163
rect 12250 9160 12256 9172
rect 11839 9132 12256 9160
rect 11839 9129 11851 9132
rect 11793 9123 11851 9129
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 13446 9160 13452 9172
rect 13407 9132 13452 9160
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 16298 9160 16304 9172
rect 16259 9132 16304 9160
rect 16298 9120 16304 9132
rect 16356 9120 16362 9172
rect 19610 9160 19616 9172
rect 19571 9132 19616 9160
rect 19610 9120 19616 9132
rect 19668 9120 19674 9172
rect 20993 9163 21051 9169
rect 20993 9129 21005 9163
rect 21039 9160 21051 9163
rect 21818 9160 21824 9172
rect 21039 9132 21824 9160
rect 21039 9129 21051 9132
rect 20993 9123 21051 9129
rect 21818 9120 21824 9132
rect 21876 9120 21882 9172
rect 11146 8916 11152 8968
rect 11204 8956 11210 8968
rect 11609 8959 11667 8965
rect 11609 8956 11621 8959
rect 11204 8928 11621 8956
rect 11204 8916 11210 8928
rect 11609 8925 11621 8928
rect 11655 8925 11667 8959
rect 11609 8919 11667 8925
rect 13265 8959 13323 8965
rect 13265 8925 13277 8959
rect 13311 8956 13323 8959
rect 13446 8956 13452 8968
rect 13311 8928 13452 8956
rect 13311 8925 13323 8928
rect 13265 8919 13323 8925
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 16485 8959 16543 8965
rect 16485 8925 16497 8959
rect 16531 8956 16543 8959
rect 16942 8956 16948 8968
rect 16531 8928 16948 8956
rect 16531 8925 16543 8928
rect 16485 8919 16543 8925
rect 16942 8916 16948 8928
rect 17000 8916 17006 8968
rect 19610 8916 19616 8968
rect 19668 8956 19674 8968
rect 20070 8956 20076 8968
rect 19668 8928 20076 8956
rect 19668 8916 19674 8928
rect 20070 8916 20076 8928
rect 20128 8956 20134 8968
rect 20257 8959 20315 8965
rect 20257 8956 20269 8959
rect 20128 8928 20269 8956
rect 20128 8916 20134 8928
rect 20257 8925 20269 8928
rect 20303 8925 20315 8959
rect 20530 8956 20536 8968
rect 20491 8928 20536 8956
rect 20257 8919 20315 8925
rect 20530 8916 20536 8928
rect 20588 8916 20594 8968
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 21177 8959 21235 8965
rect 21177 8956 21189 8959
rect 20680 8928 21189 8956
rect 20680 8916 20686 8928
rect 21177 8925 21189 8928
rect 21223 8925 21235 8959
rect 21177 8919 21235 8925
rect 14826 8820 14832 8832
rect 14787 8792 14832 8820
rect 14826 8780 14832 8792
rect 14884 8780 14890 8832
rect 17310 8780 17316 8832
rect 17368 8820 17374 8832
rect 17405 8823 17463 8829
rect 17405 8820 17417 8823
rect 17368 8792 17417 8820
rect 17368 8780 17374 8792
rect 17405 8789 17417 8792
rect 17451 8789 17463 8823
rect 20714 8820 20720 8832
rect 20675 8792 20720 8820
rect 17405 8783 17463 8789
rect 20714 8780 20720 8792
rect 20772 8780 20778 8832
rect 1104 8730 21896 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21896 8730
rect 1104 8656 21896 8678
rect 11146 8616 11152 8628
rect 11107 8588 11152 8616
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 13446 8616 13452 8628
rect 13407 8588 13452 8616
rect 13446 8576 13452 8588
rect 13504 8576 13510 8628
rect 19610 8616 19616 8628
rect 19571 8588 19616 8616
rect 19610 8576 19616 8588
rect 19668 8576 19674 8628
rect 20073 8619 20131 8625
rect 20073 8585 20085 8619
rect 20119 8616 20131 8619
rect 20622 8616 20628 8628
rect 20119 8588 20628 8616
rect 20119 8585 20131 8588
rect 20073 8579 20131 8585
rect 20622 8576 20628 8588
rect 20680 8576 20686 8628
rect 20809 8619 20867 8625
rect 20809 8585 20821 8619
rect 20855 8585 20867 8619
rect 21358 8616 21364 8628
rect 21319 8588 21364 8616
rect 20809 8579 20867 8585
rect 18690 8508 18696 8560
rect 18748 8548 18754 8560
rect 19242 8548 19248 8560
rect 18748 8520 19248 8548
rect 18748 8508 18754 8520
rect 19242 8508 19248 8520
rect 19300 8508 19306 8560
rect 9398 8480 9404 8492
rect 9359 8452 9404 8480
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 10965 8483 11023 8489
rect 10965 8449 10977 8483
rect 11011 8480 11023 8483
rect 11238 8480 11244 8492
rect 11011 8452 11244 8480
rect 11011 8449 11023 8452
rect 10965 8443 11023 8449
rect 11238 8440 11244 8452
rect 11296 8440 11302 8492
rect 11514 8480 11520 8492
rect 11475 8452 11520 8480
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 13633 8483 13691 8489
rect 13633 8449 13645 8483
rect 13679 8480 13691 8483
rect 13814 8480 13820 8492
rect 13679 8452 13820 8480
rect 13679 8449 13691 8452
rect 13633 8443 13691 8449
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 15286 8440 15292 8492
rect 15344 8480 15350 8492
rect 15473 8483 15531 8489
rect 15473 8480 15485 8483
rect 15344 8452 15485 8480
rect 15344 8440 15350 8452
rect 15473 8449 15485 8452
rect 15519 8449 15531 8483
rect 17126 8480 17132 8492
rect 17087 8452 17132 8480
rect 15473 8443 15531 8449
rect 17126 8440 17132 8452
rect 17184 8440 17190 8492
rect 18500 8483 18558 8489
rect 18500 8449 18512 8483
rect 18546 8480 18558 8483
rect 19794 8480 19800 8492
rect 18546 8452 19800 8480
rect 18546 8449 18558 8452
rect 18500 8443 18558 8449
rect 19794 8440 19800 8452
rect 19852 8440 19858 8492
rect 19889 8483 19947 8489
rect 19889 8449 19901 8483
rect 19935 8449 19947 8483
rect 19889 8443 19947 8449
rect 20533 8483 20591 8489
rect 20533 8449 20545 8483
rect 20579 8480 20591 8483
rect 20824 8480 20852 8579
rect 21358 8576 21364 8588
rect 21416 8576 21422 8628
rect 20579 8452 20852 8480
rect 20993 8483 21051 8489
rect 20579 8449 20591 8452
rect 20533 8443 20591 8449
rect 20993 8449 21005 8483
rect 21039 8480 21051 8483
rect 21082 8480 21088 8492
rect 21039 8452 21088 8480
rect 21039 8449 21051 8452
rect 20993 8443 21051 8449
rect 12437 8415 12495 8421
rect 12437 8381 12449 8415
rect 12483 8412 12495 8415
rect 12526 8412 12532 8424
rect 12483 8384 12532 8412
rect 12483 8381 12495 8384
rect 12437 8375 12495 8381
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 14458 8412 14464 8424
rect 14419 8384 14464 8412
rect 14458 8372 14464 8384
rect 14516 8372 14522 8424
rect 18230 8412 18236 8424
rect 18191 8384 18236 8412
rect 18230 8372 18236 8384
rect 18288 8372 18294 8424
rect 19904 8412 19932 8443
rect 21082 8440 21088 8452
rect 21140 8440 21146 8492
rect 21376 8412 21404 8576
rect 19904 8384 21404 8412
rect 19242 8304 19248 8356
rect 19300 8344 19306 8356
rect 20349 8347 20407 8353
rect 20349 8344 20361 8347
rect 19300 8316 20361 8344
rect 19300 8304 19306 8316
rect 20349 8313 20361 8316
rect 20395 8313 20407 8347
rect 20349 8307 20407 8313
rect 10042 8276 10048 8288
rect 10003 8248 10048 8276
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 12158 8276 12164 8288
rect 12119 8248 12164 8276
rect 12158 8236 12164 8248
rect 12216 8236 12222 8288
rect 16114 8276 16120 8288
rect 16075 8248 16120 8276
rect 16114 8236 16120 8248
rect 16172 8236 16178 8288
rect 17770 8276 17776 8288
rect 17731 8248 17776 8276
rect 17770 8236 17776 8248
rect 17828 8236 17834 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 19794 8032 19800 8084
rect 19852 8072 19858 8084
rect 19889 8075 19947 8081
rect 19889 8072 19901 8075
rect 19852 8044 19901 8072
rect 19852 8032 19858 8044
rect 19889 8041 19901 8044
rect 19935 8041 19947 8075
rect 19889 8035 19947 8041
rect 20806 8004 20812 8016
rect 20767 7976 20812 8004
rect 20806 7964 20812 7976
rect 20864 7964 20870 8016
rect 21358 7936 21364 7948
rect 20180 7908 21364 7936
rect 8386 7828 8392 7880
rect 8444 7868 8450 7880
rect 10042 7877 10048 7880
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 8444 7840 9781 7868
rect 8444 7828 8450 7840
rect 9769 7837 9781 7840
rect 9815 7837 9827 7871
rect 10036 7868 10048 7877
rect 10003 7840 10048 7868
rect 9769 7831 9827 7837
rect 10036 7831 10048 7840
rect 10042 7828 10048 7831
rect 10100 7828 10106 7880
rect 11701 7871 11759 7877
rect 11701 7837 11713 7871
rect 11747 7868 11759 7871
rect 12434 7868 12440 7880
rect 11747 7840 12440 7868
rect 11747 7837 11759 7840
rect 11701 7831 11759 7837
rect 12434 7828 12440 7840
rect 12492 7868 12498 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 12492 7840 14105 7868
rect 12492 7828 12498 7840
rect 14093 7837 14105 7840
rect 14139 7868 14151 7871
rect 15749 7871 15807 7877
rect 15749 7868 15761 7871
rect 14139 7840 15761 7868
rect 14139 7837 14151 7840
rect 14093 7831 14151 7837
rect 15749 7837 15761 7840
rect 15795 7868 15807 7871
rect 17405 7871 17463 7877
rect 17405 7868 17417 7871
rect 15795 7840 17417 7868
rect 15795 7837 15807 7840
rect 15749 7831 15807 7837
rect 17405 7837 17417 7840
rect 17451 7868 17463 7871
rect 18230 7868 18236 7880
rect 17451 7840 18236 7868
rect 17451 7837 17463 7840
rect 17405 7831 17463 7837
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 20180 7877 20208 7908
rect 21358 7896 21364 7908
rect 21416 7896 21422 7948
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 18800 7840 19257 7868
rect 11514 7760 11520 7812
rect 11572 7760 11578 7812
rect 11968 7803 12026 7809
rect 11968 7769 11980 7803
rect 12014 7800 12026 7803
rect 12158 7800 12164 7812
rect 12014 7772 12164 7800
rect 12014 7769 12026 7772
rect 11968 7763 12026 7769
rect 12158 7760 12164 7772
rect 12216 7760 12222 7812
rect 13722 7760 13728 7812
rect 13780 7800 13786 7812
rect 14338 7803 14396 7809
rect 14338 7800 14350 7803
rect 13780 7772 14350 7800
rect 13780 7760 13786 7772
rect 14338 7769 14350 7772
rect 14384 7769 14396 7803
rect 14338 7763 14396 7769
rect 16016 7803 16074 7809
rect 16016 7769 16028 7803
rect 16062 7800 16074 7803
rect 16114 7800 16120 7812
rect 16062 7772 16120 7800
rect 16062 7769 16074 7772
rect 16016 7763 16074 7769
rect 16114 7760 16120 7772
rect 16172 7760 16178 7812
rect 17672 7803 17730 7809
rect 17672 7769 17684 7803
rect 17718 7800 17730 7803
rect 17770 7800 17776 7812
rect 17718 7772 17776 7800
rect 17718 7769 17730 7772
rect 17672 7763 17730 7769
rect 17770 7760 17776 7772
rect 17828 7760 17834 7812
rect 11149 7735 11207 7741
rect 11149 7701 11161 7735
rect 11195 7732 11207 7735
rect 11532 7732 11560 7760
rect 12066 7732 12072 7744
rect 11195 7704 12072 7732
rect 11195 7701 11207 7704
rect 11149 7695 11207 7701
rect 12066 7692 12072 7704
rect 12124 7692 12130 7744
rect 13081 7735 13139 7741
rect 13081 7701 13093 7735
rect 13127 7732 13139 7735
rect 13170 7732 13176 7744
rect 13127 7704 13176 7732
rect 13127 7701 13139 7704
rect 13081 7695 13139 7701
rect 13170 7692 13176 7704
rect 13228 7692 13234 7744
rect 15286 7692 15292 7744
rect 15344 7732 15350 7744
rect 15473 7735 15531 7741
rect 15473 7732 15485 7735
rect 15344 7704 15485 7732
rect 15344 7692 15350 7704
rect 15473 7701 15485 7704
rect 15519 7701 15531 7735
rect 17126 7732 17132 7744
rect 17087 7704 17132 7732
rect 15473 7695 15531 7701
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 17586 7692 17592 7744
rect 17644 7732 17650 7744
rect 18800 7741 18828 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7837 20223 7871
rect 20165 7831 20223 7837
rect 20714 7828 20720 7880
rect 20772 7868 20778 7880
rect 20993 7871 21051 7877
rect 20993 7868 21005 7871
rect 20772 7840 21005 7868
rect 20772 7828 20778 7840
rect 20993 7837 21005 7840
rect 21039 7837 21051 7871
rect 20993 7831 21051 7837
rect 18785 7735 18843 7741
rect 18785 7732 18797 7735
rect 17644 7704 18797 7732
rect 17644 7692 17650 7704
rect 18785 7701 18797 7704
rect 18831 7701 18843 7735
rect 18785 7695 18843 7701
rect 20349 7735 20407 7741
rect 20349 7701 20361 7735
rect 20395 7732 20407 7735
rect 20714 7732 20720 7744
rect 20395 7704 20720 7732
rect 20395 7701 20407 7704
rect 20349 7695 20407 7701
rect 20714 7692 20720 7704
rect 20772 7692 20778 7744
rect 1104 7642 21896 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21896 7642
rect 1104 7568 21896 7590
rect 9398 7528 9404 7540
rect 9359 7500 9404 7528
rect 9398 7488 9404 7500
rect 9456 7488 9462 7540
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11296 7500 11529 7528
rect 11296 7488 11302 7500
rect 11517 7497 11529 7500
rect 11563 7497 11575 7531
rect 11517 7491 11575 7497
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 12526 7528 12532 7540
rect 11931 7500 12532 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 13722 7528 13728 7540
rect 13683 7500 13728 7528
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 13814 7488 13820 7540
rect 13872 7528 13878 7540
rect 14001 7531 14059 7537
rect 14001 7528 14013 7531
rect 13872 7500 14013 7528
rect 13872 7488 13878 7500
rect 14001 7497 14013 7500
rect 14047 7497 14059 7531
rect 14001 7491 14059 7497
rect 14369 7531 14427 7537
rect 14369 7497 14381 7531
rect 14415 7528 14427 7531
rect 14458 7528 14464 7540
rect 14415 7500 14464 7528
rect 14415 7497 14427 7500
rect 14369 7491 14427 7497
rect 14458 7488 14464 7500
rect 14516 7488 14522 7540
rect 15470 7528 15476 7540
rect 15431 7500 15476 7528
rect 15470 7488 15476 7500
rect 15528 7488 15534 7540
rect 16942 7528 16948 7540
rect 16903 7500 16948 7528
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17310 7528 17316 7540
rect 17271 7500 17316 7528
rect 17310 7488 17316 7500
rect 17368 7488 17374 7540
rect 17405 7531 17463 7537
rect 17405 7497 17417 7531
rect 17451 7528 17463 7531
rect 17957 7531 18015 7537
rect 17957 7528 17969 7531
rect 17451 7500 17969 7528
rect 17451 7497 17463 7500
rect 17405 7491 17463 7497
rect 17957 7497 17969 7500
rect 18003 7497 18015 7531
rect 17957 7491 18015 7497
rect 18325 7531 18383 7537
rect 18325 7497 18337 7531
rect 18371 7528 18383 7531
rect 20073 7531 20131 7537
rect 18371 7500 20024 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 8386 7460 8392 7472
rect 8036 7432 8392 7460
rect 8036 7401 8064 7432
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 13170 7420 13176 7472
rect 13228 7460 13234 7472
rect 13228 7432 15608 7460
rect 13228 7420 13234 7432
rect 8294 7401 8300 7404
rect 8021 7395 8079 7401
rect 8021 7361 8033 7395
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 8288 7355 8300 7401
rect 8352 7392 8358 7404
rect 13081 7395 13139 7401
rect 8352 7364 8388 7392
rect 8294 7352 8300 7355
rect 8352 7352 8358 7364
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 13188 7392 13216 7420
rect 13127 7364 13216 7392
rect 15381 7395 15439 7401
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 15381 7361 15393 7395
rect 15427 7361 15439 7395
rect 15381 7355 15439 7361
rect 11974 7324 11980 7336
rect 11935 7296 11980 7324
rect 11974 7284 11980 7296
rect 12032 7284 12038 7336
rect 12066 7284 12072 7336
rect 12124 7324 12130 7336
rect 14461 7327 14519 7333
rect 12124 7296 12169 7324
rect 12124 7284 12130 7296
rect 14461 7293 14473 7327
rect 14507 7293 14519 7327
rect 14461 7287 14519 7293
rect 14645 7327 14703 7333
rect 14645 7293 14657 7327
rect 14691 7324 14703 7327
rect 15286 7324 15292 7336
rect 14691 7296 15292 7324
rect 14691 7293 14703 7296
rect 14645 7287 14703 7293
rect 14476 7256 14504 7287
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 15013 7259 15071 7265
rect 15013 7256 15025 7259
rect 14476 7228 15025 7256
rect 15013 7225 15025 7228
rect 15059 7225 15071 7259
rect 15396 7256 15424 7355
rect 15580 7333 15608 7432
rect 17126 7420 17132 7472
rect 17184 7460 17190 7472
rect 17184 7432 18552 7460
rect 17184 7420 17190 7432
rect 15565 7327 15623 7333
rect 15565 7293 15577 7327
rect 15611 7293 15623 7327
rect 17586 7324 17592 7336
rect 17547 7296 17592 7324
rect 15565 7287 15623 7293
rect 17586 7284 17592 7296
rect 17644 7284 17650 7336
rect 18046 7284 18052 7336
rect 18104 7324 18110 7336
rect 18524 7333 18552 7432
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7392 19671 7395
rect 19886 7392 19892 7404
rect 19659 7364 19892 7392
rect 19659 7361 19671 7364
rect 19613 7355 19671 7361
rect 19886 7352 19892 7364
rect 19944 7352 19950 7404
rect 18417 7327 18475 7333
rect 18417 7324 18429 7327
rect 18104 7296 18429 7324
rect 18104 7284 18110 7296
rect 18417 7293 18429 7296
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 18509 7327 18567 7333
rect 18509 7293 18521 7327
rect 18555 7293 18567 7327
rect 19996 7324 20024 7500
rect 20073 7497 20085 7531
rect 20119 7497 20131 7531
rect 20073 7491 20131 7497
rect 20088 7460 20116 7491
rect 20990 7488 20996 7540
rect 21048 7528 21054 7540
rect 21177 7531 21235 7537
rect 21177 7528 21189 7531
rect 21048 7500 21189 7528
rect 21048 7488 21054 7500
rect 21177 7497 21189 7500
rect 21223 7497 21235 7531
rect 21177 7491 21235 7497
rect 20438 7460 20444 7472
rect 20088 7432 20444 7460
rect 20438 7420 20444 7432
rect 20496 7420 20502 7472
rect 20901 7463 20959 7469
rect 20901 7429 20913 7463
rect 20947 7460 20959 7463
rect 21082 7460 21088 7472
rect 20947 7432 21088 7460
rect 20947 7429 20959 7432
rect 20901 7423 20959 7429
rect 21082 7420 21088 7432
rect 21140 7420 21146 7472
rect 20533 7395 20591 7401
rect 20533 7361 20545 7395
rect 20579 7392 20591 7395
rect 21174 7392 21180 7404
rect 20579 7364 21180 7392
rect 20579 7361 20591 7364
rect 20533 7355 20591 7361
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7392 21419 7395
rect 21542 7392 21548 7404
rect 21407 7364 21548 7392
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 21542 7352 21548 7364
rect 21600 7352 21606 7404
rect 20898 7324 20904 7336
rect 19996 7296 20904 7324
rect 18509 7287 18567 7293
rect 20898 7284 20904 7296
rect 20956 7284 20962 7336
rect 21082 7256 21088 7268
rect 15396 7228 21088 7256
rect 15013 7219 15071 7225
rect 21082 7216 21088 7228
rect 21140 7216 21146 7268
rect 17862 7148 17868 7200
rect 17920 7188 17926 7200
rect 20349 7191 20407 7197
rect 20349 7188 20361 7191
rect 17920 7160 20361 7188
rect 17920 7148 17926 7160
rect 20349 7157 20361 7160
rect 20395 7157 20407 7191
rect 20349 7151 20407 7157
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 11885 6987 11943 6993
rect 11885 6953 11897 6987
rect 11931 6984 11943 6987
rect 11974 6984 11980 6996
rect 11931 6956 11980 6984
rect 11931 6953 11943 6956
rect 11885 6947 11943 6953
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 21361 6987 21419 6993
rect 21361 6953 21373 6987
rect 21407 6984 21419 6987
rect 21542 6984 21548 6996
rect 21407 6956 21548 6984
rect 21407 6953 21419 6956
rect 21361 6947 21419 6953
rect 21542 6944 21548 6956
rect 21600 6944 21606 6996
rect 20349 6919 20407 6925
rect 20349 6885 20361 6919
rect 20395 6885 20407 6919
rect 20349 6879 20407 6885
rect 9398 6808 9404 6860
rect 9456 6848 9462 6860
rect 11241 6851 11299 6857
rect 11241 6848 11253 6851
rect 9456 6820 11253 6848
rect 9456 6808 9462 6820
rect 11241 6817 11253 6820
rect 11287 6817 11299 6851
rect 11241 6811 11299 6817
rect 16390 6808 16396 6860
rect 16448 6848 16454 6860
rect 20364 6848 20392 6879
rect 16448 6820 20392 6848
rect 16448 6808 16454 6820
rect 14829 6783 14887 6789
rect 14829 6780 14841 6783
rect 12406 6752 14841 6780
rect 12406 6712 12434 6752
rect 14829 6749 14841 6752
rect 14875 6780 14887 6783
rect 15470 6780 15476 6792
rect 14875 6752 15476 6780
rect 14875 6749 14887 6752
rect 14829 6743 14887 6749
rect 15470 6740 15476 6752
rect 15528 6780 15534 6792
rect 17773 6783 17831 6789
rect 17773 6780 17785 6783
rect 15528 6752 17785 6780
rect 15528 6740 15534 6752
rect 17773 6749 17785 6752
rect 17819 6780 17831 6783
rect 18046 6780 18052 6792
rect 17819 6752 18052 6780
rect 17819 6749 17831 6752
rect 17773 6743 17831 6749
rect 18046 6740 18052 6752
rect 18104 6740 18110 6792
rect 20438 6740 20444 6792
rect 20496 6780 20502 6792
rect 20533 6783 20591 6789
rect 20533 6780 20545 6783
rect 20496 6752 20545 6780
rect 20496 6740 20502 6752
rect 20533 6749 20545 6752
rect 20579 6749 20591 6783
rect 20533 6743 20591 6749
rect 20714 6740 20720 6792
rect 20772 6780 20778 6792
rect 20993 6783 21051 6789
rect 20993 6780 21005 6783
rect 20772 6752 21005 6780
rect 20772 6740 20778 6752
rect 20993 6749 21005 6752
rect 21039 6749 21051 6783
rect 20993 6743 21051 6749
rect 20162 6712 20168 6724
rect 11440 6684 12434 6712
rect 14752 6684 20168 6712
rect 3970 6604 3976 6656
rect 4028 6644 4034 6656
rect 11440 6653 11468 6684
rect 10781 6647 10839 6653
rect 10781 6644 10793 6647
rect 4028 6616 10793 6644
rect 4028 6604 4034 6616
rect 10781 6613 10793 6616
rect 10827 6644 10839 6647
rect 11425 6647 11483 6653
rect 11425 6644 11437 6647
rect 10827 6616 11437 6644
rect 10827 6613 10839 6616
rect 10781 6607 10839 6613
rect 11425 6613 11437 6616
rect 11471 6613 11483 6647
rect 11425 6607 11483 6613
rect 11517 6647 11575 6653
rect 11517 6613 11529 6647
rect 11563 6644 11575 6647
rect 14752 6644 14780 6684
rect 20162 6672 20168 6684
rect 20220 6672 20226 6724
rect 20272 6684 20852 6712
rect 11563 6616 14780 6644
rect 11563 6613 11575 6616
rect 11517 6607 11575 6613
rect 17494 6604 17500 6656
rect 17552 6644 17558 6656
rect 20272 6644 20300 6684
rect 20824 6653 20852 6684
rect 17552 6616 20300 6644
rect 20809 6647 20867 6653
rect 17552 6604 17558 6616
rect 20809 6613 20821 6647
rect 20855 6613 20867 6647
rect 20809 6607 20867 6613
rect 1104 6554 21896 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21896 6554
rect 1104 6480 21896 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 8294 6440 8300 6452
rect 1627 6412 8300 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 20441 6443 20499 6449
rect 20441 6409 20453 6443
rect 20487 6409 20499 6443
rect 21174 6440 21180 6452
rect 21135 6412 21180 6440
rect 20441 6403 20499 6409
rect 1394 6304 1400 6316
rect 1355 6276 1400 6304
rect 1394 6264 1400 6276
rect 1452 6304 1458 6316
rect 1857 6307 1915 6313
rect 1857 6304 1869 6307
rect 1452 6276 1869 6304
rect 1452 6264 1458 6276
rect 1857 6273 1869 6276
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 19981 6307 20039 6313
rect 19981 6273 19993 6307
rect 20027 6304 20039 6307
rect 20254 6304 20260 6316
rect 20027 6276 20260 6304
rect 20027 6273 20039 6276
rect 19981 6267 20039 6273
rect 20254 6264 20260 6276
rect 20312 6264 20318 6316
rect 20456 6304 20484 6403
rect 21174 6400 21180 6412
rect 21232 6400 21238 6452
rect 20530 6332 20536 6384
rect 20588 6372 20594 6384
rect 20588 6344 21404 6372
rect 20588 6332 20594 6344
rect 21376 6313 21404 6344
rect 20901 6307 20959 6313
rect 20901 6304 20913 6307
rect 20456 6276 20913 6304
rect 20901 6273 20913 6276
rect 20947 6273 20959 6307
rect 20901 6267 20959 6273
rect 21361 6307 21419 6313
rect 21361 6273 21373 6307
rect 21407 6273 21419 6307
rect 21361 6267 21419 6273
rect 19613 6239 19671 6245
rect 19613 6205 19625 6239
rect 19659 6236 19671 6239
rect 20530 6236 20536 6248
rect 19659 6208 20536 6236
rect 19659 6205 19671 6208
rect 19613 6199 19671 6205
rect 20530 6196 20536 6208
rect 20588 6196 20594 6248
rect 14642 6128 14648 6180
rect 14700 6168 14706 6180
rect 20717 6171 20775 6177
rect 20717 6168 20729 6171
rect 14700 6140 20729 6168
rect 14700 6128 14706 6140
rect 20717 6137 20729 6140
rect 20763 6137 20775 6171
rect 20717 6131 20775 6137
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 14734 5788 14740 5840
rect 14792 5828 14798 5840
rect 20809 5831 20867 5837
rect 20809 5828 20821 5831
rect 14792 5800 20821 5828
rect 14792 5788 14798 5800
rect 20809 5797 20821 5800
rect 20855 5797 20867 5831
rect 20809 5791 20867 5797
rect 20073 5695 20131 5701
rect 20073 5661 20085 5695
rect 20119 5692 20131 5695
rect 20346 5692 20352 5704
rect 20119 5664 20352 5692
rect 20119 5661 20131 5664
rect 20073 5655 20131 5661
rect 20346 5652 20352 5664
rect 20404 5652 20410 5704
rect 20993 5627 21051 5633
rect 20993 5624 21005 5627
rect 20548 5596 21005 5624
rect 20548 5565 20576 5596
rect 20993 5593 21005 5596
rect 21039 5593 21051 5627
rect 20993 5587 21051 5593
rect 20533 5559 20591 5565
rect 20533 5525 20545 5559
rect 20579 5525 20591 5559
rect 20533 5519 20591 5525
rect 1104 5466 21896 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21896 5466
rect 1104 5392 21896 5414
rect 20714 5352 20720 5364
rect 20675 5324 20720 5352
rect 20714 5312 20720 5324
rect 20772 5312 20778 5364
rect 20898 5312 20904 5364
rect 20956 5352 20962 5364
rect 21177 5355 21235 5361
rect 21177 5352 21189 5355
rect 20956 5324 21189 5352
rect 20956 5312 20962 5324
rect 21177 5321 21189 5324
rect 21223 5321 21235 5355
rect 21177 5315 21235 5321
rect 20441 5287 20499 5293
rect 20441 5253 20453 5287
rect 20487 5284 20499 5287
rect 20622 5284 20628 5296
rect 20487 5256 20628 5284
rect 20487 5253 20499 5256
rect 20441 5247 20499 5253
rect 20622 5244 20628 5256
rect 20680 5284 20686 5296
rect 20680 5256 21404 5284
rect 20680 5244 20686 5256
rect 20898 5216 20904 5228
rect 20859 5188 20904 5216
rect 20898 5176 20904 5188
rect 20956 5176 20962 5228
rect 21376 5225 21404 5256
rect 21361 5219 21419 5225
rect 21361 5185 21373 5219
rect 21407 5185 21419 5219
rect 21361 5179 21419 5185
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 20162 4768 20168 4820
rect 20220 4808 20226 4820
rect 20257 4811 20315 4817
rect 20257 4808 20269 4811
rect 20220 4780 20269 4808
rect 20220 4768 20226 4780
rect 20257 4777 20269 4780
rect 20303 4777 20315 4811
rect 20898 4808 20904 4820
rect 20859 4780 20904 4808
rect 20257 4771 20315 4777
rect 20898 4768 20904 4780
rect 20956 4768 20962 4820
rect 21082 4768 21088 4820
rect 21140 4808 21146 4820
rect 21177 4811 21235 4817
rect 21177 4808 21189 4811
rect 21140 4780 21189 4808
rect 21140 4768 21146 4780
rect 21177 4777 21189 4780
rect 21223 4777 21235 4811
rect 21177 4771 21235 4777
rect 20438 4604 20444 4616
rect 20399 4576 20444 4604
rect 20438 4564 20444 4576
rect 20496 4564 20502 4616
rect 20714 4604 20720 4616
rect 20675 4576 20720 4604
rect 20714 4564 20720 4576
rect 20772 4564 20778 4616
rect 21358 4604 21364 4616
rect 21319 4576 21364 4604
rect 21358 4564 21364 4576
rect 21416 4564 21422 4616
rect 19981 4539 20039 4545
rect 19981 4505 19993 4539
rect 20027 4536 20039 4539
rect 20732 4536 20760 4564
rect 20027 4508 20760 4536
rect 20027 4505 20039 4508
rect 19981 4499 20039 4505
rect 1104 4378 21896 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21896 4378
rect 1104 4304 21896 4326
rect 20438 4224 20444 4276
rect 20496 4264 20502 4276
rect 20533 4267 20591 4273
rect 20533 4264 20545 4267
rect 20496 4236 20545 4264
rect 20496 4224 20502 4236
rect 20533 4233 20545 4236
rect 20579 4233 20591 4267
rect 21174 4264 21180 4276
rect 21135 4236 21180 4264
rect 20533 4227 20591 4233
rect 21174 4224 21180 4236
rect 21232 4224 21238 4276
rect 21266 4196 21272 4208
rect 19904 4168 21272 4196
rect 19904 4137 19932 4168
rect 21266 4156 21272 4168
rect 21324 4156 21330 4208
rect 19889 4131 19947 4137
rect 19889 4097 19901 4131
rect 19935 4097 19947 4131
rect 19889 4091 19947 4097
rect 20257 4131 20315 4137
rect 20257 4097 20269 4131
rect 20303 4128 20315 4131
rect 21358 4128 21364 4140
rect 20303 4100 21364 4128
rect 20303 4097 20315 4100
rect 20257 4091 20315 4097
rect 21358 4088 21364 4100
rect 21416 4088 21422 4140
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 17954 3612 17960 3664
rect 18012 3652 18018 3664
rect 19981 3655 20039 3661
rect 19981 3652 19993 3655
rect 18012 3624 19993 3652
rect 18012 3612 18018 3624
rect 19981 3621 19993 3624
rect 20027 3621 20039 3655
rect 19981 3615 20039 3621
rect 17218 3544 17224 3596
rect 17276 3584 17282 3596
rect 20809 3587 20867 3593
rect 20809 3584 20821 3587
rect 17276 3556 20821 3584
rect 17276 3544 17282 3556
rect 20809 3553 20821 3556
rect 20855 3553 20867 3587
rect 20809 3547 20867 3553
rect 19337 3519 19395 3525
rect 19337 3485 19349 3519
rect 19383 3516 19395 3519
rect 20530 3516 20536 3528
rect 19383 3488 20536 3516
rect 19383 3485 19395 3488
rect 19337 3479 19395 3485
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 19705 3451 19763 3457
rect 19705 3417 19717 3451
rect 19751 3448 19763 3451
rect 20162 3448 20168 3460
rect 19751 3420 20168 3448
rect 19751 3417 19763 3420
rect 19705 3411 19763 3417
rect 20162 3408 20168 3420
rect 20220 3408 20226 3460
rect 1104 3290 21896 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21896 3290
rect 1104 3216 21896 3238
rect 19058 3136 19064 3188
rect 19116 3176 19122 3188
rect 20073 3179 20131 3185
rect 20073 3176 20085 3179
rect 19116 3148 20085 3176
rect 19116 3136 19122 3148
rect 20073 3145 20085 3148
rect 20119 3145 20131 3179
rect 20073 3139 20131 3145
rect 18969 3111 19027 3117
rect 18969 3077 18981 3111
rect 19015 3108 19027 3111
rect 20714 3108 20720 3120
rect 19015 3080 20720 3108
rect 19015 3077 19027 3080
rect 18969 3071 19027 3077
rect 20714 3068 20720 3080
rect 20772 3068 20778 3120
rect 19058 3000 19064 3052
rect 19116 3040 19122 3052
rect 19337 3043 19395 3049
rect 19337 3040 19349 3043
rect 19116 3012 19349 3040
rect 19116 3000 19122 3012
rect 19337 3009 19349 3012
rect 19383 3040 19395 3043
rect 20165 3043 20223 3049
rect 20165 3040 20177 3043
rect 19383 3012 20177 3040
rect 19383 3009 19395 3012
rect 19337 3003 19395 3009
rect 20165 3009 20177 3012
rect 20211 3009 20223 3043
rect 21266 3040 21272 3052
rect 21227 3012 21272 3040
rect 20165 3003 20223 3009
rect 21266 3000 21272 3012
rect 21324 3000 21330 3052
rect 18601 2975 18659 2981
rect 18601 2941 18613 2975
rect 18647 2972 18659 2975
rect 21284 2972 21312 3000
rect 18647 2944 21312 2972
rect 18647 2941 18659 2944
rect 18601 2935 18659 2941
rect 15194 2864 15200 2916
rect 15252 2904 15258 2916
rect 20533 2907 20591 2913
rect 20533 2904 20545 2907
rect 15252 2876 20545 2904
rect 15252 2864 15258 2876
rect 20533 2873 20545 2876
rect 20579 2873 20591 2907
rect 20533 2867 20591 2873
rect 19610 2836 19616 2848
rect 19571 2808 19616 2836
rect 19610 2796 19616 2808
rect 19668 2796 19674 2848
rect 19702 2796 19708 2848
rect 19760 2836 19766 2848
rect 21177 2839 21235 2845
rect 21177 2836 21189 2839
rect 19760 2808 21189 2836
rect 19760 2796 19766 2808
rect 21177 2805 21189 2808
rect 21223 2805 21235 2839
rect 21177 2799 21235 2805
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 17034 2524 17040 2576
rect 17092 2564 17098 2576
rect 19981 2567 20039 2573
rect 19981 2564 19993 2567
rect 17092 2536 19993 2564
rect 17092 2524 17098 2536
rect 19981 2533 19993 2536
rect 20027 2533 20039 2567
rect 19981 2527 20039 2533
rect 18509 2499 18567 2505
rect 18509 2465 18521 2499
rect 18555 2496 18567 2499
rect 20806 2496 20812 2508
rect 18555 2468 20576 2496
rect 20767 2468 20812 2496
rect 18555 2465 18567 2468
rect 18509 2459 18567 2465
rect 20548 2440 20576 2468
rect 20806 2456 20812 2468
rect 20864 2456 20870 2508
rect 14826 2388 14832 2440
rect 14884 2428 14890 2440
rect 19429 2431 19487 2437
rect 19429 2428 19441 2431
rect 14884 2400 19441 2428
rect 14884 2388 14890 2400
rect 19429 2397 19441 2400
rect 19475 2397 19487 2431
rect 20530 2428 20536 2440
rect 20491 2400 20536 2428
rect 19429 2391 19487 2397
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 19610 2360 19616 2372
rect 19571 2332 19616 2360
rect 19610 2320 19616 2332
rect 19668 2320 19674 2372
rect 20165 2363 20223 2369
rect 20165 2360 20177 2363
rect 19996 2332 20177 2360
rect 18877 2295 18935 2301
rect 18877 2261 18889 2295
rect 18923 2292 18935 2295
rect 19242 2292 19248 2304
rect 18923 2264 19248 2292
rect 18923 2261 18935 2264
rect 18877 2255 18935 2261
rect 19242 2252 19248 2264
rect 19300 2292 19306 2304
rect 19996 2292 20024 2332
rect 20165 2329 20177 2332
rect 20211 2329 20223 2363
rect 20165 2323 20223 2329
rect 19300 2264 20024 2292
rect 19300 2252 19306 2264
rect 1104 2202 21896 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21896 2202
rect 1104 2128 21896 2150
<< via1 >>
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 3240 20544 3292 20596
rect 4436 20544 4488 20596
rect 296 20476 348 20528
rect 2412 20476 2464 20528
rect 2688 20408 2740 20460
rect 3148 20476 3200 20528
rect 4068 20476 4120 20528
rect 3240 20451 3292 20460
rect 3240 20417 3249 20451
rect 3249 20417 3283 20451
rect 3283 20417 3292 20451
rect 3240 20408 3292 20417
rect 5724 20476 5776 20528
rect 3792 20340 3844 20392
rect 5356 20408 5408 20460
rect 4252 20340 4304 20392
rect 5264 20340 5316 20392
rect 6460 20408 6512 20460
rect 8116 20476 8168 20528
rect 7932 20451 7984 20460
rect 6828 20340 6880 20392
rect 7932 20417 7941 20451
rect 7941 20417 7975 20451
rect 7975 20417 7984 20451
rect 7932 20408 7984 20417
rect 9220 20408 9272 20460
rect 9772 20408 9824 20460
rect 10324 20408 10376 20460
rect 10876 20408 10928 20460
rect 7840 20340 7892 20392
rect 8208 20340 8260 20392
rect 12624 20544 12676 20596
rect 13176 20544 13228 20596
rect 14280 20544 14332 20596
rect 15752 20544 15804 20596
rect 12900 20476 12952 20528
rect 11244 20408 11296 20460
rect 12072 20408 12124 20460
rect 13820 20476 13872 20528
rect 16028 20476 16080 20528
rect 17684 20544 17736 20596
rect 19892 20544 19944 20596
rect 20720 20544 20772 20596
rect 13452 20451 13504 20460
rect 13452 20417 13461 20451
rect 13461 20417 13495 20451
rect 13495 20417 13504 20451
rect 13452 20408 13504 20417
rect 14924 20408 14976 20460
rect 15936 20408 15988 20460
rect 16304 20451 16356 20460
rect 16304 20417 16313 20451
rect 16313 20417 16347 20451
rect 16347 20417 16356 20451
rect 16304 20408 16356 20417
rect 17500 20451 17552 20460
rect 14280 20340 14332 20392
rect 14648 20383 14700 20392
rect 14648 20349 14657 20383
rect 14657 20349 14691 20383
rect 14691 20349 14700 20383
rect 14648 20340 14700 20349
rect 17500 20417 17509 20451
rect 17509 20417 17543 20451
rect 17543 20417 17552 20451
rect 17500 20408 17552 20417
rect 18604 20451 18656 20460
rect 1676 20272 1728 20324
rect 2504 20247 2556 20256
rect 2504 20213 2513 20247
rect 2513 20213 2547 20247
rect 2547 20213 2556 20247
rect 2504 20204 2556 20213
rect 2964 20247 3016 20256
rect 2964 20213 2973 20247
rect 2973 20213 3007 20247
rect 3007 20213 3016 20247
rect 2964 20204 3016 20213
rect 3332 20204 3384 20256
rect 4068 20247 4120 20256
rect 4068 20213 4077 20247
rect 4077 20213 4111 20247
rect 4111 20213 4120 20247
rect 4068 20204 4120 20213
rect 4804 20247 4856 20256
rect 4804 20213 4813 20247
rect 4813 20213 4847 20247
rect 4847 20213 4856 20247
rect 4804 20204 4856 20213
rect 6000 20247 6052 20256
rect 6000 20213 6009 20247
rect 6009 20213 6043 20247
rect 6043 20213 6052 20247
rect 6000 20204 6052 20213
rect 17592 20340 17644 20392
rect 18604 20417 18613 20451
rect 18613 20417 18647 20451
rect 18647 20417 18656 20451
rect 18604 20408 18656 20417
rect 18512 20340 18564 20392
rect 16856 20272 16908 20324
rect 17040 20272 17092 20324
rect 20260 20408 20312 20460
rect 21640 20408 21692 20460
rect 21732 20340 21784 20392
rect 21824 20272 21876 20324
rect 6828 20204 6880 20256
rect 7380 20204 7432 20256
rect 7656 20247 7708 20256
rect 7656 20213 7665 20247
rect 7665 20213 7699 20247
rect 7699 20213 7708 20247
rect 7656 20204 7708 20213
rect 8208 20204 8260 20256
rect 8392 20204 8444 20256
rect 9680 20204 9732 20256
rect 11060 20204 11112 20256
rect 11704 20247 11756 20256
rect 11704 20213 11713 20247
rect 11713 20213 11747 20247
rect 11747 20213 11756 20247
rect 11704 20204 11756 20213
rect 11980 20247 12032 20256
rect 11980 20213 11989 20247
rect 11989 20213 12023 20247
rect 12023 20213 12032 20247
rect 11980 20204 12032 20213
rect 13820 20204 13872 20256
rect 14740 20204 14792 20256
rect 14832 20204 14884 20256
rect 16580 20204 16632 20256
rect 18236 20204 18288 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 1676 20043 1728 20052
rect 1676 20009 1685 20043
rect 1685 20009 1719 20043
rect 1719 20009 1728 20043
rect 1676 20000 1728 20009
rect 2964 19932 3016 19984
rect 1400 19864 1452 19916
rect 1492 19839 1544 19848
rect 1492 19805 1501 19839
rect 1501 19805 1535 19839
rect 1535 19805 1544 19839
rect 1492 19796 1544 19805
rect 3332 19864 3384 19916
rect 4160 19907 4212 19916
rect 2044 19796 2096 19848
rect 2596 19839 2648 19848
rect 2596 19805 2605 19839
rect 2605 19805 2639 19839
rect 2639 19805 2648 19839
rect 2596 19796 2648 19805
rect 3424 19796 3476 19848
rect 4160 19873 4169 19907
rect 4169 19873 4203 19907
rect 4203 19873 4212 19907
rect 4160 19864 4212 19873
rect 6828 20000 6880 20052
rect 7748 20000 7800 20052
rect 11244 20000 11296 20052
rect 12072 20000 12124 20052
rect 12440 20043 12492 20052
rect 12440 20009 12449 20043
rect 12449 20009 12483 20043
rect 12483 20009 12492 20043
rect 12440 20000 12492 20009
rect 13820 20000 13872 20052
rect 18788 20000 18840 20052
rect 19524 20000 19576 20052
rect 7932 19932 7984 19984
rect 6644 19839 6696 19848
rect 6644 19805 6653 19839
rect 6653 19805 6687 19839
rect 6687 19805 6696 19839
rect 6644 19796 6696 19805
rect 12900 19864 12952 19916
rect 16856 19907 16908 19916
rect 9128 19796 9180 19848
rect 10600 19839 10652 19848
rect 10600 19805 10609 19839
rect 10609 19805 10643 19839
rect 10643 19805 10652 19839
rect 10600 19796 10652 19805
rect 12256 19839 12308 19848
rect 12256 19805 12265 19839
rect 12265 19805 12299 19839
rect 12299 19805 12308 19839
rect 12256 19796 12308 19805
rect 13084 19839 13136 19848
rect 13084 19805 13093 19839
rect 13093 19805 13127 19839
rect 13127 19805 13136 19839
rect 13084 19796 13136 19805
rect 14556 19796 14608 19848
rect 14740 19839 14792 19848
rect 14740 19805 14749 19839
rect 14749 19805 14783 19839
rect 14783 19805 14792 19839
rect 14740 19796 14792 19805
rect 16856 19873 16865 19907
rect 16865 19873 16899 19907
rect 16899 19873 16908 19907
rect 16856 19864 16908 19873
rect 17316 19864 17368 19916
rect 16396 19796 16448 19848
rect 18880 19839 18932 19848
rect 18880 19805 18889 19839
rect 18889 19805 18923 19839
rect 18923 19805 18932 19839
rect 18880 19796 18932 19805
rect 19892 19796 19944 19848
rect 21916 19864 21968 19916
rect 20352 19796 20404 19848
rect 21088 19839 21140 19848
rect 21088 19805 21097 19839
rect 21097 19805 21131 19839
rect 21131 19805 21140 19839
rect 21088 19796 21140 19805
rect 2136 19703 2188 19712
rect 2136 19669 2145 19703
rect 2145 19669 2179 19703
rect 2179 19669 2188 19703
rect 2136 19660 2188 19669
rect 3332 19660 3384 19712
rect 4344 19703 4396 19712
rect 4344 19669 4353 19703
rect 4353 19669 4387 19703
rect 4387 19669 4396 19703
rect 4344 19660 4396 19669
rect 4712 19703 4764 19712
rect 4712 19669 4721 19703
rect 4721 19669 4755 19703
rect 4755 19669 4764 19703
rect 4712 19660 4764 19669
rect 5264 19771 5316 19780
rect 5264 19737 5298 19771
rect 5298 19737 5316 19771
rect 5264 19728 5316 19737
rect 6460 19728 6512 19780
rect 6736 19728 6788 19780
rect 7012 19728 7064 19780
rect 12164 19728 12216 19780
rect 15568 19728 15620 19780
rect 18052 19771 18104 19780
rect 18052 19737 18061 19771
rect 18061 19737 18095 19771
rect 18095 19737 18104 19771
rect 18052 19728 18104 19737
rect 18420 19728 18472 19780
rect 22652 19728 22704 19780
rect 5816 19660 5868 19712
rect 6552 19660 6604 19712
rect 9036 19660 9088 19712
rect 10968 19660 11020 19712
rect 13636 19660 13688 19712
rect 15200 19660 15252 19712
rect 20720 19703 20772 19712
rect 20720 19669 20729 19703
rect 20729 19669 20763 19703
rect 20763 19669 20772 19703
rect 20720 19660 20772 19669
rect 21272 19703 21324 19712
rect 21272 19669 21281 19703
rect 21281 19669 21315 19703
rect 21315 19669 21324 19703
rect 21272 19660 21324 19669
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 2596 19456 2648 19508
rect 3424 19456 3476 19508
rect 7012 19499 7064 19508
rect 7012 19465 7021 19499
rect 7021 19465 7055 19499
rect 7055 19465 7064 19499
rect 7012 19456 7064 19465
rect 3240 19388 3292 19440
rect 6736 19388 6788 19440
rect 7564 19456 7616 19508
rect 7656 19456 7708 19508
rect 9036 19499 9088 19508
rect 9036 19465 9045 19499
rect 9045 19465 9079 19499
rect 9079 19465 9088 19499
rect 9036 19456 9088 19465
rect 9680 19456 9732 19508
rect 13084 19499 13136 19508
rect 13084 19465 13093 19499
rect 13093 19465 13127 19499
rect 13127 19465 13136 19499
rect 13084 19456 13136 19465
rect 13820 19456 13872 19508
rect 1952 19320 2004 19372
rect 3424 19363 3476 19372
rect 3424 19329 3433 19363
rect 3433 19329 3467 19363
rect 3467 19329 3476 19363
rect 3424 19320 3476 19329
rect 3976 19320 4028 19372
rect 5448 19363 5500 19372
rect 5448 19329 5457 19363
rect 5457 19329 5491 19363
rect 5491 19329 5500 19363
rect 5448 19320 5500 19329
rect 6552 19320 6604 19372
rect 7288 19363 7340 19372
rect 7288 19329 7297 19363
rect 7297 19329 7331 19363
rect 7331 19329 7340 19363
rect 7288 19320 7340 19329
rect 4712 19252 4764 19304
rect 9312 19320 9364 19372
rect 9956 19320 10008 19372
rect 11980 19363 12032 19372
rect 11980 19329 12014 19363
rect 12014 19329 12032 19363
rect 11980 19320 12032 19329
rect 14740 19388 14792 19440
rect 15660 19388 15712 19440
rect 13636 19363 13688 19372
rect 13636 19329 13670 19363
rect 13670 19329 13688 19363
rect 13636 19320 13688 19329
rect 14648 19320 14700 19372
rect 5356 19184 5408 19236
rect 9680 19184 9732 19236
rect 9772 19184 9824 19236
rect 15568 19320 15620 19372
rect 19984 19456 20036 19508
rect 20076 19499 20128 19508
rect 20076 19465 20085 19499
rect 20085 19465 20119 19499
rect 20119 19465 20128 19499
rect 20076 19456 20128 19465
rect 20996 19456 21048 19508
rect 18696 19388 18748 19440
rect 17316 19363 17368 19372
rect 17316 19329 17325 19363
rect 17325 19329 17359 19363
rect 17359 19329 17368 19363
rect 17316 19320 17368 19329
rect 18420 19320 18472 19372
rect 18604 19363 18656 19372
rect 18604 19329 18613 19363
rect 18613 19329 18647 19363
rect 18647 19329 18656 19363
rect 18604 19320 18656 19329
rect 18972 19320 19024 19372
rect 19064 19320 19116 19372
rect 19616 19388 19668 19440
rect 19708 19363 19760 19372
rect 19708 19329 19717 19363
rect 19717 19329 19751 19363
rect 19751 19329 19760 19363
rect 19708 19320 19760 19329
rect 20168 19320 20220 19372
rect 20444 19320 20496 19372
rect 20904 19320 20956 19372
rect 2228 19159 2280 19168
rect 2228 19125 2237 19159
rect 2237 19125 2271 19159
rect 2271 19125 2280 19159
rect 2228 19116 2280 19125
rect 5080 19159 5132 19168
rect 5080 19125 5089 19159
rect 5089 19125 5123 19159
rect 5123 19125 5132 19159
rect 5080 19116 5132 19125
rect 7564 19116 7616 19168
rect 9864 19116 9916 19168
rect 10048 19159 10100 19168
rect 10048 19125 10057 19159
rect 10057 19125 10091 19159
rect 10091 19125 10100 19159
rect 10048 19116 10100 19125
rect 16672 19159 16724 19168
rect 16672 19125 16681 19159
rect 16681 19125 16715 19159
rect 16715 19125 16724 19159
rect 16672 19116 16724 19125
rect 17868 19116 17920 19168
rect 21364 19116 21416 19168
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 1952 18912 2004 18964
rect 3976 18912 4028 18964
rect 4344 18912 4396 18964
rect 5724 18955 5776 18964
rect 5724 18921 5733 18955
rect 5733 18921 5767 18955
rect 5767 18921 5776 18955
rect 5724 18912 5776 18921
rect 6920 18912 6972 18964
rect 7288 18912 7340 18964
rect 7840 18955 7892 18964
rect 7840 18921 7849 18955
rect 7849 18921 7883 18955
rect 7883 18921 7892 18955
rect 7840 18912 7892 18921
rect 8116 18955 8168 18964
rect 8116 18921 8125 18955
rect 8125 18921 8159 18955
rect 8159 18921 8168 18955
rect 8116 18912 8168 18921
rect 9220 18912 9272 18964
rect 13820 18912 13872 18964
rect 17776 18912 17828 18964
rect 18696 18955 18748 18964
rect 18696 18921 18705 18955
rect 18705 18921 18739 18955
rect 18739 18921 18748 18955
rect 18696 18912 18748 18921
rect 20536 18912 20588 18964
rect 21548 18912 21600 18964
rect 5448 18776 5500 18828
rect 3424 18708 3476 18760
rect 2320 18683 2372 18692
rect 2320 18649 2354 18683
rect 2354 18649 2372 18683
rect 2320 18640 2372 18649
rect 4160 18640 4212 18692
rect 6736 18844 6788 18896
rect 7196 18844 7248 18896
rect 6828 18776 6880 18828
rect 22100 18844 22152 18896
rect 12072 18776 12124 18828
rect 13084 18819 13136 18828
rect 13084 18785 13093 18819
rect 13093 18785 13127 18819
rect 13127 18785 13136 18819
rect 13084 18776 13136 18785
rect 15660 18819 15712 18828
rect 15660 18785 15669 18819
rect 15669 18785 15703 18819
rect 15703 18785 15712 18819
rect 15660 18776 15712 18785
rect 7196 18708 7248 18760
rect 10600 18708 10652 18760
rect 15200 18751 15252 18760
rect 15200 18717 15209 18751
rect 15209 18717 15243 18751
rect 15243 18717 15252 18751
rect 15200 18708 15252 18717
rect 16672 18708 16724 18760
rect 9772 18683 9824 18692
rect 9772 18649 9806 18683
rect 9806 18649 9824 18683
rect 9772 18640 9824 18649
rect 9864 18640 9916 18692
rect 11060 18640 11112 18692
rect 12808 18640 12860 18692
rect 9312 18572 9364 18624
rect 10876 18615 10928 18624
rect 10876 18581 10885 18615
rect 10885 18581 10919 18615
rect 10919 18581 10928 18615
rect 10876 18572 10928 18581
rect 11152 18615 11204 18624
rect 11152 18581 11161 18615
rect 11161 18581 11195 18615
rect 11195 18581 11204 18615
rect 11152 18572 11204 18581
rect 14556 18615 14608 18624
rect 14556 18581 14565 18615
rect 14565 18581 14599 18615
rect 14599 18581 14608 18615
rect 14556 18572 14608 18581
rect 16948 18572 17000 18624
rect 17408 18708 17460 18760
rect 18328 18708 18380 18760
rect 19984 18751 20036 18760
rect 19984 18717 19993 18751
rect 19993 18717 20027 18751
rect 20027 18717 20036 18751
rect 19984 18708 20036 18717
rect 20812 18751 20864 18760
rect 20812 18717 20821 18751
rect 20821 18717 20855 18751
rect 20855 18717 20864 18751
rect 20812 18708 20864 18717
rect 21180 18708 21232 18760
rect 21548 18640 21600 18692
rect 17960 18615 18012 18624
rect 17960 18581 17969 18615
rect 17969 18581 18003 18615
rect 18003 18581 18012 18615
rect 17960 18572 18012 18581
rect 18420 18615 18472 18624
rect 18420 18581 18429 18615
rect 18429 18581 18463 18615
rect 18463 18581 18472 18615
rect 18420 18572 18472 18581
rect 21272 18615 21324 18624
rect 21272 18581 21281 18615
rect 21281 18581 21315 18615
rect 21315 18581 21324 18615
rect 21272 18572 21324 18581
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 2044 18411 2096 18420
rect 2044 18377 2053 18411
rect 2053 18377 2087 18411
rect 2087 18377 2096 18411
rect 2044 18368 2096 18377
rect 2688 18411 2740 18420
rect 2688 18377 2697 18411
rect 2697 18377 2731 18411
rect 2731 18377 2740 18411
rect 2688 18368 2740 18377
rect 3148 18411 3200 18420
rect 3148 18377 3157 18411
rect 3157 18377 3191 18411
rect 3191 18377 3200 18411
rect 3148 18368 3200 18377
rect 4252 18411 4304 18420
rect 4252 18377 4261 18411
rect 4261 18377 4295 18411
rect 4295 18377 4304 18411
rect 4252 18368 4304 18377
rect 7196 18411 7248 18420
rect 7196 18377 7205 18411
rect 7205 18377 7239 18411
rect 7239 18377 7248 18411
rect 7196 18368 7248 18377
rect 9680 18368 9732 18420
rect 10048 18368 10100 18420
rect 11152 18368 11204 18420
rect 12164 18411 12216 18420
rect 12164 18377 12173 18411
rect 12173 18377 12207 18411
rect 12207 18377 12216 18411
rect 12164 18368 12216 18377
rect 2412 18300 2464 18352
rect 1676 18275 1728 18284
rect 1676 18241 1685 18275
rect 1685 18241 1719 18275
rect 1719 18241 1728 18275
rect 1676 18232 1728 18241
rect 5080 18232 5132 18284
rect 9864 18300 9916 18352
rect 8392 18275 8444 18284
rect 8392 18241 8426 18275
rect 8426 18241 8444 18275
rect 6552 18207 6604 18216
rect 6552 18173 6561 18207
rect 6561 18173 6595 18207
rect 6595 18173 6604 18207
rect 6552 18164 6604 18173
rect 7104 18164 7156 18216
rect 6644 18096 6696 18148
rect 8392 18232 8444 18241
rect 9956 18232 10008 18284
rect 10876 18164 10928 18216
rect 17408 18368 17460 18420
rect 18328 18411 18380 18420
rect 18328 18377 18337 18411
rect 18337 18377 18371 18411
rect 18371 18377 18380 18411
rect 18328 18368 18380 18377
rect 18880 18368 18932 18420
rect 21456 18368 21508 18420
rect 17960 18300 18012 18352
rect 15660 18164 15712 18216
rect 18696 18232 18748 18284
rect 19064 18207 19116 18216
rect 19064 18173 19073 18207
rect 19073 18173 19107 18207
rect 19107 18173 19116 18207
rect 19064 18164 19116 18173
rect 19984 18275 20036 18284
rect 19984 18241 19993 18275
rect 19993 18241 20027 18275
rect 20027 18241 20036 18275
rect 19984 18232 20036 18241
rect 18788 18096 18840 18148
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 5448 18028 5500 18080
rect 12808 18028 12860 18080
rect 14740 18028 14792 18080
rect 14924 18028 14976 18080
rect 17684 18028 17736 18080
rect 18880 18028 18932 18080
rect 20996 18232 21048 18284
rect 20628 18096 20680 18148
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 2320 17867 2372 17876
rect 2320 17833 2329 17867
rect 2329 17833 2363 17867
rect 2363 17833 2372 17867
rect 2320 17824 2372 17833
rect 4068 17824 4120 17876
rect 7104 17867 7156 17876
rect 1584 17756 1636 17808
rect 7104 17833 7113 17867
rect 7113 17833 7147 17867
rect 7147 17833 7156 17867
rect 7104 17824 7156 17833
rect 10324 17867 10376 17876
rect 10324 17833 10333 17867
rect 10333 17833 10367 17867
rect 10367 17833 10376 17867
rect 10324 17824 10376 17833
rect 19064 17824 19116 17876
rect 19984 17824 20036 17876
rect 1584 17620 1636 17672
rect 5724 17620 5776 17672
rect 6644 17688 6696 17740
rect 7380 17688 7432 17740
rect 7748 17731 7800 17740
rect 7748 17697 7757 17731
rect 7757 17697 7791 17731
rect 7791 17697 7800 17731
rect 7748 17688 7800 17697
rect 11244 17688 11296 17740
rect 18788 17756 18840 17808
rect 16948 17731 17000 17740
rect 16948 17697 16957 17731
rect 16957 17697 16991 17731
rect 16991 17697 17000 17731
rect 16948 17688 17000 17697
rect 17684 17688 17736 17740
rect 16396 17620 16448 17672
rect 17776 17663 17828 17672
rect 17776 17629 17785 17663
rect 17785 17629 17819 17663
rect 17819 17629 17828 17663
rect 17776 17620 17828 17629
rect 8024 17552 8076 17604
rect 19616 17620 19668 17672
rect 20076 17620 20128 17672
rect 3148 17527 3200 17536
rect 3148 17493 3157 17527
rect 3157 17493 3191 17527
rect 3191 17493 3200 17527
rect 3148 17484 3200 17493
rect 5632 17484 5684 17536
rect 7472 17527 7524 17536
rect 7472 17493 7481 17527
rect 7481 17493 7515 17527
rect 7515 17493 7524 17527
rect 7472 17484 7524 17493
rect 10048 17484 10100 17536
rect 12440 17484 12492 17536
rect 12808 17484 12860 17536
rect 14740 17527 14792 17536
rect 14740 17493 14749 17527
rect 14749 17493 14783 17527
rect 14783 17493 14792 17527
rect 14740 17484 14792 17493
rect 16948 17484 17000 17536
rect 18328 17484 18380 17536
rect 18788 17552 18840 17604
rect 19800 17484 19852 17536
rect 20904 17552 20956 17604
rect 20720 17527 20772 17536
rect 20720 17493 20729 17527
rect 20729 17493 20763 17527
rect 20763 17493 20772 17527
rect 20720 17484 20772 17493
rect 21272 17527 21324 17536
rect 21272 17493 21281 17527
rect 21281 17493 21315 17527
rect 21315 17493 21324 17527
rect 21272 17484 21324 17493
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 3332 17280 3384 17332
rect 5264 17280 5316 17332
rect 5448 17280 5500 17332
rect 14096 17280 14148 17332
rect 18696 17280 18748 17332
rect 18972 17323 19024 17332
rect 18972 17289 18981 17323
rect 18981 17289 19015 17323
rect 19015 17289 19024 17323
rect 18972 17280 19024 17289
rect 19616 17323 19668 17332
rect 19616 17289 19625 17323
rect 19625 17289 19659 17323
rect 19659 17289 19668 17323
rect 19616 17280 19668 17289
rect 20076 17323 20128 17332
rect 20076 17289 20085 17323
rect 20085 17289 20119 17323
rect 20119 17289 20128 17323
rect 20076 17280 20128 17289
rect 7472 17212 7524 17264
rect 12440 17212 12492 17264
rect 14188 17255 14240 17264
rect 14188 17221 14197 17255
rect 14197 17221 14231 17255
rect 14231 17221 14240 17255
rect 14188 17212 14240 17221
rect 17868 17212 17920 17264
rect 3332 17144 3384 17196
rect 5632 17187 5684 17196
rect 5632 17153 5641 17187
rect 5641 17153 5675 17187
rect 5675 17153 5684 17187
rect 5632 17144 5684 17153
rect 6552 17144 6604 17196
rect 7288 17144 7340 17196
rect 7840 17144 7892 17196
rect 9220 17187 9272 17196
rect 9220 17153 9229 17187
rect 9229 17153 9263 17187
rect 9263 17153 9272 17187
rect 9220 17144 9272 17153
rect 14464 17144 14516 17196
rect 14740 17144 14792 17196
rect 16672 17187 16724 17196
rect 16672 17153 16681 17187
rect 16681 17153 16715 17187
rect 16715 17153 16724 17187
rect 16672 17144 16724 17153
rect 18144 17144 18196 17196
rect 19524 17144 19576 17196
rect 3424 17076 3476 17128
rect 3884 17119 3936 17128
rect 3884 17085 3893 17119
rect 3893 17085 3927 17119
rect 3927 17085 3936 17119
rect 3884 17076 3936 17085
rect 9772 17076 9824 17128
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12440 17076 12492 17085
rect 13820 17076 13872 17128
rect 15476 17076 15528 17128
rect 7564 17008 7616 17060
rect 15384 17008 15436 17060
rect 1584 16983 1636 16992
rect 1584 16949 1593 16983
rect 1593 16949 1627 16983
rect 1627 16949 1636 16983
rect 1584 16940 1636 16949
rect 2964 16940 3016 16992
rect 8668 16983 8720 16992
rect 8668 16949 8677 16983
rect 8677 16949 8711 16983
rect 8711 16949 8720 16983
rect 8668 16940 8720 16949
rect 9864 16983 9916 16992
rect 9864 16949 9873 16983
rect 9873 16949 9907 16983
rect 9907 16949 9916 16983
rect 9864 16940 9916 16949
rect 19616 17008 19668 17060
rect 21088 17187 21140 17196
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 21088 17144 21140 17153
rect 17316 16983 17368 16992
rect 17316 16949 17325 16983
rect 17325 16949 17359 16983
rect 17359 16949 17368 16983
rect 17316 16940 17368 16949
rect 17776 16940 17828 16992
rect 18328 16940 18380 16992
rect 21180 16940 21232 16992
rect 21364 16940 21416 16992
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 1584 16600 1636 16652
rect 2964 16643 3016 16652
rect 2964 16609 2973 16643
rect 2973 16609 3007 16643
rect 3007 16609 3016 16643
rect 2964 16600 3016 16609
rect 3424 16600 3476 16652
rect 5724 16736 5776 16788
rect 5816 16668 5868 16720
rect 9220 16643 9272 16652
rect 3148 16532 3200 16584
rect 4804 16575 4856 16584
rect 4804 16541 4838 16575
rect 4838 16541 4856 16575
rect 4804 16532 4856 16541
rect 4068 16396 4120 16448
rect 9220 16609 9229 16643
rect 9229 16609 9263 16643
rect 9263 16609 9272 16643
rect 9220 16600 9272 16609
rect 8668 16532 8720 16584
rect 9956 16600 10008 16652
rect 10232 16600 10284 16652
rect 10600 16600 10652 16652
rect 14832 16736 14884 16788
rect 15660 16736 15712 16788
rect 16396 16736 16448 16788
rect 21088 16736 21140 16788
rect 15476 16711 15528 16720
rect 15476 16677 15485 16711
rect 15485 16677 15519 16711
rect 15519 16677 15528 16711
rect 15476 16668 15528 16677
rect 15384 16600 15436 16652
rect 16672 16643 16724 16652
rect 16672 16609 16681 16643
rect 16681 16609 16715 16643
rect 16715 16609 16724 16643
rect 16672 16600 16724 16609
rect 17040 16600 17092 16652
rect 18144 16643 18196 16652
rect 18144 16609 18153 16643
rect 18153 16609 18187 16643
rect 18187 16609 18196 16643
rect 18144 16600 18196 16609
rect 9772 16464 9824 16516
rect 6828 16439 6880 16448
rect 6828 16405 6837 16439
rect 6837 16405 6871 16439
rect 6871 16405 6880 16439
rect 6828 16396 6880 16405
rect 18420 16532 18472 16584
rect 20076 16532 20128 16584
rect 21088 16575 21140 16584
rect 11152 16464 11204 16516
rect 12716 16464 12768 16516
rect 14372 16507 14424 16516
rect 14372 16473 14406 16507
rect 14406 16473 14424 16507
rect 14372 16464 14424 16473
rect 19340 16464 19392 16516
rect 21088 16541 21097 16575
rect 21097 16541 21131 16575
rect 21131 16541 21140 16575
rect 21088 16532 21140 16541
rect 10416 16396 10468 16448
rect 12440 16396 12492 16448
rect 13820 16396 13872 16448
rect 16948 16396 17000 16448
rect 19524 16396 19576 16448
rect 19708 16439 19760 16448
rect 19708 16405 19717 16439
rect 19717 16405 19751 16439
rect 19751 16405 19760 16439
rect 19708 16396 19760 16405
rect 20352 16439 20404 16448
rect 20352 16405 20361 16439
rect 20361 16405 20395 16439
rect 20395 16405 20404 16439
rect 20352 16396 20404 16405
rect 21272 16439 21324 16448
rect 21272 16405 21281 16439
rect 21281 16405 21315 16439
rect 21315 16405 21324 16439
rect 21272 16396 21324 16405
rect 21456 16396 21508 16448
rect 21732 16396 21784 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 4068 16192 4120 16244
rect 9220 16235 9272 16244
rect 3424 16124 3476 16176
rect 6828 16124 6880 16176
rect 9220 16201 9229 16235
rect 9229 16201 9263 16235
rect 9263 16201 9272 16235
rect 9220 16192 9272 16201
rect 12716 16235 12768 16244
rect 2044 16099 2096 16108
rect 2044 16065 2078 16099
rect 2078 16065 2096 16099
rect 2044 16056 2096 16065
rect 3332 15988 3384 16040
rect 3884 15920 3936 15972
rect 6920 16099 6972 16108
rect 6920 16065 6929 16099
rect 6929 16065 6963 16099
rect 6963 16065 6972 16099
rect 10600 16124 10652 16176
rect 12716 16201 12725 16235
rect 12725 16201 12759 16235
rect 12759 16201 12768 16235
rect 12716 16192 12768 16201
rect 14372 16235 14424 16244
rect 14372 16201 14381 16235
rect 14381 16201 14415 16235
rect 14415 16201 14424 16235
rect 14372 16192 14424 16201
rect 17040 16192 17092 16244
rect 18144 16192 18196 16244
rect 19800 16192 19852 16244
rect 20076 16235 20128 16244
rect 20076 16201 20085 16235
rect 20085 16201 20119 16235
rect 20119 16201 20128 16235
rect 20076 16192 20128 16201
rect 20168 16192 20220 16244
rect 20720 16192 20772 16244
rect 20904 16192 20956 16244
rect 6920 16056 6972 16065
rect 9864 16056 9916 16108
rect 12440 16056 12492 16108
rect 13820 16056 13872 16108
rect 14832 16056 14884 16108
rect 16120 16056 16172 16108
rect 16580 16056 16632 16108
rect 17316 16124 17368 16176
rect 19340 16056 19392 16108
rect 19616 16099 19668 16108
rect 19616 16065 19625 16099
rect 19625 16065 19659 16099
rect 19659 16065 19668 16099
rect 19616 16056 19668 16065
rect 7012 15988 7064 16040
rect 7288 15988 7340 16040
rect 7104 15920 7156 15972
rect 11244 15920 11296 15972
rect 19984 16056 20036 16108
rect 20904 16056 20956 16108
rect 21364 15852 21416 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 2044 15648 2096 15700
rect 5724 15691 5776 15700
rect 5724 15657 5733 15691
rect 5733 15657 5767 15691
rect 5767 15657 5776 15691
rect 5724 15648 5776 15657
rect 8116 15648 8168 15700
rect 11152 15691 11204 15700
rect 11152 15657 11161 15691
rect 11161 15657 11195 15691
rect 11195 15657 11204 15691
rect 11152 15648 11204 15657
rect 16120 15691 16172 15700
rect 16120 15657 16129 15691
rect 16129 15657 16163 15691
rect 16163 15657 16172 15691
rect 16120 15648 16172 15657
rect 7932 15580 7984 15632
rect 19984 15648 20036 15700
rect 21088 15648 21140 15700
rect 20720 15580 20772 15632
rect 20996 15580 21048 15632
rect 2872 15487 2924 15496
rect 2872 15453 2881 15487
rect 2881 15453 2915 15487
rect 2915 15453 2924 15487
rect 6920 15512 6972 15564
rect 16580 15512 16632 15564
rect 17316 15512 17368 15564
rect 7748 15487 7800 15496
rect 2872 15444 2924 15453
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 11244 15444 11296 15496
rect 15476 15487 15528 15496
rect 15476 15453 15485 15487
rect 15485 15453 15519 15487
rect 15519 15453 15528 15487
rect 15476 15444 15528 15453
rect 17776 15487 17828 15496
rect 17776 15453 17810 15487
rect 17810 15453 17828 15487
rect 17776 15444 17828 15453
rect 20168 15487 20220 15496
rect 10324 15376 10376 15428
rect 10416 15376 10468 15428
rect 20168 15453 20177 15487
rect 20177 15453 20211 15487
rect 20211 15453 20220 15487
rect 20168 15444 20220 15453
rect 20628 15487 20680 15496
rect 20628 15453 20637 15487
rect 20637 15453 20671 15487
rect 20671 15453 20680 15487
rect 20628 15444 20680 15453
rect 21088 15487 21140 15496
rect 21088 15453 21097 15487
rect 21097 15453 21131 15487
rect 21131 15453 21140 15487
rect 21088 15444 21140 15453
rect 4252 15308 4304 15360
rect 5448 15308 5500 15360
rect 18880 15351 18932 15360
rect 18880 15317 18889 15351
rect 18889 15317 18923 15351
rect 18923 15317 18932 15351
rect 18880 15308 18932 15317
rect 21272 15351 21324 15360
rect 21272 15317 21281 15351
rect 21281 15317 21315 15351
rect 21315 15317 21324 15351
rect 21272 15308 21324 15317
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 2872 15104 2924 15156
rect 4252 15104 4304 15156
rect 7748 15147 7800 15156
rect 7748 15113 7757 15147
rect 7757 15113 7791 15147
rect 7791 15113 7800 15147
rect 7748 15104 7800 15113
rect 20168 15104 20220 15156
rect 20904 15104 20956 15156
rect 2504 15036 2556 15088
rect 5448 15036 5500 15088
rect 3240 15011 3292 15020
rect 3240 14977 3258 15011
rect 3258 14977 3292 15011
rect 3240 14968 3292 14977
rect 3424 14968 3476 15020
rect 4436 14832 4488 14884
rect 6644 15011 6696 15020
rect 6644 14977 6678 15011
rect 6678 14977 6696 15011
rect 8668 15011 8720 15020
rect 6644 14968 6696 14977
rect 8668 14977 8677 15011
rect 8677 14977 8711 15011
rect 8711 14977 8720 15011
rect 8668 14968 8720 14977
rect 9680 14968 9732 15020
rect 13084 14968 13136 15020
rect 15108 14968 15160 15020
rect 20352 15036 20404 15088
rect 12532 14943 12584 14952
rect 5264 14807 5316 14816
rect 5264 14773 5273 14807
rect 5273 14773 5307 14807
rect 5307 14773 5316 14807
rect 5264 14764 5316 14773
rect 12532 14909 12541 14943
rect 12541 14909 12575 14943
rect 12575 14909 12584 14943
rect 12532 14900 12584 14909
rect 12716 14943 12768 14952
rect 12716 14909 12725 14943
rect 12725 14909 12759 14943
rect 12759 14909 12768 14943
rect 12716 14900 12768 14909
rect 16120 14900 16172 14952
rect 7288 14764 7340 14816
rect 7472 14764 7524 14816
rect 13176 14807 13228 14816
rect 13176 14773 13185 14807
rect 13185 14773 13219 14807
rect 13219 14773 13228 14807
rect 13176 14764 13228 14773
rect 13268 14764 13320 14816
rect 21272 14807 21324 14816
rect 21272 14773 21281 14807
rect 21281 14773 21315 14807
rect 21315 14773 21324 14807
rect 21272 14764 21324 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 3240 14560 3292 14612
rect 7012 14603 7064 14612
rect 7012 14569 7021 14603
rect 7021 14569 7055 14603
rect 7055 14569 7064 14603
rect 7012 14560 7064 14569
rect 9680 14603 9732 14612
rect 9680 14569 9689 14603
rect 9689 14569 9723 14603
rect 9723 14569 9732 14603
rect 9680 14560 9732 14569
rect 7104 14492 7156 14544
rect 4436 14399 4488 14408
rect 4436 14365 4445 14399
rect 4445 14365 4479 14399
rect 4479 14365 4488 14399
rect 4436 14356 4488 14365
rect 5080 14356 5132 14408
rect 7288 14356 7340 14408
rect 12440 14560 12492 14612
rect 15108 14560 15160 14612
rect 20628 14560 20680 14612
rect 21088 14560 21140 14612
rect 7564 14467 7616 14476
rect 7564 14433 7573 14467
rect 7573 14433 7607 14467
rect 7607 14433 7616 14467
rect 7564 14424 7616 14433
rect 8668 14424 8720 14476
rect 6000 14288 6052 14340
rect 5264 14220 5316 14272
rect 8208 14356 8260 14408
rect 14832 14356 14884 14408
rect 16120 14399 16172 14408
rect 9680 14288 9732 14340
rect 9772 14220 9824 14272
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 12072 14288 12124 14340
rect 12532 14288 12584 14340
rect 13268 14220 13320 14272
rect 16120 14365 16129 14399
rect 16129 14365 16163 14399
rect 16163 14365 16172 14399
rect 16120 14356 16172 14365
rect 19708 14356 19760 14408
rect 15108 14288 15160 14340
rect 16028 14288 16080 14340
rect 20536 14288 20588 14340
rect 17040 14220 17092 14272
rect 21272 14263 21324 14272
rect 21272 14229 21281 14263
rect 21281 14229 21315 14263
rect 21315 14229 21324 14263
rect 21272 14220 21324 14229
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 4436 14016 4488 14068
rect 6644 14016 6696 14068
rect 8668 14016 8720 14068
rect 9772 14059 9824 14068
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 13084 14059 13136 14068
rect 7472 13948 7524 14000
rect 9312 13948 9364 14000
rect 5080 13923 5132 13932
rect 5080 13889 5089 13923
rect 5089 13889 5123 13923
rect 5123 13889 5132 13923
rect 5080 13880 5132 13889
rect 7104 13880 7156 13932
rect 8668 13880 8720 13932
rect 10048 13880 10100 13932
rect 7288 13812 7340 13864
rect 12348 13812 12400 13864
rect 13084 14025 13093 14059
rect 13093 14025 13127 14059
rect 13127 14025 13136 14059
rect 13084 14016 13136 14025
rect 15108 14059 15160 14068
rect 15108 14025 15117 14059
rect 15117 14025 15151 14059
rect 15151 14025 15160 14059
rect 15108 14016 15160 14025
rect 16028 14059 16080 14068
rect 13176 13948 13228 14000
rect 12808 13880 12860 13932
rect 13360 13923 13412 13932
rect 13360 13889 13369 13923
rect 13369 13889 13403 13923
rect 13403 13889 13412 13923
rect 13360 13880 13412 13889
rect 16028 14025 16037 14059
rect 16037 14025 16071 14059
rect 16071 14025 16080 14059
rect 16028 14016 16080 14025
rect 19708 14059 19760 14068
rect 19708 14025 19717 14059
rect 19717 14025 19751 14059
rect 19751 14025 19760 14059
rect 19708 14016 19760 14025
rect 17960 13948 18012 14000
rect 18880 13948 18932 14000
rect 19064 13948 19116 14000
rect 17316 13923 17368 13932
rect 17316 13889 17325 13923
rect 17325 13889 17359 13923
rect 17359 13889 17368 13923
rect 17316 13880 17368 13889
rect 18512 13880 18564 13932
rect 20628 13923 20680 13932
rect 20628 13889 20637 13923
rect 20637 13889 20671 13923
rect 20671 13889 20680 13923
rect 20628 13880 20680 13889
rect 21088 13923 21140 13932
rect 21088 13889 21097 13923
rect 21097 13889 21131 13923
rect 21131 13889 21140 13923
rect 21088 13880 21140 13889
rect 14372 13812 14424 13864
rect 14924 13855 14976 13864
rect 14924 13821 14933 13855
rect 14933 13821 14967 13855
rect 14967 13821 14976 13855
rect 14924 13812 14976 13821
rect 12900 13744 12952 13796
rect 5908 13676 5960 13728
rect 11612 13676 11664 13728
rect 11796 13676 11848 13728
rect 19984 13855 20036 13864
rect 19984 13821 19993 13855
rect 19993 13821 20027 13855
rect 20027 13821 20036 13855
rect 19984 13812 20036 13821
rect 20996 13676 21048 13728
rect 21272 13719 21324 13728
rect 21272 13685 21281 13719
rect 21281 13685 21315 13719
rect 21315 13685 21324 13719
rect 21272 13676 21324 13685
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 7012 13472 7064 13524
rect 7564 13472 7616 13524
rect 9680 13515 9732 13524
rect 9680 13481 9689 13515
rect 9689 13481 9723 13515
rect 9723 13481 9732 13515
rect 9680 13472 9732 13481
rect 12716 13472 12768 13524
rect 18512 13515 18564 13524
rect 18512 13481 18521 13515
rect 18521 13481 18555 13515
rect 18555 13481 18564 13515
rect 18512 13472 18564 13481
rect 19064 13472 19116 13524
rect 20352 13472 20404 13524
rect 21548 13472 21600 13524
rect 2228 13268 2280 13320
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 8668 13336 8720 13388
rect 9128 13336 9180 13388
rect 10324 13379 10376 13388
rect 10324 13345 10333 13379
rect 10333 13345 10367 13379
rect 10367 13345 10376 13379
rect 10324 13336 10376 13345
rect 11612 13404 11664 13456
rect 17408 13447 17460 13456
rect 17408 13413 17417 13447
rect 17417 13413 17451 13447
rect 17451 13413 17460 13447
rect 17408 13404 17460 13413
rect 11796 13268 11848 13320
rect 12900 13336 12952 13388
rect 17960 13379 18012 13388
rect 17960 13345 17969 13379
rect 17969 13345 18003 13379
rect 18003 13345 18012 13379
rect 17960 13336 18012 13345
rect 18052 13268 18104 13320
rect 19984 13268 20036 13320
rect 20076 13268 20128 13320
rect 20996 13311 21048 13320
rect 20996 13277 21005 13311
rect 21005 13277 21039 13311
rect 21039 13277 21048 13311
rect 20996 13268 21048 13277
rect 17684 13200 17736 13252
rect 21180 13200 21232 13252
rect 9588 13132 9640 13184
rect 12440 13132 12492 13184
rect 13544 13132 13596 13184
rect 17408 13132 17460 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 6000 12928 6052 12980
rect 12072 12971 12124 12980
rect 12072 12937 12081 12971
rect 12081 12937 12115 12971
rect 12115 12937 12124 12971
rect 12072 12928 12124 12937
rect 20536 12971 20588 12980
rect 10324 12860 10376 12912
rect 14832 12860 14884 12912
rect 16580 12860 16632 12912
rect 17684 12903 17736 12912
rect 17684 12869 17693 12903
rect 17693 12869 17727 12903
rect 17727 12869 17736 12903
rect 17684 12860 17736 12869
rect 20536 12937 20545 12971
rect 20545 12937 20579 12971
rect 20579 12937 20588 12971
rect 20536 12928 20588 12937
rect 20812 12971 20864 12980
rect 20812 12937 20821 12971
rect 20821 12937 20855 12971
rect 20855 12937 20864 12971
rect 20812 12928 20864 12937
rect 21364 12971 21416 12980
rect 21364 12937 21373 12971
rect 21373 12937 21407 12971
rect 21407 12937 21416 12971
rect 21364 12928 21416 12937
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 11796 12792 11848 12844
rect 12900 12792 12952 12844
rect 17316 12792 17368 12844
rect 19248 12792 19300 12844
rect 19524 12792 19576 12844
rect 17132 12767 17184 12776
rect 17132 12733 17141 12767
rect 17141 12733 17175 12767
rect 17175 12733 17184 12767
rect 17132 12724 17184 12733
rect 17224 12767 17276 12776
rect 17224 12733 17233 12767
rect 17233 12733 17267 12767
rect 17267 12733 17276 12767
rect 17224 12724 17276 12733
rect 18420 12724 18472 12776
rect 19984 12656 20036 12708
rect 20720 12656 20772 12708
rect 9588 12588 9640 12640
rect 16580 12588 16632 12640
rect 16948 12588 17000 12640
rect 18604 12588 18656 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 8300 12384 8352 12436
rect 9588 12384 9640 12436
rect 10048 12384 10100 12436
rect 12900 12427 12952 12436
rect 7932 12291 7984 12300
rect 7932 12257 7941 12291
rect 7941 12257 7975 12291
rect 7975 12257 7984 12291
rect 7932 12248 7984 12257
rect 8024 12248 8076 12300
rect 7288 12180 7340 12232
rect 8392 12180 8444 12232
rect 9496 12180 9548 12232
rect 11612 12180 11664 12232
rect 8300 12112 8352 12164
rect 11152 12112 11204 12164
rect 12900 12393 12909 12427
rect 12909 12393 12943 12427
rect 12943 12393 12952 12427
rect 12900 12384 12952 12393
rect 17132 12384 17184 12436
rect 17316 12427 17368 12436
rect 17316 12393 17325 12427
rect 17325 12393 17359 12427
rect 17359 12393 17368 12427
rect 17316 12384 17368 12393
rect 20444 12384 20496 12436
rect 21088 12384 21140 12436
rect 18420 12316 18472 12368
rect 17776 12248 17828 12300
rect 15016 12180 15068 12232
rect 16028 12223 16080 12232
rect 16028 12189 16037 12223
rect 16037 12189 16071 12223
rect 16071 12189 16080 12223
rect 16028 12180 16080 12189
rect 16580 12223 16632 12232
rect 16580 12189 16589 12223
rect 16589 12189 16623 12223
rect 16623 12189 16632 12223
rect 16580 12180 16632 12189
rect 17684 12180 17736 12232
rect 17960 12180 18012 12232
rect 18604 12180 18656 12232
rect 8668 12044 8720 12096
rect 10784 12087 10836 12096
rect 10784 12053 10793 12087
rect 10793 12053 10827 12087
rect 10827 12053 10836 12087
rect 10784 12044 10836 12053
rect 10876 12044 10928 12096
rect 14556 12044 14608 12096
rect 15476 12044 15528 12096
rect 17132 12112 17184 12164
rect 17960 12044 18012 12096
rect 18052 12044 18104 12096
rect 19064 12044 19116 12096
rect 19340 12044 19392 12096
rect 19708 12044 19760 12096
rect 20720 12180 20772 12232
rect 21364 12087 21416 12096
rect 21364 12053 21373 12087
rect 21373 12053 21407 12087
rect 21407 12053 21416 12087
rect 21364 12044 21416 12053
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 8668 11883 8720 11892
rect 8668 11849 8677 11883
rect 8677 11849 8711 11883
rect 8711 11849 8720 11883
rect 8668 11840 8720 11849
rect 10232 11840 10284 11892
rect 10876 11840 10928 11892
rect 11152 11883 11204 11892
rect 11152 11849 11161 11883
rect 11161 11849 11195 11883
rect 11195 11849 11204 11883
rect 11152 11840 11204 11849
rect 11796 11840 11848 11892
rect 12348 11840 12400 11892
rect 9956 11772 10008 11824
rect 2136 11704 2188 11756
rect 10784 11772 10836 11824
rect 9496 11636 9548 11688
rect 9956 11679 10008 11688
rect 9956 11645 9965 11679
rect 9965 11645 9999 11679
rect 9999 11645 10008 11679
rect 11336 11704 11388 11756
rect 9956 11636 10008 11645
rect 11796 11636 11848 11688
rect 14556 11840 14608 11892
rect 16948 11883 17000 11892
rect 16948 11849 16957 11883
rect 16957 11849 16991 11883
rect 16991 11849 17000 11883
rect 16948 11840 17000 11849
rect 18052 11883 18104 11892
rect 18052 11849 18061 11883
rect 18061 11849 18095 11883
rect 18095 11849 18104 11883
rect 18052 11840 18104 11849
rect 15292 11704 15344 11756
rect 15476 11747 15528 11756
rect 15476 11713 15485 11747
rect 15485 11713 15519 11747
rect 15519 11713 15528 11747
rect 17776 11772 17828 11824
rect 19892 11840 19944 11892
rect 20260 11840 20312 11892
rect 21640 11840 21692 11892
rect 15476 11704 15528 11713
rect 13176 11543 13228 11552
rect 13176 11509 13185 11543
rect 13185 11509 13219 11543
rect 13219 11509 13228 11543
rect 13176 11500 13228 11509
rect 14280 11500 14332 11552
rect 16028 11636 16080 11688
rect 17960 11704 18012 11756
rect 19156 11747 19208 11756
rect 19156 11713 19165 11747
rect 19165 11713 19199 11747
rect 19199 11713 19208 11747
rect 19156 11704 19208 11713
rect 17132 11636 17184 11688
rect 19524 11568 19576 11620
rect 15292 11500 15344 11552
rect 21180 11772 21232 11824
rect 19892 11747 19944 11756
rect 19892 11713 19901 11747
rect 19901 11713 19935 11747
rect 19935 11713 19944 11747
rect 19892 11704 19944 11713
rect 20536 11747 20588 11756
rect 20536 11713 20545 11747
rect 20545 11713 20579 11747
rect 20579 11713 20588 11747
rect 20536 11704 20588 11713
rect 20996 11747 21048 11756
rect 20996 11713 21005 11747
rect 21005 11713 21039 11747
rect 21039 11713 21048 11747
rect 20996 11704 21048 11713
rect 21180 11500 21232 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 9588 11296 9640 11348
rect 11336 11339 11388 11348
rect 7932 11160 7984 11212
rect 11336 11305 11345 11339
rect 11345 11305 11379 11339
rect 11379 11305 11388 11339
rect 11336 11296 11388 11305
rect 11796 11296 11848 11348
rect 8392 11092 8444 11144
rect 9956 11092 10008 11144
rect 11244 11092 11296 11144
rect 11980 11228 12032 11280
rect 14464 11296 14516 11348
rect 19892 11296 19944 11348
rect 20536 11339 20588 11348
rect 20536 11305 20545 11339
rect 20545 11305 20579 11339
rect 20579 11305 20588 11339
rect 20536 11296 20588 11305
rect 21916 11296 21968 11348
rect 13176 11203 13228 11212
rect 13176 11169 13185 11203
rect 13185 11169 13219 11203
rect 13219 11169 13228 11203
rect 13176 11160 13228 11169
rect 13820 11160 13872 11212
rect 15476 11228 15528 11280
rect 14464 11160 14516 11212
rect 19708 11160 19760 11212
rect 14556 11092 14608 11144
rect 19248 11135 19300 11144
rect 19248 11101 19257 11135
rect 19257 11101 19291 11135
rect 19291 11101 19300 11135
rect 19248 11092 19300 11101
rect 13544 11024 13596 11076
rect 14464 11067 14516 11076
rect 14464 11033 14473 11067
rect 14473 11033 14507 11067
rect 14507 11033 14516 11067
rect 14464 11024 14516 11033
rect 15200 11067 15252 11076
rect 15200 11033 15209 11067
rect 15209 11033 15243 11067
rect 15243 11033 15252 11067
rect 15200 11024 15252 11033
rect 17040 11024 17092 11076
rect 17684 11024 17736 11076
rect 20904 11092 20956 11144
rect 21364 11067 21416 11076
rect 21364 11033 21373 11067
rect 21373 11033 21407 11067
rect 21407 11033 21416 11067
rect 21364 11024 21416 11033
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 10048 10752 10100 10804
rect 11244 10752 11296 10804
rect 12348 10752 12400 10804
rect 15016 10795 15068 10804
rect 15016 10761 15025 10795
rect 15025 10761 15059 10795
rect 15059 10761 15068 10795
rect 15016 10752 15068 10761
rect 15476 10795 15528 10804
rect 15476 10761 15485 10795
rect 15485 10761 15519 10795
rect 15519 10761 15528 10795
rect 15476 10752 15528 10761
rect 17132 10752 17184 10804
rect 19248 10752 19300 10804
rect 20904 10795 20956 10804
rect 20904 10761 20913 10795
rect 20913 10761 20947 10795
rect 20947 10761 20956 10795
rect 20904 10752 20956 10761
rect 20996 10752 21048 10804
rect 10324 10684 10376 10736
rect 17776 10727 17828 10736
rect 17776 10693 17794 10727
rect 17794 10693 17828 10727
rect 17776 10684 17828 10693
rect 11980 10659 12032 10668
rect 11980 10625 11989 10659
rect 11989 10625 12023 10659
rect 12023 10625 12032 10659
rect 11980 10616 12032 10625
rect 15752 10616 15804 10668
rect 18880 10659 18932 10668
rect 18880 10625 18889 10659
rect 18889 10625 18923 10659
rect 18923 10625 18932 10659
rect 18880 10616 18932 10625
rect 21456 10616 21508 10668
rect 9956 10480 10008 10532
rect 12532 10548 12584 10600
rect 18512 10548 18564 10600
rect 19524 10548 19576 10600
rect 19984 10591 20036 10600
rect 19984 10557 19993 10591
rect 19993 10557 20027 10591
rect 20027 10557 20036 10591
rect 19984 10548 20036 10557
rect 8392 10412 8444 10464
rect 14280 10455 14332 10464
rect 14280 10421 14289 10455
rect 14289 10421 14323 10455
rect 14323 10421 14332 10455
rect 14280 10412 14332 10421
rect 19892 10412 19944 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 9956 10208 10008 10260
rect 11704 10072 11756 10124
rect 12440 10004 12492 10056
rect 14280 10208 14332 10260
rect 15752 10251 15804 10260
rect 15752 10217 15761 10251
rect 15761 10217 15795 10251
rect 15795 10217 15804 10251
rect 15752 10208 15804 10217
rect 17776 10208 17828 10260
rect 19524 10251 19576 10260
rect 19524 10217 19533 10251
rect 19533 10217 19567 10251
rect 19567 10217 19576 10251
rect 19524 10208 19576 10217
rect 11888 9936 11940 9988
rect 12532 9868 12584 9920
rect 13820 9936 13872 9988
rect 14556 9868 14608 9920
rect 20076 10115 20128 10124
rect 20076 10081 20085 10115
rect 20085 10081 20119 10115
rect 20119 10081 20128 10115
rect 20076 10072 20128 10081
rect 18512 10047 18564 10056
rect 18512 10013 18521 10047
rect 18521 10013 18555 10047
rect 18555 10013 18564 10047
rect 18512 10004 18564 10013
rect 19892 10047 19944 10056
rect 19892 10013 19901 10047
rect 19901 10013 19935 10047
rect 19935 10013 19944 10047
rect 19892 10004 19944 10013
rect 19984 10004 20036 10056
rect 16120 9911 16172 9920
rect 16120 9877 16129 9911
rect 16129 9877 16163 9911
rect 16163 9877 16172 9911
rect 16120 9868 16172 9877
rect 16948 9868 17000 9920
rect 17224 9868 17276 9920
rect 18052 9868 18104 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 11888 9707 11940 9716
rect 11888 9673 11897 9707
rect 11897 9673 11931 9707
rect 11931 9673 11940 9707
rect 11888 9664 11940 9673
rect 16120 9664 16172 9716
rect 19984 9664 20036 9716
rect 21456 9664 21508 9716
rect 13360 9596 13412 9648
rect 20904 9596 20956 9648
rect 12532 9571 12584 9580
rect 12532 9537 12541 9571
rect 12541 9537 12575 9571
rect 12575 9537 12584 9571
rect 12532 9528 12584 9537
rect 16304 9528 16356 9580
rect 19616 9528 19668 9580
rect 20996 9571 21048 9580
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 13820 9503 13872 9512
rect 13820 9469 13829 9503
rect 13829 9469 13863 9503
rect 13863 9469 13872 9503
rect 13820 9460 13872 9469
rect 14372 9460 14424 9512
rect 14832 9460 14884 9512
rect 18236 9460 18288 9512
rect 18512 9460 18564 9512
rect 14464 9435 14516 9444
rect 14464 9401 14473 9435
rect 14473 9401 14507 9435
rect 14507 9401 14516 9435
rect 14464 9392 14516 9401
rect 15936 9392 15988 9444
rect 21272 9392 21324 9444
rect 20536 9367 20588 9376
rect 20536 9333 20545 9367
rect 20545 9333 20579 9367
rect 20579 9333 20588 9367
rect 20536 9324 20588 9333
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 12256 9120 12308 9172
rect 13452 9163 13504 9172
rect 13452 9129 13461 9163
rect 13461 9129 13495 9163
rect 13495 9129 13504 9163
rect 13452 9120 13504 9129
rect 16304 9163 16356 9172
rect 16304 9129 16313 9163
rect 16313 9129 16347 9163
rect 16347 9129 16356 9163
rect 16304 9120 16356 9129
rect 19616 9163 19668 9172
rect 19616 9129 19625 9163
rect 19625 9129 19659 9163
rect 19659 9129 19668 9163
rect 19616 9120 19668 9129
rect 21824 9120 21876 9172
rect 11152 8916 11204 8968
rect 13452 8916 13504 8968
rect 16948 8916 17000 8968
rect 19616 8916 19668 8968
rect 20076 8916 20128 8968
rect 20536 8959 20588 8968
rect 20536 8925 20545 8959
rect 20545 8925 20579 8959
rect 20579 8925 20588 8959
rect 20536 8916 20588 8925
rect 20628 8916 20680 8968
rect 14832 8823 14884 8832
rect 14832 8789 14841 8823
rect 14841 8789 14875 8823
rect 14875 8789 14884 8823
rect 14832 8780 14884 8789
rect 17316 8780 17368 8832
rect 20720 8823 20772 8832
rect 20720 8789 20729 8823
rect 20729 8789 20763 8823
rect 20763 8789 20772 8823
rect 20720 8780 20772 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 11152 8619 11204 8628
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 13452 8619 13504 8628
rect 13452 8585 13461 8619
rect 13461 8585 13495 8619
rect 13495 8585 13504 8619
rect 13452 8576 13504 8585
rect 19616 8619 19668 8628
rect 19616 8585 19625 8619
rect 19625 8585 19659 8619
rect 19659 8585 19668 8619
rect 19616 8576 19668 8585
rect 20628 8576 20680 8628
rect 21364 8619 21416 8628
rect 18696 8508 18748 8560
rect 19248 8508 19300 8560
rect 9404 8483 9456 8492
rect 9404 8449 9413 8483
rect 9413 8449 9447 8483
rect 9447 8449 9456 8483
rect 9404 8440 9456 8449
rect 11244 8440 11296 8492
rect 11520 8483 11572 8492
rect 11520 8449 11529 8483
rect 11529 8449 11563 8483
rect 11563 8449 11572 8483
rect 11520 8440 11572 8449
rect 13820 8440 13872 8492
rect 15292 8440 15344 8492
rect 17132 8483 17184 8492
rect 17132 8449 17141 8483
rect 17141 8449 17175 8483
rect 17175 8449 17184 8483
rect 17132 8440 17184 8449
rect 19800 8440 19852 8492
rect 21364 8585 21373 8619
rect 21373 8585 21407 8619
rect 21407 8585 21416 8619
rect 21364 8576 21416 8585
rect 12532 8372 12584 8424
rect 14464 8415 14516 8424
rect 14464 8381 14473 8415
rect 14473 8381 14507 8415
rect 14507 8381 14516 8415
rect 14464 8372 14516 8381
rect 18236 8415 18288 8424
rect 18236 8381 18245 8415
rect 18245 8381 18279 8415
rect 18279 8381 18288 8415
rect 18236 8372 18288 8381
rect 21088 8440 21140 8492
rect 19248 8304 19300 8356
rect 10048 8279 10100 8288
rect 10048 8245 10057 8279
rect 10057 8245 10091 8279
rect 10091 8245 10100 8279
rect 10048 8236 10100 8245
rect 12164 8279 12216 8288
rect 12164 8245 12173 8279
rect 12173 8245 12207 8279
rect 12207 8245 12216 8279
rect 12164 8236 12216 8245
rect 16120 8279 16172 8288
rect 16120 8245 16129 8279
rect 16129 8245 16163 8279
rect 16163 8245 16172 8279
rect 16120 8236 16172 8245
rect 17776 8279 17828 8288
rect 17776 8245 17785 8279
rect 17785 8245 17819 8279
rect 17819 8245 17828 8279
rect 17776 8236 17828 8245
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 19800 8032 19852 8084
rect 20812 8007 20864 8016
rect 20812 7973 20821 8007
rect 20821 7973 20855 8007
rect 20855 7973 20864 8007
rect 20812 7964 20864 7973
rect 21364 7939 21416 7948
rect 8392 7828 8444 7880
rect 10048 7871 10100 7880
rect 10048 7837 10082 7871
rect 10082 7837 10100 7871
rect 10048 7828 10100 7837
rect 12440 7828 12492 7880
rect 18236 7828 18288 7880
rect 21364 7905 21373 7939
rect 21373 7905 21407 7939
rect 21407 7905 21416 7939
rect 21364 7896 21416 7905
rect 11520 7760 11572 7812
rect 12164 7760 12216 7812
rect 13728 7760 13780 7812
rect 16120 7760 16172 7812
rect 17776 7760 17828 7812
rect 12072 7692 12124 7744
rect 13176 7692 13228 7744
rect 15292 7692 15344 7744
rect 17132 7735 17184 7744
rect 17132 7701 17141 7735
rect 17141 7701 17175 7735
rect 17175 7701 17184 7735
rect 17132 7692 17184 7701
rect 17592 7692 17644 7744
rect 20720 7828 20772 7880
rect 20720 7692 20772 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 9404 7531 9456 7540
rect 9404 7497 9413 7531
rect 9413 7497 9447 7531
rect 9447 7497 9456 7531
rect 9404 7488 9456 7497
rect 11244 7488 11296 7540
rect 12532 7488 12584 7540
rect 13728 7531 13780 7540
rect 13728 7497 13737 7531
rect 13737 7497 13771 7531
rect 13771 7497 13780 7531
rect 13728 7488 13780 7497
rect 13820 7488 13872 7540
rect 14464 7488 14516 7540
rect 15476 7531 15528 7540
rect 15476 7497 15485 7531
rect 15485 7497 15519 7531
rect 15519 7497 15528 7531
rect 15476 7488 15528 7497
rect 16948 7531 17000 7540
rect 16948 7497 16957 7531
rect 16957 7497 16991 7531
rect 16991 7497 17000 7531
rect 16948 7488 17000 7497
rect 17316 7531 17368 7540
rect 17316 7497 17325 7531
rect 17325 7497 17359 7531
rect 17359 7497 17368 7531
rect 17316 7488 17368 7497
rect 8392 7420 8444 7472
rect 13176 7420 13228 7472
rect 8300 7395 8352 7404
rect 8300 7361 8334 7395
rect 8334 7361 8352 7395
rect 8300 7352 8352 7361
rect 11980 7327 12032 7336
rect 11980 7293 11989 7327
rect 11989 7293 12023 7327
rect 12023 7293 12032 7327
rect 11980 7284 12032 7293
rect 12072 7327 12124 7336
rect 12072 7293 12081 7327
rect 12081 7293 12115 7327
rect 12115 7293 12124 7327
rect 12072 7284 12124 7293
rect 15292 7284 15344 7336
rect 17132 7420 17184 7472
rect 17592 7327 17644 7336
rect 17592 7293 17601 7327
rect 17601 7293 17635 7327
rect 17635 7293 17644 7327
rect 17592 7284 17644 7293
rect 18052 7284 18104 7336
rect 19892 7395 19944 7404
rect 19892 7361 19901 7395
rect 19901 7361 19935 7395
rect 19935 7361 19944 7395
rect 19892 7352 19944 7361
rect 20996 7488 21048 7540
rect 20444 7420 20496 7472
rect 21088 7420 21140 7472
rect 21180 7352 21232 7404
rect 21548 7352 21600 7404
rect 20904 7284 20956 7336
rect 21088 7216 21140 7268
rect 17868 7148 17920 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 11980 6944 12032 6996
rect 21548 6944 21600 6996
rect 9404 6808 9456 6860
rect 16396 6808 16448 6860
rect 15476 6740 15528 6792
rect 18052 6740 18104 6792
rect 20444 6740 20496 6792
rect 20720 6740 20772 6792
rect 3976 6604 4028 6656
rect 20168 6672 20220 6724
rect 17500 6604 17552 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 8300 6400 8352 6452
rect 21180 6443 21232 6452
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 21180 6409 21189 6443
rect 21189 6409 21223 6443
rect 21223 6409 21232 6443
rect 21180 6400 21232 6409
rect 20536 6332 20588 6384
rect 20536 6196 20588 6248
rect 14648 6128 14700 6180
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 14740 5788 14792 5840
rect 20352 5695 20404 5704
rect 20352 5661 20361 5695
rect 20361 5661 20395 5695
rect 20395 5661 20404 5695
rect 20352 5652 20404 5661
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 20720 5355 20772 5364
rect 20720 5321 20729 5355
rect 20729 5321 20763 5355
rect 20763 5321 20772 5355
rect 20720 5312 20772 5321
rect 20904 5312 20956 5364
rect 20628 5244 20680 5296
rect 20904 5219 20956 5228
rect 20904 5185 20913 5219
rect 20913 5185 20947 5219
rect 20947 5185 20956 5219
rect 20904 5176 20956 5185
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 20168 4768 20220 4820
rect 20904 4811 20956 4820
rect 20904 4777 20913 4811
rect 20913 4777 20947 4811
rect 20947 4777 20956 4811
rect 20904 4768 20956 4777
rect 21088 4768 21140 4820
rect 20444 4607 20496 4616
rect 20444 4573 20453 4607
rect 20453 4573 20487 4607
rect 20487 4573 20496 4607
rect 20444 4564 20496 4573
rect 20720 4607 20772 4616
rect 20720 4573 20729 4607
rect 20729 4573 20763 4607
rect 20763 4573 20772 4607
rect 20720 4564 20772 4573
rect 21364 4607 21416 4616
rect 21364 4573 21373 4607
rect 21373 4573 21407 4607
rect 21407 4573 21416 4607
rect 21364 4564 21416 4573
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 20444 4224 20496 4276
rect 21180 4267 21232 4276
rect 21180 4233 21189 4267
rect 21189 4233 21223 4267
rect 21223 4233 21232 4267
rect 21180 4224 21232 4233
rect 21272 4199 21324 4208
rect 21272 4165 21281 4199
rect 21281 4165 21315 4199
rect 21315 4165 21324 4199
rect 21272 4156 21324 4165
rect 21364 4088 21416 4140
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 17960 3612 18012 3664
rect 17224 3544 17276 3596
rect 20536 3519 20588 3528
rect 20536 3485 20545 3519
rect 20545 3485 20579 3519
rect 20579 3485 20588 3519
rect 20536 3476 20588 3485
rect 20168 3451 20220 3460
rect 20168 3417 20177 3451
rect 20177 3417 20211 3451
rect 20211 3417 20220 3451
rect 20168 3408 20220 3417
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 19064 3136 19116 3188
rect 20720 3111 20772 3120
rect 20720 3077 20729 3111
rect 20729 3077 20763 3111
rect 20763 3077 20772 3111
rect 20720 3068 20772 3077
rect 19064 3000 19116 3052
rect 21272 3043 21324 3052
rect 21272 3009 21281 3043
rect 21281 3009 21315 3043
rect 21315 3009 21324 3043
rect 21272 3000 21324 3009
rect 15200 2864 15252 2916
rect 19616 2839 19668 2848
rect 19616 2805 19625 2839
rect 19625 2805 19659 2839
rect 19659 2805 19668 2839
rect 19616 2796 19668 2805
rect 19708 2796 19760 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 17040 2524 17092 2576
rect 20812 2499 20864 2508
rect 20812 2465 20821 2499
rect 20821 2465 20855 2499
rect 20855 2465 20864 2499
rect 20812 2456 20864 2465
rect 14832 2388 14884 2440
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 19616 2363 19668 2372
rect 19616 2329 19625 2363
rect 19625 2329 19659 2363
rect 19659 2329 19668 2363
rect 19616 2320 19668 2329
rect 19248 2252 19300 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
<< metal2 >>
rect 294 22200 350 23000
rect 846 22200 902 23000
rect 952 22222 1348 22250
rect 308 20534 336 22200
rect 860 22114 888 22200
rect 952 22114 980 22222
rect 860 22086 980 22114
rect 296 20528 348 20534
rect 296 20470 348 20476
rect 1320 19938 1348 22222
rect 1398 22200 1454 23000
rect 1950 22200 2006 23000
rect 2502 22200 2558 23000
rect 2792 22222 3004 22250
rect 1412 20074 1440 22200
rect 1676 20324 1728 20330
rect 1676 20266 1728 20272
rect 1412 20046 1532 20074
rect 1688 20058 1716 20266
rect 1320 19922 1440 19938
rect 1320 19916 1452 19922
rect 1320 19910 1400 19916
rect 1400 19858 1452 19864
rect 1504 19854 1532 20046
rect 1676 20052 1728 20058
rect 1676 19994 1728 20000
rect 1492 19848 1544 19854
rect 1492 19790 1544 19796
rect 1504 18170 1532 19790
rect 1964 19378 1992 22200
rect 2412 20528 2464 20534
rect 2412 20470 2464 20476
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 1952 19372 2004 19378
rect 1952 19314 2004 19320
rect 1964 18970 1992 19314
rect 1952 18964 2004 18970
rect 1952 18906 2004 18912
rect 2056 18426 2084 19790
rect 2136 19712 2188 19718
rect 2136 19654 2188 19660
rect 2044 18420 2096 18426
rect 2044 18362 2096 18368
rect 1674 18320 1730 18329
rect 1674 18255 1676 18264
rect 1728 18255 1730 18264
rect 1676 18226 1728 18232
rect 1504 18142 1624 18170
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1504 17241 1532 18022
rect 1596 17814 1624 18142
rect 1584 17808 1636 17814
rect 1584 17750 1636 17756
rect 1584 17672 1636 17678
rect 1584 17614 1636 17620
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1596 16998 1624 17614
rect 1584 16992 1636 16998
rect 1584 16934 1636 16940
rect 1596 16658 1624 16934
rect 1584 16652 1636 16658
rect 1584 16594 1636 16600
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2056 15706 2084 16050
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2148 11762 2176 19654
rect 2228 19168 2280 19174
rect 2228 19110 2280 19116
rect 2240 13326 2268 19110
rect 2320 18692 2372 18698
rect 2320 18634 2372 18640
rect 2332 17882 2360 18634
rect 2424 18358 2452 20470
rect 2516 20346 2544 22200
rect 2792 20482 2820 22222
rect 2976 22114 3004 22222
rect 3054 22200 3110 23000
rect 3606 22200 3662 23000
rect 4158 22200 4214 23000
rect 4448 22222 4660 22250
rect 3068 22114 3096 22200
rect 2976 22086 3096 22114
rect 3240 20596 3292 20602
rect 3240 20538 3292 20544
rect 2700 20466 2820 20482
rect 3148 20528 3200 20534
rect 3148 20470 3200 20476
rect 2688 20460 2820 20466
rect 2740 20454 2820 20460
rect 2688 20402 2740 20408
rect 2516 20318 2636 20346
rect 2504 20256 2556 20262
rect 2504 20198 2556 20204
rect 2412 18352 2464 18358
rect 2412 18294 2464 18300
rect 2320 17876 2372 17882
rect 2320 17818 2372 17824
rect 2516 15094 2544 20198
rect 2608 19854 2636 20318
rect 2596 19848 2648 19854
rect 2596 19790 2648 19796
rect 2608 19514 2636 19790
rect 2596 19508 2648 19514
rect 2596 19450 2648 19456
rect 2700 18426 2728 20402
rect 2964 20256 3016 20262
rect 2964 20198 3016 20204
rect 2976 19990 3004 20198
rect 2964 19984 3016 19990
rect 2964 19926 3016 19932
rect 3160 18426 3188 20470
rect 3252 20466 3280 20538
rect 3240 20460 3292 20466
rect 3240 20402 3292 20408
rect 3252 19446 3280 20402
rect 3620 20346 3648 22200
rect 4172 20618 4200 22200
rect 4080 20590 4200 20618
rect 4448 20602 4476 22222
rect 4632 22114 4660 22222
rect 4710 22200 4766 23000
rect 5262 22200 5318 23000
rect 5814 22200 5870 23000
rect 6458 22200 6514 23000
rect 6564 22222 6776 22250
rect 4724 22114 4752 22200
rect 4632 22086 4752 22114
rect 4436 20596 4488 20602
rect 4080 20534 4108 20590
rect 4436 20538 4488 20544
rect 4068 20528 4120 20534
rect 4068 20470 4120 20476
rect 5276 20398 5304 22200
rect 5828 20618 5856 22200
rect 6472 22114 6500 22200
rect 6564 22114 6592 22222
rect 6472 22086 6592 22114
rect 6148 20700 6456 20720
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20624 6456 20644
rect 5736 20590 5856 20618
rect 5736 20534 5764 20590
rect 5724 20528 5776 20534
rect 5724 20470 5776 20476
rect 5356 20460 5408 20466
rect 5356 20402 5408 20408
rect 3436 20318 3648 20346
rect 3792 20392 3844 20398
rect 4252 20392 4304 20398
rect 3844 20340 3924 20346
rect 3792 20334 3924 20340
rect 4252 20334 4304 20340
rect 5264 20392 5316 20398
rect 5264 20334 5316 20340
rect 3804 20318 3924 20334
rect 3332 20256 3384 20262
rect 3332 20198 3384 20204
rect 3344 19922 3372 20198
rect 3332 19916 3384 19922
rect 3332 19858 3384 19864
rect 3436 19854 3464 20318
rect 3549 20156 3857 20176
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20080 3857 20100
rect 3424 19848 3476 19854
rect 3424 19790 3476 19796
rect 3332 19712 3384 19718
rect 3332 19654 3384 19660
rect 3240 19440 3292 19446
rect 3240 19382 3292 19388
rect 2688 18420 2740 18426
rect 2688 18362 2740 18368
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 3148 17536 3200 17542
rect 3148 17478 3200 17484
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 2976 16658 3004 16934
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 3160 16590 3188 17478
rect 3344 17338 3372 19654
rect 3436 19514 3464 19790
rect 3424 19508 3476 19514
rect 3424 19450 3476 19456
rect 3424 19372 3476 19378
rect 3424 19314 3476 19320
rect 3436 18766 3464 19314
rect 3549 19068 3857 19088
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 18992 3857 19012
rect 3424 18760 3476 18766
rect 3424 18702 3476 18708
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3332 17196 3384 17202
rect 3332 17138 3384 17144
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3344 16046 3372 17138
rect 3436 17134 3464 18702
rect 3896 18408 3924 20318
rect 4068 20256 4120 20262
rect 4068 20198 4120 20204
rect 3976 19372 4028 19378
rect 3976 19314 4028 19320
rect 3988 18970 4016 19314
rect 3976 18964 4028 18970
rect 3976 18906 4028 18912
rect 3896 18380 4016 18408
rect 3549 17980 3857 18000
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17904 3857 17924
rect 3424 17128 3476 17134
rect 3424 17070 3476 17076
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 3436 16658 3464 17070
rect 3549 16892 3857 16912
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16816 3857 16836
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3436 16182 3464 16594
rect 3424 16176 3476 16182
rect 3424 16118 3476 16124
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 2872 15496 2924 15502
rect 2872 15438 2924 15444
rect 2884 15162 2912 15438
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 2504 15088 2556 15094
rect 2504 15030 2556 15036
rect 3436 15026 3464 16118
rect 3896 15978 3924 17070
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3549 15804 3857 15824
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15728 3857 15748
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3424 15020 3476 15026
rect 3424 14962 3476 14968
rect 3252 14618 3280 14962
rect 3549 14716 3857 14736
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14640 3857 14660
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3549 13628 3857 13648
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13552 3857 13572
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 3549 12540 3857 12560
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12464 3857 12484
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 3549 11452 3857 11472
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11376 3857 11396
rect 3549 10364 3857 10384
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10288 3857 10308
rect 3549 9276 3857 9296
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9200 3857 9220
rect 3549 8188 3857 8208
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8112 3857 8132
rect 3549 7100 3857 7120
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7024 3857 7044
rect 3988 6662 4016 18380
rect 4080 17882 4108 20198
rect 4160 19916 4212 19922
rect 4160 19858 4212 19864
rect 4172 18698 4200 19858
rect 4160 18692 4212 18698
rect 4160 18634 4212 18640
rect 4264 18426 4292 20334
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 4344 19712 4396 19718
rect 4344 19654 4396 19660
rect 4712 19712 4764 19718
rect 4712 19654 4764 19660
rect 4356 18970 4384 19654
rect 4724 19310 4752 19654
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4344 18964 4396 18970
rect 4344 18906 4396 18912
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 4816 16590 4844 20198
rect 5264 19780 5316 19786
rect 5264 19722 5316 19728
rect 5080 19168 5132 19174
rect 5080 19110 5132 19116
rect 5092 18290 5120 19110
rect 5080 18284 5132 18290
rect 5080 18226 5132 18232
rect 5276 17338 5304 19722
rect 5368 19242 5396 20402
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5356 19236 5408 19242
rect 5356 19178 5408 19184
rect 5460 18834 5488 19314
rect 5736 18970 5764 20470
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5448 18828 5500 18834
rect 5448 18770 5500 18776
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5460 17338 5488 18022
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5632 17536 5684 17542
rect 5632 17478 5684 17484
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5448 17332 5500 17338
rect 5448 17274 5500 17280
rect 5644 17202 5672 17478
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5736 16794 5764 17614
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 4804 16584 4856 16590
rect 4804 16526 4856 16532
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4080 16250 4108 16390
rect 4068 16244 4120 16250
rect 4068 16186 4120 16192
rect 5736 15706 5764 16730
rect 5828 16726 5856 19654
rect 5816 16720 5868 16726
rect 5816 16662 5868 16668
rect 6012 16574 6040 20198
rect 6472 19786 6500 20402
rect 6748 19938 6776 22222
rect 7010 22200 7066 23000
rect 7562 22200 7618 23000
rect 8114 22200 8170 23000
rect 8312 22222 8616 22250
rect 6828 20392 6880 20398
rect 7024 20346 7052 22200
rect 6880 20340 7052 20346
rect 6828 20334 7052 20340
rect 6840 20318 7052 20334
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6840 20058 6868 20198
rect 6828 20052 6880 20058
rect 6828 19994 6880 20000
rect 6748 19910 6868 19938
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6460 19780 6512 19786
rect 6460 19722 6512 19728
rect 6552 19712 6604 19718
rect 6552 19654 6604 19660
rect 6148 19612 6456 19632
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19536 6456 19556
rect 6564 19378 6592 19654
rect 6552 19372 6604 19378
rect 6552 19314 6604 19320
rect 6148 18524 6456 18544
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18448 6456 18468
rect 6552 18216 6604 18222
rect 6552 18158 6604 18164
rect 6148 17436 6456 17456
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17360 6456 17380
rect 6564 17202 6592 18158
rect 6656 18154 6684 19790
rect 6736 19780 6788 19786
rect 6736 19722 6788 19728
rect 6748 19446 6776 19722
rect 6736 19440 6788 19446
rect 6736 19382 6788 19388
rect 6748 18902 6776 19382
rect 6736 18896 6788 18902
rect 6736 18838 6788 18844
rect 6840 18834 6868 19910
rect 6932 18970 6960 20318
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7012 19780 7064 19786
rect 7012 19722 7064 19728
rect 7024 19514 7052 19722
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 7288 19372 7340 19378
rect 7288 19314 7340 19320
rect 7300 18970 7328 19314
rect 6920 18964 6972 18970
rect 6920 18906 6972 18912
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7196 18896 7248 18902
rect 7248 18844 7328 18850
rect 7196 18838 7328 18844
rect 6828 18828 6880 18834
rect 7208 18822 7328 18838
rect 6828 18770 6880 18776
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7208 18426 7236 18702
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7104 18216 7156 18222
rect 7104 18158 7156 18164
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6656 17746 6684 18090
rect 7116 17882 7144 18158
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 7300 17202 7328 18822
rect 7392 17746 7420 20198
rect 7576 19514 7604 22200
rect 8128 20534 8156 22200
rect 8116 20528 8168 20534
rect 8116 20470 8168 20476
rect 7932 20460 7984 20466
rect 7932 20402 7984 20408
rect 7840 20392 7892 20398
rect 7840 20334 7892 20340
rect 7656 20256 7708 20262
rect 7656 20198 7708 20204
rect 7668 19514 7696 20198
rect 7748 20052 7800 20058
rect 7748 19994 7800 20000
rect 7564 19508 7616 19514
rect 7564 19450 7616 19456
rect 7656 19508 7708 19514
rect 7656 19450 7708 19456
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7380 17740 7432 17746
rect 7380 17682 7432 17688
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7484 17270 7512 17478
rect 7472 17264 7524 17270
rect 7472 17206 7524 17212
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7576 17066 7604 19110
rect 7760 18850 7788 19994
rect 7852 18970 7880 20334
rect 7944 19990 7972 20402
rect 7932 19984 7984 19990
rect 7932 19926 7984 19932
rect 8128 18970 8156 20470
rect 8208 20392 8260 20398
rect 8312 20380 8340 22222
rect 8588 22114 8616 22222
rect 8666 22200 8722 23000
rect 9218 22200 9274 23000
rect 9770 22200 9826 23000
rect 10322 22200 10378 23000
rect 10874 22200 10930 23000
rect 11426 22200 11482 23000
rect 12070 22200 12126 23000
rect 12176 22222 12388 22250
rect 8680 22114 8708 22200
rect 8588 22086 8708 22114
rect 9232 20466 9260 22200
rect 9784 20466 9812 22200
rect 10336 20466 10364 22200
rect 10888 20466 10916 22200
rect 11440 20890 11468 22200
rect 12084 22114 12112 22200
rect 12176 22114 12204 22222
rect 12084 22086 12204 22114
rect 11256 20862 11468 20890
rect 11256 20466 11284 20862
rect 11346 20700 11654 20720
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20624 11654 20644
rect 9220 20460 9272 20466
rect 9220 20402 9272 20408
rect 9772 20460 9824 20466
rect 10324 20460 10376 20466
rect 9824 20420 9904 20448
rect 9772 20402 9824 20408
rect 8260 20352 8340 20380
rect 8208 20334 8260 20340
rect 8208 20256 8260 20262
rect 8208 20198 8260 20204
rect 8392 20256 8444 20262
rect 8392 20198 8444 20204
rect 7840 18964 7892 18970
rect 7840 18906 7892 18912
rect 8116 18964 8168 18970
rect 8116 18906 8168 18912
rect 7760 18822 7880 18850
rect 7748 17740 7800 17746
rect 7748 17682 7800 17688
rect 7564 17060 7616 17066
rect 7564 17002 7616 17008
rect 5920 16546 6040 16574
rect 5724 15700 5776 15706
rect 5724 15642 5776 15648
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 4264 15162 4292 15302
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 5460 15094 5488 15302
rect 5448 15088 5500 15094
rect 5448 15030 5500 15036
rect 4436 14884 4488 14890
rect 4436 14826 4488 14832
rect 4448 14414 4476 14826
rect 5264 14816 5316 14822
rect 5264 14758 5316 14764
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 5080 14408 5132 14414
rect 5080 14350 5132 14356
rect 4448 14074 4476 14350
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 5092 13938 5120 14350
rect 5276 14278 5304 14758
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5920 13734 5948 16546
rect 6828 16448 6880 16454
rect 6828 16390 6880 16396
rect 6148 16348 6456 16368
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16272 6456 16292
rect 6840 16182 6868 16390
rect 6828 16176 6880 16182
rect 6828 16118 6880 16124
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 6932 15570 6960 16050
rect 7012 16040 7064 16046
rect 7012 15982 7064 15988
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 6920 15564 6972 15570
rect 6920 15506 6972 15512
rect 6148 15260 6456 15280
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15184 6456 15204
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 6012 12986 6040 14282
rect 6148 14172 6456 14192
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14096 6456 14116
rect 6656 14074 6684 14962
rect 7024 14618 7052 15982
rect 7104 15972 7156 15978
rect 7104 15914 7156 15920
rect 7012 14612 7064 14618
rect 7012 14554 7064 14560
rect 7116 14550 7144 15914
rect 7300 14822 7328 15982
rect 7760 15502 7788 17682
rect 7852 17354 7880 18822
rect 8024 17604 8076 17610
rect 8024 17546 8076 17552
rect 8036 17490 8064 17546
rect 8036 17462 8156 17490
rect 7852 17326 8064 17354
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7852 16640 7880 17138
rect 7852 16612 7972 16640
rect 7944 15638 7972 16612
rect 7932 15632 7984 15638
rect 7932 15574 7984 15580
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7760 15162 7788 15438
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7104 14544 7156 14550
rect 7104 14486 7156 14492
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 7116 13938 7144 14486
rect 7300 14414 7328 14758
rect 7288 14408 7340 14414
rect 7288 14350 7340 14356
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7300 13870 7328 14350
rect 7484 14006 7512 14758
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7472 14000 7524 14006
rect 7472 13942 7524 13948
rect 7288 13864 7340 13870
rect 7288 13806 7340 13812
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 6148 13084 6456 13104
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13008 6456 13028
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 7024 12850 7052 13466
rect 7300 13326 7328 13806
rect 7576 13530 7604 14418
rect 7564 13524 7616 13530
rect 7564 13466 7616 13472
rect 7288 13320 7340 13326
rect 7288 13262 7340 13268
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7300 12238 7328 13262
rect 8036 12306 8064 17326
rect 8128 15706 8156 17462
rect 8116 15700 8168 15706
rect 8116 15642 8168 15648
rect 8220 14414 8248 20198
rect 8404 18290 8432 20198
rect 8747 20156 9055 20176
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20080 9055 20100
rect 9128 19848 9180 19854
rect 9128 19790 9180 19796
rect 9036 19712 9088 19718
rect 9036 19654 9088 19660
rect 9048 19514 9076 19654
rect 9036 19508 9088 19514
rect 9036 19450 9088 19456
rect 8747 19068 9055 19088
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 18992 9055 19012
rect 8392 18284 8444 18290
rect 8392 18226 8444 18232
rect 8747 17980 9055 18000
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17904 9055 17924
rect 8668 16992 8720 16998
rect 8668 16934 8720 16940
rect 8680 16590 8708 16934
rect 8747 16892 9055 16912
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16816 9055 16836
rect 8668 16584 8720 16590
rect 8668 16526 8720 16532
rect 8747 15804 9055 15824
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15728 9055 15748
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8680 14482 8708 14962
rect 8747 14716 9055 14736
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14640 9055 14660
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8208 14408 8260 14414
rect 8208 14350 8260 14356
rect 8680 14074 8708 14418
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8668 13932 8720 13938
rect 8668 13874 8720 13880
rect 8680 13394 8708 13874
rect 8747 13628 9055 13648
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13552 9055 13572
rect 9140 13394 9168 19790
rect 9232 18970 9260 20402
rect 9680 20256 9732 20262
rect 9680 20198 9732 20204
rect 9692 19514 9720 20198
rect 9680 19508 9732 19514
rect 9680 19450 9732 19456
rect 9312 19372 9364 19378
rect 9312 19314 9364 19320
rect 9220 18964 9272 18970
rect 9220 18906 9272 18912
rect 9324 18630 9352 19314
rect 9680 19236 9732 19242
rect 9680 19178 9732 19184
rect 9772 19236 9824 19242
rect 9772 19178 9824 19184
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9232 16658 9260 17138
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9232 16250 9260 16594
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 9324 14006 9352 18566
rect 9692 18426 9720 19178
rect 9784 18698 9812 19178
rect 9876 19174 9904 20420
rect 10324 20402 10376 20408
rect 10876 20460 10928 20466
rect 10876 20402 10928 20408
rect 11244 20460 11296 20466
rect 11244 20402 11296 20408
rect 12072 20460 12124 20466
rect 12072 20402 12124 20408
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 9864 19168 9916 19174
rect 9864 19110 9916 19116
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9864 18692 9916 18698
rect 9864 18634 9916 18640
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9876 18358 9904 18634
rect 9864 18352 9916 18358
rect 9864 18294 9916 18300
rect 9968 18290 9996 19314
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 10060 18426 10088 19110
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 9956 18284 10008 18290
rect 9956 18226 10008 18232
rect 9772 17128 9824 17134
rect 9772 17070 9824 17076
rect 9784 16522 9812 17070
rect 9864 16992 9916 16998
rect 9864 16934 9916 16940
rect 9772 16516 9824 16522
rect 9772 16458 9824 16464
rect 9876 16114 9904 16934
rect 9968 16658 9996 18226
rect 10336 17882 10364 20402
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 10600 19848 10652 19854
rect 10600 19790 10652 19796
rect 10612 18766 10640 19790
rect 10968 19712 11020 19718
rect 10968 19654 11020 19660
rect 10980 18873 11008 19654
rect 10966 18864 11022 18873
rect 10966 18799 11022 18808
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 9956 16652 10008 16658
rect 9956 16594 10008 16600
rect 9864 16108 9916 16114
rect 9864 16050 9916 16056
rect 9680 15020 9732 15026
rect 9680 14962 9732 14968
rect 9692 14618 9720 14962
rect 9680 14612 9732 14618
rect 9680 14554 9732 14560
rect 10060 14362 10088 17478
rect 10612 16658 10640 18702
rect 11072 18698 11100 20198
rect 11256 20058 11284 20402
rect 11704 20256 11756 20262
rect 11704 20198 11756 20204
rect 11980 20256 12032 20262
rect 11980 20198 12032 20204
rect 11244 20052 11296 20058
rect 11244 19994 11296 20000
rect 11346 19612 11654 19632
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19536 11654 19556
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 10876 18624 10928 18630
rect 10876 18566 10928 18572
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 10888 18222 10916 18566
rect 11164 18426 11192 18566
rect 11346 18524 11654 18544
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18448 11654 18468
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 10876 18216 10928 18222
rect 10876 18158 10928 18164
rect 11244 17740 11296 17746
rect 11244 17682 11296 17688
rect 10232 16652 10284 16658
rect 10232 16594 10284 16600
rect 10600 16652 10652 16658
rect 10600 16594 10652 16600
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9968 14334 10088 14362
rect 9312 14000 9364 14006
rect 9312 13942 9364 13948
rect 9692 13530 9720 14282
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9784 14074 9812 14214
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 9128 13388 9180 13394
rect 9128 13330 9180 13336
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9600 12646 9628 13126
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 8747 12540 9055 12560
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12464 9055 12484
rect 9600 12442 9628 12582
rect 9968 12458 9996 14334
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 13938 10088 14214
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9968 12442 10088 12458
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9968 12436 10100 12442
rect 9968 12430 10048 12436
rect 7932 12300 7984 12306
rect 7932 12242 7984 12248
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 7288 12232 7340 12238
rect 7288 12174 7340 12180
rect 6148 11996 6456 12016
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11920 6456 11940
rect 7944 11218 7972 12242
rect 8312 12170 8340 12378
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 9496 12232 9548 12238
rect 9496 12174 9548 12180
rect 8300 12164 8352 12170
rect 8300 12106 8352 12112
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 8404 11150 8432 12174
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8680 11898 8708 12038
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 9508 11694 9536 12174
rect 9968 11830 9996 12430
rect 10048 12378 10100 12384
rect 10244 11898 10272 16594
rect 10416 16448 10468 16454
rect 10416 16390 10468 16396
rect 10428 15434 10456 16390
rect 10612 16182 10640 16594
rect 11152 16516 11204 16522
rect 11152 16458 11204 16464
rect 10600 16176 10652 16182
rect 10600 16118 10652 16124
rect 11164 15706 11192 16458
rect 11256 15978 11284 17682
rect 11346 17436 11654 17456
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17360 11654 17380
rect 11346 16348 11654 16368
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16272 11654 16292
rect 11244 15972 11296 15978
rect 11244 15914 11296 15920
rect 11152 15700 11204 15706
rect 11152 15642 11204 15648
rect 11256 15502 11284 15914
rect 11244 15496 11296 15502
rect 11244 15438 11296 15444
rect 10324 15428 10376 15434
rect 10324 15370 10376 15376
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 10336 13394 10364 15370
rect 11346 15260 11654 15280
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15184 11654 15204
rect 11346 14172 11654 14192
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14096 11654 14116
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11624 13462 11652 13670
rect 11612 13456 11664 13462
rect 11612 13398 11664 13404
rect 10324 13388 10376 13394
rect 10324 13330 10376 13336
rect 10336 12918 10364 13330
rect 11346 13084 11654 13104
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13008 11654 13028
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 10232 11892 10284 11898
rect 10232 11834 10284 11840
rect 9956 11824 10008 11830
rect 10008 11772 10088 11778
rect 9956 11766 10088 11772
rect 9968 11750 10088 11766
rect 9496 11688 9548 11694
rect 9496 11630 9548 11636
rect 9956 11688 10008 11694
rect 9956 11630 10008 11636
rect 9508 11506 9536 11630
rect 9508 11478 9628 11506
rect 8747 11452 9055 11472
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11376 9055 11396
rect 9600 11354 9628 11478
rect 9588 11348 9640 11354
rect 9588 11290 9640 11296
rect 9968 11150 9996 11630
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 9956 11144 10008 11150
rect 9956 11086 10008 11092
rect 6148 10908 6456 10928
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10832 6456 10852
rect 8404 10470 8432 11086
rect 9968 10538 9996 11086
rect 10060 10810 10088 11750
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10336 10742 10364 12854
rect 11716 12345 11744 20198
rect 11992 19378 12020 20198
rect 12084 20058 12112 20402
rect 12072 20052 12124 20058
rect 12360 20040 12388 22222
rect 12622 22200 12678 23000
rect 13174 22200 13230 23000
rect 13726 22200 13782 23000
rect 14278 22200 14334 23000
rect 14830 22200 14886 23000
rect 15382 22200 15438 23000
rect 15488 22222 15792 22250
rect 12636 20602 12664 22200
rect 13188 20602 13216 22200
rect 12624 20596 12676 20602
rect 12624 20538 12676 20544
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 12900 20528 12952 20534
rect 12900 20470 12952 20476
rect 12440 20052 12492 20058
rect 12360 20012 12440 20040
rect 12072 19994 12124 20000
rect 12440 19994 12492 20000
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 12084 18834 12112 19994
rect 12912 19922 12940 20470
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 12900 19916 12952 19922
rect 12900 19858 12952 19864
rect 12256 19848 12308 19854
rect 12256 19790 12308 19796
rect 13084 19848 13136 19854
rect 13084 19790 13136 19796
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12176 18426 12204 19722
rect 12164 18420 12216 18426
rect 12164 18362 12216 18368
rect 12072 14340 12124 14346
rect 12072 14282 12124 14288
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11808 13326 11836 13670
rect 11796 13320 11848 13326
rect 11796 13262 11848 13268
rect 12084 12986 12112 14282
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11796 12844 11848 12850
rect 11796 12786 11848 12792
rect 11702 12336 11758 12345
rect 11702 12271 11758 12280
rect 11612 12232 11664 12238
rect 11664 12192 11744 12220
rect 11612 12174 11664 12180
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 10876 12096 10928 12102
rect 10876 12038 10928 12044
rect 10796 11830 10824 12038
rect 10888 11898 10916 12038
rect 11164 11898 11192 12106
rect 11346 11996 11654 12016
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11920 11654 11940
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 11152 11892 11204 11898
rect 11152 11834 11204 11840
rect 10784 11824 10836 11830
rect 10784 11766 10836 11772
rect 11336 11756 11388 11762
rect 11336 11698 11388 11704
rect 11348 11354 11376 11698
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 11244 11144 11296 11150
rect 11244 11086 11296 11092
rect 11256 10810 11284 11086
rect 11346 10908 11654 10928
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10832 11654 10852
rect 11244 10804 11296 10810
rect 11244 10746 11296 10752
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 9956 10532 10008 10538
rect 9956 10474 10008 10480
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 6148 9820 6456 9840
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9744 6456 9764
rect 6148 8732 6456 8752
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8656 6456 8676
rect 8404 7886 8432 10406
rect 8747 10364 9055 10384
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10288 9055 10308
rect 9968 10266 9996 10474
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 11716 10130 11744 12192
rect 11808 11898 11836 12786
rect 11796 11892 11848 11898
rect 11796 11834 11848 11840
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11808 11354 11836 11630
rect 11796 11348 11848 11354
rect 11796 11290 11848 11296
rect 11980 11280 12032 11286
rect 11980 11222 12032 11228
rect 11992 10674 12020 11222
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11346 9820 11654 9840
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9744 11654 9764
rect 11900 9722 11928 9930
rect 11888 9716 11940 9722
rect 11888 9658 11940 9664
rect 8747 9276 9055 9296
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9200 9055 9220
rect 12268 9178 12296 19790
rect 13096 19514 13124 19790
rect 13084 19508 13136 19514
rect 13084 19450 13136 19456
rect 13096 18834 13124 19450
rect 13084 18828 13136 18834
rect 13084 18770 13136 18776
rect 12808 18692 12860 18698
rect 12808 18634 12860 18640
rect 12820 18086 12848 18634
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12820 17542 12848 18022
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12808 17536 12860 17542
rect 12808 17478 12860 17484
rect 12452 17270 12480 17478
rect 12440 17264 12492 17270
rect 12440 17206 12492 17212
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12452 16454 12480 17070
rect 12716 16516 12768 16522
rect 12716 16458 12768 16464
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 16114 12480 16390
rect 12728 16250 12756 16458
rect 12716 16244 12768 16250
rect 12716 16186 12768 16192
rect 12440 16108 12492 16114
rect 12440 16050 12492 16056
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12360 11898 12388 13806
rect 12452 13190 12480 14554
rect 12544 14346 12572 14894
rect 12532 14340 12584 14346
rect 12532 14282 12584 14288
rect 12728 13530 12756 14894
rect 12820 13938 12848 17478
rect 13084 15020 13136 15026
rect 13084 14962 13136 14968
rect 13096 14074 13124 14962
rect 13176 14816 13228 14822
rect 13176 14758 13228 14764
rect 13268 14816 13320 14822
rect 13268 14758 13320 14764
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 13188 14006 13216 14758
rect 13280 14278 13308 14758
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 13176 14000 13228 14006
rect 13176 13942 13228 13948
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 12900 13796 12952 13802
rect 12900 13738 12952 13744
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12912 13394 12940 13738
rect 12900 13388 12952 13394
rect 12900 13330 12952 13336
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12912 12850 12940 13330
rect 12900 12844 12952 12850
rect 12900 12786 12952 12792
rect 12912 12442 12940 12786
rect 12900 12436 12952 12442
rect 12900 12378 12952 12384
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12360 10810 12388 11834
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13188 11218 13216 11494
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 12348 10804 12400 10810
rect 12348 10746 12400 10752
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12440 10056 12492 10062
rect 12440 9998 12492 10004
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 11152 8968 11204 8974
rect 11152 8910 11204 8916
rect 11164 8634 11192 8910
rect 11346 8732 11654 8752
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8656 11654 8676
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 11244 8492 11296 8498
rect 11244 8434 11296 8440
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 8747 8188 9055 8208
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8112 9055 8132
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 6148 7644 6456 7664
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7568 6456 7588
rect 8404 7478 8432 7822
rect 9416 7546 9444 8434
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 10060 7886 10088 8230
rect 10048 7880 10100 7886
rect 10048 7822 10100 7828
rect 11256 7546 11284 8434
rect 11532 7818 11560 8434
rect 12164 8288 12216 8294
rect 12164 8230 12216 8236
rect 12176 7818 12204 8230
rect 12452 7886 12480 9998
rect 12544 9926 12572 10542
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12544 9586 12572 9862
rect 13372 9654 13400 13874
rect 13360 9648 13412 9654
rect 13360 9590 13412 9596
rect 12532 9580 12584 9586
rect 12532 9522 12584 9528
rect 13464 9178 13492 20402
rect 13740 20040 13768 22200
rect 14292 20602 14320 22200
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 13832 20262 13860 20470
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14648 20392 14700 20398
rect 14648 20334 14700 20340
rect 13820 20256 13872 20262
rect 13820 20198 13872 20204
rect 13945 20156 14253 20176
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20080 14253 20100
rect 13820 20052 13872 20058
rect 13740 20012 13820 20040
rect 13820 19994 13872 20000
rect 13636 19712 13688 19718
rect 13636 19654 13688 19660
rect 13648 19378 13676 19654
rect 13820 19508 13872 19514
rect 13820 19450 13872 19456
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13832 18970 13860 19450
rect 13945 19068 14253 19088
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 18992 14253 19012
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13945 17980 14253 18000
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17904 14253 17924
rect 14292 17762 14320 20334
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14568 18630 14596 19790
rect 14660 19378 14688 20334
rect 14844 20262 14872 22200
rect 15396 22114 15424 22200
rect 15488 22114 15516 22222
rect 15396 22086 15516 22114
rect 15764 20602 15792 22222
rect 15934 22200 15990 23000
rect 16486 22200 16542 23000
rect 17038 22200 17094 23000
rect 17682 22200 17738 23000
rect 18234 22200 18290 23000
rect 18786 22200 18842 23000
rect 18878 22672 18934 22681
rect 18878 22607 18934 22616
rect 15948 20618 15976 22200
rect 16500 20890 16528 22200
rect 16408 20862 16528 20890
rect 15752 20596 15804 20602
rect 15948 20590 16068 20618
rect 15752 20538 15804 20544
rect 16040 20534 16068 20590
rect 16028 20528 16080 20534
rect 16028 20470 16080 20476
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 16304 20460 16356 20466
rect 16304 20402 16356 20408
rect 14740 20256 14792 20262
rect 14740 20198 14792 20204
rect 14832 20256 14884 20262
rect 14832 20198 14884 20204
rect 14752 20074 14780 20198
rect 14752 20046 14872 20074
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14752 19446 14780 19790
rect 14740 19440 14792 19446
rect 14740 19382 14792 19388
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14556 18624 14608 18630
rect 14556 18566 14608 18572
rect 14200 17734 14320 17762
rect 14094 17640 14150 17649
rect 14094 17575 14150 17584
rect 14108 17338 14136 17575
rect 14096 17332 14148 17338
rect 14096 17274 14148 17280
rect 14200 17270 14228 17734
rect 14188 17264 14240 17270
rect 14188 17206 14240 17212
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13832 16454 13860 17070
rect 13945 16892 14253 16912
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16816 14253 16836
rect 14372 16516 14424 16522
rect 14372 16458 14424 16464
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 13832 16114 13860 16390
rect 14384 16250 14412 16458
rect 14372 16244 14424 16250
rect 14372 16186 14424 16192
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13945 15804 14253 15824
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15728 14253 15748
rect 13945 14716 14253 14736
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14640 14253 14660
rect 14372 13864 14424 13870
rect 14372 13806 14424 13812
rect 13945 13628 14253 13648
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13552 14253 13572
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13556 11082 13584 13126
rect 13945 12540 14253 12560
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12464 14253 12484
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 13945 11452 14253 11472
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11376 14253 11396
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13832 9994 13860 11154
rect 14292 10470 14320 11494
rect 14280 10464 14332 10470
rect 14280 10406 14332 10412
rect 13945 10364 14253 10384
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10288 14253 10308
rect 14292 10266 14320 10406
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13832 9518 13860 9930
rect 14384 9518 14412 13806
rect 14476 11354 14504 17138
rect 14568 12434 14596 18566
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14752 17542 14780 18022
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14752 17202 14780 17478
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14844 17082 14872 20046
rect 14936 18086 14964 20402
rect 15568 19780 15620 19786
rect 15568 19722 15620 19728
rect 15200 19712 15252 19718
rect 15200 19654 15252 19660
rect 15212 18766 15240 19654
rect 15580 19378 15608 19722
rect 15660 19440 15712 19446
rect 15660 19382 15712 19388
rect 15568 19372 15620 19378
rect 15568 19314 15620 19320
rect 15672 18834 15700 19382
rect 15660 18828 15712 18834
rect 15660 18770 15712 18776
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15672 18222 15700 18770
rect 15660 18216 15712 18222
rect 15660 18158 15712 18164
rect 14924 18080 14976 18086
rect 14924 18022 14976 18028
rect 14752 17054 14872 17082
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15384 17060 15436 17066
rect 14568 12406 14688 12434
rect 14556 12096 14608 12102
rect 14556 12038 14608 12044
rect 14568 11898 14596 12038
rect 14556 11892 14608 11898
rect 14556 11834 14608 11840
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14476 11218 14504 11290
rect 14464 11212 14516 11218
rect 14464 11154 14516 11160
rect 14556 11144 14608 11150
rect 14556 11086 14608 11092
rect 14464 11076 14516 11082
rect 14464 11018 14516 11024
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 14476 9450 14504 11018
rect 14568 9926 14596 11086
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 13945 9276 14253 9296
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9200 14253 9220
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13464 8634 13492 8910
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12440 7880 12492 7886
rect 12440 7822 12492 7828
rect 11520 7812 11572 7818
rect 11520 7754 11572 7760
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 11346 7644 11654 7664
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7568 11654 7588
rect 9404 7540 9456 7546
rect 9404 7482 9456 7488
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8300 7404 8352 7410
rect 8300 7346 8352 7352
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 6148 6556 6456 6576
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6480 6456 6500
rect 8312 6458 8340 7346
rect 8747 7100 9055 7120
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7024 9055 7044
rect 9416 6866 9444 7482
rect 12084 7342 12112 7686
rect 12544 7546 12572 8366
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13176 7744 13228 7750
rect 13176 7686 13228 7692
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 13188 7478 13216 7686
rect 13740 7546 13768 7754
rect 13832 7546 13860 8434
rect 14464 8424 14516 8430
rect 14464 8366 14516 8372
rect 13945 8188 14253 8208
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8112 14253 8132
rect 14476 7546 14504 8366
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 13176 7472 13228 7478
rect 13176 7414 13228 7420
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 12072 7336 12124 7342
rect 12072 7278 12124 7284
rect 11992 7002 12020 7278
rect 13945 7100 14253 7120
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7024 14253 7044
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 11346 6556 11654 6576
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6480 11654 6500
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 1400 6316 1452 6322
rect 1400 6258 1452 6264
rect 1412 5817 1440 6258
rect 14660 6186 14688 12406
rect 14648 6180 14700 6186
rect 14648 6122 14700 6128
rect 3549 6012 3857 6032
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5936 3857 5956
rect 8747 6012 9055 6032
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5936 9055 5956
rect 13945 6012 14253 6032
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5936 14253 5956
rect 14752 5846 14780 17054
rect 15384 17002 15436 17008
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 14844 16114 14872 16730
rect 15396 16658 15424 17002
rect 15488 16726 15516 17070
rect 15672 16794 15700 18158
rect 15660 16788 15712 16794
rect 15660 16730 15712 16736
rect 15476 16720 15528 16726
rect 15476 16662 15528 16668
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14844 14414 14872 16050
rect 15488 15502 15516 16662
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15108 15020 15160 15026
rect 15108 14962 15160 14968
rect 15120 14618 15148 14962
rect 15108 14612 15160 14618
rect 15108 14554 15160 14560
rect 15120 14498 15148 14554
rect 14936 14470 15148 14498
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14844 12918 14872 14350
rect 14936 13870 14964 14470
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 15120 14074 15148 14282
rect 15108 14068 15160 14074
rect 15108 14010 15160 14016
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 15028 10810 15056 12174
rect 15476 12096 15528 12102
rect 15476 12038 15528 12044
rect 15488 11762 15516 12038
rect 15292 11756 15344 11762
rect 15292 11698 15344 11704
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15304 11558 15332 11698
rect 15292 11552 15344 11558
rect 15292 11494 15344 11500
rect 15476 11280 15528 11286
rect 15476 11222 15528 11228
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14844 8838 14872 9454
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14740 5840 14792 5846
rect 1398 5808 1454 5817
rect 14740 5782 14792 5788
rect 1398 5743 1454 5752
rect 6148 5468 6456 5488
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5392 6456 5412
rect 11346 5468 11654 5488
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5392 11654 5412
rect 3549 4924 3857 4944
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4848 3857 4868
rect 8747 4924 9055 4944
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4848 9055 4868
rect 13945 4924 14253 4944
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4848 14253 4868
rect 6148 4380 6456 4400
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4304 6456 4324
rect 11346 4380 11654 4400
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4304 11654 4324
rect 3549 3836 3857 3856
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3760 3857 3780
rect 8747 3836 9055 3856
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3760 9055 3780
rect 13945 3836 14253 3856
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3760 14253 3780
rect 6148 3292 6456 3312
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3216 6456 3236
rect 11346 3292 11654 3312
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3216 11654 3236
rect 3549 2748 3857 2768
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2672 3857 2692
rect 8747 2748 9055 2768
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2672 9055 2692
rect 13945 2748 14253 2768
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2672 14253 2692
rect 14844 2446 14872 8774
rect 15212 2922 15240 11018
rect 15488 10810 15516 11222
rect 15476 10804 15528 10810
rect 15476 10746 15528 10752
rect 15752 10668 15804 10674
rect 15752 10610 15804 10616
rect 15764 10266 15792 10610
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15948 9450 15976 20402
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16132 15706 16160 16050
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 16120 14952 16172 14958
rect 16120 14894 16172 14900
rect 16132 14414 16160 14894
rect 16120 14408 16172 14414
rect 16120 14350 16172 14356
rect 16028 14340 16080 14346
rect 16028 14282 16080 14288
rect 16040 14074 16068 14282
rect 16028 14068 16080 14074
rect 16028 14010 16080 14016
rect 16316 12434 16344 20402
rect 16408 20244 16436 20862
rect 16544 20700 16852 20720
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20624 16852 20644
rect 17052 20330 17080 22200
rect 17696 20602 17724 22200
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 17500 20460 17552 20466
rect 17500 20402 17552 20408
rect 16856 20324 16908 20330
rect 16856 20266 16908 20272
rect 17040 20324 17092 20330
rect 17040 20266 17092 20272
rect 16580 20256 16632 20262
rect 16408 20216 16580 20244
rect 16580 20198 16632 20204
rect 16868 19922 16896 20266
rect 16856 19916 16908 19922
rect 16856 19858 16908 19864
rect 17316 19916 17368 19922
rect 17316 19858 17368 19864
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16408 17678 16436 19790
rect 16544 19612 16852 19632
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19536 16852 19556
rect 17328 19378 17356 19858
rect 17316 19372 17368 19378
rect 17316 19314 17368 19320
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16684 18766 16712 19110
rect 16672 18760 16724 18766
rect 16672 18702 16724 18708
rect 17408 18760 17460 18766
rect 17408 18702 17460 18708
rect 16948 18624 17000 18630
rect 16948 18566 17000 18572
rect 16544 18524 16852 18544
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18448 16852 18468
rect 16960 17746 16988 18566
rect 17420 18426 17448 18702
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 16948 17740 17000 17746
rect 16948 17682 17000 17688
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16948 17536 17000 17542
rect 16948 17478 17000 17484
rect 16544 17436 16852 17456
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17360 16852 17380
rect 16672 17196 16724 17202
rect 16672 17138 16724 17144
rect 16396 16788 16448 16794
rect 16396 16730 16448 16736
rect 16408 16130 16436 16730
rect 16684 16658 16712 17138
rect 16672 16652 16724 16658
rect 16672 16594 16724 16600
rect 16960 16454 16988 17478
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17040 16652 17092 16658
rect 17040 16594 17092 16600
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16544 16348 16852 16368
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16272 16852 16292
rect 16408 16114 16620 16130
rect 16408 16108 16632 16114
rect 16408 16102 16580 16108
rect 16580 16050 16632 16056
rect 16592 15570 16620 16050
rect 16960 15994 16988 16390
rect 17052 16250 17080 16594
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 17328 16182 17356 16934
rect 17316 16176 17368 16182
rect 17316 16118 17368 16124
rect 16960 15966 17080 15994
rect 16580 15564 16632 15570
rect 16580 15506 16632 15512
rect 16544 15260 16852 15280
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15184 16852 15204
rect 17052 14278 17080 15966
rect 17316 15564 17368 15570
rect 17316 15506 17368 15512
rect 17040 14272 17092 14278
rect 17040 14214 17092 14220
rect 16544 14172 16852 14192
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14096 16852 14116
rect 16544 13084 16852 13104
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13008 16852 13028
rect 16580 12912 16632 12918
rect 16580 12854 16632 12860
rect 16592 12646 16620 12854
rect 16580 12640 16632 12646
rect 16580 12582 16632 12588
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16316 12406 16436 12434
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16040 11694 16068 12174
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16132 9722 16160 9862
rect 16120 9716 16172 9722
rect 16120 9658 16172 9664
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 16316 9178 16344 9522
rect 16304 9172 16356 9178
rect 16304 9114 16356 9120
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15304 7750 15332 8434
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16132 7818 16160 8230
rect 16120 7812 16172 7818
rect 16120 7754 16172 7760
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15304 7342 15332 7686
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15488 6798 15516 7482
rect 16408 6866 16436 12406
rect 16578 12336 16634 12345
rect 16578 12271 16634 12280
rect 16592 12238 16620 12271
rect 16580 12232 16632 12238
rect 16580 12174 16632 12180
rect 16544 11996 16852 12016
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11920 16852 11940
rect 16960 11898 16988 12582
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 17052 11234 17080 14214
rect 17328 13938 17356 15506
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17408 13456 17460 13462
rect 17408 13398 17460 13404
rect 17420 13190 17448 13398
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17316 12844 17368 12850
rect 17316 12786 17368 12792
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 17224 12776 17276 12782
rect 17224 12718 17276 12724
rect 17144 12442 17172 12718
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 17236 12186 17264 12718
rect 17328 12442 17356 12786
rect 17316 12436 17368 12442
rect 17316 12378 17368 12384
rect 17144 12170 17264 12186
rect 17132 12164 17264 12170
rect 17184 12158 17264 12164
rect 17132 12106 17184 12112
rect 17144 11694 17172 12106
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 16960 11206 17080 11234
rect 16544 10908 16852 10928
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10832 16852 10852
rect 16960 9926 16988 11206
rect 17040 11076 17092 11082
rect 17040 11018 17092 11024
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16544 9820 16852 9840
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9744 16852 9764
rect 16948 8968 17000 8974
rect 16948 8910 17000 8916
rect 16544 8732 16852 8752
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8656 16852 8676
rect 16544 7644 16852 7664
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7568 16852 7588
rect 16960 7546 16988 8910
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16396 6860 16448 6866
rect 16396 6802 16448 6808
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 16544 6556 16852 6576
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6480 16852 6500
rect 16544 5468 16852 5488
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5392 16852 5412
rect 16544 4380 16852 4400
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4304 16852 4324
rect 16544 3292 16852 3312
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3216 16852 3236
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 17052 2582 17080 11018
rect 17144 10810 17172 11630
rect 17132 10804 17184 10810
rect 17132 10746 17184 10752
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17144 7750 17172 8434
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17144 7478 17172 7686
rect 17132 7472 17184 7478
rect 17132 7414 17184 7420
rect 17236 3602 17264 9862
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17328 7546 17356 8774
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17512 6662 17540 20402
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17604 17082 17632 20334
rect 18248 20262 18276 22200
rect 18694 22128 18750 22137
rect 18694 22063 18750 22072
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18512 20392 18564 20398
rect 18512 20334 18564 20340
rect 18236 20256 18288 20262
rect 18236 20198 18288 20204
rect 18052 19780 18104 19786
rect 18052 19722 18104 19728
rect 18420 19780 18472 19786
rect 18420 19722 18472 19728
rect 17868 19168 17920 19174
rect 17868 19110 17920 19116
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17684 18080 17736 18086
rect 17684 18022 17736 18028
rect 17696 17746 17724 18022
rect 17684 17740 17736 17746
rect 17684 17682 17736 17688
rect 17788 17678 17816 18906
rect 17776 17672 17828 17678
rect 17776 17614 17828 17620
rect 17880 17270 17908 19110
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 18358 18000 18566
rect 17960 18352 18012 18358
rect 17960 18294 18012 18300
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17604 17054 17908 17082
rect 17776 16992 17828 16998
rect 17776 16934 17828 16940
rect 17788 15502 17816 16934
rect 17776 15496 17828 15502
rect 17776 15438 17828 15444
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17696 12918 17724 13194
rect 17684 12912 17736 12918
rect 17684 12854 17736 12860
rect 17696 12238 17724 12854
rect 17776 12300 17828 12306
rect 17776 12242 17828 12248
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17696 11082 17724 12174
rect 17788 11830 17816 12242
rect 17776 11824 17828 11830
rect 17776 11766 17828 11772
rect 17684 11076 17736 11082
rect 17684 11018 17736 11024
rect 17788 10742 17816 11766
rect 17776 10736 17828 10742
rect 17776 10678 17828 10684
rect 17788 10266 17816 10678
rect 17776 10260 17828 10266
rect 17776 10202 17828 10208
rect 17776 8288 17828 8294
rect 17776 8230 17828 8236
rect 17788 7818 17816 8230
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17604 7342 17632 7686
rect 17592 7336 17644 7342
rect 17592 7278 17644 7284
rect 17880 7206 17908 17054
rect 17960 14000 18012 14006
rect 17960 13942 18012 13948
rect 17972 13394 18000 13942
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 18064 13326 18092 19722
rect 18432 19378 18460 19722
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 18326 18864 18382 18873
rect 18326 18799 18382 18808
rect 18340 18766 18368 18799
rect 18328 18760 18380 18766
rect 18328 18702 18380 18708
rect 18420 18624 18472 18630
rect 18420 18566 18472 18572
rect 18328 18420 18380 18426
rect 18328 18362 18380 18368
rect 18340 18329 18368 18362
rect 18326 18320 18382 18329
rect 18326 18255 18382 18264
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18156 16658 18184 17138
rect 18340 16998 18368 17478
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18144 16652 18196 16658
rect 18144 16594 18196 16600
rect 18156 16250 18184 16594
rect 18432 16590 18460 18566
rect 18524 17626 18552 20334
rect 18616 19553 18644 20402
rect 18602 19544 18658 19553
rect 18708 19530 18736 22063
rect 18800 20058 18828 22200
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 18892 19854 18920 22607
rect 19338 22200 19394 23000
rect 19890 22200 19946 23000
rect 20442 22200 20498 23000
rect 20994 22200 21050 23000
rect 21546 22200 21602 23000
rect 22098 22200 22154 23000
rect 22650 22200 22706 23000
rect 19062 21312 19118 21321
rect 19062 21247 19118 21256
rect 18880 19848 18932 19854
rect 18880 19790 18932 19796
rect 18708 19502 18828 19530
rect 18602 19479 18658 19488
rect 18696 19440 18748 19446
rect 18602 19408 18658 19417
rect 18696 19382 18748 19388
rect 18602 19343 18604 19352
rect 18656 19343 18658 19352
rect 18604 19314 18656 19320
rect 18708 18970 18736 19382
rect 18696 18964 18748 18970
rect 18696 18906 18748 18912
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18524 17598 18644 17626
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18616 16402 18644 17598
rect 18708 17338 18736 18226
rect 18800 18154 18828 19502
rect 18892 18426 18920 19790
rect 19076 19378 19104 21247
rect 19352 20244 19380 22200
rect 19614 20904 19670 20913
rect 19614 20839 19670 20848
rect 19352 20216 19564 20244
rect 19143 20156 19451 20176
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20080 19451 20100
rect 19536 20058 19564 20216
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19628 19446 19656 20839
rect 19904 20602 19932 22200
rect 20456 20618 20484 22200
rect 20456 20602 20760 20618
rect 19892 20596 19944 20602
rect 20456 20596 20772 20602
rect 20456 20590 20720 20596
rect 19892 20538 19944 20544
rect 20720 20538 20772 20544
rect 20260 20460 20312 20466
rect 20260 20402 20312 20408
rect 20074 19952 20130 19961
rect 20074 19887 20130 19896
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19616 19440 19668 19446
rect 19616 19382 19668 19388
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 19064 19372 19116 19378
rect 19064 19314 19116 19320
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 18880 18420 18932 18426
rect 18880 18362 18932 18368
rect 18788 18148 18840 18154
rect 18788 18090 18840 18096
rect 18880 18080 18932 18086
rect 18880 18022 18932 18028
rect 18892 17898 18920 18022
rect 18800 17870 18920 17898
rect 18800 17814 18828 17870
rect 18788 17808 18840 17814
rect 18788 17750 18840 17756
rect 18786 17640 18842 17649
rect 18786 17575 18788 17584
rect 18840 17575 18842 17584
rect 18788 17546 18840 17552
rect 18984 17338 19012 19314
rect 19143 19068 19451 19088
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 18992 19451 19012
rect 19064 18216 19116 18222
rect 19064 18158 19116 18164
rect 19076 17882 19104 18158
rect 19143 17980 19451 18000
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17904 19451 17924
rect 19064 17876 19116 17882
rect 19064 17818 19116 17824
rect 19616 17672 19668 17678
rect 19616 17614 19668 17620
rect 19628 17338 19656 17614
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18972 17332 19024 17338
rect 18972 17274 19024 17280
rect 19616 17332 19668 17338
rect 19616 17274 19668 17280
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 19143 16892 19451 16912
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16816 19451 16836
rect 19340 16516 19392 16522
rect 19340 16458 19392 16464
rect 18616 16374 18736 16402
rect 18144 16244 18196 16250
rect 18144 16186 18196 16192
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 18524 13530 18552 13874
rect 18512 13524 18564 13530
rect 18512 13466 18564 13472
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 18420 12776 18472 12782
rect 18420 12718 18472 12724
rect 18432 12374 18460 12718
rect 18604 12640 18656 12646
rect 18604 12582 18656 12588
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18616 12238 18644 12582
rect 17960 12232 18012 12238
rect 17960 12174 18012 12180
rect 18604 12232 18656 12238
rect 18604 12174 18656 12180
rect 17972 12102 18000 12174
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 18052 12096 18104 12102
rect 18052 12038 18104 12044
rect 17972 11762 18000 12038
rect 18064 11898 18092 12038
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17972 3670 18000 11698
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18524 10062 18552 10542
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18052 9920 18104 9926
rect 18052 9862 18104 9868
rect 18064 7342 18092 9862
rect 18524 9518 18552 9998
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18512 9512 18564 9518
rect 18512 9454 18564 9460
rect 18248 8430 18276 9454
rect 18708 8566 18736 16374
rect 19352 16114 19380 16458
rect 19536 16454 19564 17138
rect 19616 17060 19668 17066
rect 19616 17002 19668 17008
rect 19524 16448 19576 16454
rect 19524 16390 19576 16396
rect 19628 16114 19656 17002
rect 19720 16454 19748 19314
rect 19800 17536 19852 17542
rect 19800 17478 19852 17484
rect 19708 16448 19760 16454
rect 19708 16390 19760 16396
rect 19812 16250 19840 17478
rect 19800 16244 19852 16250
rect 19800 16186 19852 16192
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 19143 15804 19451 15824
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15728 19451 15748
rect 18880 15360 18932 15366
rect 18880 15302 18932 15308
rect 18892 14006 18920 15302
rect 19143 14716 19451 14736
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14640 19451 14660
rect 19708 14408 19760 14414
rect 19708 14350 19760 14356
rect 19720 14074 19748 14350
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 18880 14000 18932 14006
rect 18880 13942 18932 13948
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 19076 13530 19104 13942
rect 19143 13628 19451 13648
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13552 19451 13572
rect 19064 13524 19116 13530
rect 19064 13466 19116 13472
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19260 12753 19288 12786
rect 19246 12744 19302 12753
rect 19246 12679 19302 12688
rect 19143 12540 19451 12560
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12464 19451 12484
rect 19064 12096 19116 12102
rect 19064 12038 19116 12044
rect 19340 12096 19392 12102
rect 19340 12038 19392 12044
rect 18880 10668 18932 10674
rect 18880 10610 18932 10616
rect 18892 10577 18920 10610
rect 18878 10568 18934 10577
rect 18878 10503 18934 10512
rect 18696 8560 18748 8566
rect 18696 8502 18748 8508
rect 18236 8424 18288 8430
rect 18236 8366 18288 8372
rect 18248 7886 18276 8366
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 6798 18092 7278
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 19076 3194 19104 12038
rect 19352 11778 19380 12038
rect 19168 11762 19380 11778
rect 19156 11756 19380 11762
rect 19208 11750 19380 11756
rect 19156 11698 19208 11704
rect 19536 11626 19564 12786
rect 19708 12096 19760 12102
rect 19708 12038 19760 12044
rect 19524 11620 19576 11626
rect 19524 11562 19576 11568
rect 19143 11452 19451 11472
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11376 19451 11396
rect 19720 11218 19748 12038
rect 19904 11898 19932 19790
rect 20088 19514 20116 19887
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 19996 18766 20024 19450
rect 20168 19372 20220 19378
rect 20168 19314 20220 19320
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19996 17882 20024 18226
rect 19984 17876 20036 17882
rect 19984 17818 20036 17824
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 20088 17338 20116 17614
rect 20076 17332 20128 17338
rect 20076 17274 20128 17280
rect 20076 16584 20128 16590
rect 20076 16526 20128 16532
rect 20088 16250 20116 16526
rect 20180 16250 20208 19314
rect 20076 16244 20128 16250
rect 20076 16186 20128 16192
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 19984 16108 20036 16114
rect 19984 16050 20036 16056
rect 19996 15706 20024 16050
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 20168 15496 20220 15502
rect 20168 15438 20220 15444
rect 20180 15162 20208 15438
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 19984 13864 20036 13870
rect 19984 13806 20036 13812
rect 19996 13326 20024 13806
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 20088 12866 20116 13262
rect 19996 12838 20116 12866
rect 19996 12714 20024 12838
rect 19984 12708 20036 12714
rect 19984 12650 20036 12656
rect 20272 11898 20300 20402
rect 20534 20360 20590 20369
rect 20534 20295 20590 20304
rect 20352 19848 20404 19854
rect 20352 19790 20404 19796
rect 20364 16454 20392 19790
rect 20444 19372 20496 19378
rect 20444 19314 20496 19320
rect 20352 16448 20404 16454
rect 20352 16390 20404 16396
rect 20352 15088 20404 15094
rect 20352 15030 20404 15036
rect 20364 13530 20392 15030
rect 20352 13524 20404 13530
rect 20352 13466 20404 13472
rect 20456 12442 20484 19314
rect 20548 18970 20576 20295
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20732 19417 20760 19654
rect 21008 19514 21036 22200
rect 21454 21720 21510 21729
rect 21454 21655 21510 21664
rect 21088 19848 21140 19854
rect 21088 19790 21140 19796
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 20718 19408 20774 19417
rect 20718 19343 20774 19352
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20628 18148 20680 18154
rect 20628 18090 20680 18096
rect 20640 17241 20668 18090
rect 20718 17640 20774 17649
rect 20718 17575 20774 17584
rect 20732 17542 20760 17575
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20626 17232 20682 17241
rect 20626 17167 20682 17176
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20732 15638 20760 16186
rect 20720 15632 20772 15638
rect 20720 15574 20772 15580
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20640 14618 20668 15438
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20536 14340 20588 14346
rect 20536 14282 20588 14288
rect 20548 12986 20576 14282
rect 20628 13932 20680 13938
rect 20628 13874 20680 13880
rect 20640 13025 20668 13874
rect 20626 13016 20682 13025
rect 20536 12980 20588 12986
rect 20824 12986 20852 18702
rect 20916 17610 20944 19314
rect 20996 18284 21048 18290
rect 20996 18226 21048 18232
rect 20904 17604 20956 17610
rect 20904 17546 20956 17552
rect 21008 17490 21036 18226
rect 20916 17462 21036 17490
rect 20916 16250 20944 17462
rect 21100 17354 21128 19790
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21284 19009 21312 19654
rect 21364 19168 21416 19174
rect 21364 19110 21416 19116
rect 21270 19000 21326 19009
rect 21270 18935 21326 18944
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 21008 17326 21128 17354
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20916 15162 20944 16050
rect 21008 15638 21036 17326
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21100 16794 21128 17138
rect 21192 16998 21220 18702
rect 21272 18624 21324 18630
rect 21376 18601 21404 19110
rect 21272 18566 21324 18572
rect 21362 18592 21418 18601
rect 21284 18057 21312 18566
rect 21362 18527 21418 18536
rect 21468 18426 21496 21655
rect 21560 18970 21588 22200
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21548 18964 21600 18970
rect 21548 18906 21600 18912
rect 21548 18692 21600 18698
rect 21548 18634 21600 18640
rect 21456 18420 21508 18426
rect 21456 18362 21508 18368
rect 21270 18048 21326 18057
rect 21270 17983 21326 17992
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21180 16992 21232 16998
rect 21180 16934 21232 16940
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21284 16697 21312 17478
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21270 16688 21326 16697
rect 21270 16623 21326 16632
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 21100 15706 21128 16526
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21284 15745 21312 16390
rect 21376 16289 21404 16934
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21362 16280 21418 16289
rect 21362 16215 21418 16224
rect 21364 15904 21416 15910
rect 21364 15846 21416 15852
rect 21270 15736 21326 15745
rect 21088 15700 21140 15706
rect 21270 15671 21326 15680
rect 21088 15642 21140 15648
rect 20996 15632 21048 15638
rect 20996 15574 21048 15580
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 21100 14618 21128 15438
rect 21272 15360 21324 15366
rect 21376 15337 21404 15846
rect 21272 15302 21324 15308
rect 21362 15328 21418 15337
rect 21284 14929 21312 15302
rect 21362 15263 21418 15272
rect 21270 14920 21326 14929
rect 21270 14855 21326 14864
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21284 14385 21312 14758
rect 21270 14376 21326 14385
rect 21270 14311 21326 14320
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 21284 13977 21312 14214
rect 21270 13968 21326 13977
rect 21088 13932 21140 13938
rect 21270 13903 21326 13912
rect 21088 13874 21140 13880
rect 20996 13728 21048 13734
rect 20996 13670 21048 13676
rect 21008 13326 21036 13670
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 20626 12951 20682 12960
rect 20812 12980 20864 12986
rect 20536 12922 20588 12928
rect 20812 12922 20864 12928
rect 20720 12708 20772 12714
rect 20720 12650 20772 12656
rect 20444 12436 20496 12442
rect 20444 12378 20496 12384
rect 20732 12238 20760 12650
rect 21100 12442 21128 13874
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21284 13569 21312 13670
rect 21270 13560 21326 13569
rect 21270 13495 21326 13504
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 21088 12436 21140 12442
rect 21088 12378 21140 12384
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 19892 11892 19944 11898
rect 19892 11834 19944 11840
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 21192 11830 21220 13194
rect 21362 13016 21418 13025
rect 21362 12951 21364 12960
rect 21416 12951 21418 12960
rect 21364 12922 21416 12928
rect 21468 12434 21496 16390
rect 21560 13530 21588 18634
rect 21548 13524 21600 13530
rect 21548 13466 21600 13472
rect 21284 12406 21496 12434
rect 21180 11824 21232 11830
rect 21180 11766 21232 11772
rect 19892 11756 19944 11762
rect 19892 11698 19944 11704
rect 20536 11756 20588 11762
rect 20536 11698 20588 11704
rect 20996 11756 21048 11762
rect 20996 11698 21048 11704
rect 19904 11354 19932 11698
rect 20548 11354 20576 11698
rect 19892 11348 19944 11354
rect 19892 11290 19944 11296
rect 20536 11348 20588 11354
rect 20536 11290 20588 11296
rect 20902 11248 20958 11257
rect 19708 11212 19760 11218
rect 20902 11183 20958 11192
rect 19708 11154 19760 11160
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19260 10810 19288 11086
rect 19248 10804 19300 10810
rect 19248 10746 19300 10752
rect 19524 10600 19576 10606
rect 19524 10542 19576 10548
rect 19143 10364 19451 10384
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10288 19451 10308
rect 19536 10266 19564 10542
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 19616 9580 19668 9586
rect 19616 9522 19668 9528
rect 19143 9276 19451 9296
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9200 19451 9220
rect 19628 9178 19656 9522
rect 19616 9172 19668 9178
rect 19616 9114 19668 9120
rect 19616 8968 19668 8974
rect 19616 8910 19668 8916
rect 19628 8634 19656 8910
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19248 8560 19300 8566
rect 19248 8502 19300 8508
rect 19260 8362 19288 8502
rect 19248 8356 19300 8362
rect 19248 8298 19300 8304
rect 19143 8188 19451 8208
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8112 19451 8132
rect 19143 7100 19451 7120
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7024 19451 7044
rect 19143 6012 19451 6032
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5936 19451 5956
rect 19143 4924 19451 4944
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4848 19451 4868
rect 19143 3836 19451 3856
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3760 19451 3780
rect 19064 3188 19116 3194
rect 19064 3130 19116 3136
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 17040 2576 17092 2582
rect 17040 2518 17092 2524
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 6148 2204 6456 2224
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2128 6456 2148
rect 11346 2204 11654 2224
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2128 11654 2148
rect 16544 2204 16852 2224
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2128 16852 2148
rect 19076 1057 19104 2994
rect 19720 2854 19748 11154
rect 20916 11150 20944 11183
rect 20904 11144 20956 11150
rect 20904 11086 20956 11092
rect 20916 10810 20944 11086
rect 21008 10810 21036 11698
rect 21192 11558 21220 11766
rect 21180 11552 21232 11558
rect 21180 11494 21232 11500
rect 20904 10804 20956 10810
rect 20904 10746 20956 10752
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 19984 10600 20036 10606
rect 19984 10542 20036 10548
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 10062 19932 10406
rect 19996 10062 20024 10542
rect 20076 10124 20128 10130
rect 20076 10066 20128 10072
rect 19892 10056 19944 10062
rect 19892 9998 19944 10004
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 19996 9722 20024 9998
rect 19984 9716 20036 9722
rect 19984 9658 20036 9664
rect 20088 8974 20116 10066
rect 20904 9648 20956 9654
rect 20904 9590 20956 9596
rect 20536 9376 20588 9382
rect 20536 9318 20588 9324
rect 20548 8974 20576 9318
rect 20076 8968 20128 8974
rect 20536 8968 20588 8974
rect 20076 8910 20128 8916
rect 20534 8936 20536 8945
rect 20628 8968 20680 8974
rect 20588 8936 20590 8945
rect 20628 8910 20680 8916
rect 20534 8871 20590 8880
rect 20640 8634 20668 8910
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19812 8090 19840 8434
rect 19800 8084 19852 8090
rect 19800 8026 19852 8032
rect 20732 7886 20760 8774
rect 20812 8016 20864 8022
rect 20810 7984 20812 7993
rect 20864 7984 20866 7993
rect 20810 7919 20866 7928
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20534 7576 20590 7585
rect 20534 7511 20590 7520
rect 20444 7472 20496 7478
rect 20444 7414 20496 7420
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19904 7041 19932 7346
rect 19890 7032 19946 7041
rect 19890 6967 19946 6976
rect 20456 6798 20484 7414
rect 20444 6792 20496 6798
rect 20444 6734 20496 6740
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 20180 4826 20208 6666
rect 20548 6390 20576 7511
rect 20732 6798 20760 7686
rect 20916 7426 20944 9590
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 21008 7546 21036 9522
rect 21192 9330 21220 11494
rect 21284 9450 21312 12406
rect 21364 12096 21416 12102
rect 21362 12064 21364 12073
rect 21416 12064 21418 12073
rect 21362 11999 21418 12008
rect 21652 11898 21680 20402
rect 21732 20392 21784 20398
rect 21732 20334 21784 20340
rect 21744 16454 21772 20334
rect 21824 20324 21876 20330
rect 21824 20266 21876 20272
rect 21732 16448 21784 16454
rect 21732 16390 21784 16396
rect 21640 11892 21692 11898
rect 21640 11834 21692 11840
rect 21454 11656 21510 11665
rect 21454 11591 21510 11600
rect 21364 11076 21416 11082
rect 21364 11018 21416 11024
rect 21376 10713 21404 11018
rect 21362 10704 21418 10713
rect 21468 10674 21496 11591
rect 21362 10639 21418 10648
rect 21456 10668 21508 10674
rect 21456 10610 21508 10616
rect 21468 9722 21496 10610
rect 21546 9752 21602 9761
rect 21456 9716 21508 9722
rect 21546 9687 21602 9696
rect 21456 9658 21508 9664
rect 21272 9444 21324 9450
rect 21272 9386 21324 9392
rect 21362 9344 21418 9353
rect 21192 9302 21312 9330
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21100 8401 21128 8434
rect 21086 8392 21142 8401
rect 21086 8327 21142 8336
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 21100 7478 21128 8327
rect 21088 7472 21140 7478
rect 20916 7398 21036 7426
rect 21088 7414 21140 7420
rect 20904 7336 20956 7342
rect 20904 7278 20956 7284
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20626 6624 20682 6633
rect 20626 6559 20682 6568
rect 20536 6384 20588 6390
rect 20536 6326 20588 6332
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20272 6089 20300 6258
rect 20548 6254 20576 6326
rect 20536 6248 20588 6254
rect 20536 6190 20588 6196
rect 20258 6080 20314 6089
rect 20258 6015 20314 6024
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20364 5273 20392 5646
rect 20640 5302 20668 6559
rect 20718 5400 20774 5409
rect 20916 5370 20944 7278
rect 20718 5335 20720 5344
rect 20772 5335 20774 5344
rect 20904 5364 20956 5370
rect 20720 5306 20772 5312
rect 20904 5306 20956 5312
rect 20628 5296 20680 5302
rect 20350 5264 20406 5273
rect 20628 5238 20680 5244
rect 20350 5199 20406 5208
rect 20904 5228 20956 5234
rect 20904 5170 20956 5176
rect 20916 4826 20944 5170
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 20442 4720 20498 4729
rect 20442 4655 20498 4664
rect 20456 4622 20484 4655
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20720 4616 20772 4622
rect 20720 4558 20772 4564
rect 20456 4282 20484 4558
rect 20732 4321 20760 4558
rect 20718 4312 20774 4321
rect 20444 4276 20496 4282
rect 20718 4247 20774 4256
rect 20444 4218 20496 4224
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20168 3460 20220 3466
rect 20168 3402 20220 3408
rect 19616 2848 19668 2854
rect 19616 2790 19668 2796
rect 19708 2848 19760 2854
rect 19708 2790 19760 2796
rect 19143 2748 19451 2768
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2672 19451 2692
rect 19628 2378 19656 2790
rect 19616 2372 19668 2378
rect 19616 2314 19668 2320
rect 19248 2304 19300 2310
rect 19248 2246 19300 2252
rect 19062 1048 19118 1057
rect 19062 983 19118 992
rect 19260 241 19288 2246
rect 19628 1601 19656 2314
rect 20180 2009 20208 3402
rect 20548 3369 20576 3470
rect 20534 3360 20590 3369
rect 20534 3295 20590 3304
rect 20720 3120 20772 3126
rect 20720 3062 20772 3068
rect 20536 2440 20588 2446
rect 20534 2408 20536 2417
rect 20588 2408 20590 2417
rect 20534 2343 20590 2352
rect 20166 2000 20222 2009
rect 20166 1935 20222 1944
rect 19614 1592 19670 1601
rect 19614 1527 19670 1536
rect 20732 649 20760 3062
rect 21008 2774 21036 7398
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 21088 7268 21140 7274
rect 21088 7210 21140 7216
rect 21100 4826 21128 7210
rect 21192 6458 21220 7346
rect 21180 6452 21232 6458
rect 21180 6394 21232 6400
rect 21284 6338 21312 9302
rect 21362 9279 21418 9288
rect 21376 8634 21404 9279
rect 21364 8628 21416 8634
rect 21364 8570 21416 8576
rect 21362 7984 21418 7993
rect 21362 7919 21364 7928
rect 21416 7919 21418 7928
rect 21364 7890 21416 7896
rect 21560 7410 21588 9687
rect 21836 9178 21864 20266
rect 21916 19916 21968 19922
rect 21916 19858 21968 19864
rect 21928 11354 21956 19858
rect 22112 18902 22140 22200
rect 22664 19786 22692 22200
rect 22652 19780 22704 19786
rect 22652 19722 22704 19728
rect 22100 18896 22152 18902
rect 22100 18838 22152 18844
rect 21916 11348 21968 11354
rect 21916 11290 21968 11296
rect 21824 9172 21876 9178
rect 21824 9114 21876 9120
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 21560 7002 21588 7346
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 21192 6310 21312 6338
rect 21088 4820 21140 4826
rect 21088 4762 21140 4768
rect 21192 4282 21220 6310
rect 21362 5672 21418 5681
rect 21362 5607 21418 5616
rect 21376 4622 21404 5607
rect 21364 4616 21416 4622
rect 21364 4558 21416 4564
rect 21180 4276 21232 4282
rect 21180 4218 21232 4224
rect 21272 4208 21324 4214
rect 21272 4150 21324 4156
rect 21284 3913 21312 4150
rect 21376 4146 21404 4558
rect 21364 4140 21416 4146
rect 21364 4082 21416 4088
rect 21270 3904 21326 3913
rect 21270 3839 21326 3848
rect 21272 3052 21324 3058
rect 21272 2994 21324 3000
rect 21284 2961 21312 2994
rect 21270 2952 21326 2961
rect 21270 2887 21326 2896
rect 20824 2746 21036 2774
rect 20824 2514 20852 2746
rect 20812 2508 20864 2514
rect 20812 2450 20864 2456
rect 20718 640 20774 649
rect 20718 575 20774 584
rect 19246 232 19302 241
rect 19246 167 19302 176
<< via2 >>
rect 1674 18284 1730 18320
rect 1674 18264 1676 18284
rect 1676 18264 1728 18284
rect 1728 18264 1730 18284
rect 1490 17176 1546 17232
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 10966 18808 11022 18864
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 11702 12280 11758 12336
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 18878 22616 18934 22672
rect 14094 17584 14150 17640
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 1398 5752 1454 5808
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16578 12280 16634 12336
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 18694 22072 18750 22128
rect 18326 18808 18382 18864
rect 18326 18264 18382 18320
rect 18602 19488 18658 19544
rect 19062 21256 19118 21312
rect 18602 19372 18658 19408
rect 18602 19352 18604 19372
rect 18604 19352 18656 19372
rect 18656 19352 18658 19372
rect 19614 20848 19670 20904
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 20074 19896 20130 19952
rect 18786 17604 18842 17640
rect 18786 17584 18788 17604
rect 18788 17584 18840 17604
rect 18840 17584 18842 17604
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19246 12688 19302 12744
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 18878 10512 18934 10568
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 20534 20304 20590 20360
rect 21454 21664 21510 21720
rect 20718 19352 20774 19408
rect 20718 17584 20774 17640
rect 20626 17176 20682 17232
rect 20626 12960 20682 13016
rect 21270 18944 21326 19000
rect 21362 18536 21418 18592
rect 21270 17992 21326 18048
rect 21270 16632 21326 16688
rect 21362 16224 21418 16280
rect 21270 15680 21326 15736
rect 21362 15272 21418 15328
rect 21270 14864 21326 14920
rect 21270 14320 21326 14376
rect 21270 13912 21326 13968
rect 21270 13504 21326 13560
rect 21362 12980 21418 13016
rect 21362 12960 21364 12980
rect 21364 12960 21416 12980
rect 21416 12960 21418 12980
rect 20902 11192 20958 11248
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 20534 8916 20536 8936
rect 20536 8916 20588 8936
rect 20588 8916 20590 8936
rect 20534 8880 20590 8916
rect 20810 7964 20812 7984
rect 20812 7964 20864 7984
rect 20864 7964 20866 7984
rect 20810 7928 20866 7964
rect 20534 7520 20590 7576
rect 19890 6976 19946 7032
rect 21362 12044 21364 12064
rect 21364 12044 21416 12064
rect 21416 12044 21418 12064
rect 21362 12008 21418 12044
rect 21454 11600 21510 11656
rect 21362 10648 21418 10704
rect 21546 9696 21602 9752
rect 21086 8336 21142 8392
rect 20626 6568 20682 6624
rect 20258 6024 20314 6080
rect 20718 5364 20774 5400
rect 20718 5344 20720 5364
rect 20720 5344 20772 5364
rect 20772 5344 20774 5364
rect 20350 5208 20406 5264
rect 20442 4664 20498 4720
rect 20718 4256 20774 4312
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 19062 992 19118 1048
rect 20534 3304 20590 3360
rect 20534 2388 20536 2408
rect 20536 2388 20588 2408
rect 20588 2388 20590 2408
rect 20534 2352 20590 2388
rect 20166 1944 20222 2000
rect 19614 1536 19670 1592
rect 21362 9288 21418 9344
rect 21362 7948 21418 7984
rect 21362 7928 21364 7948
rect 21364 7928 21416 7948
rect 21416 7928 21418 7948
rect 21362 5616 21418 5672
rect 21270 3848 21326 3904
rect 21270 2896 21326 2952
rect 20718 584 20774 640
rect 19246 176 19302 232
<< metal3 >>
rect 18873 22674 18939 22677
rect 22200 22674 23000 22704
rect 18873 22672 23000 22674
rect 18873 22616 18878 22672
rect 18934 22616 23000 22672
rect 18873 22614 23000 22616
rect 18873 22611 18939 22614
rect 22200 22584 23000 22614
rect 22200 22266 23000 22296
rect 18830 22206 23000 22266
rect 18689 22130 18755 22133
rect 18830 22130 18890 22206
rect 22200 22176 23000 22206
rect 18689 22128 18890 22130
rect 18689 22072 18694 22128
rect 18750 22072 18890 22128
rect 18689 22070 18890 22072
rect 18689 22067 18755 22070
rect 21449 21722 21515 21725
rect 22200 21722 23000 21752
rect 21449 21720 23000 21722
rect 21449 21664 21454 21720
rect 21510 21664 23000 21720
rect 21449 21662 23000 21664
rect 21449 21659 21515 21662
rect 22200 21632 23000 21662
rect 19057 21314 19123 21317
rect 22200 21314 23000 21344
rect 19057 21312 23000 21314
rect 19057 21256 19062 21312
rect 19118 21256 23000 21312
rect 19057 21254 23000 21256
rect 19057 21251 19123 21254
rect 22200 21224 23000 21254
rect 19609 20906 19675 20909
rect 22200 20906 23000 20936
rect 19609 20904 23000 20906
rect 19609 20848 19614 20904
rect 19670 20848 23000 20904
rect 19609 20846 23000 20848
rect 19609 20843 19675 20846
rect 22200 20816 23000 20846
rect 6142 20704 6462 20705
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 20639 6462 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 16538 20704 16858 20705
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 20639 16858 20640
rect 20529 20362 20595 20365
rect 22200 20362 23000 20392
rect 20529 20360 23000 20362
rect 20529 20304 20534 20360
rect 20590 20304 23000 20360
rect 20529 20302 23000 20304
rect 20529 20299 20595 20302
rect 22200 20272 23000 20302
rect 3543 20160 3863 20161
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 20095 3863 20096
rect 8741 20160 9061 20161
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 20095 9061 20096
rect 13939 20160 14259 20161
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 20095 14259 20096
rect 19137 20160 19457 20161
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 20095 19457 20096
rect 20069 19954 20135 19957
rect 22200 19954 23000 19984
rect 20069 19952 23000 19954
rect 20069 19896 20074 19952
rect 20130 19896 23000 19952
rect 20069 19894 23000 19896
rect 20069 19891 20135 19894
rect 22200 19864 23000 19894
rect 6142 19616 6462 19617
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 19551 6462 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 16538 19616 16858 19617
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 19551 16858 19552
rect 18597 19546 18663 19549
rect 18822 19546 18828 19548
rect 18597 19544 18828 19546
rect 18597 19488 18602 19544
rect 18658 19488 18828 19544
rect 18597 19486 18828 19488
rect 18597 19483 18663 19486
rect 18822 19484 18828 19486
rect 18892 19484 18898 19548
rect 18597 19412 18663 19413
rect 18597 19408 18644 19412
rect 18708 19410 18714 19412
rect 20713 19410 20779 19413
rect 22200 19410 23000 19440
rect 18597 19352 18602 19408
rect 18597 19348 18644 19352
rect 18708 19350 18754 19410
rect 20713 19408 23000 19410
rect 20713 19352 20718 19408
rect 20774 19352 23000 19408
rect 20713 19350 23000 19352
rect 18708 19348 18714 19350
rect 18597 19347 18663 19348
rect 20713 19347 20779 19350
rect 22200 19320 23000 19350
rect 3543 19072 3863 19073
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 19007 3863 19008
rect 8741 19072 9061 19073
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 19007 9061 19008
rect 13939 19072 14259 19073
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 19007 14259 19008
rect 19137 19072 19457 19073
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 19007 19457 19008
rect 21265 19002 21331 19005
rect 22200 19002 23000 19032
rect 21265 19000 23000 19002
rect 21265 18944 21270 19000
rect 21326 18944 23000 19000
rect 21265 18942 23000 18944
rect 21265 18939 21331 18942
rect 22200 18912 23000 18942
rect 10961 18866 11027 18869
rect 18321 18866 18387 18869
rect 10961 18864 18387 18866
rect 10961 18808 10966 18864
rect 11022 18808 18326 18864
rect 18382 18808 18387 18864
rect 10961 18806 18387 18808
rect 10961 18803 11027 18806
rect 18321 18803 18387 18806
rect 21357 18594 21423 18597
rect 22200 18594 23000 18624
rect 21357 18592 23000 18594
rect 21357 18536 21362 18592
rect 21418 18536 23000 18592
rect 21357 18534 23000 18536
rect 21357 18531 21423 18534
rect 6142 18528 6462 18529
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 18463 6462 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 16538 18528 16858 18529
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 22200 18504 23000 18534
rect 16538 18463 16858 18464
rect 1669 18322 1735 18325
rect 18321 18322 18387 18325
rect 1669 18320 18387 18322
rect 1669 18264 1674 18320
rect 1730 18264 18326 18320
rect 18382 18264 18387 18320
rect 1669 18262 18387 18264
rect 1669 18259 1735 18262
rect 18321 18259 18387 18262
rect 21265 18050 21331 18053
rect 22200 18050 23000 18080
rect 21265 18048 23000 18050
rect 21265 17992 21270 18048
rect 21326 17992 23000 18048
rect 21265 17990 23000 17992
rect 21265 17987 21331 17990
rect 3543 17984 3863 17985
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 17919 3863 17920
rect 8741 17984 9061 17985
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 17919 9061 17920
rect 13939 17984 14259 17985
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 17919 14259 17920
rect 19137 17984 19457 17985
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 22200 17960 23000 17990
rect 19137 17919 19457 17920
rect 14089 17642 14155 17645
rect 18781 17642 18847 17645
rect 14089 17640 18847 17642
rect 14089 17584 14094 17640
rect 14150 17584 18786 17640
rect 18842 17584 18847 17640
rect 14089 17582 18847 17584
rect 14089 17579 14155 17582
rect 18781 17579 18847 17582
rect 20713 17642 20779 17645
rect 22200 17642 23000 17672
rect 20713 17640 23000 17642
rect 20713 17584 20718 17640
rect 20774 17584 23000 17640
rect 20713 17582 23000 17584
rect 20713 17579 20779 17582
rect 22200 17552 23000 17582
rect 6142 17440 6462 17441
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 17375 6462 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 16538 17440 16858 17441
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 17375 16858 17376
rect 0 17234 800 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 800 17174
rect 1485 17171 1551 17174
rect 20621 17234 20687 17237
rect 22200 17234 23000 17264
rect 20621 17232 23000 17234
rect 20621 17176 20626 17232
rect 20682 17176 23000 17232
rect 20621 17174 23000 17176
rect 20621 17171 20687 17174
rect 22200 17144 23000 17174
rect 3543 16896 3863 16897
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 16831 3863 16832
rect 8741 16896 9061 16897
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 16831 9061 16832
rect 13939 16896 14259 16897
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 16831 14259 16832
rect 19137 16896 19457 16897
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 16831 19457 16832
rect 21265 16690 21331 16693
rect 22200 16690 23000 16720
rect 21265 16688 23000 16690
rect 21265 16632 21270 16688
rect 21326 16632 23000 16688
rect 21265 16630 23000 16632
rect 21265 16627 21331 16630
rect 22200 16600 23000 16630
rect 6142 16352 6462 16353
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 16287 6462 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 16538 16352 16858 16353
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 16287 16858 16288
rect 21357 16282 21423 16285
rect 22200 16282 23000 16312
rect 21357 16280 23000 16282
rect 21357 16224 21362 16280
rect 21418 16224 23000 16280
rect 21357 16222 23000 16224
rect 21357 16219 21423 16222
rect 22200 16192 23000 16222
rect 3543 15808 3863 15809
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 15743 3863 15744
rect 8741 15808 9061 15809
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 15743 9061 15744
rect 13939 15808 14259 15809
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 15743 14259 15744
rect 19137 15808 19457 15809
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 15743 19457 15744
rect 21265 15738 21331 15741
rect 22200 15738 23000 15768
rect 21265 15736 23000 15738
rect 21265 15680 21270 15736
rect 21326 15680 23000 15736
rect 21265 15678 23000 15680
rect 21265 15675 21331 15678
rect 22200 15648 23000 15678
rect 21357 15330 21423 15333
rect 22200 15330 23000 15360
rect 21357 15328 23000 15330
rect 21357 15272 21362 15328
rect 21418 15272 23000 15328
rect 21357 15270 23000 15272
rect 21357 15267 21423 15270
rect 6142 15264 6462 15265
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 15199 6462 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 16538 15264 16858 15265
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 22200 15240 23000 15270
rect 16538 15199 16858 15200
rect 21265 14922 21331 14925
rect 22200 14922 23000 14952
rect 21265 14920 23000 14922
rect 21265 14864 21270 14920
rect 21326 14864 23000 14920
rect 21265 14862 23000 14864
rect 21265 14859 21331 14862
rect 22200 14832 23000 14862
rect 3543 14720 3863 14721
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 14655 3863 14656
rect 8741 14720 9061 14721
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 14655 9061 14656
rect 13939 14720 14259 14721
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 14655 14259 14656
rect 19137 14720 19457 14721
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 14655 19457 14656
rect 21265 14378 21331 14381
rect 22200 14378 23000 14408
rect 21265 14376 23000 14378
rect 21265 14320 21270 14376
rect 21326 14320 23000 14376
rect 21265 14318 23000 14320
rect 21265 14315 21331 14318
rect 22200 14288 23000 14318
rect 6142 14176 6462 14177
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 14111 6462 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 16538 14176 16858 14177
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 14111 16858 14112
rect 21265 13970 21331 13973
rect 22200 13970 23000 14000
rect 21265 13968 23000 13970
rect 21265 13912 21270 13968
rect 21326 13912 23000 13968
rect 21265 13910 23000 13912
rect 21265 13907 21331 13910
rect 22200 13880 23000 13910
rect 3543 13632 3863 13633
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 13567 3863 13568
rect 8741 13632 9061 13633
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 13567 9061 13568
rect 13939 13632 14259 13633
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 13567 14259 13568
rect 19137 13632 19457 13633
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 13567 19457 13568
rect 21265 13562 21331 13565
rect 22200 13562 23000 13592
rect 21265 13560 23000 13562
rect 21265 13504 21270 13560
rect 21326 13504 23000 13560
rect 21265 13502 23000 13504
rect 21265 13499 21331 13502
rect 22200 13472 23000 13502
rect 6142 13088 6462 13089
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 13023 6462 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 16538 13088 16858 13089
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 13023 16858 13024
rect 20621 13018 20687 13021
rect 21357 13018 21423 13021
rect 22200 13018 23000 13048
rect 20621 13016 23000 13018
rect 20621 12960 20626 13016
rect 20682 12960 21362 13016
rect 21418 12960 23000 13016
rect 20621 12958 23000 12960
rect 20621 12955 20687 12958
rect 21357 12955 21423 12958
rect 22200 12928 23000 12958
rect 19241 12746 19307 12749
rect 19241 12744 19626 12746
rect 19241 12688 19246 12744
rect 19302 12688 19626 12744
rect 19241 12686 19626 12688
rect 19241 12683 19307 12686
rect 19566 12610 19626 12686
rect 22200 12610 23000 12640
rect 19566 12550 23000 12610
rect 3543 12544 3863 12545
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 12479 3863 12480
rect 8741 12544 9061 12545
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 12479 9061 12480
rect 13939 12544 14259 12545
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 12479 14259 12480
rect 19137 12544 19457 12545
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 22200 12520 23000 12550
rect 19137 12479 19457 12480
rect 11697 12338 11763 12341
rect 16573 12338 16639 12341
rect 11697 12336 16639 12338
rect 11697 12280 11702 12336
rect 11758 12280 16578 12336
rect 16634 12280 16639 12336
rect 11697 12278 16639 12280
rect 11697 12275 11763 12278
rect 16573 12275 16639 12278
rect 21357 12066 21423 12069
rect 22200 12066 23000 12096
rect 21357 12064 23000 12066
rect 21357 12008 21362 12064
rect 21418 12008 23000 12064
rect 21357 12006 23000 12008
rect 21357 12003 21423 12006
rect 6142 12000 6462 12001
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 11935 6462 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 16538 12000 16858 12001
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 22200 11976 23000 12006
rect 16538 11935 16858 11936
rect 21449 11658 21515 11661
rect 22200 11658 23000 11688
rect 21449 11656 23000 11658
rect 21449 11600 21454 11656
rect 21510 11600 23000 11656
rect 21449 11598 23000 11600
rect 21449 11595 21515 11598
rect 22200 11568 23000 11598
rect 3543 11456 3863 11457
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 11391 3863 11392
rect 8741 11456 9061 11457
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 11391 9061 11392
rect 13939 11456 14259 11457
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 11391 14259 11392
rect 19137 11456 19457 11457
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 11391 19457 11392
rect 20897 11250 20963 11253
rect 22200 11250 23000 11280
rect 20897 11248 23000 11250
rect 20897 11192 20902 11248
rect 20958 11192 23000 11248
rect 20897 11190 23000 11192
rect 20897 11187 20963 11190
rect 22200 11160 23000 11190
rect 6142 10912 6462 10913
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 10847 6462 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 16538 10912 16858 10913
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 10847 16858 10848
rect 21357 10706 21423 10709
rect 22200 10706 23000 10736
rect 21357 10704 23000 10706
rect 21357 10648 21362 10704
rect 21418 10648 23000 10704
rect 21357 10646 23000 10648
rect 21357 10643 21423 10646
rect 22200 10616 23000 10646
rect 18873 10570 18939 10573
rect 18873 10568 19626 10570
rect 18873 10512 18878 10568
rect 18934 10512 19626 10568
rect 18873 10510 19626 10512
rect 18873 10507 18939 10510
rect 3543 10368 3863 10369
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 10303 3863 10304
rect 8741 10368 9061 10369
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 10303 9061 10304
rect 13939 10368 14259 10369
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 10303 14259 10304
rect 19137 10368 19457 10369
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 10303 19457 10304
rect 19566 10298 19626 10510
rect 22200 10298 23000 10328
rect 19566 10238 23000 10298
rect 22200 10208 23000 10238
rect 6142 9824 6462 9825
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 9759 6462 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 16538 9824 16858 9825
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 9759 16858 9760
rect 21541 9754 21607 9757
rect 22200 9754 23000 9784
rect 21541 9752 23000 9754
rect 21541 9696 21546 9752
rect 21602 9696 23000 9752
rect 21541 9694 23000 9696
rect 21541 9691 21607 9694
rect 22200 9664 23000 9694
rect 21357 9346 21423 9349
rect 22200 9346 23000 9376
rect 21357 9344 23000 9346
rect 21357 9288 21362 9344
rect 21418 9288 23000 9344
rect 21357 9286 23000 9288
rect 21357 9283 21423 9286
rect 3543 9280 3863 9281
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 9215 3863 9216
rect 8741 9280 9061 9281
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 9215 9061 9216
rect 13939 9280 14259 9281
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 9215 14259 9216
rect 19137 9280 19457 9281
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 22200 9256 23000 9286
rect 19137 9215 19457 9216
rect 20529 8938 20595 8941
rect 22200 8938 23000 8968
rect 20529 8936 23000 8938
rect 20529 8880 20534 8936
rect 20590 8880 23000 8936
rect 20529 8878 23000 8880
rect 20529 8875 20595 8878
rect 22200 8848 23000 8878
rect 6142 8736 6462 8737
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 8671 6462 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 16538 8736 16858 8737
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 8671 16858 8672
rect 21081 8394 21147 8397
rect 22200 8394 23000 8424
rect 21081 8392 23000 8394
rect 21081 8336 21086 8392
rect 21142 8336 23000 8392
rect 21081 8334 23000 8336
rect 21081 8331 21147 8334
rect 22200 8304 23000 8334
rect 3543 8192 3863 8193
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 8127 3863 8128
rect 8741 8192 9061 8193
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 8127 9061 8128
rect 13939 8192 14259 8193
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 8127 14259 8128
rect 19137 8192 19457 8193
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 8127 19457 8128
rect 18822 7924 18828 7988
rect 18892 7986 18898 7988
rect 20805 7986 20871 7989
rect 18892 7984 20871 7986
rect 18892 7928 20810 7984
rect 20866 7928 20871 7984
rect 18892 7926 20871 7928
rect 18892 7924 18898 7926
rect 20805 7923 20871 7926
rect 21357 7986 21423 7989
rect 22200 7986 23000 8016
rect 21357 7984 23000 7986
rect 21357 7928 21362 7984
rect 21418 7928 23000 7984
rect 21357 7926 23000 7928
rect 21357 7923 21423 7926
rect 22200 7896 23000 7926
rect 6142 7648 6462 7649
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 7583 6462 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 16538 7648 16858 7649
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 7583 16858 7584
rect 20529 7578 20595 7581
rect 22200 7578 23000 7608
rect 20529 7576 23000 7578
rect 20529 7520 20534 7576
rect 20590 7520 23000 7576
rect 20529 7518 23000 7520
rect 20529 7515 20595 7518
rect 22200 7488 23000 7518
rect 3543 7104 3863 7105
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 7039 3863 7040
rect 8741 7104 9061 7105
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 7039 9061 7040
rect 13939 7104 14259 7105
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 7039 14259 7040
rect 19137 7104 19457 7105
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 7039 19457 7040
rect 19885 7034 19951 7037
rect 22200 7034 23000 7064
rect 19885 7032 23000 7034
rect 19885 6976 19890 7032
rect 19946 6976 23000 7032
rect 19885 6974 23000 6976
rect 19885 6971 19951 6974
rect 22200 6944 23000 6974
rect 20621 6626 20687 6629
rect 22200 6626 23000 6656
rect 20621 6624 23000 6626
rect 20621 6568 20626 6624
rect 20682 6568 23000 6624
rect 20621 6566 23000 6568
rect 20621 6563 20687 6566
rect 6142 6560 6462 6561
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 6495 6462 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 16538 6560 16858 6561
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 22200 6536 23000 6566
rect 16538 6495 16858 6496
rect 20253 6082 20319 6085
rect 22200 6082 23000 6112
rect 20253 6080 23000 6082
rect 20253 6024 20258 6080
rect 20314 6024 23000 6080
rect 20253 6022 23000 6024
rect 20253 6019 20319 6022
rect 3543 6016 3863 6017
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 5951 3863 5952
rect 8741 6016 9061 6017
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 5951 9061 5952
rect 13939 6016 14259 6017
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 5951 14259 5952
rect 19137 6016 19457 6017
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 22200 5992 23000 6022
rect 19137 5951 19457 5952
rect 0 5810 800 5840
rect 1393 5810 1459 5813
rect 0 5808 1459 5810
rect 0 5752 1398 5808
rect 1454 5752 1459 5808
rect 0 5750 1459 5752
rect 0 5720 800 5750
rect 1393 5747 1459 5750
rect 21357 5674 21423 5677
rect 22200 5674 23000 5704
rect 21357 5672 23000 5674
rect 21357 5616 21362 5672
rect 21418 5616 23000 5672
rect 21357 5614 23000 5616
rect 21357 5611 21423 5614
rect 22200 5584 23000 5614
rect 6142 5472 6462 5473
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 5407 6462 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 16538 5472 16858 5473
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 5407 16858 5408
rect 18638 5340 18644 5404
rect 18708 5402 18714 5404
rect 20713 5402 20779 5405
rect 18708 5400 20779 5402
rect 18708 5344 20718 5400
rect 20774 5344 20779 5400
rect 18708 5342 20779 5344
rect 18708 5340 18714 5342
rect 20713 5339 20779 5342
rect 20345 5266 20411 5269
rect 22200 5266 23000 5296
rect 20345 5264 23000 5266
rect 20345 5208 20350 5264
rect 20406 5208 23000 5264
rect 20345 5206 23000 5208
rect 20345 5203 20411 5206
rect 22200 5176 23000 5206
rect 3543 4928 3863 4929
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 4863 3863 4864
rect 8741 4928 9061 4929
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 4863 9061 4864
rect 13939 4928 14259 4929
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 4863 14259 4864
rect 19137 4928 19457 4929
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 4863 19457 4864
rect 20437 4722 20503 4725
rect 22200 4722 23000 4752
rect 20437 4720 23000 4722
rect 20437 4664 20442 4720
rect 20498 4664 23000 4720
rect 20437 4662 23000 4664
rect 20437 4659 20503 4662
rect 22200 4632 23000 4662
rect 6142 4384 6462 4385
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 4319 6462 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 16538 4384 16858 4385
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 4319 16858 4320
rect 20713 4314 20779 4317
rect 22200 4314 23000 4344
rect 20713 4312 23000 4314
rect 20713 4256 20718 4312
rect 20774 4256 23000 4312
rect 20713 4254 23000 4256
rect 20713 4251 20779 4254
rect 22200 4224 23000 4254
rect 21265 3906 21331 3909
rect 22200 3906 23000 3936
rect 21265 3904 23000 3906
rect 21265 3848 21270 3904
rect 21326 3848 23000 3904
rect 21265 3846 23000 3848
rect 21265 3843 21331 3846
rect 3543 3840 3863 3841
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 3775 3863 3776
rect 8741 3840 9061 3841
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 3775 9061 3776
rect 13939 3840 14259 3841
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 3775 14259 3776
rect 19137 3840 19457 3841
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 22200 3816 23000 3846
rect 19137 3775 19457 3776
rect 20529 3362 20595 3365
rect 22200 3362 23000 3392
rect 20529 3360 23000 3362
rect 20529 3304 20534 3360
rect 20590 3304 23000 3360
rect 20529 3302 23000 3304
rect 20529 3299 20595 3302
rect 6142 3296 6462 3297
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 3231 6462 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 16538 3296 16858 3297
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 22200 3272 23000 3302
rect 16538 3231 16858 3232
rect 21265 2954 21331 2957
rect 22200 2954 23000 2984
rect 21265 2952 23000 2954
rect 21265 2896 21270 2952
rect 21326 2896 23000 2952
rect 21265 2894 23000 2896
rect 21265 2891 21331 2894
rect 22200 2864 23000 2894
rect 3543 2752 3863 2753
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2687 3863 2688
rect 8741 2752 9061 2753
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2687 9061 2688
rect 13939 2752 14259 2753
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2687 14259 2688
rect 19137 2752 19457 2753
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2687 19457 2688
rect 20529 2410 20595 2413
rect 22200 2410 23000 2440
rect 20529 2408 23000 2410
rect 20529 2352 20534 2408
rect 20590 2352 23000 2408
rect 20529 2350 23000 2352
rect 20529 2347 20595 2350
rect 22200 2320 23000 2350
rect 6142 2208 6462 2209
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2143 6462 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 16538 2208 16858 2209
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2143 16858 2144
rect 20161 2002 20227 2005
rect 22200 2002 23000 2032
rect 20161 2000 23000 2002
rect 20161 1944 20166 2000
rect 20222 1944 23000 2000
rect 20161 1942 23000 1944
rect 20161 1939 20227 1942
rect 22200 1912 23000 1942
rect 19609 1594 19675 1597
rect 22200 1594 23000 1624
rect 19609 1592 23000 1594
rect 19609 1536 19614 1592
rect 19670 1536 23000 1592
rect 19609 1534 23000 1536
rect 19609 1531 19675 1534
rect 22200 1504 23000 1534
rect 19057 1050 19123 1053
rect 22200 1050 23000 1080
rect 19057 1048 23000 1050
rect 19057 992 19062 1048
rect 19118 992 23000 1048
rect 19057 990 23000 992
rect 19057 987 19123 990
rect 22200 960 23000 990
rect 20713 642 20779 645
rect 22200 642 23000 672
rect 20713 640 23000 642
rect 20713 584 20718 640
rect 20774 584 23000 640
rect 20713 582 23000 584
rect 20713 579 20779 582
rect 22200 552 23000 582
rect 19241 234 19307 237
rect 22200 234 23000 264
rect 19241 232 23000 234
rect 19241 176 19246 232
rect 19302 176 23000 232
rect 19241 174 23000 176
rect 19241 171 19307 174
rect 22200 144 23000 174
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 18828 19484 18892 19548
rect 18644 19408 18708 19412
rect 18644 19352 18658 19408
rect 18658 19352 18708 19408
rect 18644 19348 18708 19352
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 18828 7924 18892 7988
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 18644 5340 18708 5404
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 18827 19548 18893 19549
rect 18827 19484 18828 19548
rect 18892 19484 18893 19548
rect 18827 19483 18893 19484
rect 18643 19412 18709 19413
rect 18643 19348 18644 19412
rect 18708 19348 18709 19412
rect 18643 19347 18709 19348
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 18646 5405 18706 19347
rect 18830 7989 18890 19483
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 18827 7988 18893 7989
rect 18827 7924 18828 7988
rect 18892 7924 18893 7988
rect 18827 7923 18893 7924
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 18643 5404 18709 5405
rect 18643 5340 18644 5404
rect 18708 5340 18709 5404
rect 18643 5339 18709 5340
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2024 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 20056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 20608 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 18676 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 20976 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 19228 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 20700 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 20148 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 20332 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 20056 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 20516 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 19688 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 19688 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform 1 0 21252 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 20976 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 7544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 6256 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 6716 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 8280 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 7912 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 8096 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 9108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 10396 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 2760 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 1840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 1840 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 2760 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 3220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 3220 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 2852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 4324 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 5796 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 18584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 18676 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 19412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 19964 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 19044 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 19780 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 19780 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 3588 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17664 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 18308 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 18768 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 19504 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15088 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12604 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 14720 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14720 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 16744 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11040 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10212 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12512 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_6.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 16744 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 10120 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_10.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5152 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_12.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4232 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_14.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5244 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_18.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12512 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14720 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_22.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17480 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_26.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_28.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8280 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_30.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10028 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 16560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17756 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output84_A
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output86_A
timestamp 1649977179
transform 1 0 14536 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 19780 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_181 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_187
timestamp 1649977179
transform 1 0 18308 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_190 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1649977179
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_203
timestamp 1649977179
transform 1 0 19780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_181 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_191
timestamp 1649977179
transform 1 0 18676 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_195
timestamp 1649977179
transform 1 0 19044 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_199
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_203
timestamp 1649977179
transform 1 0 19780 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1649977179
transform 1 0 20332 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_215
timestamp 1649977179
transform 1 0 20884 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1649977179
transform 1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_199
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_203
timestamp 1649977179
transform 1 0 19780 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_201
timestamp 1649977179
transform 1 0 19596 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_209
timestamp 1649977179
transform 1 0 20332 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_213
timestamp 1649977179
transform 1 0 20700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1649977179
transform 1 0 21436 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_203
timestamp 1649977179
transform 1 0 19780 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_206
timestamp 1649977179
transform 1 0 20056 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_211
timestamp 1649977179
transform 1 0 20516 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_216
timestamp 1649977179
transform 1 0 20976 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_211
timestamp 1649977179
transform 1 0 20516 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_216
timestamp 1649977179
transform 1 0 20976 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_221
timestamp 1649977179
transform 1 0 21436 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_207
timestamp 1649977179
transform 1 0 20148 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1649977179
transform 1 0 20608 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_218
timestamp 1649977179
transform 1 0 21160 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_222
timestamp 1649977179
transform 1 0 21528 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1649977179
transform 1 0 1656 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_10
timestamp 1649977179
transform 1 0 2024 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_22
timestamp 1649977179
transform 1 0 3128 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_34
timestamp 1649977179
transform 1 0 4232 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_46
timestamp 1649977179
transform 1 0 5336 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_199
timestamp 1649977179
transform 1 0 19412 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_202
timestamp 1649977179
transform 1 0 19688 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_206
timestamp 1649977179
transform 1 0 20056 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_211
timestamp 1649977179
transform 1 0 20516 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_216
timestamp 1649977179
transform 1 0 20976 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_107
timestamp 1649977179
transform 1 0 10948 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_118
timestamp 1649977179
transform 1 0 11960 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_130
timestamp 1649977179
transform 1 0 13064 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_151
timestamp 1649977179
transform 1 0 14996 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_163
timestamp 1649977179
transform 1 0 16100 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_175
timestamp 1649977179
transform 1 0 17204 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_183
timestamp 1649977179
transform 1 0 17940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_212
timestamp 1649977179
transform 1 0 20608 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_217
timestamp 1649977179
transform 1 0 21068 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_91
timestamp 1649977179
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1649977179
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_122
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_138
timestamp 1649977179
transform 1 0 13800 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_160
timestamp 1649977179
transform 1 0 15824 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_192
timestamp 1649977179
transform 1 0 18768 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_202
timestamp 1649977179
transform 1 0 19688 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_207
timestamp 1649977179
transform 1 0 20148 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_212
timestamp 1649977179
transform 1 0 20608 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_216
timestamp 1649977179
transform 1 0 20976 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1649977179
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1649977179
transform 1 0 9660 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_110
timestamp 1649977179
transform 1 0 11224 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_114
timestamp 1649977179
transform 1 0 11592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_131
timestamp 1649977179
transform 1 0 13156 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_157
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_175
timestamp 1649977179
transform 1 0 17204 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_193
timestamp 1649977179
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_205
timestamp 1649977179
transform 1 0 19964 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_210
timestamp 1649977179
transform 1 0 20424 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_217
timestamp 1649977179
transform 1 0 21068 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_89
timestamp 1649977179
transform 1 0 9292 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_98
timestamp 1649977179
transform 1 0 10120 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_106
timestamp 1649977179
transform 1 0 10856 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_121
timestamp 1649977179
transform 1 0 12236 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_126
timestamp 1649977179
transform 1 0 12696 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_11_148
timestamp 1649977179
transform 1 0 14720 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_173
timestamp 1649977179
transform 1 0 17020 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_182
timestamp 1649977179
transform 1 0 17848 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_202
timestamp 1649977179
transform 1 0 19688 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_207
timestamp 1649977179
transform 1 0 20148 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_212
timestamp 1649977179
transform 1 0 20608 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_113
timestamp 1649977179
transform 1 0 11500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_117
timestamp 1649977179
transform 1 0 11868 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_129
timestamp 1649977179
transform 1 0 12972 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_147
timestamp 1649977179
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_150
timestamp 1649977179
transform 1 0 14904 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_162
timestamp 1649977179
transform 1 0 16008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_168
timestamp 1649977179
transform 1 0 16560 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_176
timestamp 1649977179
transform 1 0 17296 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_180
timestamp 1649977179
transform 1 0 17664 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1649977179
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_214
timestamp 1649977179
transform 1 0 20792 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_219
timestamp 1649977179
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_146
timestamp 1649977179
transform 1 0 14536 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_150
timestamp 1649977179
transform 1 0 14904 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_157
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_165
timestamp 1649977179
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_189
timestamp 1649977179
transform 1 0 18492 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_208
timestamp 1649977179
transform 1 0 20240 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_212
timestamp 1649977179
transform 1 0 20608 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_114
timestamp 1649977179
transform 1 0 11592 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_132
timestamp 1649977179
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_157
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_168
timestamp 1649977179
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_172
timestamp 1649977179
transform 1 0 16928 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_190
timestamp 1649977179
transform 1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_219
timestamp 1649977179
transform 1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_15_101
timestamp 1649977179
transform 1 0 10396 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1649977179
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_122
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_126
timestamp 1649977179
transform 1 0 12696 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_160
timestamp 1649977179
transform 1 0 15824 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_185
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_191
timestamp 1649977179
transform 1 0 18676 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_196
timestamp 1649977179
transform 1 0 19136 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_207
timestamp 1649977179
transform 1 0 20148 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_212
timestamp 1649977179
transform 1 0 20608 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_216
timestamp 1649977179
transform 1 0 20976 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_101
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_112
timestamp 1649977179
transform 1 0 11408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_117
timestamp 1649977179
transform 1 0 11868 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_123
timestamp 1649977179
transform 1 0 12420 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_127
timestamp 1649977179
transform 1 0 12788 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_150
timestamp 1649977179
transform 1 0 14904 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_154
timestamp 1649977179
transform 1 0 15272 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_166
timestamp 1649977179
transform 1 0 16376 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_178
timestamp 1649977179
transform 1 0 17480 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_190
timestamp 1649977179
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_200
timestamp 1649977179
transform 1 0 19504 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_207
timestamp 1649977179
transform 1 0 20148 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_212
timestamp 1649977179
transform 1 0 20608 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_217
timestamp 1649977179
transform 1 0 21068 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_77
timestamp 1649977179
transform 1 0 8188 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_99
timestamp 1649977179
transform 1 0 10212 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_122
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_130
timestamp 1649977179
transform 1 0 13064 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_147
timestamp 1649977179
transform 1 0 14628 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_157
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1649977179
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_178
timestamp 1649977179
transform 1 0 17480 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_189
timestamp 1649977179
transform 1 0 18492 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1649977179
transform 1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_212
timestamp 1649977179
transform 1 0 20608 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_87
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_106
timestamp 1649977179
transform 1 0 10856 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_110
timestamp 1649977179
transform 1 0 11224 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_129
timestamp 1649977179
transform 1 0 12972 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 1649977179
transform 1 0 13708 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_144
timestamp 1649977179
transform 1 0 14352 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_163
timestamp 1649977179
transform 1 0 16100 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_174
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_185
timestamp 1649977179
transform 1 0 18124 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_190
timestamp 1649977179
transform 1 0 18584 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1649977179
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_202
timestamp 1649977179
transform 1 0 19688 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_207
timestamp 1649977179
transform 1 0 20148 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1649977179
transform 1 0 20608 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_217
timestamp 1649977179
transform 1 0 21068 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_65
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_77
timestamp 1649977179
transform 1 0 8188 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_89
timestamp 1649977179
transform 1 0 9292 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_101
timestamp 1649977179
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1649977179
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_117
timestamp 1649977179
transform 1 0 11868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_127
timestamp 1649977179
transform 1 0 12788 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_178
timestamp 1649977179
transform 1 0 17480 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_182
timestamp 1649977179
transform 1 0 17848 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_186
timestamp 1649977179
transform 1 0 18216 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_19_197
timestamp 1649977179
transform 1 0 19228 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_202
timestamp 1649977179
transform 1 0 19688 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_207
timestamp 1649977179
transform 1 0 20148 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_212
timestamp 1649977179
transform 1 0 20608 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1649977179
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_49
timestamp 1649977179
transform 1 0 5612 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_68
timestamp 1649977179
transform 1 0 7360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1649977179
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_94
timestamp 1649977179
transform 1 0 9752 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_98
timestamp 1649977179
transform 1 0 10120 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_120
timestamp 1649977179
transform 1 0 12144 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_131
timestamp 1649977179
transform 1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_135
timestamp 1649977179
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_179
timestamp 1649977179
transform 1 0 17572 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_190
timestamp 1649977179
transform 1 0 18584 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_206
timestamp 1649977179
transform 1 0 20056 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_212
timestamp 1649977179
transform 1 0 20608 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_217
timestamp 1649977179
transform 1 0 21068 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_44
timestamp 1649977179
transform 1 0 5152 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_87
timestamp 1649977179
transform 1 0 9108 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_103
timestamp 1649977179
transform 1 0 10580 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1649977179
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_115
timestamp 1649977179
transform 1 0 11684 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_121
timestamp 1649977179
transform 1 0 12236 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_131
timestamp 1649977179
transform 1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_135
timestamp 1649977179
transform 1 0 13524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_139
timestamp 1649977179
transform 1 0 13892 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_147
timestamp 1649977179
transform 1 0 14628 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_157
timestamp 1649977179
transform 1 0 15548 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1649977179
transform 1 0 16100 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_175
timestamp 1649977179
transform 1 0 17204 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_192
timestamp 1649977179
transform 1 0 18768 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_203
timestamp 1649977179
transform 1 0 19780 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_208
timestamp 1649977179
transform 1 0 20240 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_215
timestamp 1649977179
transform 1 0 20884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1649977179
transform 1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_37
timestamp 1649977179
transform 1 0 4508 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_45
timestamp 1649977179
transform 1 0 5244 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_62
timestamp 1649977179
transform 1 0 6808 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_73
timestamp 1649977179
transform 1 0 7820 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_94
timestamp 1649977179
transform 1 0 9752 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_113
timestamp 1649977179
transform 1 0 11500 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1649977179
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_157
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_168
timestamp 1649977179
transform 1 0 16560 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_172
timestamp 1649977179
transform 1 0 16928 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_184
timestamp 1649977179
transform 1 0 18032 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_205
timestamp 1649977179
transform 1 0 19964 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1649977179
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_23_42
timestamp 1649977179
transform 1 0 4968 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_46
timestamp 1649977179
transform 1 0 5336 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_73
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_83
timestamp 1649977179
transform 1 0 8740 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_89
timestamp 1649977179
transform 1 0 9292 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_121
timestamp 1649977179
transform 1 0 12236 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_132
timestamp 1649977179
transform 1 0 13248 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_140
timestamp 1649977179
transform 1 0 13984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_23_150
timestamp 1649977179
transform 1 0 14904 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_23_159
timestamp 1649977179
transform 1 0 15732 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_209
timestamp 1649977179
transform 1 0 20332 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_215
timestamp 1649977179
transform 1 0 20884 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1649977179
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_11
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_20
timestamp 1649977179
transform 1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_38
timestamp 1649977179
transform 1 0 4600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_43
timestamp 1649977179
transform 1 0 5060 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_70
timestamp 1649977179
transform 1 0 7544 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_80
timestamp 1649977179
transform 1 0 8464 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_117
timestamp 1649977179
transform 1 0 11868 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_129
timestamp 1649977179
transform 1 0 12972 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_137
timestamp 1649977179
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_164
timestamp 1649977179
transform 1 0 16192 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_176
timestamp 1649977179
transform 1 0 17296 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1649977179
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_201
timestamp 1649977179
transform 1 0 19596 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_205
timestamp 1649977179
transform 1 0 19964 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1649977179
transform 1 0 20424 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1649977179
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_23
timestamp 1649977179
transform 1 0 3220 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_33
timestamp 1649977179
transform 1 0 4140 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_45
timestamp 1649977179
transform 1 0 5244 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1649977179
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_68
timestamp 1649977179
transform 1 0 7360 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_72
timestamp 1649977179
transform 1 0 7728 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_89
timestamp 1649977179
transform 1 0 9292 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1649977179
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_127
timestamp 1649977179
transform 1 0 12788 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_135
timestamp 1649977179
transform 1 0 13524 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_145
timestamp 1649977179
transform 1 0 14444 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_185
timestamp 1649977179
transform 1 0 18124 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_197
timestamp 1649977179
transform 1 0 19228 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_202
timestamp 1649977179
transform 1 0 19688 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_207
timestamp 1649977179
transform 1 0 20148 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_211
timestamp 1649977179
transform 1 0 20516 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1649977179
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1649977179
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_32
timestamp 1649977179
transform 1 0 4048 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_36
timestamp 1649977179
transform 1 0 4416 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_63
timestamp 1649977179
transform 1 0 6900 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_71
timestamp 1649977179
transform 1 0 7636 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_96
timestamp 1649977179
transform 1 0 9936 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_101
timestamp 1649977179
transform 1 0 10396 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_120
timestamp 1649977179
transform 1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1649977179
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_157
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_176
timestamp 1649977179
transform 1 0 17296 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_180
timestamp 1649977179
transform 1 0 17664 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1649977179
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_200
timestamp 1649977179
transform 1 0 19504 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_205
timestamp 1649977179
transform 1 0 19964 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1649977179
transform 1 0 20424 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1649977179
transform 1 0 20884 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_21
timestamp 1649977179
transform 1 0 3036 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_32
timestamp 1649977179
transform 1 0 4048 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_27_36
timestamp 1649977179
transform 1 0 4416 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_27_50
timestamp 1649977179
transform 1 0 5704 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_84
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_96
timestamp 1649977179
transform 1 0 9936 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_101
timestamp 1649977179
transform 1 0 10396 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_121
timestamp 1649977179
transform 1 0 12236 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_131
timestamp 1649977179
transform 1 0 13156 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_136
timestamp 1649977179
transform 1 0 13616 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_148
timestamp 1649977179
transform 1 0 14720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_159
timestamp 1649977179
transform 1 0 15732 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_164
timestamp 1649977179
transform 1 0 16192 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_177
timestamp 1649977179
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_182
timestamp 1649977179
transform 1 0 17848 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_192
timestamp 1649977179
transform 1 0 18768 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_197
timestamp 1649977179
transform 1 0 19228 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_202
timestamp 1649977179
transform 1 0 19688 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_207
timestamp 1649977179
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_212
timestamp 1649977179
transform 1 0 20608 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_216
timestamp 1649977179
transform 1 0 20976 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1649977179
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_14
timestamp 1649977179
transform 1 0 2392 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_18
timestamp 1649977179
transform 1 0 2760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_25
timestamp 1649977179
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_57
timestamp 1649977179
transform 1 0 6348 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_74
timestamp 1649977179
transform 1 0 7912 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_78
timestamp 1649977179
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_101
timestamp 1649977179
transform 1 0 10396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_122
timestamp 1649977179
transform 1 0 12328 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_126
timestamp 1649977179
transform 1 0 12696 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1649977179
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_147
timestamp 1649977179
transform 1 0 14628 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_150
timestamp 1649977179
transform 1 0 14904 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_162
timestamp 1649977179
transform 1 0 16008 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp 1649977179
transform 1 0 16560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_179
timestamp 1649977179
transform 1 0 17572 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_184
timestamp 1649977179
transform 1 0 18032 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1649977179
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_200
timestamp 1649977179
transform 1 0 19504 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_205
timestamp 1649977179
transform 1 0 19964 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1649977179
transform 1 0 20884 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_11
timestamp 1649977179
transform 1 0 2116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_18
timestamp 1649977179
transform 1 0 2760 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_23
timestamp 1649977179
transform 1 0 3220 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_35
timestamp 1649977179
transform 1 0 4324 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_43
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_67
timestamp 1649977179
transform 1 0 7268 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_72
timestamp 1649977179
transform 1 0 7728 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_92
timestamp 1649977179
transform 1 0 9568 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_96
timestamp 1649977179
transform 1 0 9936 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_99
timestamp 1649977179
transform 1 0 10212 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1649977179
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_121
timestamp 1649977179
transform 1 0 12236 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_127
timestamp 1649977179
transform 1 0 12788 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_139
timestamp 1649977179
transform 1 0 13892 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_151
timestamp 1649977179
transform 1 0 14996 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_156
timestamp 1649977179
transform 1 0 15456 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_162
timestamp 1649977179
transform 1 0 16008 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_188
timestamp 1649977179
transform 1 0 18400 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_199
timestamp 1649977179
transform 1 0 19412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_203
timestamp 1649977179
transform 1 0 19780 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_209
timestamp 1649977179
transform 1 0 20332 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1649977179
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_8
timestamp 1649977179
transform 1 0 1840 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1649977179
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_37
timestamp 1649977179
transform 1 0 4508 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_43
timestamp 1649977179
transform 1 0 5060 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_47
timestamp 1649977179
transform 1 0 5428 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_51
timestamp 1649977179
transform 1 0 5796 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_56
timestamp 1649977179
transform 1 0 6256 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_61
timestamp 1649977179
transform 1 0 6716 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_66
timestamp 1649977179
transform 1 0 7176 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_70
timestamp 1649977179
transform 1 0 7544 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_74
timestamp 1649977179
transform 1 0 7912 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_78
timestamp 1649977179
transform 1 0 8280 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1649977179
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_89
timestamp 1649977179
transform 1 0 9292 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_107
timestamp 1649977179
transform 1 0 10948 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_112
timestamp 1649977179
transform 1 0 11408 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_125
timestamp 1649977179
transform 1 0 12604 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_144
timestamp 1649977179
transform 1 0 14352 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_148
timestamp 1649977179
transform 1 0 14720 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1649977179
transform 1 0 15088 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_156
timestamp 1649977179
transform 1 0 15456 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_174
timestamp 1649977179
transform 1 0 17112 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_184
timestamp 1649977179
transform 1 0 18032 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1649977179
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_203
timestamp 1649977179
transform 1 0 19780 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1649977179
transform 1 0 20884 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_8
timestamp 1649977179
transform 1 0 1840 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_13
timestamp 1649977179
transform 1 0 2300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_19
timestamp 1649977179
transform 1 0 2852 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_23
timestamp 1649977179
transform 1 0 3220 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_41
timestamp 1649977179
transform 1 0 4876 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1649977179
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_65
timestamp 1649977179
transform 1 0 7084 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_70
timestamp 1649977179
transform 1 0 7544 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_76
timestamp 1649977179
transform 1 0 8096 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_87
timestamp 1649977179
transform 1 0 9108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_98
timestamp 1649977179
transform 1 0 10120 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1649977179
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_131
timestamp 1649977179
transform 1 0 13156 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_159
timestamp 1649977179
transform 1 0 15732 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1649977179
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_177
timestamp 1649977179
transform 1 0 17388 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_182
timestamp 1649977179
transform 1 0 17848 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_186
timestamp 1649977179
transform 1 0 18216 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_191
timestamp 1649977179
transform 1 0 18676 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1649977179
transform 1 0 19228 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1649977179
transform 1 0 19780 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_215
timestamp 1649977179
transform 1 0 20884 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_12
timestamp 1649977179
transform 1 0 2208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_19
timestamp 1649977179
transform 1 0 2852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1649977179
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_40
timestamp 1649977179
transform 1 0 4784 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_58
timestamp 1649977179
transform 1 0 6440 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_76
timestamp 1649977179
transform 1 0 8096 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1649977179
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_94
timestamp 1649977179
transform 1 0 9752 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_98
timestamp 1649977179
transform 1 0 10120 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_101
timestamp 1649977179
transform 1 0 10396 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_119
timestamp 1649977179
transform 1 0 12052 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_125
timestamp 1649977179
transform 1 0 12604 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_129
timestamp 1649977179
transform 1 0 12972 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1649977179
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_145
timestamp 1649977179
transform 1 0 14444 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_164
timestamp 1649977179
transform 1 0 16192 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_175
timestamp 1649977179
transform 1 0 17204 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_180
timestamp 1649977179
transform 1 0 17664 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1649977179
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_201
timestamp 1649977179
transform 1 0 19596 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_207
timestamp 1649977179
transform 1 0 20148 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1649977179
transform 1 0 20884 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_9
timestamp 1649977179
transform 1 0 1932 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_16
timestamp 1649977179
transform 1 0 2576 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_21
timestamp 1649977179
transform 1 0 3036 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_26
timestamp 1649977179
transform 1 0 3496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_33
timestamp 1649977179
transform 1 0 4140 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_38
timestamp 1649977179
transform 1 0 4600 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_48
timestamp 1649977179
transform 1 0 5520 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1649977179
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_62
timestamp 1649977179
transform 1 0 6808 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_67
timestamp 1649977179
transform 1 0 7268 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_72
timestamp 1649977179
transform 1 0 7728 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_82
timestamp 1649977179
transform 1 0 8648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_87
timestamp 1649977179
transform 1 0 9108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_92
timestamp 1649977179
transform 1 0 9568 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_98
timestamp 1649977179
transform 1 0 10120 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_104
timestamp 1649977179
transform 1 0 10672 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1649977179
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_116
timestamp 1649977179
transform 1 0 11776 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_126
timestamp 1649977179
transform 1 0 12696 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_132
timestamp 1649977179
transform 1 0 13248 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_138
timestamp 1649977179
transform 1 0 13800 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_143
timestamp 1649977179
transform 1 0 14260 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_154
timestamp 1649977179
transform 1 0 15272 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_160
timestamp 1649977179
transform 1 0 15824 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_166
timestamp 1649977179
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_173
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1649977179
transform 1 0 17572 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_185
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1649977179
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_195
timestamp 1649977179
transform 1 0 19044 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_201
timestamp 1649977179
transform 1 0 19596 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_207
timestamp 1649977179
transform 1 0 20148 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_213
timestamp 1649977179
transform 1 0 20700 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_219
timestamp 1649977179
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _48_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21068 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1649977179
transform -1 0 20608 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1649977179
transform -1 0 20608 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1649977179
transform -1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1649977179
transform -1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1649977179
transform -1 0 20424 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1649977179
transform -1 0 20884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1649977179
transform -1 0 18952 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1649977179
transform -1 0 19964 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1649977179
transform -1 0 20148 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1649977179
transform -1 0 18492 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1649977179
transform -1 0 19964 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1649977179
transform -1 0 20884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1649977179
transform -1 0 20424 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1649977179
transform 1 0 20608 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1649977179
transform -1 0 16192 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1649977179
transform 1 0 19688 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform 1 0 18952 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform -1 0 18032 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform -1 0 19504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform -1 0 11868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _69_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21160 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform -1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform 1 0 20700 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform 1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform 1 0 20332 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1649977179
transform 1 0 20792 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1649977179
transform 1 0 20332 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1649977179
transform 1 0 20792 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp 1649977179
transform 1 0 20976 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp 1649977179
transform 1 0 20792 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp 1649977179
transform 1 0 19688 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1649977179
transform 1 0 20792 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1649977179
transform 1 0 20332 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _83_
timestamp 1649977179
transform 1 0 20792 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _84_
timestamp 1649977179
transform -1 0 20608 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _85_
timestamp 1649977179
transform 1 0 20792 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _86_
timestamp 1649977179
transform 1 0 20792 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _87_
timestamp 1649977179
transform 1 0 20700 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_right_track_0.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12144 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_mem_right_track_0.prog_clk
timestamp 1649977179
transform -1 0 9660 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_mem_right_track_0.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_mem_right_track_0.prog_clk
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_mem_right_track_0.prog_clk
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9200 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1649977179
transform 1 0 10488 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1649977179
transform -1 0 4508 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1649977179
transform 1 0 7728 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1649977179
transform 1 0 12052 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1649977179
transform -1 0 12696 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1649977179
transform 1 0 17296 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1649977179
transform 1 0 10304 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1649977179
transform 1 0 14996 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1649977179
transform -1 0 7452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1649977179
transform 1 0 13064 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1649977179
transform 1 0 15456 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1649977179
transform 1 0 17112 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1649977179
transform -1 0 18768 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1649977179
transform 1 0 15456 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1649977179
transform -1 0 4508 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1649977179
transform -1 0 17388 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1649977179
transform 1 0 6164 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1649977179
transform -1 0 4140 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1649977179
transform -1 0 7084 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1649977179
transform 1 0 13064 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1649977179
transform -1 0 11868 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1649977179
transform -1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1649977179
transform 1 0 9384 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1649977179
transform 1 0 20516 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1649977179
transform -1 0 12788 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1649977179
transform 1 0 7912 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1649977179
transform -1 0 5520 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1649977179
transform -1 0 15548 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1649977179
transform -1 0 2944 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1649977179
transform -1 0 12604 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1649977179
transform 1 0 1656 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1649977179
transform -1 0 8740 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1649977179
transform -1 0 14904 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1649977179
transform -1 0 5704 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 20976 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 20792 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 21160 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 19136 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 20148 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 20608 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform 1 0 21160 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 20148 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 19688 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform 1 0 20240 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 20516 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform 1 0 21160 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 20148 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform 1 0 21160 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 20424 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform 1 0 20792 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 2208 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 7544 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 6072 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 6808 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform -1 0 7268 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 7728 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 9568 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 10120 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform -1 0 10672 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform -1 0 11224 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform -1 0 11776 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 2300 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 2852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 2576 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 3496 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 3036 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform -1 0 3496 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 4140 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform -1 0 4600 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20516 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1649977179
transform -1 0 21436 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1649977179
transform 1 0 20516 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1649977179
transform -1 0 21436 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1649977179
transform -1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1649977179
transform -1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1649977179
transform -1 0 20332 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform -1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform -1 0 20332 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1649977179
transform 1 0 1564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18584 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16100 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14628 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13248 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11592 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9384 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11500 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12052 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11500 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7636 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5152 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3588 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3036 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2024 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 3404 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4508 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7820 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9752 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10672 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12328 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14904 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17480 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17296 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7360 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 5336 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6348 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4968 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6624 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8096 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9476 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10580 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11684 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 13340 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14720 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15640 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16928 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8004 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9752 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11684 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15732 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18216 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18768 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17112 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17296 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 18676 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_0.mux_l2_in_1__106 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18308 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17664 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20148 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13800 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 14536 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15732 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_2.mux_l2_in_1__112
timestamp 1649977179
transform -1 0 15548 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14996 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14352 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9384 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9200 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_4.mux_l2_in_1__99
timestamp 1649977179
transform 1 0 11592 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 11408 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11868 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13156 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13156 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13248 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_6.mux_l2_in_1__100
timestamp 1649977179
transform -1 0 15732 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15732 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_8.mux_l1_in_1__101
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9752 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9660 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4140 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_10.mux_l2_in_0__107
timestamp 1649977179
transform 1 0 4784 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20332 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3220 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_12.mux_l2_in_0__108
timestamp 1649977179
transform 1 0 3128 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 3496 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4784 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5060 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_14.mux_l2_in_0__109
timestamp 1649977179
transform -1 0 5060 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5060 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_16.mux_l2_in_0__110
timestamp 1649977179
transform 1 0 10120 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9936 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10396 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_18.mux_l2_in_0__111
timestamp 1649977179
transform 1 0 13340 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13156 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20332 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14720 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_20.mux_l2_in_0__113
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15732 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19412 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17296 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_22.mux_l2_in_0__114
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18768 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19688 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18584 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_24.mux_l1_in_1__115
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 19780 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20332 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6992 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7360 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_26.mux_l2_in_0__116
timestamp 1649977179
transform 1 0 7268 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20148 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_28.mux_l2_in_0__93
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7268 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7176 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9108 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_30.mux_l2_in_0__94
timestamp 1649977179
transform -1 0 8648 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18676 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10120 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_32.mux_l2_in_0__95
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18492 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12604 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_34.mux_l2_in_0__96
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13800 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17848 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15272 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_36.mux_l2_in_0__97
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16376 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15456 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17572 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18584 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_38.mux_l2_in_0__98
timestamp 1649977179
transform -1 0 17848 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16376 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11960 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_0.mux_l2_in_0__102
timestamp 1649977179
transform 1 0 12420 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11224 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14996 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_4.mux_l2_in_0__104
timestamp 1649977179
transform 1 0 14444 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13984 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17940 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_8.mux_l2_in_0__105
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16928 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19504 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_24.mux_l2_in_0__103
timestamp 1649977179
transform 1 0 20332 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19320 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output52 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform 1 0 21068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform 1 0 21068 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform 1 0 20516 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform -1 0 20332 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform 1 0 19964 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform -1 0 19780 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform 1 0 20516 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 21068 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform 1 0 21068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 20516 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 20148 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform -1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 20148 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 20884 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 20884 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 19780 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform -1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 13248 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform 1 0 13432 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 14444 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform -1 0 15824 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform -1 0 16376 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform -1 0 17020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18952 0 1 19584
box -38 -48 1142 592
<< labels >>
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 0 nsew ground input
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 0 nsew ground input
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 0 nsew ground input
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 1 nsew power input
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 1 nsew power input
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 1 nsew power input
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 1 nsew power input
rlabel metal3 s 0 5720 800 5840 6 ccff_head
port 2 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 ccff_tail
port 3 nsew signal tristate
rlabel metal3 s 22200 4224 23000 4344 6 chanx_right_in[0]
port 4 nsew signal input
rlabel metal3 s 22200 8848 23000 8968 6 chanx_right_in[10]
port 5 nsew signal input
rlabel metal3 s 22200 9256 23000 9376 6 chanx_right_in[11]
port 6 nsew signal input
rlabel metal3 s 22200 9664 23000 9784 6 chanx_right_in[12]
port 7 nsew signal input
rlabel metal3 s 22200 10208 23000 10328 6 chanx_right_in[13]
port 8 nsew signal input
rlabel metal3 s 22200 10616 23000 10736 6 chanx_right_in[14]
port 9 nsew signal input
rlabel metal3 s 22200 11160 23000 11280 6 chanx_right_in[15]
port 10 nsew signal input
rlabel metal3 s 22200 11568 23000 11688 6 chanx_right_in[16]
port 11 nsew signal input
rlabel metal3 s 22200 11976 23000 12096 6 chanx_right_in[17]
port 12 nsew signal input
rlabel metal3 s 22200 12520 23000 12640 6 chanx_right_in[18]
port 13 nsew signal input
rlabel metal3 s 22200 12928 23000 13048 6 chanx_right_in[19]
port 14 nsew signal input
rlabel metal3 s 22200 4632 23000 4752 6 chanx_right_in[1]
port 15 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[2]
port 16 nsew signal input
rlabel metal3 s 22200 5584 23000 5704 6 chanx_right_in[3]
port 17 nsew signal input
rlabel metal3 s 22200 5992 23000 6112 6 chanx_right_in[4]
port 18 nsew signal input
rlabel metal3 s 22200 6536 23000 6656 6 chanx_right_in[5]
port 19 nsew signal input
rlabel metal3 s 22200 6944 23000 7064 6 chanx_right_in[6]
port 20 nsew signal input
rlabel metal3 s 22200 7488 23000 7608 6 chanx_right_in[7]
port 21 nsew signal input
rlabel metal3 s 22200 7896 23000 8016 6 chanx_right_in[8]
port 22 nsew signal input
rlabel metal3 s 22200 8304 23000 8424 6 chanx_right_in[9]
port 23 nsew signal input
rlabel metal3 s 22200 13472 23000 13592 6 chanx_right_out[0]
port 24 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[10]
port 25 nsew signal tristate
rlabel metal3 s 22200 18504 23000 18624 6 chanx_right_out[11]
port 26 nsew signal tristate
rlabel metal3 s 22200 18912 23000 19032 6 chanx_right_out[12]
port 27 nsew signal tristate
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[13]
port 28 nsew signal tristate
rlabel metal3 s 22200 19864 23000 19984 6 chanx_right_out[14]
port 29 nsew signal tristate
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[15]
port 30 nsew signal tristate
rlabel metal3 s 22200 20816 23000 20936 6 chanx_right_out[16]
port 31 nsew signal tristate
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[17]
port 32 nsew signal tristate
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[18]
port 33 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 chanx_right_out[19]
port 34 nsew signal tristate
rlabel metal3 s 22200 13880 23000 14000 6 chanx_right_out[1]
port 35 nsew signal tristate
rlabel metal3 s 22200 14288 23000 14408 6 chanx_right_out[2]
port 36 nsew signal tristate
rlabel metal3 s 22200 14832 23000 14952 6 chanx_right_out[3]
port 37 nsew signal tristate
rlabel metal3 s 22200 15240 23000 15360 6 chanx_right_out[4]
port 38 nsew signal tristate
rlabel metal3 s 22200 15648 23000 15768 6 chanx_right_out[5]
port 39 nsew signal tristate
rlabel metal3 s 22200 16192 23000 16312 6 chanx_right_out[6]
port 40 nsew signal tristate
rlabel metal3 s 22200 16600 23000 16720 6 chanx_right_out[7]
port 41 nsew signal tristate
rlabel metal3 s 22200 17144 23000 17264 6 chanx_right_out[8]
port 42 nsew signal tristate
rlabel metal3 s 22200 17552 23000 17672 6 chanx_right_out[9]
port 43 nsew signal tristate
rlabel metal2 s 846 22200 902 23000 6 chany_top_in[0]
port 44 nsew signal input
rlabel metal2 s 6458 22200 6514 23000 6 chany_top_in[10]
port 45 nsew signal input
rlabel metal2 s 7010 22200 7066 23000 6 chany_top_in[11]
port 46 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[12]
port 47 nsew signal input
rlabel metal2 s 8114 22200 8170 23000 6 chany_top_in[13]
port 48 nsew signal input
rlabel metal2 s 8666 22200 8722 23000 6 chany_top_in[14]
port 49 nsew signal input
rlabel metal2 s 9218 22200 9274 23000 6 chany_top_in[15]
port 50 nsew signal input
rlabel metal2 s 9770 22200 9826 23000 6 chany_top_in[16]
port 51 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[17]
port 52 nsew signal input
rlabel metal2 s 10874 22200 10930 23000 6 chany_top_in[18]
port 53 nsew signal input
rlabel metal2 s 11426 22200 11482 23000 6 chany_top_in[19]
port 54 nsew signal input
rlabel metal2 s 1398 22200 1454 23000 6 chany_top_in[1]
port 55 nsew signal input
rlabel metal2 s 1950 22200 2006 23000 6 chany_top_in[2]
port 56 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 chany_top_in[3]
port 57 nsew signal input
rlabel metal2 s 3054 22200 3110 23000 6 chany_top_in[4]
port 58 nsew signal input
rlabel metal2 s 3606 22200 3662 23000 6 chany_top_in[5]
port 59 nsew signal input
rlabel metal2 s 4158 22200 4214 23000 6 chany_top_in[6]
port 60 nsew signal input
rlabel metal2 s 4710 22200 4766 23000 6 chany_top_in[7]
port 61 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[8]
port 62 nsew signal input
rlabel metal2 s 5814 22200 5870 23000 6 chany_top_in[9]
port 63 nsew signal input
rlabel metal2 s 12070 22200 12126 23000 6 chany_top_out[0]
port 64 nsew signal tristate
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 65 nsew signal tristate
rlabel metal2 s 18234 22200 18290 23000 6 chany_top_out[11]
port 66 nsew signal tristate
rlabel metal2 s 18786 22200 18842 23000 6 chany_top_out[12]
port 67 nsew signal tristate
rlabel metal2 s 19338 22200 19394 23000 6 chany_top_out[13]
port 68 nsew signal tristate
rlabel metal2 s 19890 22200 19946 23000 6 chany_top_out[14]
port 69 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[15]
port 70 nsew signal tristate
rlabel metal2 s 20994 22200 21050 23000 6 chany_top_out[16]
port 71 nsew signal tristate
rlabel metal2 s 21546 22200 21602 23000 6 chany_top_out[17]
port 72 nsew signal tristate
rlabel metal2 s 22098 22200 22154 23000 6 chany_top_out[18]
port 73 nsew signal tristate
rlabel metal2 s 22650 22200 22706 23000 6 chany_top_out[19]
port 74 nsew signal tristate
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_out[1]
port 75 nsew signal tristate
rlabel metal2 s 13174 22200 13230 23000 6 chany_top_out[2]
port 76 nsew signal tristate
rlabel metal2 s 13726 22200 13782 23000 6 chany_top_out[3]
port 77 nsew signal tristate
rlabel metal2 s 14278 22200 14334 23000 6 chany_top_out[4]
port 78 nsew signal tristate
rlabel metal2 s 14830 22200 14886 23000 6 chany_top_out[5]
port 79 nsew signal tristate
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[6]
port 80 nsew signal tristate
rlabel metal2 s 15934 22200 15990 23000 6 chany_top_out[7]
port 81 nsew signal tristate
rlabel metal2 s 16486 22200 16542 23000 6 chany_top_out[8]
port 82 nsew signal tristate
rlabel metal2 s 17038 22200 17094 23000 6 chany_top_out[9]
port 83 nsew signal tristate
rlabel metal3 s 22200 22584 23000 22704 6 prog_clk_0_E_in
port 84 nsew signal input
rlabel metal3 s 22200 2320 23000 2440 6 right_bottom_grid_pin_11_
port 85 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_13_
port 86 nsew signal input
rlabel metal3 s 22200 3272 23000 3392 6 right_bottom_grid_pin_15_
port 87 nsew signal input
rlabel metal3 s 22200 3816 23000 3936 6 right_bottom_grid_pin_17_
port 88 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_1_
port 89 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_3_
port 90 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_5_
port 91 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_7_
port 92 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_9_
port 93 nsew signal input
rlabel metal2 s 294 22200 350 23000 6 top_left_grid_pin_1_
port 94 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
