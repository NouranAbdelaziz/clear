magic
tech sky130A
magscale 1 2
timestamp 1650633435
<< viali >>
rect 5273 14025 5307 14059
rect 18061 14025 18095 14059
rect 18429 14025 18463 14059
rect 13093 13957 13127 13991
rect 14013 13957 14047 13991
rect 15577 13957 15611 13991
rect 16497 13957 16531 13991
rect 16865 13957 16899 13991
rect 4905 13889 4939 13923
rect 13277 13889 13311 13923
rect 13645 13889 13679 13923
rect 14105 13889 14139 13923
rect 17877 13889 17911 13923
rect 18245 13889 18279 13923
rect 4629 13821 4663 13855
rect 4813 13821 4847 13855
rect 6929 13821 6963 13855
rect 15485 13821 15519 13855
rect 16773 13821 16807 13855
rect 17049 13821 17083 13855
rect 6009 13685 6043 13719
rect 9781 13685 9815 13719
rect 14749 13685 14783 13719
rect 3893 13481 3927 13515
rect 5089 13481 5123 13515
rect 12541 13481 12575 13515
rect 16589 13481 16623 13515
rect 4261 13413 4295 13447
rect 6009 13413 6043 13447
rect 10517 13413 10551 13447
rect 15899 13413 15933 13447
rect 4445 13345 4479 13379
rect 5733 13345 5767 13379
rect 6561 13345 6595 13379
rect 9413 13345 9447 13379
rect 9597 13345 9631 13379
rect 11621 13345 11655 13379
rect 4721 13277 4755 13311
rect 6469 13277 6503 13311
rect 8401 13277 8435 13311
rect 9781 13277 9815 13311
rect 11345 13277 11379 13311
rect 13921 13277 13955 13311
rect 15209 13277 15243 13311
rect 15796 13277 15830 13311
rect 18061 13277 18095 13311
rect 4077 13209 4111 13243
rect 4629 13209 4663 13243
rect 5549 13209 5583 13243
rect 8134 13209 8168 13243
rect 8493 13209 8527 13243
rect 13676 13209 13710 13243
rect 16773 13209 16807 13243
rect 5181 13141 5215 13175
rect 5641 13141 5675 13175
rect 6377 13141 6411 13175
rect 6929 13141 6963 13175
rect 7021 13141 7055 13175
rect 8953 13141 8987 13175
rect 9321 13141 9355 13175
rect 10425 13141 10459 13175
rect 14565 13141 14599 13175
rect 17693 13141 17727 13175
rect 1593 12937 1627 12971
rect 2697 12937 2731 12971
rect 4353 12937 4387 12971
rect 4629 12937 4663 12971
rect 4997 12937 5031 12971
rect 5457 12937 5491 12971
rect 8493 12937 8527 12971
rect 13553 12937 13587 12971
rect 13737 12937 13771 12971
rect 18061 12937 18095 12971
rect 18429 12937 18463 12971
rect 10066 12869 10100 12903
rect 12440 12869 12474 12903
rect 14850 12869 14884 12903
rect 2513 12801 2547 12835
rect 3056 12801 3090 12835
rect 5825 12801 5859 12835
rect 7582 12801 7616 12835
rect 7849 12801 7883 12835
rect 8033 12801 8067 12835
rect 10425 12801 10459 12835
rect 15117 12801 15151 12835
rect 15761 12801 15795 12835
rect 17969 12801 18003 12835
rect 2789 12733 2823 12767
rect 5089 12733 5123 12767
rect 5181 12733 5215 12767
rect 5917 12733 5951 12767
rect 6009 12733 6043 12767
rect 8217 12733 8251 12767
rect 8401 12733 8435 12767
rect 10333 12733 10367 12767
rect 12173 12733 12207 12767
rect 15853 12733 15887 12767
rect 15945 12733 15979 12767
rect 18153 12733 18187 12767
rect 1869 12665 1903 12699
rect 6469 12665 6503 12699
rect 8953 12665 8987 12699
rect 1961 12597 1995 12631
rect 2145 12597 2179 12631
rect 4169 12597 4203 12631
rect 4537 12597 4571 12631
rect 8861 12597 8895 12631
rect 11069 12597 11103 12631
rect 15393 12597 15427 12631
rect 17325 12597 17359 12631
rect 17601 12597 17635 12631
rect 2329 12393 2363 12427
rect 5365 12393 5399 12427
rect 6193 12393 6227 12427
rect 8769 12393 8803 12427
rect 16037 12393 16071 12427
rect 5181 12325 5215 12359
rect 7113 12325 7147 12359
rect 10977 12325 11011 12359
rect 13921 12325 13955 12359
rect 15853 12325 15887 12359
rect 5917 12257 5951 12291
rect 6837 12257 6871 12291
rect 7389 12257 7423 12291
rect 9229 12257 9263 12291
rect 9873 12257 9907 12291
rect 10701 12257 10735 12291
rect 13369 12257 13403 12291
rect 14749 12257 14783 12291
rect 15393 12257 15427 12291
rect 15485 12257 15519 12291
rect 17693 12257 17727 12291
rect 1685 12189 1719 12223
rect 2973 12189 3007 12223
rect 3801 12189 3835 12223
rect 6561 12189 6595 12223
rect 7656 12189 7690 12223
rect 10517 12189 10551 12223
rect 12357 12189 12391 12223
rect 13461 12189 13495 12223
rect 14473 12189 14507 12223
rect 17417 12189 17451 12223
rect 17877 12189 17911 12223
rect 2421 12121 2455 12155
rect 2605 12121 2639 12155
rect 2881 12121 2915 12155
rect 4068 12121 4102 12155
rect 7205 12121 7239 12155
rect 9689 12121 9723 12155
rect 12090 12121 12124 12155
rect 13093 12121 13127 12155
rect 13553 12121 13587 12155
rect 17172 12121 17206 12155
rect 18337 12121 18371 12155
rect 1501 12053 1535 12087
rect 1777 12053 1811 12087
rect 1961 12053 1995 12087
rect 3617 12053 3651 12087
rect 5733 12053 5767 12087
rect 5825 12053 5859 12087
rect 6653 12053 6687 12087
rect 9321 12053 9355 12087
rect 9781 12053 9815 12087
rect 10149 12053 10183 12087
rect 10609 12053 10643 12087
rect 14105 12053 14139 12087
rect 14565 12053 14599 12087
rect 14933 12053 14967 12087
rect 15301 12053 15335 12087
rect 17785 12053 17819 12087
rect 18245 12053 18279 12087
rect 2513 11849 2547 11883
rect 6377 11849 6411 11883
rect 7205 11849 7239 11883
rect 8493 11849 8527 11883
rect 9413 11849 9447 11883
rect 9781 11849 9815 11883
rect 10241 11849 10275 11883
rect 10609 11849 10643 11883
rect 11897 11849 11931 11883
rect 12541 11849 12575 11883
rect 13737 11849 13771 11883
rect 14197 11849 14231 11883
rect 15209 11849 15243 11883
rect 15577 11849 15611 11883
rect 15669 11849 15703 11883
rect 16681 11849 16715 11883
rect 17509 11849 17543 11883
rect 3065 11781 3099 11815
rect 3525 11781 3559 11815
rect 3985 11781 4019 11815
rect 4344 11781 4378 11815
rect 6193 11781 6227 11815
rect 8585 11781 8619 11815
rect 10149 11781 10183 11815
rect 13645 11781 13679 11815
rect 16221 11781 16255 11815
rect 17141 11781 17175 11815
rect 1501 11713 1535 11747
rect 2973 11713 3007 11747
rect 5549 11713 5583 11747
rect 6745 11713 6779 11747
rect 7573 11713 7607 11747
rect 9321 11713 9355 11747
rect 10977 11713 11011 11747
rect 11989 11713 12023 11747
rect 14565 11713 14599 11747
rect 15025 11713 15059 11747
rect 16037 11713 16071 11747
rect 17049 11713 17083 11747
rect 17877 11713 17911 11747
rect 17969 11713 18003 11747
rect 18337 11713 18371 11747
rect 2145 11645 2179 11679
rect 3249 11645 3283 11679
rect 4077 11645 4111 11679
rect 6837 11645 6871 11679
rect 7021 11645 7055 11679
rect 7665 11645 7699 11679
rect 7757 11645 7791 11679
rect 8769 11645 8803 11679
rect 9597 11645 9631 11679
rect 10333 11645 10367 11679
rect 11069 11645 11103 11679
rect 11161 11645 11195 11679
rect 12081 11645 12115 11679
rect 13553 11645 13587 11679
rect 14657 11645 14691 11679
rect 14749 11645 14783 11679
rect 15761 11645 15795 11679
rect 17325 11645 17359 11679
rect 18061 11645 18095 11679
rect 8953 11577 8987 11611
rect 11529 11577 11563 11611
rect 16497 11577 16531 11611
rect 2237 11509 2271 11543
rect 2605 11509 2639 11543
rect 3801 11509 3835 11543
rect 5457 11509 5491 11543
rect 8125 11509 8159 11543
rect 12357 11509 12391 11543
rect 13001 11509 13035 11543
rect 13277 11509 13311 11543
rect 14105 11509 14139 11543
rect 6193 11305 6227 11339
rect 8769 11305 8803 11339
rect 9413 11305 9447 11339
rect 9597 11305 9631 11339
rect 11161 11305 11195 11339
rect 16313 11305 16347 11339
rect 18337 11305 18371 11339
rect 4169 11237 4203 11271
rect 7573 11237 7607 11271
rect 12357 11237 12391 11271
rect 13185 11237 13219 11271
rect 3801 11169 3835 11203
rect 6009 11169 6043 11203
rect 7205 11169 7239 11203
rect 8125 11169 8159 11203
rect 11805 11169 11839 11203
rect 12909 11169 12943 11203
rect 13645 11169 13679 11203
rect 13737 11169 13771 11203
rect 14933 11169 14967 11203
rect 2145 11101 2179 11135
rect 3617 11101 3651 11135
rect 5733 11101 5767 11135
rect 10977 11101 11011 11135
rect 11621 11101 11655 11135
rect 12725 11101 12759 11135
rect 14197 11101 14231 11135
rect 16405 11101 16439 11135
rect 18061 11101 18095 11135
rect 1501 11033 1535 11067
rect 3372 11033 3406 11067
rect 5466 11033 5500 11067
rect 6469 11033 6503 11067
rect 7021 11033 7055 11067
rect 7389 11033 7423 11067
rect 7941 11033 7975 11067
rect 8033 11033 8067 11067
rect 8401 11033 8435 11067
rect 9229 11033 9263 11067
rect 10710 11033 10744 11067
rect 12265 11033 12299 11067
rect 13553 11033 13587 11067
rect 15200 11033 15234 11067
rect 17816 11033 17850 11067
rect 2237 10965 2271 10999
rect 4353 10965 4387 10999
rect 6561 10965 6595 10999
rect 6929 10965 6963 10999
rect 9045 10965 9079 10999
rect 11529 10965 11563 10999
rect 11989 10965 12023 10999
rect 12817 10965 12851 10999
rect 14841 10965 14875 10999
rect 16681 10965 16715 10999
rect 18153 10965 18187 10999
rect 3249 10761 3283 10795
rect 4353 10761 4387 10795
rect 4721 10761 4755 10795
rect 5181 10761 5215 10795
rect 6653 10761 6687 10795
rect 7113 10761 7147 10795
rect 8585 10761 8619 10795
rect 10793 10761 10827 10795
rect 16681 10761 16715 10795
rect 17969 10761 18003 10795
rect 18337 10761 18371 10795
rect 2522 10693 2556 10727
rect 5089 10693 5123 10727
rect 11069 10693 11103 10727
rect 17141 10693 17175 10727
rect 4261 10625 4295 10659
rect 6193 10625 6227 10659
rect 6745 10625 6779 10659
rect 7205 10625 7239 10659
rect 7472 10625 7506 10659
rect 8677 10625 8711 10659
rect 8944 10625 8978 10659
rect 10149 10625 10183 10659
rect 11161 10625 11195 10659
rect 11529 10625 11563 10659
rect 11785 10625 11819 10659
rect 13001 10625 13035 10659
rect 13257 10625 13291 10659
rect 15597 10625 15631 10659
rect 15853 10625 15887 10659
rect 17049 10625 17083 10659
rect 17877 10625 17911 10659
rect 2789 10557 2823 10591
rect 3341 10557 3375 10591
rect 3525 10557 3559 10591
rect 4445 10557 4479 10591
rect 5273 10557 5307 10591
rect 6561 10557 6595 10591
rect 17233 10557 17267 10591
rect 18061 10557 18095 10591
rect 3801 10489 3835 10523
rect 1409 10421 1443 10455
rect 2881 10421 2915 10455
rect 3893 10421 3927 10455
rect 5549 10421 5583 10455
rect 10057 10421 10091 10455
rect 12909 10421 12943 10455
rect 14381 10421 14415 10455
rect 14473 10421 14507 10455
rect 15945 10421 15979 10455
rect 16405 10421 16439 10455
rect 17509 10421 17543 10455
rect 1593 10217 1627 10251
rect 4077 10217 4111 10251
rect 6745 10217 6779 10251
rect 7665 10217 7699 10251
rect 9413 10217 9447 10251
rect 13093 10217 13127 10251
rect 1777 10149 1811 10183
rect 7573 10149 7607 10183
rect 9321 10149 9355 10183
rect 15485 10149 15519 10183
rect 18061 10149 18095 10183
rect 2605 10081 2639 10115
rect 3341 10081 3375 10115
rect 3525 10081 3559 10115
rect 3801 10081 3835 10115
rect 4997 10081 5031 10115
rect 7389 10081 7423 10115
rect 8217 10081 8251 10115
rect 10241 10081 10275 10115
rect 12173 10081 12207 10115
rect 12449 10081 12483 10115
rect 13737 10081 13771 10115
rect 16129 10081 16163 10115
rect 16957 10081 16991 10115
rect 17877 10081 17911 10115
rect 1961 10013 1995 10047
rect 2421 10013 2455 10047
rect 4261 10013 4295 10047
rect 4905 10013 4939 10047
rect 5273 10013 5307 10047
rect 7113 10013 7147 10047
rect 10425 10013 10459 10047
rect 12633 10013 12667 10047
rect 14105 10013 14139 10047
rect 15945 10013 15979 10047
rect 17601 10013 17635 10047
rect 18245 10013 18279 10047
rect 3249 9945 3283 9979
rect 4813 9945 4847 9979
rect 8033 9945 8067 9979
rect 9965 9945 9999 9979
rect 14372 9945 14406 9979
rect 16773 9945 16807 9979
rect 17693 9945 17727 9979
rect 18521 9945 18555 9979
rect 2053 9877 2087 9911
rect 2513 9877 2547 9911
rect 2881 9877 2915 9911
rect 4445 9877 4479 9911
rect 8125 9877 8159 9911
rect 8585 9877 8619 9911
rect 8769 9877 8803 9911
rect 9045 9877 9079 9911
rect 9597 9877 9631 9911
rect 10057 9877 10091 9911
rect 12541 9877 12575 9911
rect 13001 9877 13035 9911
rect 13461 9877 13495 9911
rect 13553 9877 13587 9911
rect 15577 9877 15611 9911
rect 16037 9877 16071 9911
rect 16405 9877 16439 9911
rect 16865 9877 16899 9911
rect 17233 9877 17267 9911
rect 3341 9673 3375 9707
rect 5365 9673 5399 9707
rect 7757 9673 7791 9707
rect 8401 9673 8435 9707
rect 11253 9673 11287 9707
rect 18245 9673 18279 9707
rect 4997 9605 5031 9639
rect 15516 9605 15550 9639
rect 16497 9605 16531 9639
rect 18337 9605 18371 9639
rect 1869 9537 1903 9571
rect 1961 9537 1995 9571
rect 2228 9537 2262 9571
rect 3433 9537 3467 9571
rect 3689 9537 3723 9571
rect 5825 9537 5859 9571
rect 6377 9537 6411 9571
rect 6644 9537 6678 9571
rect 9229 9537 9263 9571
rect 10802 9537 10836 9571
rect 11069 9537 11103 9571
rect 12173 9537 12207 9571
rect 13001 9537 13035 9571
rect 13829 9537 13863 9571
rect 15761 9537 15795 9571
rect 15853 9537 15887 9571
rect 17132 9537 17166 9571
rect 5641 9469 5675 9503
rect 5733 9469 5767 9503
rect 8493 9469 8527 9503
rect 8677 9469 8711 9503
rect 9045 9469 9079 9503
rect 9137 9469 9171 9503
rect 11897 9469 11931 9503
rect 12081 9469 12115 9503
rect 13093 9469 13127 9503
rect 13277 9469 13311 9503
rect 13921 9469 13955 9503
rect 14013 9469 14047 9503
rect 16865 9469 16899 9503
rect 12633 9401 12667 9435
rect 13461 9401 13495 9435
rect 1409 9333 1443 9367
rect 1685 9333 1719 9367
rect 4813 9333 4847 9367
rect 5181 9333 5215 9367
rect 6193 9333 6227 9367
rect 7849 9333 7883 9367
rect 8033 9333 8067 9367
rect 9597 9333 9631 9367
rect 9689 9333 9723 9367
rect 11621 9333 11655 9367
rect 12541 9333 12575 9367
rect 14381 9333 14415 9367
rect 16681 9333 16715 9367
rect 4353 9129 4387 9163
rect 6561 9129 6595 9163
rect 10425 9129 10459 9163
rect 12265 9129 12299 9163
rect 14105 9129 14139 9163
rect 17601 9129 17635 9163
rect 6653 9061 6687 9095
rect 9045 9061 9079 9095
rect 12357 9061 12391 9095
rect 15761 9061 15795 9095
rect 2513 8993 2547 9027
rect 2605 8993 2639 9027
rect 2973 8993 3007 9027
rect 3157 8993 3191 9027
rect 4997 8993 5031 9027
rect 5181 8993 5215 9027
rect 10057 8993 10091 9027
rect 10241 8993 10275 9027
rect 10977 8993 11011 9027
rect 11713 8993 11747 9027
rect 14565 8993 14599 9027
rect 14657 8993 14691 9027
rect 15577 8993 15611 9027
rect 18153 8993 18187 9027
rect 1961 8925 1995 8959
rect 2421 8925 2455 8959
rect 3249 8925 3283 8959
rect 4077 8925 4111 8959
rect 5448 8925 5482 8959
rect 8033 8925 8067 8959
rect 8125 8925 8159 8959
rect 9965 8925 9999 8959
rect 13737 8925 13771 8959
rect 16129 8925 16163 8959
rect 17969 8925 18003 8959
rect 18429 8925 18463 8959
rect 1685 8857 1719 8891
rect 4721 8857 4755 8891
rect 7788 8857 7822 8891
rect 8769 8857 8803 8891
rect 10885 8857 10919 8891
rect 11805 8857 11839 8891
rect 13492 8857 13526 8891
rect 15301 8857 15335 8891
rect 16396 8857 16430 8891
rect 2053 8789 2087 8823
rect 3617 8789 3651 8823
rect 3893 8789 3927 8823
rect 4169 8789 4203 8823
rect 4813 8789 4847 8823
rect 9229 8789 9263 8823
rect 9413 8789 9447 8823
rect 9597 8789 9631 8823
rect 10793 8789 10827 8823
rect 11253 8789 11287 8823
rect 11897 8789 11931 8823
rect 13829 8789 13863 8823
rect 14473 8789 14507 8823
rect 14933 8789 14967 8823
rect 15393 8789 15427 8823
rect 15945 8789 15979 8823
rect 17509 8789 17543 8823
rect 18061 8789 18095 8823
rect 2973 8585 3007 8619
rect 3433 8585 3467 8619
rect 4813 8585 4847 8619
rect 6653 8585 6687 8619
rect 7113 8585 7147 8619
rect 8125 8585 8159 8619
rect 10885 8585 10919 8619
rect 12909 8585 12943 8619
rect 13737 8585 13771 8619
rect 14105 8585 14139 8619
rect 14657 8585 14691 8619
rect 15117 8585 15151 8619
rect 15485 8585 15519 8619
rect 15853 8585 15887 8619
rect 16405 8585 16439 8619
rect 3341 8517 3375 8551
rect 4169 8517 4203 8551
rect 9597 8517 9631 8551
rect 13277 8517 13311 8551
rect 14197 8517 14231 8551
rect 16926 8517 16960 8551
rect 2533 8449 2567 8483
rect 5926 8449 5960 8483
rect 6193 8449 6227 8483
rect 7021 8449 7055 8483
rect 9249 8449 9283 8483
rect 11796 8449 11830 8483
rect 13369 8449 13403 8483
rect 15025 8449 15059 8483
rect 15945 8449 15979 8483
rect 16681 8449 16715 8483
rect 18153 8449 18187 8483
rect 2789 8381 2823 8415
rect 3617 8381 3651 8415
rect 4261 8381 4295 8415
rect 4353 8381 4387 8415
rect 7297 8381 7331 8415
rect 7849 8381 7883 8415
rect 9505 8381 9539 8415
rect 11529 8381 11563 8415
rect 13093 8381 13127 8415
rect 14013 8381 14047 8415
rect 15301 8381 15335 8415
rect 16129 8381 16163 8415
rect 1409 8313 1443 8347
rect 6469 8313 6503 8347
rect 7573 8313 7607 8347
rect 8033 8313 8067 8347
rect 18061 8313 18095 8347
rect 18337 8313 18371 8347
rect 3801 8245 3835 8279
rect 4721 8245 4755 8279
rect 14565 8245 14599 8279
rect 4169 8041 4203 8075
rect 11069 8041 11103 8075
rect 12541 8041 12575 8075
rect 12909 8041 12943 8075
rect 16957 8041 16991 8075
rect 18245 8041 18279 8075
rect 1961 7973 1995 8007
rect 4997 7973 5031 8007
rect 9137 7973 9171 8007
rect 10149 7973 10183 8007
rect 13001 7973 13035 8007
rect 15485 7973 15519 8007
rect 2421 7905 2455 7939
rect 2513 7905 2547 7939
rect 3525 7905 3559 7939
rect 4813 7905 4847 7939
rect 7757 7905 7791 7939
rect 8401 7905 8435 7939
rect 8585 7905 8619 7939
rect 9505 7905 9539 7939
rect 9689 7905 9723 7939
rect 10333 7905 10367 7939
rect 11529 7905 11563 7939
rect 11713 7905 11747 7939
rect 13369 7905 13403 7939
rect 14289 7905 14323 7939
rect 14381 7905 14415 7939
rect 17601 7905 17635 7939
rect 17785 7905 17819 7939
rect 18337 7905 18371 7939
rect 1869 7837 1903 7871
rect 2329 7837 2363 7871
rect 4077 7837 4111 7871
rect 4537 7837 4571 7871
rect 6377 7837 6411 7871
rect 6745 7837 6779 7871
rect 7481 7837 7515 7871
rect 9781 7837 9815 7871
rect 10609 7837 10643 7871
rect 11897 7837 11931 7871
rect 1593 7769 1627 7803
rect 3249 7769 3283 7803
rect 6110 7769 6144 7803
rect 6837 7769 6871 7803
rect 8309 7769 8343 7803
rect 11437 7769 11471 7803
rect 13553 7769 13587 7803
rect 14933 7769 14967 7803
rect 15669 7769 15703 7803
rect 17877 7769 17911 7803
rect 2881 7701 2915 7735
rect 3341 7701 3375 7735
rect 3893 7701 3927 7735
rect 4629 7701 4663 7735
rect 6561 7701 6595 7735
rect 7113 7701 7147 7735
rect 7573 7701 7607 7735
rect 7941 7701 7975 7735
rect 9321 7701 9355 7735
rect 10517 7701 10551 7735
rect 10977 7701 11011 7735
rect 12725 7701 12759 7735
rect 13461 7701 13495 7735
rect 13921 7701 13955 7735
rect 14473 7701 14507 7735
rect 14841 7701 14875 7735
rect 15301 7701 15335 7735
rect 1501 7497 1535 7531
rect 4997 7497 5031 7531
rect 6929 7497 6963 7531
rect 8493 7497 8527 7531
rect 11897 7497 11931 7531
rect 12357 7497 12391 7531
rect 12817 7497 12851 7531
rect 13185 7497 13219 7531
rect 13645 7497 13679 7531
rect 14289 7497 14323 7531
rect 16773 7497 16807 7531
rect 17509 7497 17543 7531
rect 18429 7497 18463 7531
rect 2789 7429 2823 7463
rect 4353 7429 4387 7463
rect 5733 7429 5767 7463
rect 9628 7429 9662 7463
rect 14657 7429 14691 7463
rect 1685 7361 1719 7395
rect 2145 7361 2179 7395
rect 4445 7361 4479 7395
rect 5825 7361 5859 7395
rect 6653 7361 6687 7395
rect 7297 7361 7331 7395
rect 7757 7361 7791 7395
rect 9873 7361 9907 7395
rect 9965 7361 9999 7395
rect 10232 7361 10266 7395
rect 12725 7361 12759 7395
rect 13553 7361 13587 7395
rect 15117 7361 15151 7395
rect 15384 7361 15418 7395
rect 17417 7361 17451 7395
rect 18153 7361 18187 7395
rect 18245 7361 18279 7395
rect 1961 7293 1995 7327
rect 2053 7293 2087 7327
rect 4813 7293 4847 7327
rect 4905 7293 4939 7327
rect 5641 7293 5675 7327
rect 7389 7293 7423 7327
rect 7481 7293 7515 7327
rect 11621 7293 11655 7327
rect 11805 7293 11839 7327
rect 12909 7293 12943 7327
rect 13737 7293 13771 7327
rect 14013 7293 14047 7327
rect 14749 7293 14783 7327
rect 14933 7293 14967 7327
rect 11345 7225 11379 7259
rect 2513 7157 2547 7191
rect 5365 7157 5399 7191
rect 6193 7157 6227 7191
rect 6469 7157 6503 7191
rect 6745 7157 6779 7191
rect 8401 7157 8435 7191
rect 12265 7157 12299 7191
rect 16497 7157 16531 7191
rect 6561 6953 6595 6987
rect 9965 6953 9999 6987
rect 11529 6953 11563 6987
rect 12725 6953 12759 6987
rect 16865 6953 16899 6987
rect 17417 6953 17451 6987
rect 12633 6885 12667 6919
rect 6193 6817 6227 6851
rect 6285 6817 6319 6851
rect 7205 6817 7239 6851
rect 9045 6817 9079 6851
rect 9781 6817 9815 6851
rect 11345 6817 11379 6851
rect 12173 6817 12207 6851
rect 13369 6817 13403 6851
rect 16129 6817 16163 6851
rect 16405 6817 16439 6851
rect 1593 6749 1627 6783
rect 3525 6749 3559 6783
rect 3893 6749 3927 6783
rect 5641 6749 5675 6783
rect 7021 6749 7055 6783
rect 8769 6749 8803 6783
rect 12449 6749 12483 6783
rect 13093 6749 13127 6783
rect 13553 6749 13587 6783
rect 13829 6749 13863 6783
rect 14105 6749 14139 6783
rect 15945 6749 15979 6783
rect 16957 6749 16991 6783
rect 17509 6749 17543 6783
rect 17877 6749 17911 6783
rect 18245 6749 18279 6783
rect 1838 6681 1872 6715
rect 3249 6681 3283 6715
rect 4160 6681 4194 6715
rect 8524 6681 8558 6715
rect 9321 6681 9355 6715
rect 11100 6681 11134 6715
rect 14350 6681 14384 6715
rect 16589 6681 16623 6715
rect 1501 6613 1535 6647
rect 2973 6613 3007 6647
rect 5273 6613 5307 6647
rect 5457 6613 5491 6647
rect 5733 6613 5767 6647
rect 6101 6613 6135 6647
rect 6929 6613 6963 6647
rect 7389 6613 7423 6647
rect 9229 6613 9263 6647
rect 9689 6613 9723 6647
rect 11897 6613 11931 6647
rect 11989 6613 12023 6647
rect 13185 6613 13219 6647
rect 15485 6613 15519 6647
rect 15577 6613 15611 6647
rect 16037 6613 16071 6647
rect 17141 6613 17175 6647
rect 17693 6613 17727 6647
rect 18061 6613 18095 6647
rect 18429 6613 18463 6647
rect 2237 6409 2271 6443
rect 4629 6409 4663 6443
rect 4997 6409 5031 6443
rect 5457 6409 5491 6443
rect 5825 6409 5859 6443
rect 7849 6409 7883 6443
rect 8217 6409 8251 6443
rect 8677 6409 8711 6443
rect 9045 6409 9079 6443
rect 11805 6409 11839 6443
rect 11989 6409 12023 6443
rect 12817 6409 12851 6443
rect 13277 6409 13311 6443
rect 14473 6409 14507 6443
rect 14933 6409 14967 6443
rect 17049 6409 17083 6443
rect 18429 6409 18463 6443
rect 2329 6341 2363 6375
rect 3902 6341 3936 6375
rect 5089 6341 5123 6375
rect 11529 6341 11563 6375
rect 14105 6341 14139 6375
rect 16037 6341 16071 6375
rect 16865 6341 16899 6375
rect 1869 6273 1903 6307
rect 4537 6273 4571 6307
rect 5917 6273 5951 6307
rect 6377 6273 6411 6307
rect 6644 6273 6678 6307
rect 9781 6273 9815 6307
rect 10997 6273 11031 6307
rect 11253 6273 11287 6307
rect 12357 6273 12391 6307
rect 13185 6273 13219 6307
rect 14013 6273 14047 6307
rect 14841 6273 14875 6307
rect 15301 6273 15335 6307
rect 15945 6273 15979 6307
rect 17509 6273 17543 6307
rect 17877 6273 17911 6307
rect 18245 6273 18279 6307
rect 1685 6205 1719 6239
rect 2145 6205 2179 6239
rect 4169 6205 4203 6239
rect 5181 6205 5215 6239
rect 6101 6205 6135 6239
rect 8309 6205 8343 6239
rect 8401 6205 8435 6239
rect 9137 6205 9171 6239
rect 9321 6205 9355 6239
rect 12449 6205 12483 6239
rect 12633 6205 12667 6239
rect 13369 6205 13403 6239
rect 14197 6205 14231 6239
rect 15025 6205 15059 6239
rect 16313 6205 16347 6239
rect 16773 6205 16807 6239
rect 17785 6205 17819 6239
rect 2697 6137 2731 6171
rect 13645 6137 13679 6171
rect 16497 6137 16531 6171
rect 18061 6137 18095 6171
rect 2789 6069 2823 6103
rect 4353 6069 4387 6103
rect 7757 6069 7791 6103
rect 9597 6069 9631 6103
rect 9873 6069 9907 6103
rect 17325 6069 17359 6103
rect 1593 5865 1627 5899
rect 6745 5865 6779 5899
rect 10885 5865 10919 5899
rect 16405 5865 16439 5899
rect 17325 5865 17359 5899
rect 17785 5865 17819 5899
rect 5181 5797 5215 5831
rect 14933 5797 14967 5831
rect 4537 5729 4571 5763
rect 8493 5729 8527 5763
rect 8953 5729 8987 5763
rect 14657 5729 14691 5763
rect 15485 5729 15519 5763
rect 2717 5661 2751 5695
rect 2973 5661 3007 5695
rect 3525 5661 3559 5695
rect 4353 5661 4387 5695
rect 4813 5661 4847 5695
rect 5273 5661 5307 5695
rect 9209 5661 9243 5695
rect 12173 5661 12207 5695
rect 12265 5661 12299 5695
rect 14473 5661 14507 5695
rect 15761 5661 15795 5695
rect 17877 5661 17911 5695
rect 18245 5661 18279 5695
rect 3249 5593 3283 5627
rect 4077 5593 4111 5627
rect 8226 5593 8260 5627
rect 12532 5593 12566 5627
rect 13829 5593 13863 5627
rect 1501 5525 1535 5559
rect 4721 5525 4755 5559
rect 7113 5525 7147 5559
rect 8769 5525 8803 5559
rect 10333 5525 10367 5559
rect 13645 5525 13679 5559
rect 14105 5525 14139 5559
rect 14565 5525 14599 5559
rect 15301 5525 15335 5559
rect 15393 5525 15427 5559
rect 16497 5525 16531 5559
rect 17509 5525 17543 5559
rect 18061 5525 18095 5559
rect 18429 5525 18463 5559
rect 2237 5321 2271 5355
rect 4997 5321 5031 5355
rect 5365 5321 5399 5355
rect 5917 5321 5951 5355
rect 7021 5321 7055 5355
rect 7481 5321 7515 5355
rect 9045 5321 9079 5355
rect 9597 5321 9631 5355
rect 9965 5321 9999 5355
rect 10057 5321 10091 5355
rect 10425 5321 10459 5355
rect 10885 5321 10919 5355
rect 13001 5321 13035 5355
rect 13829 5321 13863 5355
rect 15577 5321 15611 5355
rect 16037 5321 16071 5355
rect 16313 5321 16347 5355
rect 16497 5321 16531 5355
rect 16681 5321 16715 5355
rect 16865 5321 16899 5355
rect 17693 5321 17727 5355
rect 18429 5321 18463 5355
rect 2605 5253 2639 5287
rect 4537 5253 4571 5287
rect 5825 5253 5859 5287
rect 7389 5253 7423 5287
rect 10793 5253 10827 5287
rect 11253 5253 11287 5287
rect 11796 5253 11830 5287
rect 15945 5253 15979 5287
rect 1685 5185 1719 5219
rect 2145 5185 2179 5219
rect 6929 5185 6963 5219
rect 8217 5185 8251 5219
rect 9137 5185 9171 5219
rect 13369 5185 13403 5219
rect 13461 5185 13495 5219
rect 14372 5185 14406 5219
rect 17877 5185 17911 5219
rect 18245 5185 18279 5219
rect 2329 5117 2363 5151
rect 4721 5117 4755 5151
rect 4905 5117 4939 5151
rect 6009 5117 6043 5151
rect 6745 5117 6779 5151
rect 7573 5117 7607 5151
rect 8309 5117 8343 5151
rect 8493 5117 8527 5151
rect 8953 5117 8987 5151
rect 10241 5117 10275 5151
rect 10977 5117 11011 5151
rect 11529 5117 11563 5151
rect 13645 5117 13679 5151
rect 14105 5117 14139 5151
rect 1501 5049 1535 5083
rect 5457 5049 5491 5083
rect 12909 5049 12943 5083
rect 15485 5049 15519 5083
rect 1777 4981 1811 5015
rect 3893 4981 3927 5015
rect 7849 4981 7883 5015
rect 9505 4981 9539 5015
rect 18061 4981 18095 5015
rect 3893 4777 3927 4811
rect 13921 4777 13955 4811
rect 16681 4777 16715 4811
rect 17693 4777 17727 4811
rect 14933 4709 14967 4743
rect 17233 4709 17267 4743
rect 1593 4641 1627 4675
rect 1685 4641 1719 4675
rect 6837 4641 6871 4675
rect 7389 4641 7423 4675
rect 11621 4641 11655 4675
rect 12173 4641 12207 4675
rect 13093 4641 13127 4675
rect 14657 4641 14691 4675
rect 15485 4641 15519 4675
rect 17509 4641 17543 4675
rect 1777 4573 1811 4607
rect 2237 4573 2271 4607
rect 3985 4573 4019 4607
rect 6570 4573 6604 4607
rect 7205 4573 7239 4607
rect 9045 4573 9079 4607
rect 10710 4573 10744 4607
rect 10977 4573 11011 4607
rect 13277 4573 13311 4607
rect 15761 4573 15795 4607
rect 17877 4573 17911 4607
rect 2504 4505 2538 4539
rect 4252 4505 4286 4539
rect 7634 4505 7668 4539
rect 9321 4505 9355 4539
rect 11437 4505 11471 4539
rect 11897 4505 11931 4539
rect 12909 4505 12943 4539
rect 14473 4505 14507 4539
rect 15301 4505 15335 4539
rect 16497 4505 16531 4539
rect 18429 4505 18463 4539
rect 2145 4437 2179 4471
rect 3617 4437 3651 4471
rect 5365 4437 5399 4471
rect 5457 4437 5491 4471
rect 7021 4437 7055 4471
rect 8769 4437 8803 4471
rect 9597 4437 9631 4471
rect 11069 4437 11103 4471
rect 11529 4437 11563 4471
rect 12449 4437 12483 4471
rect 12817 4437 12851 4471
rect 14105 4437 14139 4471
rect 14565 4437 14599 4471
rect 15393 4437 15427 4471
rect 16405 4437 16439 4471
rect 16865 4437 16899 4471
rect 17049 4437 17083 4471
rect 18061 4437 18095 4471
rect 18337 4437 18371 4471
rect 2145 4233 2179 4267
rect 2605 4233 2639 4267
rect 5365 4233 5399 4267
rect 8033 4233 8067 4267
rect 8401 4233 8435 4267
rect 8769 4233 8803 4267
rect 10057 4233 10091 4267
rect 13461 4233 13495 4267
rect 15117 4233 15151 4267
rect 15485 4233 15519 4267
rect 16313 4233 16347 4267
rect 16957 4233 16991 4267
rect 17325 4233 17359 4267
rect 2237 4165 2271 4199
rect 3718 4165 3752 4199
rect 5825 4165 5859 4199
rect 17969 4165 18003 4199
rect 1685 4097 1719 4131
rect 4261 4097 4295 4131
rect 4537 4097 4571 4131
rect 4905 4097 4939 4131
rect 4997 4097 5031 4131
rect 7593 4097 7627 4131
rect 7849 4097 7883 4131
rect 8217 4097 8251 4131
rect 9505 4097 9539 4131
rect 10885 4097 10919 4131
rect 11785 4097 11819 4131
rect 13277 4097 13311 4131
rect 13645 4097 13679 4131
rect 13912 4097 13946 4131
rect 16129 4097 16163 4131
rect 18337 4097 18371 4131
rect 2421 4029 2455 4063
rect 3985 4029 4019 4063
rect 4721 4029 4755 4063
rect 5917 4029 5951 4063
rect 6009 4029 6043 4063
rect 8861 4029 8895 4063
rect 8953 4029 8987 4063
rect 10149 4029 10183 4063
rect 10333 4029 10367 4063
rect 10977 4029 11011 4063
rect 11069 4029 11103 4063
rect 11529 4029 11563 4063
rect 13093 4029 13127 4063
rect 15577 4029 15611 4063
rect 15669 4029 15703 4063
rect 15945 4029 15979 4063
rect 16773 4029 16807 4063
rect 17785 4029 17819 4063
rect 1501 3961 1535 3995
rect 1777 3961 1811 3995
rect 5457 3961 5491 3995
rect 9321 3961 9355 3995
rect 10517 3961 10551 3995
rect 17601 3961 17635 3995
rect 6469 3893 6503 3927
rect 9689 3893 9723 3927
rect 12909 3893 12943 3927
rect 15025 3893 15059 3927
rect 17141 3893 17175 3927
rect 17509 3893 17543 3927
rect 18245 3893 18279 3927
rect 3617 3689 3651 3723
rect 4629 3689 4663 3723
rect 7941 3689 7975 3723
rect 8953 3689 8987 3723
rect 9781 3689 9815 3723
rect 10057 3689 10091 3723
rect 10885 3689 10919 3723
rect 13921 3689 13955 3723
rect 14841 3689 14875 3723
rect 15577 3689 15611 3723
rect 15669 3689 15703 3723
rect 15853 3689 15887 3723
rect 16865 3689 16899 3723
rect 2881 3621 2915 3655
rect 4537 3621 4571 3655
rect 11805 3621 11839 3655
rect 16221 3621 16255 3655
rect 17693 3621 17727 3655
rect 18429 3621 18463 3655
rect 3985 3553 4019 3587
rect 4077 3553 4111 3587
rect 5089 3553 5123 3587
rect 5273 3553 5307 3587
rect 8493 3553 8527 3587
rect 9413 3553 9447 3587
rect 9597 3553 9631 3587
rect 10701 3553 10735 3587
rect 11437 3553 11471 3587
rect 14289 3553 14323 3587
rect 14381 3553 14415 3587
rect 16037 3553 16071 3587
rect 1501 3485 1535 3519
rect 2973 3485 3007 3519
rect 4997 3485 5031 3519
rect 7849 3485 7883 3519
rect 9321 3485 9355 3519
rect 10425 3485 10459 3519
rect 10517 3485 10551 3519
rect 11989 3485 12023 3519
rect 12173 3485 12207 3519
rect 13737 3485 13771 3519
rect 14933 3485 14967 3519
rect 17141 3485 17175 3519
rect 17325 3485 17359 3519
rect 17509 3485 17543 3519
rect 17877 3485 17911 3519
rect 18245 3485 18279 3519
rect 1768 3417 1802 3451
rect 5457 3417 5491 3451
rect 7481 3417 7515 3451
rect 11253 3417 11287 3451
rect 12440 3417 12474 3451
rect 16405 3417 16439 3451
rect 16589 3417 16623 3451
rect 16957 3417 16991 3451
rect 4169 3349 4203 3383
rect 6193 3349 6227 3383
rect 7665 3349 7699 3383
rect 8309 3349 8343 3383
rect 8401 3349 8435 3383
rect 11345 3349 11379 3383
rect 13553 3349 13587 3383
rect 14473 3349 14507 3383
rect 18061 3349 18095 3383
rect 1501 3145 1535 3179
rect 3065 3145 3099 3179
rect 4537 3145 4571 3179
rect 7021 3145 7055 3179
rect 10149 3145 10183 3179
rect 10885 3145 10919 3179
rect 11253 3145 11287 3179
rect 11989 3145 12023 3179
rect 13461 3145 13495 3179
rect 4353 3077 4387 3111
rect 7849 3077 7883 3111
rect 12633 3077 12667 3111
rect 16221 3077 16255 3111
rect 1685 3009 1719 3043
rect 2145 3009 2179 3043
rect 4721 3009 4755 3043
rect 4813 3009 4847 3043
rect 5080 3009 5114 3043
rect 6929 3009 6963 3043
rect 7389 3009 7423 3043
rect 7481 3009 7515 3043
rect 10057 3009 10091 3043
rect 10793 3009 10827 3043
rect 11897 3009 11931 3043
rect 12357 3009 12391 3043
rect 14749 3009 14783 3043
rect 14841 3009 14875 3043
rect 15393 3009 15427 3043
rect 15945 3009 15979 3043
rect 16957 3009 16991 3043
rect 17141 3009 17175 3043
rect 17509 3009 17543 3043
rect 17877 3009 17911 3043
rect 18245 3009 18279 3043
rect 1869 2941 1903 2975
rect 2053 2941 2087 2975
rect 6745 2941 6779 2975
rect 7573 2941 7607 2975
rect 10241 2941 10275 2975
rect 10609 2941 10643 2975
rect 12081 2941 12115 2975
rect 15117 2941 15151 2975
rect 15577 2941 15611 2975
rect 16773 2873 16807 2907
rect 2513 2805 2547 2839
rect 6193 2805 6227 2839
rect 9137 2805 9171 2839
rect 9689 2805 9723 2839
rect 11529 2805 11563 2839
rect 17325 2805 17359 2839
rect 17693 2805 17727 2839
rect 18061 2805 18095 2839
rect 18429 2805 18463 2839
rect 2881 2601 2915 2635
rect 5089 2601 5123 2635
rect 6193 2601 6227 2635
rect 10609 2601 10643 2635
rect 11529 2601 11563 2635
rect 13921 2601 13955 2635
rect 16221 2601 16255 2635
rect 16405 2601 16439 2635
rect 16957 2601 16991 2635
rect 6561 2533 6595 2567
rect 9689 2533 9723 2567
rect 13001 2533 13035 2567
rect 2145 2465 2179 2499
rect 2329 2465 2363 2499
rect 3341 2465 3375 2499
rect 3525 2465 3559 2499
rect 4169 2465 4203 2499
rect 4353 2465 4387 2499
rect 5825 2465 5859 2499
rect 7113 2465 7147 2499
rect 8217 2465 8251 2499
rect 9045 2465 9079 2499
rect 9229 2465 9263 2499
rect 9965 2465 9999 2499
rect 11161 2465 11195 2499
rect 12081 2465 12115 2499
rect 14197 2465 14231 2499
rect 15209 2465 15243 2499
rect 16037 2465 16071 2499
rect 1961 2397 1995 2431
rect 2421 2397 2455 2431
rect 5549 2397 5583 2431
rect 6469 2397 6503 2431
rect 6929 2397 6963 2431
rect 7665 2397 7699 2431
rect 8769 2397 8803 2431
rect 10057 2397 10091 2431
rect 12357 2397 12391 2431
rect 13093 2397 13127 2431
rect 14381 2397 14415 2431
rect 14933 2397 14967 2431
rect 15485 2397 15519 2431
rect 17693 2397 17727 2431
rect 18061 2397 18095 2431
rect 1685 2329 1719 2363
rect 3985 2329 4019 2363
rect 4445 2329 4479 2363
rect 10149 2329 10183 2363
rect 11069 2329 11103 2363
rect 11989 2329 12023 2363
rect 15761 2329 15795 2363
rect 17417 2329 17451 2363
rect 18429 2329 18463 2363
rect 2789 2261 2823 2295
rect 3249 2261 3283 2295
rect 4813 2261 4847 2295
rect 5181 2261 5215 2295
rect 5641 2261 5675 2295
rect 7021 2261 7055 2295
rect 7481 2261 7515 2295
rect 9321 2261 9355 2295
rect 10517 2261 10551 2295
rect 10977 2261 11011 2295
rect 11897 2261 11931 2295
rect 13737 2261 13771 2295
rect 14473 2261 14507 2295
rect 14841 2261 14875 2295
rect 16681 2261 16715 2295
rect 17049 2261 17083 2295
rect 17233 2261 17267 2295
rect 17877 2261 17911 2295
rect 18245 2261 18279 2295
<< metal1 >>
rect 3694 15376 3700 15428
rect 3752 15416 3758 15428
rect 7466 15416 7472 15428
rect 3752 15388 7472 15416
rect 3752 15376 3758 15388
rect 7466 15376 7472 15388
rect 7524 15376 7530 15428
rect 13170 15308 13176 15360
rect 13228 15348 13234 15360
rect 18046 15348 18052 15360
rect 13228 15320 18052 15348
rect 13228 15308 13234 15320
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 3510 15172 3516 15224
rect 3568 15212 3574 15224
rect 9214 15212 9220 15224
rect 3568 15184 9220 15212
rect 3568 15172 3574 15184
rect 9214 15172 9220 15184
rect 9272 15172 9278 15224
rect 13262 15172 13268 15224
rect 13320 15212 13326 15224
rect 15194 15212 15200 15224
rect 13320 15184 15200 15212
rect 13320 15172 13326 15184
rect 15194 15172 15200 15184
rect 15252 15172 15258 15224
rect 1104 14714 18860 14736
rect 1104 14662 3174 14714
rect 3226 14662 3238 14714
rect 3290 14662 3302 14714
rect 3354 14662 3366 14714
rect 3418 14662 3430 14714
rect 3482 14662 7622 14714
rect 7674 14662 7686 14714
rect 7738 14662 7750 14714
rect 7802 14662 7814 14714
rect 7866 14662 7878 14714
rect 7930 14662 12070 14714
rect 12122 14662 12134 14714
rect 12186 14662 12198 14714
rect 12250 14662 12262 14714
rect 12314 14662 12326 14714
rect 12378 14662 16518 14714
rect 16570 14662 16582 14714
rect 16634 14662 16646 14714
rect 16698 14662 16710 14714
rect 16762 14662 16774 14714
rect 16826 14662 18860 14714
rect 1104 14640 18860 14662
rect 3786 14424 3792 14476
rect 3844 14464 3850 14476
rect 10502 14464 10508 14476
rect 3844 14436 10508 14464
rect 3844 14424 3850 14436
rect 10502 14424 10508 14436
rect 10560 14424 10566 14476
rect 10594 14424 10600 14476
rect 10652 14464 10658 14476
rect 15286 14464 15292 14476
rect 10652 14436 15292 14464
rect 10652 14424 10658 14436
rect 15286 14424 15292 14436
rect 15344 14424 15350 14476
rect 1118 14356 1124 14408
rect 1176 14396 1182 14408
rect 13078 14396 13084 14408
rect 1176 14368 13084 14396
rect 1176 14356 1182 14368
rect 13078 14356 13084 14368
rect 13136 14356 13142 14408
rect 5534 14288 5540 14340
rect 5592 14328 5598 14340
rect 18046 14328 18052 14340
rect 5592 14300 18052 14328
rect 5592 14288 5598 14300
rect 18046 14288 18052 14300
rect 18104 14288 18110 14340
rect 4062 14220 4068 14272
rect 4120 14260 4126 14272
rect 7190 14260 7196 14272
rect 4120 14232 7196 14260
rect 4120 14220 4126 14232
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 7558 14220 7564 14272
rect 7616 14260 7622 14272
rect 15654 14260 15660 14272
rect 7616 14232 15660 14260
rect 7616 14220 7622 14232
rect 15654 14220 15660 14232
rect 15712 14220 15718 14272
rect 1104 14170 18860 14192
rect 1104 14118 5398 14170
rect 5450 14118 5462 14170
rect 5514 14118 5526 14170
rect 5578 14118 5590 14170
rect 5642 14118 5654 14170
rect 5706 14118 9846 14170
rect 9898 14118 9910 14170
rect 9962 14118 9974 14170
rect 10026 14118 10038 14170
rect 10090 14118 10102 14170
rect 10154 14118 14294 14170
rect 14346 14118 14358 14170
rect 14410 14118 14422 14170
rect 14474 14118 14486 14170
rect 14538 14118 14550 14170
rect 14602 14118 18860 14170
rect 1104 14096 18860 14118
rect 3878 14016 3884 14068
rect 3936 14056 3942 14068
rect 5261 14059 5319 14065
rect 3936 14028 5120 14056
rect 3936 14016 3942 14028
rect 2130 13948 2136 14000
rect 2188 13988 2194 14000
rect 4982 13988 4988 14000
rect 2188 13960 4988 13988
rect 2188 13948 2194 13960
rect 4982 13948 4988 13960
rect 5040 13948 5046 14000
rect 4890 13920 4896 13932
rect 4851 13892 4896 13920
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 5092 13920 5120 14028
rect 5261 14025 5273 14059
rect 5307 14056 5319 14059
rect 10962 14056 10968 14068
rect 5307 14028 10968 14056
rect 5307 14025 5319 14028
rect 5261 14019 5319 14025
rect 10962 14016 10968 14028
rect 11020 14016 11026 14068
rect 15194 14056 15200 14068
rect 12406 14028 15200 14056
rect 5166 13948 5172 14000
rect 5224 13988 5230 14000
rect 7558 13988 7564 14000
rect 5224 13960 7564 13988
rect 5224 13948 5230 13960
rect 7558 13948 7564 13960
rect 7616 13948 7622 14000
rect 12406 13988 12434 14028
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 18046 14056 18052 14068
rect 16500 14028 17724 14056
rect 18007 14028 18052 14056
rect 13078 13988 13084 14000
rect 7659 13960 12434 13988
rect 13039 13960 13084 13988
rect 7659 13920 7687 13960
rect 13078 13948 13084 13960
rect 13136 13988 13142 14000
rect 14001 13991 14059 13997
rect 13136 13960 13308 13988
rect 13136 13948 13142 13960
rect 13280 13929 13308 13960
rect 14001 13957 14013 13991
rect 14047 13988 14059 13991
rect 14182 13988 14188 14000
rect 14047 13960 14188 13988
rect 14047 13957 14059 13960
rect 14001 13951 14059 13957
rect 14182 13948 14188 13960
rect 14240 13988 14246 14000
rect 15102 13988 15108 14000
rect 14240 13960 15108 13988
rect 14240 13948 14246 13960
rect 15102 13948 15108 13960
rect 15160 13988 15166 14000
rect 16500 13997 16528 14028
rect 15565 13991 15623 13997
rect 15565 13988 15577 13991
rect 15160 13960 15577 13988
rect 15160 13948 15166 13960
rect 15565 13957 15577 13960
rect 15611 13957 15623 13991
rect 15565 13951 15623 13957
rect 16485 13991 16543 13997
rect 16485 13957 16497 13991
rect 16531 13957 16543 13991
rect 16485 13951 16543 13957
rect 16853 13991 16911 13997
rect 16853 13957 16865 13991
rect 16899 13988 16911 13991
rect 16942 13988 16948 14000
rect 16899 13960 16948 13988
rect 16899 13957 16911 13960
rect 16853 13951 16911 13957
rect 16942 13948 16948 13960
rect 17000 13948 17006 14000
rect 17696 13988 17724 14028
rect 18046 14016 18052 14028
rect 18104 14016 18110 14068
rect 18417 14059 18475 14065
rect 18417 14025 18429 14059
rect 18463 14056 18475 14059
rect 18506 14056 18512 14068
rect 18463 14028 18512 14056
rect 18463 14025 18475 14028
rect 18417 14019 18475 14025
rect 18506 14016 18512 14028
rect 18564 14016 18570 14068
rect 18782 13988 18788 14000
rect 17696 13960 18788 13988
rect 18782 13948 18788 13960
rect 18840 13948 18846 14000
rect 5092 13892 7687 13920
rect 13265 13923 13323 13929
rect 13265 13889 13277 13923
rect 13311 13889 13323 13923
rect 13630 13920 13636 13932
rect 13591 13892 13636 13920
rect 13265 13883 13323 13889
rect 13630 13880 13636 13892
rect 13688 13880 13694 13932
rect 14093 13923 14151 13929
rect 14093 13889 14105 13923
rect 14139 13889 14151 13923
rect 17862 13920 17868 13932
rect 17823 13892 17868 13920
rect 14093 13883 14151 13889
rect 4617 13855 4675 13861
rect 4617 13821 4629 13855
rect 4663 13821 4675 13855
rect 4798 13852 4804 13864
rect 4759 13824 4804 13852
rect 4617 13815 4675 13821
rect 4632 13784 4660 13815
rect 4798 13812 4804 13824
rect 4856 13812 4862 13864
rect 6914 13852 6920 13864
rect 6827 13824 6920 13852
rect 6914 13812 6920 13824
rect 6972 13852 6978 13864
rect 13446 13852 13452 13864
rect 6972 13824 13452 13852
rect 6972 13812 6978 13824
rect 13446 13812 13452 13824
rect 13504 13812 13510 13864
rect 13538 13812 13544 13864
rect 13596 13852 13602 13864
rect 14108 13852 14136 13883
rect 17862 13880 17868 13892
rect 17920 13880 17926 13932
rect 18046 13880 18052 13932
rect 18104 13920 18110 13932
rect 18233 13923 18291 13929
rect 18233 13920 18245 13923
rect 18104 13892 18245 13920
rect 18104 13880 18110 13892
rect 18233 13889 18245 13892
rect 18279 13889 18291 13923
rect 18233 13883 18291 13889
rect 13596 13824 14136 13852
rect 15473 13855 15531 13861
rect 13596 13812 13602 13824
rect 15473 13821 15485 13855
rect 15519 13852 15531 13855
rect 16761 13855 16819 13861
rect 15519 13824 16574 13852
rect 15519 13821 15531 13824
rect 15473 13815 15531 13821
rect 5166 13784 5172 13796
rect 4632 13756 5172 13784
rect 5166 13744 5172 13756
rect 5224 13744 5230 13796
rect 6932 13784 6960 13812
rect 15562 13784 15568 13796
rect 5276 13756 6960 13784
rect 7024 13756 15568 13784
rect 4430 13676 4436 13728
rect 4488 13716 4494 13728
rect 5276 13716 5304 13756
rect 4488 13688 5304 13716
rect 4488 13676 4494 13688
rect 5810 13676 5816 13728
rect 5868 13716 5874 13728
rect 5997 13719 6055 13725
rect 5997 13716 6009 13719
rect 5868 13688 6009 13716
rect 5868 13676 5874 13688
rect 5997 13685 6009 13688
rect 6043 13685 6055 13719
rect 5997 13679 6055 13685
rect 6086 13676 6092 13728
rect 6144 13716 6150 13728
rect 7024 13716 7052 13756
rect 15562 13744 15568 13756
rect 15620 13744 15626 13796
rect 16546 13784 16574 13824
rect 16761 13821 16773 13855
rect 16807 13852 16819 13855
rect 16850 13852 16856 13864
rect 16807 13824 16856 13852
rect 16807 13821 16819 13824
rect 16761 13815 16819 13821
rect 16850 13812 16856 13824
rect 16908 13812 16914 13864
rect 17034 13852 17040 13864
rect 16995 13824 17040 13852
rect 17034 13812 17040 13824
rect 17092 13812 17098 13864
rect 17126 13784 17132 13796
rect 16546 13756 17132 13784
rect 17126 13744 17132 13756
rect 17184 13744 17190 13796
rect 6144 13688 7052 13716
rect 6144 13676 6150 13688
rect 9398 13676 9404 13728
rect 9456 13716 9462 13728
rect 9769 13719 9827 13725
rect 9769 13716 9781 13719
rect 9456 13688 9781 13716
rect 9456 13676 9462 13688
rect 9769 13685 9781 13688
rect 9815 13716 9827 13719
rect 10594 13716 10600 13728
rect 9815 13688 10600 13716
rect 9815 13685 9827 13688
rect 9769 13679 9827 13685
rect 10594 13676 10600 13688
rect 10652 13676 10658 13728
rect 14734 13716 14740 13728
rect 14695 13688 14740 13716
rect 14734 13676 14740 13688
rect 14792 13676 14798 13728
rect 1104 13626 18860 13648
rect 1104 13574 3174 13626
rect 3226 13574 3238 13626
rect 3290 13574 3302 13626
rect 3354 13574 3366 13626
rect 3418 13574 3430 13626
rect 3482 13574 7622 13626
rect 7674 13574 7686 13626
rect 7738 13574 7750 13626
rect 7802 13574 7814 13626
rect 7866 13574 7878 13626
rect 7930 13574 12070 13626
rect 12122 13574 12134 13626
rect 12186 13574 12198 13626
rect 12250 13574 12262 13626
rect 12314 13574 12326 13626
rect 12378 13574 16518 13626
rect 16570 13574 16582 13626
rect 16634 13574 16646 13626
rect 16698 13574 16710 13626
rect 16762 13574 16774 13626
rect 16826 13574 18860 13626
rect 1104 13552 18860 13574
rect 3878 13512 3884 13524
rect 3839 13484 3884 13512
rect 3878 13472 3884 13484
rect 3936 13472 3942 13524
rect 4890 13472 4896 13524
rect 4948 13512 4954 13524
rect 5077 13515 5135 13521
rect 5077 13512 5089 13515
rect 4948 13484 5089 13512
rect 4948 13472 4954 13484
rect 5077 13481 5089 13484
rect 5123 13481 5135 13515
rect 8478 13512 8484 13524
rect 5077 13475 5135 13481
rect 5368 13484 8484 13512
rect 3970 13404 3976 13456
rect 4028 13444 4034 13456
rect 4249 13447 4307 13453
rect 4249 13444 4261 13447
rect 4028 13416 4261 13444
rect 4028 13404 4034 13416
rect 4249 13413 4261 13416
rect 4295 13444 4307 13447
rect 5258 13444 5264 13456
rect 4295 13416 5264 13444
rect 4295 13413 4307 13416
rect 4249 13407 4307 13413
rect 5258 13404 5264 13416
rect 5316 13404 5322 13456
rect 4433 13379 4491 13385
rect 4433 13345 4445 13379
rect 4479 13345 4491 13379
rect 4433 13339 4491 13345
rect 4154 13268 4160 13320
rect 4212 13308 4218 13320
rect 4448 13308 4476 13339
rect 4614 13336 4620 13388
rect 4672 13376 4678 13388
rect 5368 13376 5396 13484
rect 8478 13472 8484 13484
rect 8536 13472 8542 13524
rect 10226 13472 10232 13524
rect 10284 13512 10290 13524
rect 12529 13515 12587 13521
rect 12529 13512 12541 13515
rect 10284 13484 12541 13512
rect 10284 13472 10290 13484
rect 12529 13481 12541 13484
rect 12575 13512 12587 13515
rect 13630 13512 13636 13524
rect 12575 13484 13636 13512
rect 12575 13481 12587 13484
rect 12529 13475 12587 13481
rect 13630 13472 13636 13484
rect 13688 13472 13694 13524
rect 16577 13515 16635 13521
rect 16577 13481 16589 13515
rect 16623 13512 16635 13515
rect 16850 13512 16856 13524
rect 16623 13484 16856 13512
rect 16623 13481 16635 13484
rect 16577 13475 16635 13481
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 5997 13447 6055 13453
rect 5997 13444 6009 13447
rect 4672 13348 5396 13376
rect 5552 13416 6009 13444
rect 4672 13336 4678 13348
rect 4212 13280 4476 13308
rect 4709 13311 4767 13317
rect 4212 13268 4218 13280
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 5552 13308 5580 13416
rect 5997 13413 6009 13416
rect 6043 13413 6055 13447
rect 10502 13444 10508 13456
rect 10463 13416 10508 13444
rect 5997 13407 6055 13413
rect 10502 13404 10508 13416
rect 10560 13404 10566 13456
rect 15887 13447 15945 13453
rect 15887 13413 15899 13447
rect 15933 13444 15945 13447
rect 16942 13444 16948 13456
rect 15933 13416 16948 13444
rect 15933 13413 15945 13416
rect 15887 13407 15945 13413
rect 16942 13404 16948 13416
rect 17000 13404 17006 13456
rect 5718 13376 5724 13388
rect 5679 13348 5724 13376
rect 5718 13336 5724 13348
rect 5776 13336 5782 13388
rect 6546 13376 6552 13388
rect 6507 13348 6552 13376
rect 6546 13336 6552 13348
rect 6604 13336 6610 13388
rect 8478 13336 8484 13388
rect 8536 13376 8542 13388
rect 9398 13376 9404 13388
rect 8536 13348 9404 13376
rect 8536 13336 8542 13348
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 9585 13379 9643 13385
rect 9585 13345 9597 13379
rect 9631 13376 9643 13379
rect 9674 13376 9680 13388
rect 9631 13348 9680 13376
rect 9631 13345 9643 13348
rect 9585 13339 9643 13345
rect 9674 13336 9680 13348
rect 9732 13336 9738 13388
rect 11609 13379 11667 13385
rect 11609 13345 11621 13379
rect 11655 13376 11667 13379
rect 11882 13376 11888 13388
rect 11655 13348 11888 13376
rect 11655 13345 11667 13348
rect 11609 13339 11667 13345
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 15102 13336 15108 13388
rect 15160 13376 15166 13388
rect 15160 13348 15332 13376
rect 15160 13336 15166 13348
rect 4755 13280 5580 13308
rect 6457 13311 6515 13317
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 6457 13277 6469 13311
rect 6503 13308 6515 13311
rect 6914 13308 6920 13320
rect 6503 13280 6920 13308
rect 6503 13277 6515 13280
rect 6457 13271 6515 13277
rect 6914 13268 6920 13280
rect 6972 13268 6978 13320
rect 7834 13268 7840 13320
rect 7892 13308 7898 13320
rect 8389 13311 8447 13317
rect 8389 13308 8401 13311
rect 7892 13280 8401 13308
rect 7892 13268 7898 13280
rect 8389 13277 8401 13280
rect 8435 13277 8447 13311
rect 8389 13271 8447 13277
rect 9030 13268 9036 13320
rect 9088 13308 9094 13320
rect 9769 13311 9827 13317
rect 9769 13308 9781 13311
rect 9088 13280 9781 13308
rect 9088 13268 9094 13280
rect 9769 13277 9781 13280
rect 9815 13277 9827 13311
rect 9769 13271 9827 13277
rect 10962 13268 10968 13320
rect 11020 13308 11026 13320
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 11020 13280 11345 13308
rect 11020 13268 11026 13280
rect 11333 13277 11345 13280
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 12158 13268 12164 13320
rect 12216 13308 12222 13320
rect 13909 13311 13967 13317
rect 13909 13308 13921 13311
rect 12216 13280 13921 13308
rect 12216 13268 12222 13280
rect 13909 13277 13921 13280
rect 13955 13277 13967 13311
rect 15194 13308 15200 13320
rect 15155 13280 15200 13308
rect 13909 13271 13967 13277
rect 15194 13268 15200 13280
rect 15252 13268 15258 13320
rect 15304 13308 15332 13348
rect 15784 13311 15842 13317
rect 15784 13308 15796 13311
rect 15304 13280 15796 13308
rect 15784 13277 15796 13280
rect 15830 13277 15842 13311
rect 18046 13308 18052 13320
rect 18007 13280 18052 13308
rect 15784 13271 15842 13277
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 4065 13243 4123 13249
rect 4065 13209 4077 13243
rect 4111 13240 4123 13243
rect 4617 13243 4675 13249
rect 4111 13212 4568 13240
rect 4111 13209 4123 13212
rect 4065 13203 4123 13209
rect 1946 13132 1952 13184
rect 2004 13172 2010 13184
rect 3878 13172 3884 13184
rect 2004 13144 3884 13172
rect 2004 13132 2010 13144
rect 3878 13132 3884 13144
rect 3936 13132 3942 13184
rect 4540 13172 4568 13212
rect 4617 13209 4629 13243
rect 4663 13240 4675 13243
rect 4663 13212 5212 13240
rect 4663 13209 4675 13212
rect 4617 13203 4675 13209
rect 4890 13172 4896 13184
rect 4540 13144 4896 13172
rect 4890 13132 4896 13144
rect 4948 13132 4954 13184
rect 5184 13181 5212 13212
rect 5258 13200 5264 13252
rect 5316 13240 5322 13252
rect 5537 13243 5595 13249
rect 5537 13240 5549 13243
rect 5316 13212 5549 13240
rect 5316 13200 5322 13212
rect 5537 13209 5549 13212
rect 5583 13240 5595 13243
rect 5583 13212 7236 13240
rect 5583 13209 5595 13212
rect 5537 13203 5595 13209
rect 5169 13175 5227 13181
rect 5169 13141 5181 13175
rect 5215 13141 5227 13175
rect 5169 13135 5227 13141
rect 5629 13175 5687 13181
rect 5629 13141 5641 13175
rect 5675 13172 5687 13175
rect 5810 13172 5816 13184
rect 5675 13144 5816 13172
rect 5675 13141 5687 13144
rect 5629 13135 5687 13141
rect 5810 13132 5816 13144
rect 5868 13132 5874 13184
rect 6362 13172 6368 13184
rect 6323 13144 6368 13172
rect 6362 13132 6368 13144
rect 6420 13132 6426 13184
rect 6914 13172 6920 13184
rect 6875 13144 6920 13172
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 7006 13132 7012 13184
rect 7064 13172 7070 13184
rect 7208 13172 7236 13212
rect 8018 13200 8024 13252
rect 8076 13240 8082 13252
rect 8122 13243 8180 13249
rect 8122 13240 8134 13243
rect 8076 13212 8134 13240
rect 8076 13200 8082 13212
rect 8122 13209 8134 13212
rect 8168 13240 8180 13243
rect 8481 13243 8539 13249
rect 8481 13240 8493 13243
rect 8168 13212 8493 13240
rect 8168 13209 8180 13212
rect 8122 13203 8180 13209
rect 8481 13209 8493 13212
rect 8527 13209 8539 13243
rect 13664 13243 13722 13249
rect 8481 13203 8539 13209
rect 8588 13212 13584 13240
rect 8588 13172 8616 13212
rect 8938 13172 8944 13184
rect 7064 13144 7109 13172
rect 7208 13144 8616 13172
rect 8899 13144 8944 13172
rect 7064 13132 7070 13144
rect 8938 13132 8944 13144
rect 8996 13132 9002 13184
rect 9306 13172 9312 13184
rect 9267 13144 9312 13172
rect 9306 13132 9312 13144
rect 9364 13132 9370 13184
rect 10410 13172 10416 13184
rect 10371 13144 10416 13172
rect 10410 13132 10416 13144
rect 10468 13132 10474 13184
rect 13556 13172 13584 13212
rect 13664 13209 13676 13243
rect 13710 13240 13722 13243
rect 14734 13240 14740 13252
rect 13710 13212 14740 13240
rect 13710 13209 13722 13212
rect 13664 13203 13722 13209
rect 14734 13200 14740 13212
rect 14792 13200 14798 13252
rect 16761 13243 16819 13249
rect 16761 13209 16773 13243
rect 16807 13240 16819 13243
rect 17126 13240 17132 13252
rect 16807 13212 17132 13240
rect 16807 13209 16819 13212
rect 16761 13203 16819 13209
rect 17126 13200 17132 13212
rect 17184 13240 17190 13252
rect 18690 13240 18696 13252
rect 17184 13212 18696 13240
rect 17184 13200 17190 13212
rect 18690 13200 18696 13212
rect 18748 13200 18754 13252
rect 13998 13172 14004 13184
rect 13556 13144 14004 13172
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 14553 13175 14611 13181
rect 14553 13141 14565 13175
rect 14599 13172 14611 13175
rect 15286 13172 15292 13184
rect 14599 13144 15292 13172
rect 14599 13141 14611 13144
rect 14553 13135 14611 13141
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 17218 13132 17224 13184
rect 17276 13172 17282 13184
rect 17681 13175 17739 13181
rect 17681 13172 17693 13175
rect 17276 13144 17693 13172
rect 17276 13132 17282 13144
rect 17681 13141 17693 13144
rect 17727 13172 17739 13175
rect 17862 13172 17868 13184
rect 17727 13144 17868 13172
rect 17727 13141 17739 13144
rect 17681 13135 17739 13141
rect 17862 13132 17868 13144
rect 17920 13132 17926 13184
rect 1104 13082 18860 13104
rect 1104 13030 5398 13082
rect 5450 13030 5462 13082
rect 5514 13030 5526 13082
rect 5578 13030 5590 13082
rect 5642 13030 5654 13082
rect 5706 13030 9846 13082
rect 9898 13030 9910 13082
rect 9962 13030 9974 13082
rect 10026 13030 10038 13082
rect 10090 13030 10102 13082
rect 10154 13030 14294 13082
rect 14346 13030 14358 13082
rect 14410 13030 14422 13082
rect 14474 13030 14486 13082
rect 14538 13030 14550 13082
rect 14602 13030 18860 13082
rect 1104 13008 18860 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 2685 12971 2743 12977
rect 2685 12937 2697 12971
rect 2731 12968 2743 12971
rect 4341 12971 4399 12977
rect 2731 12940 4016 12968
rect 2731 12937 2743 12940
rect 2685 12931 2743 12937
rect 3878 12900 3884 12912
rect 2746 12872 3884 12900
rect 2501 12835 2559 12841
rect 2501 12801 2513 12835
rect 2547 12832 2559 12835
rect 2746 12832 2774 12872
rect 3878 12860 3884 12872
rect 3936 12860 3942 12912
rect 3988 12900 4016 12940
rect 4341 12937 4353 12971
rect 4387 12968 4399 12971
rect 4430 12968 4436 12980
rect 4387 12940 4436 12968
rect 4387 12937 4399 12940
rect 4341 12931 4399 12937
rect 4430 12928 4436 12940
rect 4488 12928 4494 12980
rect 4617 12971 4675 12977
rect 4617 12937 4629 12971
rect 4663 12968 4675 12971
rect 4798 12968 4804 12980
rect 4663 12940 4804 12968
rect 4663 12937 4675 12940
rect 4617 12931 4675 12937
rect 4798 12928 4804 12940
rect 4856 12928 4862 12980
rect 4985 12971 5043 12977
rect 4985 12937 4997 12971
rect 5031 12968 5043 12971
rect 5445 12971 5503 12977
rect 5445 12968 5457 12971
rect 5031 12940 5457 12968
rect 5031 12937 5043 12940
rect 4985 12931 5043 12937
rect 5445 12937 5457 12940
rect 5491 12937 5503 12971
rect 5445 12931 5503 12937
rect 5810 12928 5816 12980
rect 5868 12968 5874 12980
rect 8481 12971 8539 12977
rect 5868 12940 8156 12968
rect 5868 12928 5874 12940
rect 8128 12912 8156 12940
rect 8481 12937 8493 12971
rect 8527 12968 8539 12971
rect 8938 12968 8944 12980
rect 8527 12940 8944 12968
rect 8527 12937 8539 12940
rect 8481 12931 8539 12937
rect 8938 12928 8944 12940
rect 8996 12928 9002 12980
rect 13078 12968 13084 12980
rect 9048 12940 13084 12968
rect 4706 12900 4712 12912
rect 3988 12872 4712 12900
rect 4706 12860 4712 12872
rect 4764 12860 4770 12912
rect 7374 12860 7380 12912
rect 7432 12900 7438 12912
rect 7432 12872 7788 12900
rect 7432 12860 7438 12872
rect 2547 12804 2774 12832
rect 3044 12835 3102 12841
rect 2547 12801 2559 12804
rect 2501 12795 2559 12801
rect 3044 12801 3056 12835
rect 3090 12832 3102 12835
rect 5810 12832 5816 12844
rect 3090 12804 5580 12832
rect 5723 12804 5816 12832
rect 3090 12801 3102 12804
rect 3044 12795 3102 12801
rect 2774 12724 2780 12776
rect 2832 12764 2838 12776
rect 4614 12764 4620 12776
rect 2832 12736 2877 12764
rect 4356 12736 4620 12764
rect 2832 12724 2838 12736
rect 1857 12699 1915 12705
rect 1857 12665 1869 12699
rect 1903 12696 1915 12699
rect 4356 12696 4384 12736
rect 4614 12724 4620 12736
rect 4672 12724 4678 12776
rect 5074 12764 5080 12776
rect 5035 12736 5080 12764
rect 5074 12724 5080 12736
rect 5132 12724 5138 12776
rect 5169 12767 5227 12773
rect 5169 12733 5181 12767
rect 5215 12733 5227 12767
rect 5169 12727 5227 12733
rect 5184 12696 5212 12727
rect 1903 12668 2774 12696
rect 1903 12665 1915 12668
rect 1857 12659 1915 12665
rect 1946 12628 1952 12640
rect 1907 12600 1952 12628
rect 1946 12588 1952 12600
rect 2004 12588 2010 12640
rect 2130 12628 2136 12640
rect 2091 12600 2136 12628
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 2746 12628 2774 12668
rect 3988 12668 4384 12696
rect 4448 12668 5212 12696
rect 5552 12696 5580 12804
rect 5810 12792 5816 12804
rect 5868 12832 5874 12844
rect 6086 12832 6092 12844
rect 5868 12804 6092 12832
rect 5868 12792 5874 12804
rect 6086 12792 6092 12804
rect 6144 12792 6150 12844
rect 7006 12792 7012 12844
rect 7064 12832 7070 12844
rect 7570 12835 7628 12841
rect 7570 12832 7582 12835
rect 7064 12804 7582 12832
rect 7064 12792 7070 12804
rect 7570 12801 7582 12804
rect 7616 12801 7628 12835
rect 7760 12832 7788 12872
rect 8110 12860 8116 12912
rect 8168 12900 8174 12912
rect 9048 12900 9076 12940
rect 13078 12928 13084 12940
rect 13136 12928 13142 12980
rect 13538 12968 13544 12980
rect 13499 12940 13544 12968
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 13725 12971 13783 12977
rect 13725 12937 13737 12971
rect 13771 12937 13783 12971
rect 13725 12931 13783 12937
rect 18049 12971 18107 12977
rect 18049 12937 18061 12971
rect 18095 12968 18107 12971
rect 18138 12968 18144 12980
rect 18095 12940 18144 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 8168 12872 9076 12900
rect 8168 12860 8174 12872
rect 9674 12860 9680 12912
rect 9732 12900 9738 12912
rect 10054 12903 10112 12909
rect 10054 12900 10066 12903
rect 9732 12872 10066 12900
rect 9732 12860 9738 12872
rect 10054 12869 10066 12872
rect 10100 12869 10112 12903
rect 10962 12900 10968 12912
rect 10054 12863 10112 12869
rect 10152 12872 10968 12900
rect 7834 12832 7840 12844
rect 7747 12804 7840 12832
rect 7570 12795 7628 12801
rect 7834 12792 7840 12804
rect 7892 12792 7898 12844
rect 8021 12835 8079 12841
rect 8021 12801 8033 12835
rect 8067 12832 8079 12835
rect 10152 12832 10180 12872
rect 10962 12860 10968 12872
rect 11020 12860 11026 12912
rect 12428 12903 12486 12909
rect 12428 12869 12440 12903
rect 12474 12900 12486 12903
rect 13740 12900 13768 12931
rect 18138 12928 18144 12940
rect 18196 12968 18202 12980
rect 18417 12971 18475 12977
rect 18417 12968 18429 12971
rect 18196 12940 18429 12968
rect 18196 12928 18202 12940
rect 18417 12937 18429 12940
rect 18463 12937 18475 12971
rect 18417 12931 18475 12937
rect 13814 12900 13820 12912
rect 12474 12872 13820 12900
rect 12474 12869 12486 12872
rect 12428 12863 12486 12869
rect 13814 12860 13820 12872
rect 13872 12860 13878 12912
rect 14826 12860 14832 12912
rect 14884 12909 14890 12912
rect 14884 12900 14896 12909
rect 14884 12872 15332 12900
rect 14884 12863 14896 12872
rect 14884 12860 14890 12863
rect 8067 12804 10180 12832
rect 8067 12801 8079 12804
rect 8021 12795 8079 12801
rect 5902 12764 5908 12776
rect 5863 12736 5908 12764
rect 5902 12724 5908 12736
rect 5960 12724 5966 12776
rect 5997 12767 6055 12773
rect 5997 12733 6009 12767
rect 6043 12733 6055 12767
rect 5997 12727 6055 12733
rect 5718 12696 5724 12708
rect 5552 12668 5724 12696
rect 3988 12628 4016 12668
rect 4154 12628 4160 12640
rect 2746 12600 4016 12628
rect 4115 12600 4160 12628
rect 4154 12588 4160 12600
rect 4212 12628 4218 12640
rect 4448 12628 4476 12668
rect 5718 12656 5724 12668
rect 5776 12696 5782 12708
rect 6012 12696 6040 12727
rect 6457 12699 6515 12705
rect 6457 12696 6469 12699
rect 5776 12668 6469 12696
rect 5776 12656 5782 12668
rect 6457 12665 6469 12668
rect 6503 12696 6515 12699
rect 6546 12696 6552 12708
rect 6503 12668 6552 12696
rect 6503 12665 6515 12668
rect 6457 12659 6515 12665
rect 6546 12656 6552 12668
rect 6604 12656 6610 12708
rect 4212 12600 4476 12628
rect 4212 12588 4218 12600
rect 4522 12588 4528 12640
rect 4580 12628 4586 12640
rect 5810 12628 5816 12640
rect 4580 12600 5816 12628
rect 4580 12588 4586 12600
rect 5810 12588 5816 12600
rect 5868 12588 5874 12640
rect 7098 12588 7104 12640
rect 7156 12628 7162 12640
rect 8036 12628 8064 12795
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 10413 12835 10471 12841
rect 10413 12832 10425 12835
rect 10284 12804 10425 12832
rect 10284 12792 10290 12804
rect 10413 12801 10425 12804
rect 10459 12801 10471 12835
rect 14550 12832 14556 12844
rect 10413 12795 10471 12801
rect 14108 12804 14556 12832
rect 8205 12767 8263 12773
rect 8205 12733 8217 12767
rect 8251 12733 8263 12767
rect 8386 12764 8392 12776
rect 8347 12736 8392 12764
rect 8205 12727 8263 12733
rect 8220 12696 8248 12727
rect 8386 12724 8392 12736
rect 8444 12724 8450 12776
rect 10321 12767 10379 12773
rect 10321 12733 10333 12767
rect 10367 12764 10379 12767
rect 12158 12764 12164 12776
rect 10367 12736 12164 12764
rect 10367 12733 10379 12736
rect 10321 12727 10379 12733
rect 12158 12724 12164 12736
rect 12216 12724 12222 12776
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 14108 12764 14136 12804
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 15010 12792 15016 12844
rect 15068 12832 15074 12844
rect 15105 12835 15163 12841
rect 15105 12832 15117 12835
rect 15068 12804 15117 12832
rect 15068 12792 15074 12804
rect 15105 12801 15117 12804
rect 15151 12801 15163 12835
rect 15105 12795 15163 12801
rect 13872 12736 14136 12764
rect 13872 12724 13878 12736
rect 8941 12699 8999 12705
rect 8941 12696 8953 12699
rect 8220 12668 8953 12696
rect 8941 12665 8953 12668
rect 8987 12696 8999 12699
rect 9030 12696 9036 12708
rect 8987 12668 9036 12696
rect 8987 12665 8999 12668
rect 8941 12659 8999 12665
rect 9030 12656 9036 12668
rect 9088 12656 9094 12708
rect 15304 12696 15332 12872
rect 15749 12835 15807 12841
rect 15749 12801 15761 12835
rect 15795 12832 15807 12835
rect 17494 12832 17500 12844
rect 15795 12804 17500 12832
rect 15795 12801 15807 12804
rect 15749 12795 15807 12801
rect 17494 12792 17500 12804
rect 17552 12792 17558 12844
rect 17957 12835 18015 12841
rect 17957 12801 17969 12835
rect 18003 12832 18015 12835
rect 18322 12832 18328 12844
rect 18003 12804 18328 12832
rect 18003 12801 18015 12804
rect 17957 12795 18015 12801
rect 18322 12792 18328 12804
rect 18380 12792 18386 12844
rect 15838 12764 15844 12776
rect 15799 12736 15844 12764
rect 15838 12724 15844 12736
rect 15896 12724 15902 12776
rect 15933 12767 15991 12773
rect 15933 12733 15945 12767
rect 15979 12733 15991 12767
rect 15933 12727 15991 12733
rect 15948 12696 15976 12727
rect 18138 12724 18144 12776
rect 18196 12764 18202 12776
rect 18196 12736 18241 12764
rect 18196 12724 18202 12736
rect 17770 12696 17776 12708
rect 15304 12668 15976 12696
rect 17328 12668 17776 12696
rect 8846 12628 8852 12640
rect 7156 12600 8064 12628
rect 8807 12600 8852 12628
rect 7156 12588 7162 12600
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 9048 12628 9076 12656
rect 9582 12628 9588 12640
rect 9048 12600 9588 12628
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 11054 12628 11060 12640
rect 11015 12600 11060 12628
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 11790 12588 11796 12640
rect 11848 12628 11854 12640
rect 15102 12628 15108 12640
rect 11848 12600 15108 12628
rect 11848 12588 11854 12600
rect 15102 12588 15108 12600
rect 15160 12588 15166 12640
rect 15378 12628 15384 12640
rect 15339 12600 15384 12628
rect 15378 12588 15384 12600
rect 15436 12588 15442 12640
rect 17034 12588 17040 12640
rect 17092 12628 17098 12640
rect 17328 12637 17356 12668
rect 17770 12656 17776 12668
rect 17828 12656 17834 12708
rect 17313 12631 17371 12637
rect 17313 12628 17325 12631
rect 17092 12600 17325 12628
rect 17092 12588 17098 12600
rect 17313 12597 17325 12600
rect 17359 12597 17371 12631
rect 17586 12628 17592 12640
rect 17547 12600 17592 12628
rect 17313 12591 17371 12597
rect 17586 12588 17592 12600
rect 17644 12588 17650 12640
rect 1104 12538 18860 12560
rect 1104 12486 3174 12538
rect 3226 12486 3238 12538
rect 3290 12486 3302 12538
rect 3354 12486 3366 12538
rect 3418 12486 3430 12538
rect 3482 12486 7622 12538
rect 7674 12486 7686 12538
rect 7738 12486 7750 12538
rect 7802 12486 7814 12538
rect 7866 12486 7878 12538
rect 7930 12486 12070 12538
rect 12122 12486 12134 12538
rect 12186 12486 12198 12538
rect 12250 12486 12262 12538
rect 12314 12486 12326 12538
rect 12378 12486 16518 12538
rect 16570 12486 16582 12538
rect 16634 12486 16646 12538
rect 16698 12486 16710 12538
rect 16762 12486 16774 12538
rect 16826 12486 18860 12538
rect 1104 12464 18860 12486
rect 2317 12427 2375 12433
rect 2317 12393 2329 12427
rect 2363 12424 2375 12427
rect 4798 12424 4804 12436
rect 2363 12396 4804 12424
rect 2363 12393 2375 12396
rect 2317 12387 2375 12393
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 5074 12384 5080 12436
rect 5132 12424 5138 12436
rect 5353 12427 5411 12433
rect 5353 12424 5365 12427
rect 5132 12396 5365 12424
rect 5132 12384 5138 12396
rect 5353 12393 5365 12396
rect 5399 12393 5411 12427
rect 5353 12387 5411 12393
rect 5902 12384 5908 12436
rect 5960 12424 5966 12436
rect 6181 12427 6239 12433
rect 6181 12424 6193 12427
rect 5960 12396 6193 12424
rect 5960 12384 5966 12396
rect 6181 12393 6193 12396
rect 6227 12393 6239 12427
rect 8754 12424 8760 12436
rect 8667 12396 8760 12424
rect 6181 12387 6239 12393
rect 8754 12384 8760 12396
rect 8812 12424 8818 12436
rect 10226 12424 10232 12436
rect 8812 12396 10232 12424
rect 8812 12384 8818 12396
rect 10226 12384 10232 12396
rect 10284 12384 10290 12436
rect 14734 12424 14740 12436
rect 13372 12396 14740 12424
rect 5166 12356 5172 12368
rect 5127 12328 5172 12356
rect 5166 12316 5172 12328
rect 5224 12316 5230 12368
rect 7101 12359 7159 12365
rect 7101 12356 7113 12359
rect 6104 12328 7113 12356
rect 2608 12260 3924 12288
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12220 1731 12223
rect 2314 12220 2320 12232
rect 1719 12192 2320 12220
rect 1719 12189 1731 12192
rect 1673 12183 1731 12189
rect 2314 12180 2320 12192
rect 2372 12180 2378 12232
rect 2608 12164 2636 12260
rect 2958 12220 2964 12232
rect 2919 12192 2964 12220
rect 2958 12180 2964 12192
rect 3016 12180 3022 12232
rect 3786 12220 3792 12232
rect 3747 12192 3792 12220
rect 3786 12180 3792 12192
rect 3844 12180 3850 12232
rect 3896 12220 3924 12260
rect 5718 12248 5724 12300
rect 5776 12288 5782 12300
rect 5905 12291 5963 12297
rect 5905 12288 5917 12291
rect 5776 12260 5917 12288
rect 5776 12248 5782 12260
rect 5905 12257 5917 12260
rect 5951 12257 5963 12291
rect 5905 12251 5963 12257
rect 6104 12220 6132 12328
rect 7101 12325 7113 12328
rect 7147 12356 7159 12359
rect 7190 12356 7196 12368
rect 7147 12328 7196 12356
rect 7147 12325 7159 12328
rect 7101 12319 7159 12325
rect 7190 12316 7196 12328
rect 7248 12316 7254 12368
rect 9674 12316 9680 12368
rect 9732 12356 9738 12368
rect 10965 12359 11023 12365
rect 10965 12356 10977 12359
rect 9732 12328 10977 12356
rect 9732 12316 9738 12328
rect 6825 12291 6883 12297
rect 6825 12257 6837 12291
rect 6871 12288 6883 12291
rect 7006 12288 7012 12300
rect 6871 12260 7012 12288
rect 6871 12257 6883 12260
rect 6825 12251 6883 12257
rect 7006 12248 7012 12260
rect 7064 12248 7070 12300
rect 7374 12288 7380 12300
rect 7335 12260 7380 12288
rect 7374 12248 7380 12260
rect 7432 12248 7438 12300
rect 9217 12291 9275 12297
rect 9217 12257 9229 12291
rect 9263 12288 9275 12291
rect 9306 12288 9312 12300
rect 9263 12260 9312 12288
rect 9263 12257 9275 12260
rect 9217 12251 9275 12257
rect 9306 12248 9312 12260
rect 9364 12248 9370 12300
rect 9582 12248 9588 12300
rect 9640 12288 9646 12300
rect 10704 12297 10732 12328
rect 10965 12325 10977 12328
rect 11011 12325 11023 12359
rect 10965 12319 11023 12325
rect 13372 12297 13400 12396
rect 14734 12384 14740 12396
rect 14792 12424 14798 12436
rect 16025 12427 16083 12433
rect 16025 12424 16037 12427
rect 14792 12396 16037 12424
rect 14792 12384 14798 12396
rect 16025 12393 16037 12396
rect 16071 12393 16083 12427
rect 16025 12387 16083 12393
rect 13909 12359 13967 12365
rect 13909 12325 13921 12359
rect 13955 12325 13967 12359
rect 13909 12319 13967 12325
rect 9861 12291 9919 12297
rect 9861 12288 9873 12291
rect 9640 12260 9873 12288
rect 9640 12248 9646 12260
rect 9861 12257 9873 12260
rect 9907 12257 9919 12291
rect 9861 12251 9919 12257
rect 10689 12291 10747 12297
rect 10689 12257 10701 12291
rect 10735 12257 10747 12291
rect 10689 12251 10747 12257
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12257 13415 12291
rect 13924 12288 13952 12319
rect 14550 12316 14556 12368
rect 14608 12356 14614 12368
rect 15841 12359 15899 12365
rect 14608 12328 15516 12356
rect 14608 12316 14614 12328
rect 14752 12297 14780 12328
rect 14737 12291 14795 12297
rect 13924 12260 14504 12288
rect 13357 12251 13415 12257
rect 3896 12192 6132 12220
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12220 6607 12223
rect 7098 12220 7104 12232
rect 6595 12192 7104 12220
rect 6595 12189 6607 12192
rect 6549 12183 6607 12189
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 7644 12223 7702 12229
rect 7644 12189 7656 12223
rect 7690 12220 7702 12223
rect 10410 12220 10416 12232
rect 7690 12192 10416 12220
rect 7690 12189 7702 12192
rect 7644 12183 7702 12189
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 10502 12180 10508 12232
rect 10560 12220 10566 12232
rect 11330 12220 11336 12232
rect 10560 12192 11336 12220
rect 10560 12180 10566 12192
rect 11330 12180 11336 12192
rect 11388 12180 11394 12232
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12220 12403 12223
rect 12434 12220 12440 12232
rect 12391 12192 12440 12220
rect 12391 12189 12403 12192
rect 12345 12183 12403 12189
rect 12434 12180 12440 12192
rect 12492 12220 12498 12232
rect 12986 12220 12992 12232
rect 12492 12192 12992 12220
rect 12492 12180 12498 12192
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 13446 12220 13452 12232
rect 13407 12192 13452 12220
rect 13446 12180 13452 12192
rect 13504 12180 13510 12232
rect 14476 12229 14504 12260
rect 14737 12257 14749 12291
rect 14783 12257 14795 12291
rect 15378 12288 15384 12300
rect 15339 12260 15384 12288
rect 14737 12251 14795 12257
rect 15378 12248 15384 12260
rect 15436 12248 15442 12300
rect 15488 12297 15516 12328
rect 15841 12325 15853 12359
rect 15887 12356 15899 12359
rect 15930 12356 15936 12368
rect 15887 12328 15936 12356
rect 15887 12325 15899 12328
rect 15841 12319 15899 12325
rect 15930 12316 15936 12328
rect 15988 12316 15994 12368
rect 15473 12291 15531 12297
rect 15473 12257 15485 12291
rect 15519 12257 15531 12291
rect 15473 12251 15531 12257
rect 17681 12291 17739 12297
rect 17681 12257 17693 12291
rect 17727 12288 17739 12291
rect 18138 12288 18144 12300
rect 17727 12260 18144 12288
rect 17727 12257 17739 12260
rect 17681 12251 17739 12257
rect 18138 12248 18144 12260
rect 18196 12248 18202 12300
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12189 14519 12223
rect 14461 12183 14519 12189
rect 14918 12180 14924 12232
rect 14976 12220 14982 12232
rect 17402 12220 17408 12232
rect 14976 12192 17408 12220
rect 14976 12180 14982 12192
rect 17402 12180 17408 12192
rect 17460 12180 17466 12232
rect 17770 12180 17776 12232
rect 17828 12220 17834 12232
rect 17865 12223 17923 12229
rect 17865 12220 17877 12223
rect 17828 12192 17877 12220
rect 17828 12180 17834 12192
rect 17865 12189 17877 12192
rect 17911 12189 17923 12223
rect 17865 12183 17923 12189
rect 2038 12112 2044 12164
rect 2096 12152 2102 12164
rect 2409 12155 2467 12161
rect 2409 12152 2421 12155
rect 2096 12124 2421 12152
rect 2096 12112 2102 12124
rect 2409 12121 2421 12124
rect 2455 12121 2467 12155
rect 2590 12152 2596 12164
rect 2551 12124 2596 12152
rect 2409 12115 2467 12121
rect 2590 12112 2596 12124
rect 2648 12112 2654 12164
rect 2869 12155 2927 12161
rect 2869 12121 2881 12155
rect 2915 12152 2927 12155
rect 4056 12155 4114 12161
rect 2915 12124 4016 12152
rect 2915 12121 2927 12124
rect 2869 12115 2927 12121
rect 1486 12084 1492 12096
rect 1447 12056 1492 12084
rect 1486 12044 1492 12056
rect 1544 12044 1550 12096
rect 1762 12084 1768 12096
rect 1723 12056 1768 12084
rect 1762 12044 1768 12056
rect 1820 12044 1826 12096
rect 1946 12084 1952 12096
rect 1907 12056 1952 12084
rect 1946 12044 1952 12056
rect 2004 12044 2010 12096
rect 3602 12084 3608 12096
rect 3563 12056 3608 12084
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 3988 12084 4016 12124
rect 4056 12121 4068 12155
rect 4102 12152 4114 12155
rect 4154 12152 4160 12164
rect 4102 12124 4160 12152
rect 4102 12121 4114 12124
rect 4056 12115 4114 12121
rect 4154 12112 4160 12124
rect 4212 12112 4218 12164
rect 4246 12112 4252 12164
rect 4304 12152 4310 12164
rect 4522 12152 4528 12164
rect 4304 12124 4528 12152
rect 4304 12112 4310 12124
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 6730 12112 6736 12164
rect 6788 12152 6794 12164
rect 7193 12155 7251 12161
rect 7193 12152 7205 12155
rect 6788 12124 7205 12152
rect 6788 12112 6794 12124
rect 7193 12121 7205 12124
rect 7239 12152 7251 12155
rect 9490 12152 9496 12164
rect 7239 12124 9496 12152
rect 7239 12121 7251 12124
rect 7193 12115 7251 12121
rect 9490 12112 9496 12124
rect 9548 12112 9554 12164
rect 9677 12155 9735 12161
rect 9677 12121 9689 12155
rect 9723 12152 9735 12155
rect 12078 12155 12136 12161
rect 9723 12124 10180 12152
rect 9723 12121 9735 12124
rect 9677 12115 9735 12121
rect 5258 12084 5264 12096
rect 3988 12056 5264 12084
rect 5258 12044 5264 12056
rect 5316 12044 5322 12096
rect 5718 12084 5724 12096
rect 5679 12056 5724 12084
rect 5718 12044 5724 12056
rect 5776 12044 5782 12096
rect 5813 12087 5871 12093
rect 5813 12053 5825 12087
rect 5859 12084 5871 12087
rect 6546 12084 6552 12096
rect 5859 12056 6552 12084
rect 5859 12053 5871 12056
rect 5813 12047 5871 12053
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 6641 12087 6699 12093
rect 6641 12053 6653 12087
rect 6687 12084 6699 12087
rect 6822 12084 6828 12096
rect 6687 12056 6828 12084
rect 6687 12053 6699 12056
rect 6641 12047 6699 12053
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 8938 12044 8944 12096
rect 8996 12084 9002 12096
rect 9309 12087 9367 12093
rect 9309 12084 9321 12087
rect 8996 12056 9321 12084
rect 8996 12044 9002 12056
rect 9309 12053 9321 12056
rect 9355 12053 9367 12087
rect 9309 12047 9367 12053
rect 9766 12044 9772 12096
rect 9824 12084 9830 12096
rect 10152 12093 10180 12124
rect 12078 12121 12090 12155
rect 12124 12121 12136 12155
rect 12078 12115 12136 12121
rect 13081 12155 13139 12161
rect 13081 12121 13093 12155
rect 13127 12152 13139 12155
rect 13541 12155 13599 12161
rect 13541 12152 13553 12155
rect 13127 12124 13553 12152
rect 13127 12121 13139 12124
rect 13081 12115 13139 12121
rect 13541 12121 13553 12124
rect 13587 12121 13599 12155
rect 13541 12115 13599 12121
rect 10137 12087 10195 12093
rect 9824 12056 9869 12084
rect 9824 12044 9830 12056
rect 10137 12053 10149 12087
rect 10183 12053 10195 12087
rect 10137 12047 10195 12053
rect 10594 12044 10600 12096
rect 10652 12084 10658 12096
rect 10652 12056 10697 12084
rect 10652 12044 10658 12056
rect 10778 12044 10784 12096
rect 10836 12084 10842 12096
rect 11514 12084 11520 12096
rect 10836 12056 11520 12084
rect 10836 12044 10842 12056
rect 11514 12044 11520 12056
rect 11572 12044 11578 12096
rect 11698 12044 11704 12096
rect 11756 12084 11762 12096
rect 12084 12084 12112 12115
rect 14182 12112 14188 12164
rect 14240 12152 14246 12164
rect 17160 12155 17218 12161
rect 14240 12124 14504 12152
rect 14240 12112 14246 12124
rect 14090 12084 14096 12096
rect 11756 12056 12112 12084
rect 14051 12056 14096 12084
rect 11756 12044 11762 12056
rect 14090 12044 14096 12056
rect 14148 12044 14154 12096
rect 14476 12084 14504 12124
rect 17160 12121 17172 12155
rect 17206 12152 17218 12155
rect 17310 12152 17316 12164
rect 17206 12124 17316 12152
rect 17206 12121 17218 12124
rect 17160 12115 17218 12121
rect 17310 12112 17316 12124
rect 17368 12112 17374 12164
rect 18325 12155 18383 12161
rect 18325 12152 18337 12155
rect 17788 12124 18337 12152
rect 14553 12087 14611 12093
rect 14553 12084 14565 12087
rect 14476 12056 14565 12084
rect 14553 12053 14565 12056
rect 14599 12053 14611 12087
rect 14553 12047 14611 12053
rect 14642 12044 14648 12096
rect 14700 12084 14706 12096
rect 14921 12087 14979 12093
rect 14921 12084 14933 12087
rect 14700 12056 14933 12084
rect 14700 12044 14706 12056
rect 14921 12053 14933 12056
rect 14967 12053 14979 12087
rect 14921 12047 14979 12053
rect 15194 12044 15200 12096
rect 15252 12084 15258 12096
rect 15289 12087 15347 12093
rect 15289 12084 15301 12087
rect 15252 12056 15301 12084
rect 15252 12044 15258 12056
rect 15289 12053 15301 12056
rect 15335 12053 15347 12087
rect 15289 12047 15347 12053
rect 16482 12044 16488 12096
rect 16540 12084 16546 12096
rect 17788 12093 17816 12124
rect 18325 12121 18337 12124
rect 18371 12152 18383 12155
rect 18414 12152 18420 12164
rect 18371 12124 18420 12152
rect 18371 12121 18383 12124
rect 18325 12115 18383 12121
rect 18414 12112 18420 12124
rect 18472 12112 18478 12164
rect 17773 12087 17831 12093
rect 17773 12084 17785 12087
rect 16540 12056 17785 12084
rect 16540 12044 16546 12056
rect 17773 12053 17785 12056
rect 17819 12053 17831 12087
rect 17773 12047 17831 12053
rect 17862 12044 17868 12096
rect 17920 12084 17926 12096
rect 18233 12087 18291 12093
rect 18233 12084 18245 12087
rect 17920 12056 18245 12084
rect 17920 12044 17926 12056
rect 18233 12053 18245 12056
rect 18279 12053 18291 12087
rect 18233 12047 18291 12053
rect 1104 11994 18860 12016
rect 1104 11942 5398 11994
rect 5450 11942 5462 11994
rect 5514 11942 5526 11994
rect 5578 11942 5590 11994
rect 5642 11942 5654 11994
rect 5706 11942 9846 11994
rect 9898 11942 9910 11994
rect 9962 11942 9974 11994
rect 10026 11942 10038 11994
rect 10090 11942 10102 11994
rect 10154 11942 14294 11994
rect 14346 11942 14358 11994
rect 14410 11942 14422 11994
rect 14474 11942 14486 11994
rect 14538 11942 14550 11994
rect 14602 11942 18860 11994
rect 1104 11920 18860 11942
rect 2501 11883 2559 11889
rect 2501 11849 2513 11883
rect 2547 11880 2559 11883
rect 2682 11880 2688 11892
rect 2547 11852 2688 11880
rect 2547 11849 2559 11852
rect 2501 11843 2559 11849
rect 2682 11840 2688 11852
rect 2740 11880 2746 11892
rect 4246 11880 4252 11892
rect 2740 11852 4252 11880
rect 2740 11840 2746 11852
rect 4246 11840 4252 11852
rect 4304 11840 4310 11892
rect 5718 11840 5724 11892
rect 5776 11880 5782 11892
rect 6365 11883 6423 11889
rect 6365 11880 6377 11883
rect 5776 11852 6377 11880
rect 5776 11840 5782 11852
rect 6365 11849 6377 11852
rect 6411 11849 6423 11883
rect 6365 11843 6423 11849
rect 6546 11840 6552 11892
rect 6604 11880 6610 11892
rect 7193 11883 7251 11889
rect 7193 11880 7205 11883
rect 6604 11852 7205 11880
rect 6604 11840 6610 11852
rect 7193 11849 7205 11852
rect 7239 11849 7251 11883
rect 7193 11843 7251 11849
rect 7650 11840 7656 11892
rect 7708 11880 7714 11892
rect 8481 11883 8539 11889
rect 7708 11852 8432 11880
rect 7708 11840 7714 11852
rect 1670 11772 1676 11824
rect 1728 11812 1734 11824
rect 1946 11812 1952 11824
rect 1728 11784 1952 11812
rect 1728 11772 1734 11784
rect 1946 11772 1952 11784
rect 2004 11812 2010 11824
rect 3053 11815 3111 11821
rect 3053 11812 3065 11815
rect 2004 11784 3065 11812
rect 2004 11772 2010 11784
rect 3053 11781 3065 11784
rect 3099 11812 3111 11815
rect 3510 11812 3516 11824
rect 3099 11784 3516 11812
rect 3099 11781 3111 11784
rect 3053 11775 3111 11781
rect 3510 11772 3516 11784
rect 3568 11772 3574 11824
rect 3973 11815 4031 11821
rect 3973 11781 3985 11815
rect 4019 11812 4031 11815
rect 4062 11812 4068 11824
rect 4019 11784 4068 11812
rect 4019 11781 4031 11784
rect 3973 11775 4031 11781
rect 4062 11772 4068 11784
rect 4120 11772 4126 11824
rect 4332 11815 4390 11821
rect 4332 11781 4344 11815
rect 4378 11812 4390 11815
rect 6181 11815 6239 11821
rect 6181 11812 6193 11815
rect 4378 11784 6193 11812
rect 4378 11781 4390 11784
rect 4332 11775 4390 11781
rect 6181 11781 6193 11784
rect 6227 11781 6239 11815
rect 6181 11775 6239 11781
rect 6840 11784 8340 11812
rect 1489 11747 1547 11753
rect 1489 11713 1501 11747
rect 1535 11744 1547 11747
rect 1578 11744 1584 11756
rect 1535 11716 1584 11744
rect 1535 11713 1547 11716
rect 1489 11707 1547 11713
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11744 3019 11747
rect 3694 11744 3700 11756
rect 3007 11716 3700 11744
rect 3007 11713 3019 11716
rect 2961 11707 3019 11713
rect 3694 11704 3700 11716
rect 3752 11704 3758 11756
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 4764 11716 5120 11744
rect 4764 11704 4770 11716
rect 2133 11679 2191 11685
rect 2133 11645 2145 11679
rect 2179 11676 2191 11679
rect 2222 11676 2228 11688
rect 2179 11648 2228 11676
rect 2179 11645 2191 11648
rect 2133 11639 2191 11645
rect 2222 11636 2228 11648
rect 2280 11636 2286 11688
rect 3237 11679 3295 11685
rect 3237 11645 3249 11679
rect 3283 11676 3295 11679
rect 3510 11676 3516 11688
rect 3283 11648 3516 11676
rect 3283 11645 3295 11648
rect 3237 11639 3295 11645
rect 3510 11636 3516 11648
rect 3568 11636 3574 11688
rect 3786 11636 3792 11688
rect 3844 11676 3850 11688
rect 4062 11676 4068 11688
rect 3844 11648 4068 11676
rect 3844 11636 3850 11648
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 5092 11676 5120 11716
rect 5166 11704 5172 11756
rect 5224 11744 5230 11756
rect 5537 11747 5595 11753
rect 5537 11744 5549 11747
rect 5224 11716 5549 11744
rect 5224 11704 5230 11716
rect 5537 11713 5549 11716
rect 5583 11713 5595 11747
rect 6730 11744 6736 11756
rect 6643 11716 6736 11744
rect 5537 11707 5595 11713
rect 6656 11676 6684 11716
rect 6730 11704 6736 11716
rect 6788 11704 6794 11756
rect 6840 11688 6868 11784
rect 7561 11747 7619 11753
rect 7561 11744 7573 11747
rect 6932 11716 7573 11744
rect 6822 11676 6828 11688
rect 5092 11648 6684 11676
rect 6783 11648 6828 11676
rect 6822 11636 6828 11648
rect 6880 11636 6886 11688
rect 6730 11568 6736 11620
rect 6788 11608 6794 11620
rect 6932 11608 6960 11716
rect 7561 11713 7573 11716
rect 7607 11744 7619 11747
rect 8202 11744 8208 11756
rect 7607 11716 8208 11744
rect 7607 11713 7619 11716
rect 7561 11707 7619 11713
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 7006 11636 7012 11688
rect 7064 11676 7070 11688
rect 7064 11648 7157 11676
rect 7064 11636 7070 11648
rect 7190 11636 7196 11688
rect 7248 11676 7254 11688
rect 7650 11676 7656 11688
rect 7248 11648 7656 11676
rect 7248 11636 7254 11648
rect 7650 11636 7656 11648
rect 7708 11636 7714 11688
rect 7745 11679 7803 11685
rect 7745 11645 7757 11679
rect 7791 11645 7803 11679
rect 7745 11639 7803 11645
rect 6788 11580 6960 11608
rect 7024 11608 7052 11636
rect 7760 11608 7788 11639
rect 7024 11580 7788 11608
rect 6788 11568 6794 11580
rect 2038 11500 2044 11552
rect 2096 11540 2102 11552
rect 2225 11543 2283 11549
rect 2225 11540 2237 11543
rect 2096 11512 2237 11540
rect 2096 11500 2102 11512
rect 2225 11509 2237 11512
rect 2271 11509 2283 11543
rect 2225 11503 2283 11509
rect 2498 11500 2504 11552
rect 2556 11540 2562 11552
rect 2593 11543 2651 11549
rect 2593 11540 2605 11543
rect 2556 11512 2605 11540
rect 2556 11500 2562 11512
rect 2593 11509 2605 11512
rect 2639 11509 2651 11543
rect 3786 11540 3792 11552
rect 3747 11512 3792 11540
rect 2593 11503 2651 11509
rect 3786 11500 3792 11512
rect 3844 11500 3850 11552
rect 5442 11540 5448 11552
rect 5403 11512 5448 11540
rect 5442 11500 5448 11512
rect 5500 11500 5506 11552
rect 7190 11500 7196 11552
rect 7248 11540 7254 11552
rect 8113 11543 8171 11549
rect 8113 11540 8125 11543
rect 7248 11512 8125 11540
rect 7248 11500 7254 11512
rect 8113 11509 8125 11512
rect 8159 11509 8171 11543
rect 8312 11540 8340 11784
rect 8404 11744 8432 11852
rect 8481 11849 8493 11883
rect 8527 11880 8539 11883
rect 8846 11880 8852 11892
rect 8527 11852 8852 11880
rect 8527 11849 8539 11852
rect 8481 11843 8539 11849
rect 8846 11840 8852 11852
rect 8904 11840 8910 11892
rect 9398 11880 9404 11892
rect 9359 11852 9404 11880
rect 9398 11840 9404 11852
rect 9456 11840 9462 11892
rect 9766 11880 9772 11892
rect 9727 11852 9772 11880
rect 9766 11840 9772 11852
rect 9824 11840 9830 11892
rect 10229 11883 10287 11889
rect 10229 11849 10241 11883
rect 10275 11880 10287 11883
rect 10597 11883 10655 11889
rect 10597 11880 10609 11883
rect 10275 11852 10609 11880
rect 10275 11849 10287 11852
rect 10229 11843 10287 11849
rect 10597 11849 10609 11852
rect 10643 11849 10655 11883
rect 10597 11843 10655 11849
rect 10778 11840 10784 11892
rect 10836 11840 10842 11892
rect 11882 11880 11888 11892
rect 11843 11852 11888 11880
rect 11882 11840 11888 11852
rect 11940 11880 11946 11892
rect 12526 11880 12532 11892
rect 11940 11852 12532 11880
rect 11940 11840 11946 11852
rect 12526 11840 12532 11852
rect 12584 11840 12590 11892
rect 13725 11883 13783 11889
rect 13725 11849 13737 11883
rect 13771 11880 13783 11883
rect 14090 11880 14096 11892
rect 13771 11852 14096 11880
rect 13771 11849 13783 11852
rect 13725 11843 13783 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14182 11840 14188 11892
rect 14240 11880 14246 11892
rect 15194 11880 15200 11892
rect 14240 11852 14285 11880
rect 15155 11852 15200 11880
rect 14240 11840 14246 11852
rect 15194 11840 15200 11852
rect 15252 11840 15258 11892
rect 15562 11880 15568 11892
rect 15523 11852 15568 11880
rect 15562 11840 15568 11852
rect 15620 11840 15626 11892
rect 15657 11883 15715 11889
rect 15657 11849 15669 11883
rect 15703 11880 15715 11883
rect 16669 11883 16727 11889
rect 16669 11880 16681 11883
rect 15703 11852 16681 11880
rect 15703 11849 15715 11852
rect 15657 11843 15715 11849
rect 16669 11849 16681 11852
rect 16715 11849 16727 11883
rect 17494 11880 17500 11892
rect 17455 11852 17500 11880
rect 16669 11843 16727 11849
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 8573 11815 8631 11821
rect 8573 11781 8585 11815
rect 8619 11812 8631 11815
rect 8938 11812 8944 11824
rect 8619 11784 8944 11812
rect 8619 11781 8631 11784
rect 8573 11775 8631 11781
rect 8938 11772 8944 11784
rect 8996 11772 9002 11824
rect 10137 11815 10195 11821
rect 10137 11781 10149 11815
rect 10183 11812 10195 11815
rect 10796 11812 10824 11840
rect 10183 11784 10824 11812
rect 13633 11815 13691 11821
rect 10183 11781 10195 11784
rect 10137 11775 10195 11781
rect 13633 11781 13645 11815
rect 13679 11812 13691 11815
rect 14642 11812 14648 11824
rect 13679 11784 14648 11812
rect 13679 11781 13691 11784
rect 13633 11775 13691 11781
rect 14642 11772 14648 11784
rect 14700 11772 14706 11824
rect 15470 11772 15476 11824
rect 15528 11812 15534 11824
rect 16114 11812 16120 11824
rect 15528 11784 16120 11812
rect 15528 11772 15534 11784
rect 16114 11772 16120 11784
rect 16172 11812 16178 11824
rect 16209 11815 16267 11821
rect 16209 11812 16221 11815
rect 16172 11784 16221 11812
rect 16172 11772 16178 11784
rect 16209 11781 16221 11784
rect 16255 11781 16267 11815
rect 17126 11812 17132 11824
rect 17087 11784 17132 11812
rect 16209 11775 16267 11781
rect 17126 11772 17132 11784
rect 17184 11772 17190 11824
rect 8404 11716 8984 11744
rect 8754 11676 8760 11688
rect 8715 11648 8760 11676
rect 8754 11636 8760 11648
rect 8812 11636 8818 11688
rect 8956 11676 8984 11716
rect 9030 11704 9036 11756
rect 9088 11744 9094 11756
rect 9214 11744 9220 11756
rect 9088 11716 9220 11744
rect 9088 11704 9094 11716
rect 9214 11704 9220 11716
rect 9272 11744 9278 11756
rect 9309 11747 9367 11753
rect 9309 11744 9321 11747
rect 9272 11716 9321 11744
rect 9272 11704 9278 11716
rect 9309 11713 9321 11716
rect 9355 11713 9367 11747
rect 9309 11707 9367 11713
rect 9490 11704 9496 11756
rect 9548 11744 9554 11756
rect 10502 11744 10508 11756
rect 9548 11716 10508 11744
rect 9548 11704 9554 11716
rect 10502 11704 10508 11716
rect 10560 11704 10566 11756
rect 10778 11704 10784 11756
rect 10836 11744 10842 11756
rect 10965 11747 11023 11753
rect 10965 11744 10977 11747
rect 10836 11716 10977 11744
rect 10836 11704 10842 11716
rect 10965 11713 10977 11716
rect 11011 11713 11023 11747
rect 10965 11707 11023 11713
rect 11977 11747 12035 11753
rect 11977 11713 11989 11747
rect 12023 11744 12035 11747
rect 12023 11716 12388 11744
rect 12023 11713 12035 11716
rect 11977 11707 12035 11713
rect 9585 11679 9643 11685
rect 8956 11648 9076 11676
rect 8386 11568 8392 11620
rect 8444 11608 8450 11620
rect 8941 11611 8999 11617
rect 8941 11608 8953 11611
rect 8444 11580 8953 11608
rect 8444 11568 8450 11580
rect 8941 11577 8953 11580
rect 8987 11577 8999 11611
rect 9048 11608 9076 11648
rect 9585 11645 9597 11679
rect 9631 11676 9643 11679
rect 9674 11676 9680 11688
rect 9631 11648 9680 11676
rect 9631 11645 9643 11648
rect 9585 11639 9643 11645
rect 9674 11636 9680 11648
rect 9732 11676 9738 11688
rect 10321 11679 10379 11685
rect 10321 11676 10333 11679
rect 9732 11648 10333 11676
rect 9732 11636 9738 11648
rect 10321 11645 10333 11648
rect 10367 11645 10379 11679
rect 10321 11639 10379 11645
rect 10410 11636 10416 11688
rect 10468 11676 10474 11688
rect 10870 11676 10876 11688
rect 10468 11648 10876 11676
rect 10468 11636 10474 11648
rect 10870 11636 10876 11648
rect 10928 11676 10934 11688
rect 11057 11679 11115 11685
rect 11057 11676 11069 11679
rect 10928 11648 11069 11676
rect 10928 11636 10934 11648
rect 11057 11645 11069 11648
rect 11103 11645 11115 11679
rect 11057 11639 11115 11645
rect 11149 11679 11207 11685
rect 11149 11645 11161 11679
rect 11195 11676 11207 11679
rect 11698 11676 11704 11688
rect 11195 11648 11704 11676
rect 11195 11645 11207 11648
rect 11149 11639 11207 11645
rect 10134 11608 10140 11620
rect 9048 11580 10140 11608
rect 8941 11571 8999 11577
rect 10134 11568 10140 11580
rect 10192 11568 10198 11620
rect 10226 11568 10232 11620
rect 10284 11608 10290 11620
rect 11164 11608 11192 11639
rect 11698 11636 11704 11648
rect 11756 11676 11762 11688
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11756 11648 12081 11676
rect 11756 11636 11762 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 11514 11608 11520 11620
rect 10284 11580 11192 11608
rect 11475 11580 11520 11608
rect 10284 11568 10290 11580
rect 11514 11568 11520 11580
rect 11572 11568 11578 11620
rect 12360 11608 12388 11716
rect 13078 11704 13084 11756
rect 13136 11744 13142 11756
rect 13136 11716 13952 11744
rect 13136 11704 13142 11716
rect 13538 11676 13544 11688
rect 13499 11648 13544 11676
rect 13538 11636 13544 11648
rect 13596 11636 13602 11688
rect 13924 11676 13952 11716
rect 13998 11704 14004 11756
rect 14056 11744 14062 11756
rect 14553 11747 14611 11753
rect 14553 11744 14565 11747
rect 14056 11716 14565 11744
rect 14056 11704 14062 11716
rect 14553 11713 14565 11716
rect 14599 11744 14611 11747
rect 15013 11747 15071 11753
rect 15013 11744 15025 11747
rect 14599 11716 15025 11744
rect 14599 11713 14611 11716
rect 14553 11707 14611 11713
rect 15013 11713 15025 11716
rect 15059 11713 15071 11747
rect 15013 11707 15071 11713
rect 15562 11704 15568 11756
rect 15620 11744 15626 11756
rect 16025 11747 16083 11753
rect 16025 11744 16037 11747
rect 15620 11716 16037 11744
rect 15620 11704 15626 11716
rect 16025 11713 16037 11716
rect 16071 11713 16083 11747
rect 16025 11707 16083 11713
rect 16850 11704 16856 11756
rect 16908 11744 16914 11756
rect 17037 11747 17095 11753
rect 17037 11744 17049 11747
rect 16908 11716 17049 11744
rect 16908 11704 16914 11716
rect 17037 11713 17049 11716
rect 17083 11713 17095 11747
rect 17770 11744 17776 11756
rect 17037 11707 17095 11713
rect 17135 11716 17776 11744
rect 14645 11679 14703 11685
rect 14645 11676 14657 11679
rect 13924 11648 14657 11676
rect 14645 11645 14657 11648
rect 14691 11645 14703 11679
rect 14645 11639 14703 11645
rect 14458 11608 14464 11620
rect 12360 11580 14464 11608
rect 12360 11549 12388 11580
rect 14458 11568 14464 11580
rect 14516 11568 14522 11620
rect 14660 11608 14688 11639
rect 14734 11636 14740 11688
rect 14792 11676 14798 11688
rect 15749 11679 15807 11685
rect 15749 11676 15761 11679
rect 14792 11648 15761 11676
rect 14792 11636 14798 11648
rect 15749 11645 15761 11648
rect 15795 11645 15807 11679
rect 15749 11639 15807 11645
rect 16206 11636 16212 11688
rect 16264 11676 16270 11688
rect 17135 11676 17163 11716
rect 17770 11704 17776 11716
rect 17828 11744 17834 11756
rect 17865 11747 17923 11753
rect 17865 11744 17877 11747
rect 17828 11716 17877 11744
rect 17828 11704 17834 11716
rect 17865 11713 17877 11716
rect 17911 11713 17923 11747
rect 17865 11707 17923 11713
rect 17957 11747 18015 11753
rect 17957 11713 17969 11747
rect 18003 11744 18015 11747
rect 18325 11747 18383 11753
rect 18325 11744 18337 11747
rect 18003 11716 18337 11744
rect 18003 11713 18015 11716
rect 17957 11707 18015 11713
rect 17310 11676 17316 11688
rect 16264 11648 17163 11676
rect 17271 11648 17316 11676
rect 16264 11636 16270 11648
rect 17310 11636 17316 11648
rect 17368 11636 17374 11688
rect 18049 11679 18107 11685
rect 18049 11645 18061 11679
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 15470 11608 15476 11620
rect 14660 11580 15476 11608
rect 15470 11568 15476 11580
rect 15528 11568 15534 11620
rect 16114 11568 16120 11620
rect 16172 11608 16178 11620
rect 16485 11611 16543 11617
rect 16485 11608 16497 11611
rect 16172 11580 16497 11608
rect 16172 11568 16178 11580
rect 16485 11577 16497 11580
rect 16531 11608 16543 11611
rect 17126 11608 17132 11620
rect 16531 11580 17132 11608
rect 16531 11577 16543 11580
rect 16485 11571 16543 11577
rect 17126 11568 17132 11580
rect 17184 11568 17190 11620
rect 17328 11608 17356 11636
rect 18064 11608 18092 11639
rect 17328 11580 18092 11608
rect 12345 11543 12403 11549
rect 12345 11540 12357 11543
rect 8312 11512 12357 11540
rect 8113 11503 8171 11509
rect 12345 11509 12357 11512
rect 12391 11509 12403 11543
rect 12345 11503 12403 11509
rect 12989 11543 13047 11549
rect 12989 11509 13001 11543
rect 13035 11540 13047 11543
rect 13078 11540 13084 11552
rect 13035 11512 13084 11540
rect 13035 11509 13047 11512
rect 12989 11503 13047 11509
rect 13078 11500 13084 11512
rect 13136 11500 13142 11552
rect 13262 11540 13268 11552
rect 13223 11512 13268 11540
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 14090 11540 14096 11552
rect 14051 11512 14096 11540
rect 14090 11500 14096 11512
rect 14148 11500 14154 11552
rect 16390 11500 16396 11552
rect 16448 11540 16454 11552
rect 18156 11540 18184 11716
rect 18325 11713 18337 11716
rect 18371 11713 18383 11747
rect 18325 11707 18383 11713
rect 16448 11512 18184 11540
rect 16448 11500 16454 11512
rect 1104 11450 18860 11472
rect 1104 11398 3174 11450
rect 3226 11398 3238 11450
rect 3290 11398 3302 11450
rect 3354 11398 3366 11450
rect 3418 11398 3430 11450
rect 3482 11398 7622 11450
rect 7674 11398 7686 11450
rect 7738 11398 7750 11450
rect 7802 11398 7814 11450
rect 7866 11398 7878 11450
rect 7930 11398 12070 11450
rect 12122 11398 12134 11450
rect 12186 11398 12198 11450
rect 12250 11398 12262 11450
rect 12314 11398 12326 11450
rect 12378 11398 16518 11450
rect 16570 11398 16582 11450
rect 16634 11398 16646 11450
rect 16698 11398 16710 11450
rect 16762 11398 16774 11450
rect 16826 11398 18860 11450
rect 1104 11376 18860 11398
rect 2038 11296 2044 11348
rect 2096 11336 2102 11348
rect 6181 11339 6239 11345
rect 6181 11336 6193 11339
rect 2096 11308 6193 11336
rect 2096 11296 2102 11308
rect 6181 11305 6193 11308
rect 6227 11336 6239 11339
rect 6822 11336 6828 11348
rect 6227 11308 6828 11336
rect 6227 11305 6239 11308
rect 6181 11299 6239 11305
rect 6822 11296 6828 11308
rect 6880 11296 6886 11348
rect 7466 11296 7472 11348
rect 7524 11336 7530 11348
rect 8757 11339 8815 11345
rect 7524 11308 7972 11336
rect 7524 11296 7530 11308
rect 7944 11280 7972 11308
rect 8757 11305 8769 11339
rect 8803 11336 8815 11339
rect 8846 11336 8852 11348
rect 8803 11308 8852 11336
rect 8803 11305 8815 11308
rect 8757 11299 8815 11305
rect 8846 11296 8852 11308
rect 8904 11296 8910 11348
rect 9398 11336 9404 11348
rect 9359 11308 9404 11336
rect 9398 11296 9404 11308
rect 9456 11296 9462 11348
rect 9585 11339 9643 11345
rect 9585 11305 9597 11339
rect 9631 11336 9643 11339
rect 10226 11336 10232 11348
rect 9631 11308 10232 11336
rect 9631 11305 9643 11308
rect 9585 11299 9643 11305
rect 10226 11296 10232 11308
rect 10284 11296 10290 11348
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 11149 11339 11207 11345
rect 11149 11336 11161 11339
rect 10652 11308 11161 11336
rect 10652 11296 10658 11308
rect 11149 11305 11161 11308
rect 11195 11305 11207 11339
rect 11149 11299 11207 11305
rect 11698 11296 11704 11348
rect 11756 11336 11762 11348
rect 11756 11308 12112 11336
rect 11756 11296 11762 11308
rect 4154 11268 4160 11280
rect 4115 11240 4160 11268
rect 4154 11228 4160 11240
rect 4212 11268 4218 11280
rect 4338 11268 4344 11280
rect 4212 11240 4344 11268
rect 4212 11228 4218 11240
rect 4338 11228 4344 11240
rect 4396 11228 4402 11280
rect 6270 11228 6276 11280
rect 6328 11268 6334 11280
rect 6328 11240 6592 11268
rect 6328 11228 6334 11240
rect 3694 11160 3700 11212
rect 3752 11200 3758 11212
rect 3789 11203 3847 11209
rect 3789 11200 3801 11203
rect 3752 11172 3801 11200
rect 3752 11160 3758 11172
rect 3789 11169 3801 11172
rect 3835 11169 3847 11203
rect 3789 11163 3847 11169
rect 3878 11160 3884 11212
rect 3936 11200 3942 11212
rect 5997 11203 6055 11209
rect 3936 11172 4752 11200
rect 3936 11160 3942 11172
rect 2133 11135 2191 11141
rect 2133 11101 2145 11135
rect 2179 11101 2191 11135
rect 2133 11095 2191 11101
rect 1489 11067 1547 11073
rect 1489 11033 1501 11067
rect 1535 11064 1547 11067
rect 1946 11064 1952 11076
rect 1535 11036 1952 11064
rect 1535 11033 1547 11036
rect 1489 11027 1547 11033
rect 1946 11024 1952 11036
rect 2004 11024 2010 11076
rect 2148 11064 2176 11095
rect 2774 11092 2780 11144
rect 2832 11132 2838 11144
rect 3605 11135 3663 11141
rect 3605 11132 3617 11135
rect 2832 11104 3617 11132
rect 2832 11092 2838 11104
rect 3605 11101 3617 11104
rect 3651 11132 3663 11135
rect 4062 11132 4068 11144
rect 3651 11104 4068 11132
rect 3651 11101 3663 11104
rect 3605 11095 3663 11101
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 4724 11132 4752 11172
rect 5997 11169 6009 11203
rect 6043 11200 6055 11203
rect 6362 11200 6368 11212
rect 6043 11172 6368 11200
rect 6043 11169 6055 11172
rect 5997 11163 6055 11169
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 6564 11200 6592 11240
rect 6638 11228 6644 11280
rect 6696 11268 6702 11280
rect 7561 11271 7619 11277
rect 7561 11268 7573 11271
rect 6696 11240 7573 11268
rect 6696 11228 6702 11240
rect 7561 11237 7573 11240
rect 7607 11237 7619 11271
rect 7561 11231 7619 11237
rect 7926 11228 7932 11280
rect 7984 11268 7990 11280
rect 9214 11268 9220 11280
rect 7984 11240 9220 11268
rect 7984 11228 7990 11240
rect 9214 11228 9220 11240
rect 9272 11228 9278 11280
rect 6730 11200 6736 11212
rect 6564 11172 6736 11200
rect 6730 11160 6736 11172
rect 6788 11200 6794 11212
rect 7193 11203 7251 11209
rect 6788 11172 7144 11200
rect 6788 11160 6794 11172
rect 5721 11135 5779 11141
rect 4724 11104 5672 11132
rect 2958 11064 2964 11076
rect 2148 11036 2964 11064
rect 2958 11024 2964 11036
rect 3016 11024 3022 11076
rect 3360 11067 3418 11073
rect 3360 11033 3372 11067
rect 3406 11064 3418 11067
rect 3510 11064 3516 11076
rect 3406 11036 3516 11064
rect 3406 11033 3418 11036
rect 3360 11027 3418 11033
rect 3510 11024 3516 11036
rect 3568 11064 3574 11076
rect 3568 11036 4384 11064
rect 3568 11024 3574 11036
rect 2225 10999 2283 11005
rect 2225 10965 2237 10999
rect 2271 10996 2283 10999
rect 2498 10996 2504 11008
rect 2271 10968 2504 10996
rect 2271 10965 2283 10968
rect 2225 10959 2283 10965
rect 2498 10956 2504 10968
rect 2556 10956 2562 11008
rect 4356 11005 4384 11036
rect 4982 11024 4988 11076
rect 5040 11064 5046 11076
rect 5442 11064 5448 11076
rect 5500 11073 5506 11076
rect 5040 11036 5448 11064
rect 5040 11024 5046 11036
rect 5442 11024 5448 11036
rect 5500 11027 5512 11073
rect 5644 11064 5672 11104
rect 5721 11101 5733 11135
rect 5767 11132 5779 11135
rect 6822 11132 6828 11144
rect 5767 11104 6828 11132
rect 5767 11101 5779 11104
rect 5721 11095 5779 11101
rect 6822 11092 6828 11104
rect 6880 11092 6886 11144
rect 6086 11064 6092 11076
rect 5644 11036 6092 11064
rect 5500 11024 5506 11027
rect 6086 11024 6092 11036
rect 6144 11024 6150 11076
rect 6454 11064 6460 11076
rect 6415 11036 6460 11064
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 7006 11064 7012 11076
rect 6967 11036 7012 11064
rect 7006 11024 7012 11036
rect 7064 11024 7070 11076
rect 7116 11064 7144 11172
rect 7193 11169 7205 11203
rect 7239 11169 7251 11203
rect 8110 11200 8116 11212
rect 8071 11172 8116 11200
rect 7193 11163 7251 11169
rect 7208 11132 7236 11163
rect 8110 11160 8116 11172
rect 8168 11160 8174 11212
rect 8202 11160 8208 11212
rect 8260 11200 8266 11212
rect 9950 11200 9956 11212
rect 8260 11172 9956 11200
rect 8260 11160 8266 11172
rect 9950 11160 9956 11172
rect 10008 11160 10014 11212
rect 11238 11160 11244 11212
rect 11296 11200 11302 11212
rect 11793 11203 11851 11209
rect 11296 11172 11652 11200
rect 11296 11160 11302 11172
rect 11624 11144 11652 11172
rect 11793 11169 11805 11203
rect 11839 11200 11851 11203
rect 12084 11200 12112 11308
rect 14458 11296 14464 11348
rect 14516 11336 14522 11348
rect 16301 11339 16359 11345
rect 14516 11308 15884 11336
rect 14516 11296 14522 11308
rect 12345 11271 12403 11277
rect 12345 11237 12357 11271
rect 12391 11268 12403 11271
rect 12618 11268 12624 11280
rect 12391 11240 12624 11268
rect 12391 11237 12403 11240
rect 12345 11231 12403 11237
rect 12618 11228 12624 11240
rect 12676 11228 12682 11280
rect 13173 11271 13231 11277
rect 13173 11268 13185 11271
rect 12728 11240 13185 11268
rect 11839 11172 12112 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 8570 11132 8576 11144
rect 7208 11104 8576 11132
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 10965 11135 11023 11141
rect 10965 11101 10977 11135
rect 11011 11132 11023 11135
rect 11514 11132 11520 11144
rect 11011 11104 11520 11132
rect 11011 11101 11023 11104
rect 10965 11095 11023 11101
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 11606 11092 11612 11144
rect 11664 11132 11670 11144
rect 12728 11141 12756 11240
rect 13173 11237 13185 11240
rect 13219 11237 13231 11271
rect 15856 11268 15884 11308
rect 16301 11305 16313 11339
rect 16347 11336 16359 11339
rect 17310 11336 17316 11348
rect 16347 11308 17316 11336
rect 16347 11305 16359 11308
rect 16301 11299 16359 11305
rect 17310 11296 17316 11308
rect 17368 11296 17374 11348
rect 17770 11296 17776 11348
rect 17828 11336 17834 11348
rect 18325 11339 18383 11345
rect 18325 11336 18337 11339
rect 17828 11308 18337 11336
rect 17828 11296 17834 11308
rect 18325 11305 18337 11308
rect 18371 11305 18383 11339
rect 18325 11299 18383 11305
rect 16390 11268 16396 11280
rect 15856 11240 16396 11268
rect 13173 11231 13231 11237
rect 16390 11228 16396 11240
rect 16448 11228 16454 11280
rect 12894 11200 12900 11212
rect 12855 11172 12900 11200
rect 12894 11160 12900 11172
rect 12952 11160 12958 11212
rect 13262 11160 13268 11212
rect 13320 11200 13326 11212
rect 13633 11203 13691 11209
rect 13633 11200 13645 11203
rect 13320 11172 13645 11200
rect 13320 11160 13326 11172
rect 13633 11169 13645 11172
rect 13679 11169 13691 11203
rect 13633 11163 13691 11169
rect 13722 11160 13728 11212
rect 13780 11200 13786 11212
rect 14918 11200 14924 11212
rect 13780 11172 13825 11200
rect 14879 11172 14924 11200
rect 13780 11160 13786 11172
rect 14918 11160 14924 11172
rect 14976 11160 14982 11212
rect 12713 11135 12771 11141
rect 11664 11104 11757 11132
rect 11664 11092 11670 11104
rect 12713 11101 12725 11135
rect 12759 11101 12771 11135
rect 12713 11095 12771 11101
rect 14090 11092 14096 11144
rect 14148 11132 14154 11144
rect 14185 11135 14243 11141
rect 14185 11132 14197 11135
rect 14148 11104 14197 11132
rect 14148 11092 14154 11104
rect 14185 11101 14197 11104
rect 14231 11101 14243 11135
rect 16393 11135 16451 11141
rect 16393 11132 16405 11135
rect 14185 11095 14243 11101
rect 14936 11104 16405 11132
rect 7377 11067 7435 11073
rect 7377 11064 7389 11067
rect 7116 11036 7389 11064
rect 7377 11033 7389 11036
rect 7423 11033 7435 11067
rect 7926 11064 7932 11076
rect 7887 11036 7932 11064
rect 7377 11027 7435 11033
rect 7926 11024 7932 11036
rect 7984 11024 7990 11076
rect 8021 11067 8079 11073
rect 8021 11033 8033 11067
rect 8067 11033 8079 11067
rect 8021 11027 8079 11033
rect 4341 10999 4399 11005
rect 4341 10965 4353 10999
rect 4387 10965 4399 10999
rect 4341 10959 4399 10965
rect 4614 10956 4620 11008
rect 4672 10996 4678 11008
rect 5074 10996 5080 11008
rect 4672 10968 5080 10996
rect 4672 10956 4678 10968
rect 5074 10956 5080 10968
rect 5132 10956 5138 11008
rect 6546 10996 6552 11008
rect 6507 10968 6552 10996
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 6914 10996 6920 11008
rect 6875 10968 6920 10996
rect 6914 10956 6920 10968
rect 6972 10956 6978 11008
rect 8036 10996 8064 11027
rect 8202 11024 8208 11076
rect 8260 11064 8266 11076
rect 8389 11067 8447 11073
rect 8389 11064 8401 11067
rect 8260 11036 8401 11064
rect 8260 11024 8266 11036
rect 8389 11033 8401 11036
rect 8435 11033 8447 11067
rect 9214 11064 9220 11076
rect 9175 11036 9220 11064
rect 8389 11027 8447 11033
rect 9214 11024 9220 11036
rect 9272 11024 9278 11076
rect 10686 11064 10692 11076
rect 10744 11073 10750 11076
rect 10656 11036 10692 11064
rect 10686 11024 10692 11036
rect 10744 11027 10756 11073
rect 12250 11064 12256 11076
rect 11532 11036 12256 11064
rect 10744 11024 10750 11027
rect 8294 10996 8300 11008
rect 8036 10968 8300 10996
rect 8294 10956 8300 10968
rect 8352 10996 8358 11008
rect 8846 10996 8852 11008
rect 8352 10968 8852 10996
rect 8352 10956 8358 10968
rect 8846 10956 8852 10968
rect 8904 10956 8910 11008
rect 9030 10996 9036 11008
rect 8991 10968 9036 10996
rect 9030 10956 9036 10968
rect 9088 10956 9094 11008
rect 11532 11005 11560 11036
rect 12250 11024 12256 11036
rect 12308 11024 12314 11076
rect 13541 11067 13599 11073
rect 13541 11033 13553 11067
rect 13587 11064 13599 11067
rect 14936 11064 14964 11104
rect 16393 11101 16405 11104
rect 16439 11101 16451 11135
rect 16393 11095 16451 11101
rect 17402 11092 17408 11144
rect 17460 11132 17466 11144
rect 18049 11135 18107 11141
rect 18049 11132 18061 11135
rect 17460 11104 18061 11132
rect 17460 11092 17466 11104
rect 18049 11101 18061 11104
rect 18095 11101 18107 11135
rect 18049 11095 18107 11101
rect 18138 11092 18144 11144
rect 18196 11092 18202 11144
rect 13587 11036 14964 11064
rect 15188 11067 15246 11073
rect 13587 11033 13599 11036
rect 13541 11027 13599 11033
rect 15188 11033 15200 11067
rect 15234 11064 15246 11067
rect 15286 11064 15292 11076
rect 15234 11036 15292 11064
rect 15234 11033 15246 11036
rect 15188 11027 15246 11033
rect 15286 11024 15292 11036
rect 15344 11024 15350 11076
rect 17804 11067 17862 11073
rect 17804 11033 17816 11067
rect 17850 11064 17862 11067
rect 18156 11064 18184 11092
rect 17850 11036 18184 11064
rect 17850 11033 17862 11036
rect 17804 11027 17862 11033
rect 11517 10999 11575 11005
rect 11517 10965 11529 10999
rect 11563 10965 11575 10999
rect 11517 10959 11575 10965
rect 11882 10956 11888 11008
rect 11940 10996 11946 11008
rect 11977 10999 12035 11005
rect 11977 10996 11989 10999
rect 11940 10968 11989 10996
rect 11940 10956 11946 10968
rect 11977 10965 11989 10968
rect 12023 10965 12035 10999
rect 12802 10996 12808 11008
rect 12763 10968 12808 10996
rect 11977 10959 12035 10965
rect 12802 10956 12808 10968
rect 12860 10956 12866 11008
rect 14826 10996 14832 11008
rect 14787 10968 14832 10996
rect 14826 10956 14832 10968
rect 14884 10956 14890 11008
rect 16666 10996 16672 11008
rect 16627 10968 16672 10996
rect 16666 10956 16672 10968
rect 16724 10956 16730 11008
rect 16850 10956 16856 11008
rect 16908 10996 16914 11008
rect 17678 10996 17684 11008
rect 16908 10968 17684 10996
rect 16908 10956 16914 10968
rect 17678 10956 17684 10968
rect 17736 10996 17742 11008
rect 18141 10999 18199 11005
rect 18141 10996 18153 10999
rect 17736 10968 18153 10996
rect 17736 10956 17742 10968
rect 18141 10965 18153 10968
rect 18187 10965 18199 10999
rect 18141 10959 18199 10965
rect 1104 10906 18860 10928
rect 1104 10854 5398 10906
rect 5450 10854 5462 10906
rect 5514 10854 5526 10906
rect 5578 10854 5590 10906
rect 5642 10854 5654 10906
rect 5706 10854 9846 10906
rect 9898 10854 9910 10906
rect 9962 10854 9974 10906
rect 10026 10854 10038 10906
rect 10090 10854 10102 10906
rect 10154 10854 14294 10906
rect 14346 10854 14358 10906
rect 14410 10854 14422 10906
rect 14474 10854 14486 10906
rect 14538 10854 14550 10906
rect 14602 10854 18860 10906
rect 1104 10832 18860 10854
rect 3237 10795 3295 10801
rect 3237 10761 3249 10795
rect 3283 10792 3295 10795
rect 4154 10792 4160 10804
rect 3283 10764 4160 10792
rect 3283 10761 3295 10764
rect 3237 10755 3295 10761
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4341 10795 4399 10801
rect 4341 10761 4353 10795
rect 4387 10792 4399 10795
rect 4709 10795 4767 10801
rect 4709 10792 4721 10795
rect 4387 10764 4721 10792
rect 4387 10761 4399 10764
rect 4341 10755 4399 10761
rect 4709 10761 4721 10764
rect 4755 10761 4767 10795
rect 4709 10755 4767 10761
rect 4798 10752 4804 10804
rect 4856 10792 4862 10804
rect 5169 10795 5227 10801
rect 5169 10792 5181 10795
rect 4856 10764 5181 10792
rect 4856 10752 4862 10764
rect 5169 10761 5181 10764
rect 5215 10792 5227 10795
rect 6362 10792 6368 10804
rect 5215 10764 6368 10792
rect 5215 10761 5227 10764
rect 5169 10755 5227 10761
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 6638 10792 6644 10804
rect 6599 10764 6644 10792
rect 6638 10752 6644 10764
rect 6696 10752 6702 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7101 10795 7159 10801
rect 7101 10792 7113 10795
rect 6972 10764 7113 10792
rect 6972 10752 6978 10764
rect 7101 10761 7113 10764
rect 7147 10761 7159 10795
rect 8294 10792 8300 10804
rect 7101 10755 7159 10761
rect 7208 10764 8300 10792
rect 2498 10684 2504 10736
rect 2556 10733 2562 10736
rect 2556 10724 2568 10733
rect 2556 10696 2601 10724
rect 2556 10687 2568 10696
rect 2556 10684 2562 10687
rect 4614 10684 4620 10736
rect 4672 10724 4678 10736
rect 4890 10724 4896 10736
rect 4672 10696 4896 10724
rect 4672 10684 4678 10696
rect 4890 10684 4896 10696
rect 4948 10724 4954 10736
rect 5077 10727 5135 10733
rect 5077 10724 5089 10727
rect 4948 10696 5089 10724
rect 4948 10684 4954 10696
rect 5077 10693 5089 10696
rect 5123 10724 5135 10727
rect 6454 10724 6460 10736
rect 5123 10696 6460 10724
rect 5123 10693 5135 10696
rect 5077 10687 5135 10693
rect 6454 10684 6460 10696
rect 6512 10684 6518 10736
rect 7208 10724 7236 10764
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 8570 10792 8576 10804
rect 8531 10764 8576 10792
rect 8570 10752 8576 10764
rect 8628 10792 8634 10804
rect 8628 10764 10180 10792
rect 8628 10752 8634 10764
rect 6656 10696 7236 10724
rect 6656 10668 6684 10696
rect 7374 10684 7380 10736
rect 7432 10724 7438 10736
rect 7432 10696 8708 10724
rect 7432 10684 7438 10696
rect 4154 10616 4160 10668
rect 4212 10656 4218 10668
rect 4249 10659 4307 10665
rect 4249 10656 4261 10659
rect 4212 10628 4261 10656
rect 4212 10616 4218 10628
rect 4249 10625 4261 10628
rect 4295 10656 4307 10659
rect 4338 10656 4344 10668
rect 4295 10628 4344 10656
rect 4295 10625 4307 10628
rect 4249 10619 4307 10625
rect 4338 10616 4344 10628
rect 4396 10616 4402 10668
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 6181 10659 6239 10665
rect 6181 10656 6193 10659
rect 5960 10628 6193 10656
rect 5960 10616 5966 10628
rect 6181 10625 6193 10628
rect 6227 10625 6239 10659
rect 6181 10619 6239 10625
rect 6638 10616 6644 10668
rect 6696 10616 6702 10668
rect 6733 10659 6791 10665
rect 6733 10625 6745 10659
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 2832 10560 2877 10588
rect 2832 10548 2838 10560
rect 3050 10548 3056 10600
rect 3108 10588 3114 10600
rect 3329 10591 3387 10597
rect 3329 10588 3341 10591
rect 3108 10560 3341 10588
rect 3108 10548 3114 10560
rect 3329 10557 3341 10560
rect 3375 10557 3387 10591
rect 3510 10588 3516 10600
rect 3471 10560 3516 10588
rect 3329 10551 3387 10557
rect 3510 10548 3516 10560
rect 3568 10588 3574 10600
rect 4433 10591 4491 10597
rect 4433 10588 4445 10591
rect 3568 10560 4445 10588
rect 3568 10548 3574 10560
rect 4433 10557 4445 10560
rect 4479 10557 4491 10591
rect 4433 10551 4491 10557
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10557 5319 10591
rect 5261 10551 5319 10557
rect 6549 10591 6607 10597
rect 6549 10557 6561 10591
rect 6595 10557 6607 10591
rect 6748 10588 6776 10619
rect 6822 10616 6828 10668
rect 6880 10656 6886 10668
rect 7193 10659 7251 10665
rect 7193 10656 7205 10659
rect 6880 10628 7205 10656
rect 6880 10616 6886 10628
rect 7193 10625 7205 10628
rect 7239 10656 7251 10659
rect 7392 10656 7420 10684
rect 7466 10665 7472 10668
rect 7239 10628 7420 10656
rect 7239 10625 7251 10628
rect 7193 10619 7251 10625
rect 7460 10619 7472 10665
rect 7524 10656 7530 10668
rect 8680 10665 8708 10696
rect 10152 10665 10180 10764
rect 10686 10752 10692 10804
rect 10744 10792 10750 10804
rect 10781 10795 10839 10801
rect 10781 10792 10793 10795
rect 10744 10764 10793 10792
rect 10744 10752 10750 10764
rect 10781 10761 10793 10764
rect 10827 10761 10839 10795
rect 11146 10792 11152 10804
rect 10781 10755 10839 10761
rect 11072 10764 11152 10792
rect 11072 10733 11100 10764
rect 11146 10752 11152 10764
rect 11204 10752 11210 10804
rect 15378 10792 15384 10804
rect 11256 10764 15384 10792
rect 11057 10727 11115 10733
rect 11057 10693 11069 10727
rect 11103 10693 11115 10727
rect 11057 10687 11115 10693
rect 8665 10659 8723 10665
rect 7524 10628 7560 10656
rect 7466 10616 7472 10619
rect 7524 10616 7530 10628
rect 8665 10625 8677 10659
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 8932 10659 8990 10665
rect 8932 10625 8944 10659
rect 8978 10656 8990 10659
rect 10137 10659 10195 10665
rect 8978 10628 9996 10656
rect 8978 10625 8990 10628
rect 8932 10619 8990 10625
rect 7098 10588 7104 10600
rect 6748 10560 7104 10588
rect 6549 10551 6607 10557
rect 3786 10520 3792 10532
rect 3699 10492 3792 10520
rect 3786 10480 3792 10492
rect 3844 10520 3850 10532
rect 4798 10520 4804 10532
rect 3844 10492 4804 10520
rect 3844 10480 3850 10492
rect 4798 10480 4804 10492
rect 4856 10480 4862 10532
rect 4982 10480 4988 10532
rect 5040 10520 5046 10532
rect 5276 10520 5304 10551
rect 5040 10492 5304 10520
rect 5040 10480 5046 10492
rect 1397 10455 1455 10461
rect 1397 10421 1409 10455
rect 1443 10452 1455 10455
rect 1578 10452 1584 10464
rect 1443 10424 1584 10452
rect 1443 10421 1455 10424
rect 1397 10415 1455 10421
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 2498 10412 2504 10464
rect 2556 10452 2562 10464
rect 2869 10455 2927 10461
rect 2869 10452 2881 10455
rect 2556 10424 2881 10452
rect 2556 10412 2562 10424
rect 2869 10421 2881 10424
rect 2915 10421 2927 10455
rect 3878 10452 3884 10464
rect 3839 10424 3884 10452
rect 2869 10415 2927 10421
rect 3878 10412 3884 10424
rect 3936 10412 3942 10464
rect 5537 10455 5595 10461
rect 5537 10421 5549 10455
rect 5583 10452 5595 10455
rect 5718 10452 5724 10464
rect 5583 10424 5724 10452
rect 5583 10421 5595 10424
rect 5537 10415 5595 10421
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 6564 10452 6592 10551
rect 7098 10548 7104 10560
rect 7156 10548 7162 10600
rect 9968 10588 9996 10628
rect 10137 10625 10149 10659
rect 10183 10625 10195 10659
rect 10137 10619 10195 10625
rect 10870 10616 10876 10668
rect 10928 10656 10934 10668
rect 11149 10659 11207 10665
rect 11149 10656 11161 10659
rect 10928 10628 11161 10656
rect 10928 10616 10934 10628
rect 11149 10625 11161 10628
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 11054 10588 11060 10600
rect 9968 10560 11060 10588
rect 11054 10548 11060 10560
rect 11112 10548 11118 10600
rect 11256 10520 11284 10764
rect 15378 10752 15384 10764
rect 15436 10752 15442 10804
rect 15838 10752 15844 10804
rect 15896 10792 15902 10804
rect 16669 10795 16727 10801
rect 16669 10792 16681 10795
rect 15896 10764 16681 10792
rect 15896 10752 15902 10764
rect 16669 10761 16681 10764
rect 16715 10761 16727 10795
rect 16669 10755 16727 10761
rect 17862 10752 17868 10804
rect 17920 10792 17926 10804
rect 17957 10795 18015 10801
rect 17957 10792 17969 10795
rect 17920 10764 17969 10792
rect 17920 10752 17926 10764
rect 17957 10761 17969 10764
rect 18003 10761 18015 10795
rect 18322 10792 18328 10804
rect 18283 10764 18328 10792
rect 17957 10755 18015 10761
rect 18322 10752 18328 10764
rect 18380 10752 18386 10804
rect 12710 10684 12716 10736
rect 12768 10724 12774 10736
rect 12768 10696 14872 10724
rect 12768 10684 12774 10696
rect 11514 10656 11520 10668
rect 11475 10628 11520 10656
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 11773 10659 11831 10665
rect 11773 10656 11785 10659
rect 11624 10628 11785 10656
rect 11624 10588 11652 10628
rect 11773 10625 11785 10628
rect 11819 10625 11831 10659
rect 12986 10656 12992 10668
rect 12947 10628 12992 10656
rect 11773 10619 11831 10625
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13245 10659 13303 10665
rect 13245 10656 13257 10659
rect 13096 10628 13257 10656
rect 9646 10492 11284 10520
rect 11532 10560 11652 10588
rect 7466 10452 7472 10464
rect 6564 10424 7472 10452
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 9646 10452 9674 10492
rect 10042 10452 10048 10464
rect 8352 10424 9674 10452
rect 10003 10424 10048 10452
rect 8352 10412 8358 10424
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 11532 10452 11560 10560
rect 12526 10548 12532 10600
rect 12584 10588 12590 10600
rect 12894 10588 12900 10600
rect 12584 10560 12900 10588
rect 12584 10548 12590 10560
rect 12894 10548 12900 10560
rect 12952 10588 12958 10600
rect 13096 10588 13124 10628
rect 13245 10625 13257 10628
rect 13291 10625 13303 10659
rect 14844 10656 14872 10696
rect 14918 10684 14924 10736
rect 14976 10724 14982 10736
rect 14976 10696 15884 10724
rect 14976 10684 14982 10696
rect 15286 10656 15292 10668
rect 14844 10628 15292 10656
rect 13245 10619 13303 10625
rect 15286 10616 15292 10628
rect 15344 10616 15350 10668
rect 15856 10665 15884 10696
rect 16298 10684 16304 10736
rect 16356 10724 16362 10736
rect 17129 10727 17187 10733
rect 17129 10724 17141 10727
rect 16356 10696 17141 10724
rect 16356 10684 16362 10696
rect 17129 10693 17141 10696
rect 17175 10693 17187 10727
rect 17129 10687 17187 10693
rect 15585 10659 15643 10665
rect 15585 10625 15597 10659
rect 15631 10656 15643 10659
rect 15841 10659 15899 10665
rect 15631 10628 15792 10656
rect 15631 10625 15643 10628
rect 15585 10619 15643 10625
rect 12952 10560 13124 10588
rect 15764 10588 15792 10628
rect 15841 10625 15853 10659
rect 15887 10625 15899 10659
rect 15841 10619 15899 10625
rect 16850 10616 16856 10668
rect 16908 10656 16914 10668
rect 17037 10659 17095 10665
rect 17037 10656 17049 10659
rect 16908 10628 17049 10656
rect 16908 10616 16914 10628
rect 17037 10625 17049 10628
rect 17083 10625 17095 10659
rect 17310 10656 17316 10668
rect 17037 10619 17095 10625
rect 17236 10628 17316 10656
rect 16666 10588 16672 10600
rect 15764 10560 16672 10588
rect 12952 10548 12958 10560
rect 16666 10548 16672 10560
rect 16724 10588 16730 10600
rect 16942 10588 16948 10600
rect 16724 10560 16948 10588
rect 16724 10548 16730 10560
rect 16942 10548 16948 10560
rect 17000 10548 17006 10600
rect 17236 10597 17264 10628
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 17586 10616 17592 10668
rect 17644 10656 17650 10668
rect 17865 10659 17923 10665
rect 17865 10656 17877 10659
rect 17644 10628 17877 10656
rect 17644 10616 17650 10628
rect 17865 10625 17877 10628
rect 17911 10625 17923 10659
rect 17865 10619 17923 10625
rect 17221 10591 17279 10597
rect 17221 10557 17233 10591
rect 17267 10557 17279 10591
rect 18049 10591 18107 10597
rect 18049 10588 18061 10591
rect 17221 10551 17279 10557
rect 17328 10560 18061 10588
rect 16960 10520 16988 10548
rect 17328 10520 17356 10560
rect 18049 10557 18061 10560
rect 18095 10557 18107 10591
rect 18049 10551 18107 10557
rect 12452 10492 13032 10520
rect 16960 10492 17356 10520
rect 12452 10452 12480 10492
rect 11532 10424 12480 10452
rect 12526 10412 12532 10464
rect 12584 10452 12590 10464
rect 12897 10455 12955 10461
rect 12897 10452 12909 10455
rect 12584 10424 12909 10452
rect 12584 10412 12590 10424
rect 12897 10421 12909 10424
rect 12943 10421 12955 10455
rect 13004 10452 13032 10492
rect 13722 10452 13728 10464
rect 13004 10424 13728 10452
rect 12897 10415 12955 10421
rect 13722 10412 13728 10424
rect 13780 10412 13786 10464
rect 14090 10412 14096 10464
rect 14148 10452 14154 10464
rect 14369 10455 14427 10461
rect 14369 10452 14381 10455
rect 14148 10424 14381 10452
rect 14148 10412 14154 10424
rect 14369 10421 14381 10424
rect 14415 10421 14427 10455
rect 14369 10415 14427 10421
rect 14461 10455 14519 10461
rect 14461 10421 14473 10455
rect 14507 10452 14519 10455
rect 15194 10452 15200 10464
rect 14507 10424 15200 10452
rect 14507 10421 14519 10424
rect 14461 10415 14519 10421
rect 15194 10412 15200 10424
rect 15252 10412 15258 10464
rect 15470 10412 15476 10464
rect 15528 10452 15534 10464
rect 15654 10452 15660 10464
rect 15528 10424 15660 10452
rect 15528 10412 15534 10424
rect 15654 10412 15660 10424
rect 15712 10452 15718 10464
rect 15933 10455 15991 10461
rect 15933 10452 15945 10455
rect 15712 10424 15945 10452
rect 15712 10412 15718 10424
rect 15933 10421 15945 10424
rect 15979 10421 15991 10455
rect 15933 10415 15991 10421
rect 16298 10412 16304 10464
rect 16356 10452 16362 10464
rect 16393 10455 16451 10461
rect 16393 10452 16405 10455
rect 16356 10424 16405 10452
rect 16356 10412 16362 10424
rect 16393 10421 16405 10424
rect 16439 10421 16451 10455
rect 17494 10452 17500 10464
rect 17455 10424 17500 10452
rect 16393 10415 16451 10421
rect 17494 10412 17500 10424
rect 17552 10412 17558 10464
rect 1104 10362 18860 10384
rect 1104 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 3430 10362
rect 3482 10310 7622 10362
rect 7674 10310 7686 10362
rect 7738 10310 7750 10362
rect 7802 10310 7814 10362
rect 7866 10310 7878 10362
rect 7930 10310 12070 10362
rect 12122 10310 12134 10362
rect 12186 10310 12198 10362
rect 12250 10310 12262 10362
rect 12314 10310 12326 10362
rect 12378 10310 16518 10362
rect 16570 10310 16582 10362
rect 16634 10310 16646 10362
rect 16698 10310 16710 10362
rect 16762 10310 16774 10362
rect 16826 10310 18860 10362
rect 1104 10288 18860 10310
rect 1581 10251 1639 10257
rect 1581 10217 1593 10251
rect 1627 10248 1639 10251
rect 3050 10248 3056 10260
rect 1627 10220 3056 10248
rect 1627 10217 1639 10220
rect 1581 10211 1639 10217
rect 106 10140 112 10192
rect 164 10180 170 10192
rect 1765 10183 1823 10189
rect 1765 10180 1777 10183
rect 164 10152 1777 10180
rect 164 10140 170 10152
rect 1765 10149 1777 10152
rect 1811 10149 1823 10183
rect 1765 10143 1823 10149
rect 1964 10053 1992 10220
rect 3050 10208 3056 10220
rect 3108 10248 3114 10260
rect 4065 10251 4123 10257
rect 4065 10248 4077 10251
rect 3108 10220 4077 10248
rect 3108 10208 3114 10220
rect 4065 10217 4077 10220
rect 4111 10248 4123 10251
rect 6638 10248 6644 10260
rect 4111 10220 6644 10248
rect 4111 10217 4123 10220
rect 4065 10211 4123 10217
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 6733 10251 6791 10257
rect 6733 10217 6745 10251
rect 6779 10248 6791 10251
rect 6822 10248 6828 10260
rect 6779 10220 6828 10248
rect 6779 10217 6791 10220
rect 6733 10211 6791 10217
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 7098 10208 7104 10260
rect 7156 10248 7162 10260
rect 7653 10251 7711 10257
rect 7653 10248 7665 10251
rect 7156 10220 7665 10248
rect 7156 10208 7162 10220
rect 7653 10217 7665 10220
rect 7699 10217 7711 10251
rect 9398 10248 9404 10260
rect 7653 10211 7711 10217
rect 7760 10220 9404 10248
rect 7760 10192 7788 10220
rect 9398 10208 9404 10220
rect 9456 10208 9462 10260
rect 10962 10208 10968 10260
rect 11020 10248 11026 10260
rect 12710 10248 12716 10260
rect 11020 10220 12716 10248
rect 11020 10208 11026 10220
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 12802 10208 12808 10260
rect 12860 10248 12866 10260
rect 13081 10251 13139 10257
rect 13081 10248 13093 10251
rect 12860 10220 13093 10248
rect 12860 10208 12866 10220
rect 13081 10217 13093 10220
rect 13127 10217 13139 10251
rect 13081 10211 13139 10217
rect 4338 10180 4344 10192
rect 3344 10152 4344 10180
rect 2590 10112 2596 10124
rect 2551 10084 2596 10112
rect 2590 10072 2596 10084
rect 2648 10072 2654 10124
rect 3344 10121 3372 10152
rect 4338 10140 4344 10152
rect 4396 10140 4402 10192
rect 7558 10180 7564 10192
rect 6748 10152 7564 10180
rect 6748 10124 6776 10152
rect 7558 10140 7564 10152
rect 7616 10140 7622 10192
rect 7742 10140 7748 10192
rect 7800 10140 7806 10192
rect 9306 10180 9312 10192
rect 9219 10152 9312 10180
rect 9306 10140 9312 10152
rect 9364 10180 9370 10192
rect 11790 10180 11796 10192
rect 9364 10152 11796 10180
rect 9364 10140 9370 10152
rect 11790 10140 11796 10152
rect 11848 10140 11854 10192
rect 12986 10180 12992 10192
rect 12176 10152 12992 10180
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10081 3387 10115
rect 3510 10112 3516 10124
rect 3471 10084 3516 10112
rect 3329 10075 3387 10081
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 3789 10115 3847 10121
rect 3789 10081 3801 10115
rect 3835 10112 3847 10115
rect 4154 10112 4160 10124
rect 3835 10084 4160 10112
rect 3835 10081 3847 10084
rect 3789 10075 3847 10081
rect 4154 10072 4160 10084
rect 4212 10112 4218 10124
rect 4614 10112 4620 10124
rect 4212 10084 4620 10112
rect 4212 10072 4218 10084
rect 4614 10072 4620 10084
rect 4672 10072 4678 10124
rect 4982 10112 4988 10124
rect 4943 10084 4988 10112
rect 4982 10072 4988 10084
rect 5040 10072 5046 10124
rect 6730 10072 6736 10124
rect 6788 10072 6794 10124
rect 7377 10115 7435 10121
rect 7377 10081 7389 10115
rect 7423 10112 7435 10115
rect 8018 10112 8024 10124
rect 7423 10084 8024 10112
rect 7423 10081 7435 10084
rect 7377 10075 7435 10081
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 8110 10072 8116 10124
rect 8168 10112 8174 10124
rect 8205 10115 8263 10121
rect 8205 10112 8217 10115
rect 8168 10084 8217 10112
rect 8168 10072 8174 10084
rect 8205 10081 8217 10084
rect 8251 10081 8263 10115
rect 8205 10075 8263 10081
rect 10042 10072 10048 10124
rect 10100 10112 10106 10124
rect 10229 10115 10287 10121
rect 10229 10112 10241 10115
rect 10100 10084 10241 10112
rect 10100 10072 10106 10084
rect 10229 10081 10241 10084
rect 10275 10112 10287 10115
rect 10778 10112 10784 10124
rect 10275 10084 10784 10112
rect 10275 10081 10287 10084
rect 10229 10075 10287 10081
rect 10778 10072 10784 10084
rect 10836 10072 10842 10124
rect 11514 10072 11520 10124
rect 11572 10112 11578 10124
rect 11974 10112 11980 10124
rect 11572 10084 11980 10112
rect 11572 10072 11578 10084
rect 11974 10072 11980 10084
rect 12032 10112 12038 10124
rect 12176 10121 12204 10152
rect 12986 10140 12992 10152
rect 13044 10140 13050 10192
rect 14090 10180 14096 10192
rect 13556 10152 14096 10180
rect 12161 10115 12219 10121
rect 12161 10112 12173 10115
rect 12032 10084 12173 10112
rect 12032 10072 12038 10084
rect 12161 10081 12173 10084
rect 12207 10081 12219 10115
rect 12161 10075 12219 10081
rect 12437 10115 12495 10121
rect 12437 10081 12449 10115
rect 12483 10112 12495 10115
rect 13556 10112 13584 10152
rect 14090 10140 14096 10152
rect 14148 10140 14154 10192
rect 15473 10183 15531 10189
rect 15473 10149 15485 10183
rect 15519 10180 15531 10183
rect 15838 10180 15844 10192
rect 15519 10152 15844 10180
rect 15519 10149 15531 10152
rect 15473 10143 15531 10149
rect 15838 10140 15844 10152
rect 15896 10140 15902 10192
rect 16850 10140 16856 10192
rect 16908 10180 16914 10192
rect 18049 10183 18107 10189
rect 18049 10180 18061 10183
rect 16908 10152 18061 10180
rect 16908 10140 16914 10152
rect 18049 10149 18061 10152
rect 18095 10149 18107 10183
rect 18049 10143 18107 10149
rect 13722 10112 13728 10124
rect 12483 10084 13584 10112
rect 13683 10084 13728 10112
rect 12483 10081 12495 10084
rect 12437 10075 12495 10081
rect 13722 10072 13728 10084
rect 13780 10072 13786 10124
rect 15194 10072 15200 10124
rect 15252 10112 15258 10124
rect 16117 10115 16175 10121
rect 16117 10112 16129 10115
rect 15252 10084 16129 10112
rect 15252 10072 15258 10084
rect 16117 10081 16129 10084
rect 16163 10081 16175 10115
rect 16942 10112 16948 10124
rect 16903 10084 16948 10112
rect 16117 10075 16175 10081
rect 16942 10072 16948 10084
rect 17000 10072 17006 10124
rect 17865 10115 17923 10121
rect 17865 10081 17877 10115
rect 17911 10112 17923 10115
rect 18138 10112 18144 10124
rect 17911 10084 18144 10112
rect 17911 10081 17923 10084
rect 17865 10075 17923 10081
rect 18138 10072 18144 10084
rect 18196 10072 18202 10124
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10013 2007 10047
rect 1949 10007 2007 10013
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 3878 10044 3884 10056
rect 2455 10016 3884 10044
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 3878 10004 3884 10016
rect 3936 10004 3942 10056
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 4249 10047 4307 10053
rect 4249 10044 4261 10047
rect 4120 10016 4261 10044
rect 4120 10004 4126 10016
rect 4249 10013 4261 10016
rect 4295 10044 4307 10047
rect 4890 10044 4896 10056
rect 4295 10016 4896 10044
rect 4295 10013 4307 10016
rect 4249 10007 4307 10013
rect 4890 10004 4896 10016
rect 4948 10004 4954 10056
rect 5258 10044 5264 10056
rect 5219 10016 5264 10044
rect 5258 10004 5264 10016
rect 5316 10044 5322 10056
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 5316 10016 7113 10044
rect 5316 10004 5322 10016
rect 7101 10013 7113 10016
rect 7147 10044 7159 10047
rect 10413 10047 10471 10053
rect 10413 10044 10425 10047
rect 7147 10016 10425 10044
rect 7147 10013 7159 10016
rect 7101 10007 7159 10013
rect 10413 10013 10425 10016
rect 10459 10044 10471 10047
rect 10870 10044 10876 10056
rect 10459 10016 10876 10044
rect 10459 10013 10471 10016
rect 10413 10007 10471 10013
rect 10870 10004 10876 10016
rect 10928 10004 10934 10056
rect 12618 10044 12624 10056
rect 12579 10016 12624 10044
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 14093 10047 14151 10053
rect 14093 10013 14105 10047
rect 14139 10044 14151 10047
rect 14918 10044 14924 10056
rect 14139 10016 14924 10044
rect 14139 10013 14151 10016
rect 14093 10007 14151 10013
rect 14918 10004 14924 10016
rect 14976 10004 14982 10056
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10044 15991 10047
rect 17494 10044 17500 10056
rect 15979 10016 17500 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 17494 10004 17500 10016
rect 17552 10004 17558 10056
rect 17589 10047 17647 10053
rect 17589 10013 17601 10047
rect 17635 10044 17647 10047
rect 17954 10044 17960 10056
rect 17635 10016 17960 10044
rect 17635 10013 17647 10016
rect 17589 10007 17647 10013
rect 17954 10004 17960 10016
rect 18012 10044 18018 10056
rect 18233 10047 18291 10053
rect 18233 10044 18245 10047
rect 18012 10016 18245 10044
rect 18012 10004 18018 10016
rect 18233 10013 18245 10016
rect 18279 10013 18291 10047
rect 18233 10007 18291 10013
rect 2682 9936 2688 9988
rect 2740 9976 2746 9988
rect 3237 9979 3295 9985
rect 2740 9948 3004 9976
rect 2740 9936 2746 9948
rect 2041 9911 2099 9917
rect 2041 9877 2053 9911
rect 2087 9908 2099 9911
rect 2130 9908 2136 9920
rect 2087 9880 2136 9908
rect 2087 9877 2099 9880
rect 2041 9871 2099 9877
rect 2130 9868 2136 9880
rect 2188 9868 2194 9920
rect 2501 9911 2559 9917
rect 2501 9877 2513 9911
rect 2547 9908 2559 9911
rect 2869 9911 2927 9917
rect 2869 9908 2881 9911
rect 2547 9880 2881 9908
rect 2547 9877 2559 9880
rect 2501 9871 2559 9877
rect 2869 9877 2881 9880
rect 2915 9877 2927 9911
rect 2976 9908 3004 9948
rect 3237 9945 3249 9979
rect 3283 9976 3295 9979
rect 4801 9979 4859 9985
rect 3283 9948 4476 9976
rect 3283 9945 3295 9948
rect 3237 9939 3295 9945
rect 3326 9908 3332 9920
rect 2976 9880 3332 9908
rect 2869 9871 2927 9877
rect 3326 9868 3332 9880
rect 3384 9868 3390 9920
rect 4448 9917 4476 9948
rect 4801 9945 4813 9979
rect 4847 9976 4859 9979
rect 5994 9976 6000 9988
rect 4847 9948 6000 9976
rect 4847 9945 4859 9948
rect 4801 9939 4859 9945
rect 5994 9936 6000 9948
rect 6052 9936 6058 9988
rect 8021 9979 8079 9985
rect 8021 9945 8033 9979
rect 8067 9976 8079 9979
rect 8202 9976 8208 9988
rect 8067 9948 8208 9976
rect 8067 9945 8079 9948
rect 8021 9939 8079 9945
rect 8202 9936 8208 9948
rect 8260 9936 8266 9988
rect 9398 9936 9404 9988
rect 9456 9976 9462 9988
rect 9953 9979 10011 9985
rect 9456 9948 9720 9976
rect 9456 9936 9462 9948
rect 4433 9911 4491 9917
rect 4433 9877 4445 9911
rect 4479 9877 4491 9911
rect 4433 9871 4491 9877
rect 4890 9868 4896 9920
rect 4948 9908 4954 9920
rect 7742 9908 7748 9920
rect 4948 9880 7748 9908
rect 4948 9868 4954 9880
rect 7742 9868 7748 9880
rect 7800 9868 7806 9920
rect 8113 9911 8171 9917
rect 8113 9877 8125 9911
rect 8159 9908 8171 9911
rect 8573 9911 8631 9917
rect 8573 9908 8585 9911
rect 8159 9880 8585 9908
rect 8159 9877 8171 9880
rect 8113 9871 8171 9877
rect 8573 9877 8585 9880
rect 8619 9908 8631 9911
rect 8662 9908 8668 9920
rect 8619 9880 8668 9908
rect 8619 9877 8631 9880
rect 8573 9871 8631 9877
rect 8662 9868 8668 9880
rect 8720 9868 8726 9920
rect 8757 9911 8815 9917
rect 8757 9877 8769 9911
rect 8803 9908 8815 9911
rect 8846 9908 8852 9920
rect 8803 9880 8852 9908
rect 8803 9877 8815 9880
rect 8757 9871 8815 9877
rect 8846 9868 8852 9880
rect 8904 9868 8910 9920
rect 9030 9908 9036 9920
rect 8991 9880 9036 9908
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 9582 9908 9588 9920
rect 9543 9880 9588 9908
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 9692 9908 9720 9948
rect 9953 9945 9965 9979
rect 9999 9976 10011 9979
rect 10226 9976 10232 9988
rect 9999 9948 10232 9976
rect 9999 9945 10011 9948
rect 9953 9939 10011 9945
rect 10226 9936 10232 9948
rect 10284 9936 10290 9988
rect 14182 9976 14188 9988
rect 12084 9948 14188 9976
rect 10045 9911 10103 9917
rect 10045 9908 10057 9911
rect 9692 9880 10057 9908
rect 10045 9877 10057 9880
rect 10091 9908 10103 9911
rect 12084 9908 12112 9948
rect 14182 9936 14188 9948
rect 14240 9936 14246 9988
rect 14360 9979 14418 9985
rect 14360 9945 14372 9979
rect 14406 9976 14418 9979
rect 14826 9976 14832 9988
rect 14406 9948 14832 9976
rect 14406 9945 14418 9948
rect 14360 9939 14418 9945
rect 14826 9936 14832 9948
rect 14884 9936 14890 9988
rect 16761 9979 16819 9985
rect 16761 9945 16773 9979
rect 16807 9976 16819 9979
rect 17681 9979 17739 9985
rect 16807 9948 17264 9976
rect 16807 9945 16819 9948
rect 16761 9939 16819 9945
rect 10091 9880 12112 9908
rect 10091 9877 10103 9880
rect 10045 9871 10103 9877
rect 12342 9868 12348 9920
rect 12400 9908 12406 9920
rect 12529 9911 12587 9917
rect 12529 9908 12541 9911
rect 12400 9880 12541 9908
rect 12400 9868 12406 9880
rect 12529 9877 12541 9880
rect 12575 9877 12587 9911
rect 12986 9908 12992 9920
rect 12947 9880 12992 9908
rect 12529 9871 12587 9877
rect 12986 9868 12992 9880
rect 13044 9868 13050 9920
rect 13078 9868 13084 9920
rect 13136 9908 13142 9920
rect 13354 9908 13360 9920
rect 13136 9880 13360 9908
rect 13136 9868 13142 9880
rect 13354 9868 13360 9880
rect 13412 9908 13418 9920
rect 13449 9911 13507 9917
rect 13449 9908 13461 9911
rect 13412 9880 13461 9908
rect 13412 9868 13418 9880
rect 13449 9877 13461 9880
rect 13495 9877 13507 9911
rect 13449 9871 13507 9877
rect 13538 9868 13544 9920
rect 13596 9908 13602 9920
rect 15470 9908 15476 9920
rect 13596 9880 15476 9908
rect 13596 9868 13602 9880
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 15565 9911 15623 9917
rect 15565 9877 15577 9911
rect 15611 9908 15623 9911
rect 15746 9908 15752 9920
rect 15611 9880 15752 9908
rect 15611 9877 15623 9880
rect 15565 9871 15623 9877
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 16025 9911 16083 9917
rect 16025 9877 16037 9911
rect 16071 9908 16083 9911
rect 16393 9911 16451 9917
rect 16393 9908 16405 9911
rect 16071 9880 16405 9908
rect 16071 9877 16083 9880
rect 16025 9871 16083 9877
rect 16393 9877 16405 9880
rect 16439 9877 16451 9911
rect 16393 9871 16451 9877
rect 16853 9911 16911 9917
rect 16853 9877 16865 9911
rect 16899 9908 16911 9911
rect 17126 9908 17132 9920
rect 16899 9880 17132 9908
rect 16899 9877 16911 9880
rect 16853 9871 16911 9877
rect 17126 9868 17132 9880
rect 17184 9868 17190 9920
rect 17236 9917 17264 9948
rect 17681 9945 17693 9979
rect 17727 9976 17739 9979
rect 18509 9979 18567 9985
rect 18509 9976 18521 9979
rect 17727 9948 18521 9976
rect 17727 9945 17739 9948
rect 17681 9939 17739 9945
rect 18509 9945 18521 9948
rect 18555 9976 18567 9979
rect 18598 9976 18604 9988
rect 18555 9948 18604 9976
rect 18555 9945 18567 9948
rect 18509 9939 18567 9945
rect 18598 9936 18604 9948
rect 18656 9936 18662 9988
rect 17221 9911 17279 9917
rect 17221 9877 17233 9911
rect 17267 9877 17279 9911
rect 17221 9871 17279 9877
rect 1104 9818 18860 9840
rect 1104 9766 5398 9818
rect 5450 9766 5462 9818
rect 5514 9766 5526 9818
rect 5578 9766 5590 9818
rect 5642 9766 5654 9818
rect 5706 9766 9846 9818
rect 9898 9766 9910 9818
rect 9962 9766 9974 9818
rect 10026 9766 10038 9818
rect 10090 9766 10102 9818
rect 10154 9766 14294 9818
rect 14346 9766 14358 9818
rect 14410 9766 14422 9818
rect 14474 9766 14486 9818
rect 14538 9766 14550 9818
rect 14602 9766 18860 9818
rect 1104 9744 18860 9766
rect 1670 9664 1676 9716
rect 1728 9704 1734 9716
rect 3329 9707 3387 9713
rect 1728 9676 1900 9704
rect 1728 9664 1734 9676
rect 1872 9577 1900 9676
rect 3329 9673 3341 9707
rect 3375 9673 3387 9707
rect 3329 9667 3387 9673
rect 5353 9707 5411 9713
rect 5353 9673 5365 9707
rect 5399 9704 5411 9707
rect 5994 9704 6000 9716
rect 5399 9676 6000 9704
rect 5399 9673 5411 9676
rect 5353 9667 5411 9673
rect 2774 9636 2780 9648
rect 1964 9608 2780 9636
rect 1964 9577 1992 9608
rect 2774 9596 2780 9608
rect 2832 9596 2838 9648
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 3344 9636 3372 9667
rect 5994 9664 6000 9676
rect 6052 9664 6058 9716
rect 7374 9704 7380 9716
rect 6288 9676 7380 9704
rect 3016 9608 3372 9636
rect 4985 9639 5043 9645
rect 3016 9596 3022 9608
rect 4985 9605 4997 9639
rect 5031 9636 5043 9639
rect 5074 9636 5080 9648
rect 5031 9608 5080 9636
rect 5031 9605 5043 9608
rect 4985 9599 5043 9605
rect 5074 9596 5080 9608
rect 5132 9636 5138 9648
rect 6288 9636 6316 9676
rect 7374 9664 7380 9676
rect 7432 9664 7438 9716
rect 7466 9664 7472 9716
rect 7524 9704 7530 9716
rect 7745 9707 7803 9713
rect 7745 9704 7757 9707
rect 7524 9676 7757 9704
rect 7524 9664 7530 9676
rect 7745 9673 7757 9676
rect 7791 9673 7803 9707
rect 7745 9667 7803 9673
rect 8389 9707 8447 9713
rect 8389 9673 8401 9707
rect 8435 9704 8447 9707
rect 9582 9704 9588 9716
rect 8435 9676 9588 9704
rect 8435 9673 8447 9676
rect 8389 9667 8447 9673
rect 9582 9664 9588 9676
rect 9640 9664 9646 9716
rect 10226 9664 10232 9716
rect 10284 9704 10290 9716
rect 11241 9707 11299 9713
rect 11241 9704 11253 9707
rect 10284 9676 11253 9704
rect 10284 9664 10290 9676
rect 11241 9673 11253 9676
rect 11287 9704 11299 9707
rect 14642 9704 14648 9716
rect 11287 9676 14648 9704
rect 11287 9673 11299 9676
rect 11241 9667 11299 9673
rect 14642 9664 14648 9676
rect 14700 9664 14706 9716
rect 14918 9664 14924 9716
rect 14976 9704 14982 9716
rect 14976 9676 15424 9704
rect 14976 9664 14982 9676
rect 6822 9636 6828 9648
rect 5132 9608 6316 9636
rect 6380 9608 6828 9636
rect 5132 9596 5138 9608
rect 2222 9577 2228 9580
rect 1857 9571 1915 9577
rect 1857 9537 1869 9571
rect 1903 9537 1915 9571
rect 1857 9531 1915 9537
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9537 2007 9571
rect 2216 9568 2228 9577
rect 2183 9540 2228 9568
rect 1949 9531 2007 9537
rect 2216 9531 2228 9540
rect 2222 9528 2228 9531
rect 2280 9528 2286 9580
rect 2792 9568 2820 9596
rect 3421 9571 3479 9577
rect 3421 9568 3433 9571
rect 2792 9540 3433 9568
rect 3421 9537 3433 9540
rect 3467 9537 3479 9571
rect 3677 9571 3735 9577
rect 3677 9568 3689 9571
rect 3421 9531 3479 9537
rect 3528 9540 3689 9568
rect 3528 9500 3556 9540
rect 3677 9537 3689 9540
rect 3723 9537 3735 9571
rect 3677 9531 3735 9537
rect 4890 9528 4896 9580
rect 4948 9568 4954 9580
rect 5166 9568 5172 9580
rect 4948 9540 5172 9568
rect 4948 9528 4954 9540
rect 5166 9528 5172 9540
rect 5224 9568 5230 9580
rect 5813 9571 5871 9577
rect 5813 9568 5825 9571
rect 5224 9540 5825 9568
rect 5224 9528 5230 9540
rect 5813 9537 5825 9540
rect 5859 9537 5871 9571
rect 5813 9531 5871 9537
rect 6178 9528 6184 9580
rect 6236 9568 6242 9580
rect 6380 9577 6408 9608
rect 6822 9596 6828 9608
rect 6880 9596 6886 9648
rect 7282 9596 7288 9648
rect 7340 9636 7346 9648
rect 8938 9636 8944 9648
rect 7340 9608 8944 9636
rect 7340 9596 7346 9608
rect 8938 9596 8944 9608
rect 8996 9596 9002 9648
rect 12526 9636 12532 9648
rect 9048 9608 10824 9636
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 6236 9540 6377 9568
rect 6236 9528 6242 9540
rect 6365 9537 6377 9540
rect 6411 9537 6423 9571
rect 6632 9571 6690 9577
rect 6632 9568 6644 9571
rect 6365 9531 6423 9537
rect 6472 9540 6644 9568
rect 3252 9472 3556 9500
rect 5629 9503 5687 9509
rect 1302 9324 1308 9376
rect 1360 9364 1366 9376
rect 1397 9367 1455 9373
rect 1397 9364 1409 9367
rect 1360 9336 1409 9364
rect 1360 9324 1366 9336
rect 1397 9333 1409 9336
rect 1443 9364 1455 9367
rect 1486 9364 1492 9376
rect 1443 9336 1492 9364
rect 1443 9333 1455 9336
rect 1397 9327 1455 9333
rect 1486 9324 1492 9336
rect 1544 9324 1550 9376
rect 1670 9364 1676 9376
rect 1631 9336 1676 9364
rect 1670 9324 1676 9336
rect 1728 9324 1734 9376
rect 1946 9324 1952 9376
rect 2004 9364 2010 9376
rect 3252 9364 3280 9472
rect 5629 9469 5641 9503
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 5721 9503 5779 9509
rect 5721 9469 5733 9503
rect 5767 9500 5779 9503
rect 5994 9500 6000 9512
rect 5767 9472 6000 9500
rect 5767 9469 5779 9472
rect 5721 9463 5779 9469
rect 5644 9432 5672 9463
rect 5994 9460 6000 9472
rect 6052 9460 6058 9512
rect 6472 9500 6500 9540
rect 6632 9537 6644 9540
rect 6678 9568 6690 9571
rect 6914 9568 6920 9580
rect 6678 9540 6920 9568
rect 6678 9537 6690 9540
rect 6632 9531 6690 9537
rect 6914 9528 6920 9540
rect 6972 9568 6978 9580
rect 8110 9568 8116 9580
rect 6972 9540 8116 9568
rect 6972 9528 6978 9540
rect 8110 9528 8116 9540
rect 8168 9528 8174 9580
rect 8478 9500 8484 9512
rect 6104 9472 6500 9500
rect 8439 9472 8484 9500
rect 6104 9432 6132 9472
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 9048 9509 9076 9608
rect 10796 9580 10824 9608
rect 11900 9608 12532 9636
rect 9217 9571 9275 9577
rect 9217 9537 9229 9571
rect 9263 9568 9275 9571
rect 9306 9568 9312 9580
rect 9263 9540 9312 9568
rect 9263 9537 9275 9540
rect 9217 9531 9275 9537
rect 9306 9528 9312 9540
rect 9364 9528 9370 9580
rect 10778 9528 10784 9580
rect 10836 9577 10842 9580
rect 10836 9568 10848 9577
rect 11057 9571 11115 9577
rect 10836 9540 10881 9568
rect 10836 9531 10848 9540
rect 11057 9537 11069 9571
rect 11103 9537 11115 9571
rect 11057 9531 11115 9537
rect 10836 9528 10842 9531
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9469 8723 9503
rect 8665 9463 8723 9469
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9469 9091 9503
rect 9033 9463 9091 9469
rect 5644 9404 6132 9432
rect 8680 9432 8708 9463
rect 9122 9460 9128 9512
rect 9180 9500 9186 9512
rect 9180 9472 9225 9500
rect 9180 9460 9186 9472
rect 11072 9432 11100 9531
rect 11900 9509 11928 9608
rect 12526 9596 12532 9608
rect 12584 9596 12590 9648
rect 12710 9596 12716 9648
rect 12768 9636 12774 9648
rect 12768 9608 13308 9636
rect 12768 9596 12774 9608
rect 12161 9571 12219 9577
rect 12161 9537 12173 9571
rect 12207 9568 12219 9571
rect 12207 9540 12756 9568
rect 12207 9537 12219 9540
rect 12161 9531 12219 9537
rect 11885 9503 11943 9509
rect 11885 9469 11897 9503
rect 11931 9469 11943 9503
rect 12066 9500 12072 9512
rect 12027 9472 12072 9500
rect 11885 9463 11943 9469
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 11974 9432 11980 9444
rect 8680 9404 9720 9432
rect 11072 9404 11980 9432
rect 2004 9336 3280 9364
rect 2004 9324 2010 9336
rect 4062 9324 4068 9376
rect 4120 9364 4126 9376
rect 4801 9367 4859 9373
rect 4801 9364 4813 9367
rect 4120 9336 4813 9364
rect 4120 9324 4126 9336
rect 4801 9333 4813 9336
rect 4847 9333 4859 9367
rect 5166 9364 5172 9376
rect 5127 9336 5172 9364
rect 4801 9327 4859 9333
rect 5166 9324 5172 9336
rect 5224 9324 5230 9376
rect 6181 9367 6239 9373
rect 6181 9333 6193 9367
rect 6227 9364 6239 9367
rect 7098 9364 7104 9376
rect 6227 9336 7104 9364
rect 6227 9333 6239 9336
rect 6181 9327 6239 9333
rect 7098 9324 7104 9336
rect 7156 9324 7162 9376
rect 7374 9324 7380 9376
rect 7432 9364 7438 9376
rect 7837 9367 7895 9373
rect 7837 9364 7849 9367
rect 7432 9336 7849 9364
rect 7432 9324 7438 9336
rect 7837 9333 7849 9336
rect 7883 9333 7895 9367
rect 7837 9327 7895 9333
rect 8021 9367 8079 9373
rect 8021 9333 8033 9367
rect 8067 9364 8079 9367
rect 8386 9364 8392 9376
rect 8067 9336 8392 9364
rect 8067 9333 8079 9336
rect 8021 9327 8079 9333
rect 8386 9324 8392 9336
rect 8444 9324 8450 9376
rect 8846 9324 8852 9376
rect 8904 9364 8910 9376
rect 9122 9364 9128 9376
rect 8904 9336 9128 9364
rect 8904 9324 8910 9336
rect 9122 9324 9128 9336
rect 9180 9324 9186 9376
rect 9582 9364 9588 9376
rect 9543 9336 9588 9364
rect 9582 9324 9588 9336
rect 9640 9324 9646 9376
rect 9692 9373 9720 9404
rect 11974 9392 11980 9404
rect 12032 9392 12038 9444
rect 12342 9392 12348 9444
rect 12400 9392 12406 9444
rect 12621 9435 12679 9441
rect 12621 9401 12633 9435
rect 12667 9432 12679 9435
rect 12728 9432 12756 9540
rect 12802 9528 12808 9580
rect 12860 9568 12866 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12860 9540 13001 9568
rect 12860 9528 12866 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13280 9568 13308 9608
rect 13722 9596 13728 9648
rect 13780 9636 13786 9648
rect 13780 9608 14228 9636
rect 13780 9596 13786 9608
rect 13740 9568 13768 9596
rect 13280 9540 13768 9568
rect 13817 9571 13875 9577
rect 13078 9500 13084 9512
rect 13039 9472 13084 9500
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 13280 9509 13308 9540
rect 13817 9537 13829 9571
rect 13863 9568 13875 9571
rect 14090 9568 14096 9580
rect 13863 9540 14096 9568
rect 13863 9537 13875 9540
rect 13817 9531 13875 9537
rect 14090 9528 14096 9540
rect 14148 9528 14154 9580
rect 13265 9503 13323 9509
rect 13265 9469 13277 9503
rect 13311 9469 13323 9503
rect 13265 9463 13323 9469
rect 13722 9460 13728 9512
rect 13780 9500 13786 9512
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13780 9472 13921 9500
rect 13780 9460 13786 9472
rect 13909 9469 13921 9472
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 14001 9503 14059 9509
rect 14001 9469 14013 9503
rect 14047 9500 14059 9503
rect 14200 9500 14228 9608
rect 15396 9568 15424 9676
rect 18138 9664 18144 9716
rect 18196 9704 18202 9716
rect 18233 9707 18291 9713
rect 18233 9704 18245 9707
rect 18196 9676 18245 9704
rect 18196 9664 18202 9676
rect 18233 9673 18245 9676
rect 18279 9673 18291 9707
rect 18233 9667 18291 9673
rect 15504 9639 15562 9645
rect 15504 9605 15516 9639
rect 15550 9636 15562 9639
rect 16485 9639 16543 9645
rect 16485 9636 16497 9639
rect 15550 9608 16497 9636
rect 15550 9605 15562 9608
rect 15504 9599 15562 9605
rect 16485 9605 16497 9608
rect 16531 9605 16543 9639
rect 16485 9599 16543 9605
rect 17954 9596 17960 9648
rect 18012 9636 18018 9648
rect 18325 9639 18383 9645
rect 18325 9636 18337 9639
rect 18012 9608 18337 9636
rect 18012 9596 18018 9608
rect 18325 9605 18337 9608
rect 18371 9605 18383 9639
rect 18325 9599 18383 9605
rect 15749 9571 15807 9577
rect 15749 9568 15761 9571
rect 15396 9540 15761 9568
rect 15749 9537 15761 9540
rect 15795 9537 15807 9571
rect 15749 9531 15807 9537
rect 14047 9472 14228 9500
rect 15764 9500 15792 9531
rect 15838 9528 15844 9580
rect 15896 9568 15902 9580
rect 17120 9571 17178 9577
rect 15896 9540 15941 9568
rect 15896 9528 15902 9540
rect 17120 9537 17132 9571
rect 17166 9568 17178 9571
rect 17494 9568 17500 9580
rect 17166 9540 17500 9568
rect 17166 9537 17178 9540
rect 17120 9531 17178 9537
rect 17494 9528 17500 9540
rect 17552 9528 17558 9580
rect 16850 9500 16856 9512
rect 15764 9472 16856 9500
rect 14047 9469 14059 9472
rect 14001 9463 14059 9469
rect 16850 9460 16856 9472
rect 16908 9460 16914 9512
rect 13446 9432 13452 9444
rect 12667 9404 12756 9432
rect 13407 9404 13452 9432
rect 12667 9401 12679 9404
rect 12621 9395 12679 9401
rect 13446 9392 13452 9404
rect 13504 9392 13510 9444
rect 16758 9432 16764 9444
rect 16684 9404 16764 9432
rect 9677 9367 9735 9373
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 10134 9364 10140 9376
rect 9723 9336 10140 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 10928 9336 11621 9364
rect 10928 9324 10934 9336
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 12360 9364 12388 9392
rect 12529 9367 12587 9373
rect 12529 9364 12541 9367
rect 12360 9336 12541 9364
rect 11609 9327 11667 9333
rect 12529 9333 12541 9336
rect 12575 9333 12587 9367
rect 12529 9327 12587 9333
rect 14369 9367 14427 9373
rect 14369 9333 14381 9367
rect 14415 9364 14427 9367
rect 15378 9364 15384 9376
rect 14415 9336 15384 9364
rect 14415 9333 14427 9336
rect 14369 9327 14427 9333
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 16206 9324 16212 9376
rect 16264 9364 16270 9376
rect 16684 9373 16712 9404
rect 16758 9392 16764 9404
rect 16816 9392 16822 9444
rect 16669 9367 16727 9373
rect 16669 9364 16681 9367
rect 16264 9336 16681 9364
rect 16264 9324 16270 9336
rect 16669 9333 16681 9336
rect 16715 9333 16727 9367
rect 16669 9327 16727 9333
rect 1104 9274 18860 9296
rect 1104 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 3430 9274
rect 3482 9222 7622 9274
rect 7674 9222 7686 9274
rect 7738 9222 7750 9274
rect 7802 9222 7814 9274
rect 7866 9222 7878 9274
rect 7930 9222 12070 9274
rect 12122 9222 12134 9274
rect 12186 9222 12198 9274
rect 12250 9222 12262 9274
rect 12314 9222 12326 9274
rect 12378 9222 16518 9274
rect 16570 9222 16582 9274
rect 16634 9222 16646 9274
rect 16698 9222 16710 9274
rect 16762 9222 16774 9274
rect 16826 9222 18860 9274
rect 1104 9200 18860 9222
rect 4154 9160 4160 9172
rect 1964 9132 4160 9160
rect 1964 8965 1992 9132
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 4338 9160 4344 9172
rect 4299 9132 4344 9160
rect 4338 9120 4344 9132
rect 4396 9120 4402 9172
rect 6549 9163 6607 9169
rect 6549 9129 6561 9163
rect 6595 9160 6607 9163
rect 7282 9160 7288 9172
rect 6595 9132 7288 9160
rect 6595 9129 6607 9132
rect 6549 9123 6607 9129
rect 7282 9120 7288 9132
rect 7340 9160 7346 9172
rect 7340 9132 8156 9160
rect 7340 9120 7346 9132
rect 2774 9052 2780 9104
rect 2832 9092 2838 9104
rect 6641 9095 6699 9101
rect 2832 9064 5212 9092
rect 2832 9052 2838 9064
rect 2498 9024 2504 9036
rect 2459 8996 2504 9024
rect 2498 8984 2504 8996
rect 2556 8984 2562 9036
rect 2590 8984 2596 9036
rect 2648 9024 2654 9036
rect 2958 9024 2964 9036
rect 2648 8996 2693 9024
rect 2919 8996 2964 9024
rect 2648 8984 2654 8996
rect 2958 8984 2964 8996
rect 3016 8984 3022 9036
rect 3145 9027 3203 9033
rect 3145 8993 3157 9027
rect 3191 9024 3203 9027
rect 3510 9024 3516 9036
rect 3191 8996 3516 9024
rect 3191 8993 3203 8996
rect 3145 8987 3203 8993
rect 3510 8984 3516 8996
rect 3568 8984 3574 9036
rect 4982 9024 4988 9036
rect 4943 8996 4988 9024
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 5184 9033 5212 9064
rect 6641 9061 6653 9095
rect 6687 9092 6699 9095
rect 6914 9092 6920 9104
rect 6687 9064 6920 9092
rect 6687 9061 6699 9064
rect 6641 9055 6699 9061
rect 6914 9052 6920 9064
rect 6972 9052 6978 9104
rect 5169 9027 5227 9033
rect 5169 8993 5181 9027
rect 5215 8993 5227 9027
rect 5169 8987 5227 8993
rect 1949 8959 2007 8965
rect 1949 8925 1961 8959
rect 1995 8925 2007 8959
rect 2406 8956 2412 8968
rect 2367 8928 2412 8956
rect 1949 8919 2007 8925
rect 2406 8916 2412 8928
rect 2464 8916 2470 8968
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8956 3295 8959
rect 3694 8956 3700 8968
rect 3283 8928 3700 8956
rect 3283 8925 3295 8928
rect 3237 8919 3295 8925
rect 3694 8916 3700 8928
rect 3752 8916 3758 8968
rect 3970 8916 3976 8968
rect 4028 8956 4034 8968
rect 4065 8959 4123 8965
rect 4065 8956 4077 8959
rect 4028 8928 4077 8956
rect 4028 8916 4034 8928
rect 4065 8925 4077 8928
rect 4111 8925 4123 8959
rect 4065 8919 4123 8925
rect 5436 8959 5494 8965
rect 5436 8925 5448 8959
rect 5482 8956 5494 8959
rect 5718 8956 5724 8968
rect 5482 8928 5724 8956
rect 5482 8925 5494 8928
rect 5436 8919 5494 8925
rect 5718 8916 5724 8928
rect 5776 8916 5782 8968
rect 6178 8916 6184 8968
rect 6236 8956 6242 8968
rect 8128 8965 8156 9132
rect 8478 9120 8484 9172
rect 8536 9160 8542 9172
rect 10413 9163 10471 9169
rect 10413 9160 10425 9163
rect 8536 9132 10425 9160
rect 8536 9120 8542 9132
rect 10413 9129 10425 9132
rect 10459 9129 10471 9163
rect 10413 9123 10471 9129
rect 12253 9163 12311 9169
rect 12253 9129 12265 9163
rect 12299 9160 12311 9163
rect 13078 9160 13084 9172
rect 12299 9132 13084 9160
rect 12299 9129 12311 9132
rect 12253 9123 12311 9129
rect 13078 9120 13084 9132
rect 13136 9120 13142 9172
rect 14090 9160 14096 9172
rect 14051 9132 14096 9160
rect 14090 9120 14096 9132
rect 14148 9120 14154 9172
rect 15764 9132 17080 9160
rect 8938 9052 8944 9104
rect 8996 9092 9002 9104
rect 9033 9095 9091 9101
rect 9033 9092 9045 9095
rect 8996 9064 9045 9092
rect 8996 9052 9002 9064
rect 9033 9061 9045 9064
rect 9079 9061 9091 9095
rect 9033 9055 9091 9061
rect 8021 8959 8079 8965
rect 8021 8956 8033 8959
rect 6236 8928 8033 8956
rect 6236 8916 6242 8928
rect 8021 8925 8033 8928
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 8113 8959 8171 8965
rect 8113 8925 8125 8959
rect 8159 8925 8171 8959
rect 9048 8956 9076 9055
rect 9398 9052 9404 9104
rect 9456 9092 9462 9104
rect 10502 9092 10508 9104
rect 9456 9064 10508 9092
rect 9456 9052 9462 9064
rect 10502 9052 10508 9064
rect 10560 9052 10566 9104
rect 12345 9095 12403 9101
rect 12345 9061 12357 9095
rect 12391 9092 12403 9095
rect 12710 9092 12716 9104
rect 12391 9064 12716 9092
rect 12391 9061 12403 9064
rect 12345 9055 12403 9061
rect 12710 9052 12716 9064
rect 12768 9052 12774 9104
rect 15654 9092 15660 9104
rect 14568 9064 15660 9092
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 10045 9027 10103 9033
rect 10045 9024 10057 9027
rect 9640 8996 10057 9024
rect 9640 8984 9646 8996
rect 10045 8993 10057 8996
rect 10091 8993 10103 9027
rect 10226 9024 10232 9036
rect 10187 8996 10232 9024
rect 10045 8987 10103 8993
rect 10226 8984 10232 8996
rect 10284 8984 10290 9036
rect 10778 8984 10784 9036
rect 10836 9024 10842 9036
rect 10965 9027 11023 9033
rect 10965 9024 10977 9027
rect 10836 8996 10977 9024
rect 10836 8984 10842 8996
rect 10965 8993 10977 8996
rect 11011 8993 11023 9027
rect 10965 8987 11023 8993
rect 11701 9027 11759 9033
rect 11701 8993 11713 9027
rect 11747 9024 11759 9027
rect 11747 8996 11928 9024
rect 11747 8993 11759 8996
rect 11701 8987 11759 8993
rect 9950 8956 9956 8968
rect 9048 8928 9956 8956
rect 8113 8919 8171 8925
rect 9950 8916 9956 8928
rect 10008 8916 10014 8968
rect 1673 8891 1731 8897
rect 1673 8857 1685 8891
rect 1719 8888 1731 8891
rect 2590 8888 2596 8900
rect 1719 8860 2596 8888
rect 1719 8857 1731 8860
rect 1673 8851 1731 8857
rect 2590 8848 2596 8860
rect 2648 8848 2654 8900
rect 4709 8891 4767 8897
rect 4709 8857 4721 8891
rect 4755 8888 4767 8891
rect 5074 8888 5080 8900
rect 4755 8860 5080 8888
rect 4755 8857 4767 8860
rect 4709 8851 4767 8857
rect 5074 8848 5080 8860
rect 5132 8848 5138 8900
rect 6914 8848 6920 8900
rect 6972 8888 6978 8900
rect 7374 8888 7380 8900
rect 6972 8860 7380 8888
rect 6972 8848 6978 8860
rect 7374 8848 7380 8860
rect 7432 8848 7438 8900
rect 7776 8891 7834 8897
rect 7776 8857 7788 8891
rect 7822 8888 7834 8891
rect 8757 8891 8815 8897
rect 8757 8888 8769 8891
rect 7822 8860 8769 8888
rect 7822 8857 7834 8860
rect 7776 8851 7834 8857
rect 8757 8857 8769 8860
rect 8803 8857 8815 8891
rect 10873 8891 10931 8897
rect 10873 8888 10885 8891
rect 8757 8851 8815 8857
rect 9232 8860 10885 8888
rect 2038 8820 2044 8832
rect 1999 8792 2044 8820
rect 2038 8780 2044 8792
rect 2096 8780 2102 8832
rect 3418 8780 3424 8832
rect 3476 8820 3482 8832
rect 3605 8823 3663 8829
rect 3605 8820 3617 8823
rect 3476 8792 3617 8820
rect 3476 8780 3482 8792
rect 3605 8789 3617 8792
rect 3651 8789 3663 8823
rect 3605 8783 3663 8789
rect 3786 8780 3792 8832
rect 3844 8820 3850 8832
rect 3881 8823 3939 8829
rect 3881 8820 3893 8823
rect 3844 8792 3893 8820
rect 3844 8780 3850 8792
rect 3881 8789 3893 8792
rect 3927 8789 3939 8823
rect 3881 8783 3939 8789
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 4157 8823 4215 8829
rect 4157 8820 4169 8823
rect 4028 8792 4169 8820
rect 4028 8780 4034 8792
rect 4157 8789 4169 8792
rect 4203 8789 4215 8823
rect 4157 8783 4215 8789
rect 4801 8823 4859 8829
rect 4801 8789 4813 8823
rect 4847 8820 4859 8823
rect 6822 8820 6828 8832
rect 4847 8792 6828 8820
rect 4847 8789 4859 8792
rect 4801 8783 4859 8789
rect 6822 8780 6828 8792
rect 6880 8820 6886 8832
rect 9232 8829 9260 8860
rect 10873 8857 10885 8860
rect 10919 8888 10931 8891
rect 11330 8888 11336 8900
rect 10919 8860 11336 8888
rect 10919 8857 10931 8860
rect 10873 8851 10931 8857
rect 11330 8848 11336 8860
rect 11388 8848 11394 8900
rect 11698 8848 11704 8900
rect 11756 8888 11762 8900
rect 11793 8891 11851 8897
rect 11793 8888 11805 8891
rect 11756 8860 11805 8888
rect 11756 8848 11762 8860
rect 11793 8857 11805 8860
rect 11839 8857 11851 8891
rect 11900 8888 11928 8996
rect 14182 8984 14188 9036
rect 14240 9024 14246 9036
rect 14568 9033 14596 9064
rect 15654 9052 15660 9064
rect 15712 9092 15718 9104
rect 15764 9101 15792 9132
rect 15749 9095 15807 9101
rect 15749 9092 15761 9095
rect 15712 9064 15761 9092
rect 15712 9052 15718 9064
rect 15749 9061 15761 9064
rect 15795 9061 15807 9095
rect 17052 9092 17080 9132
rect 17126 9120 17132 9172
rect 17184 9160 17190 9172
rect 17589 9163 17647 9169
rect 17589 9160 17601 9163
rect 17184 9132 17601 9160
rect 17184 9120 17190 9132
rect 17589 9129 17601 9132
rect 17635 9129 17647 9163
rect 17589 9123 17647 9129
rect 17052 9064 17172 9092
rect 15749 9055 15807 9061
rect 14553 9027 14611 9033
rect 14553 9024 14565 9027
rect 14240 8996 14565 9024
rect 14240 8984 14246 8996
rect 14553 8993 14565 8996
rect 14599 8993 14611 9027
rect 14553 8987 14611 8993
rect 14645 9027 14703 9033
rect 14645 8993 14657 9027
rect 14691 8993 14703 9027
rect 14645 8987 14703 8993
rect 15565 9027 15623 9033
rect 15565 8993 15577 9027
rect 15611 9024 15623 9027
rect 15838 9024 15844 9036
rect 15611 8996 15844 9024
rect 15611 8993 15623 8996
rect 15565 8987 15623 8993
rect 11974 8916 11980 8968
rect 12032 8956 12038 8968
rect 13725 8959 13783 8965
rect 13725 8956 13737 8959
rect 12032 8928 13737 8956
rect 12032 8916 12038 8928
rect 13725 8925 13737 8928
rect 13771 8925 13783 8959
rect 13725 8919 13783 8925
rect 12894 8888 12900 8900
rect 11900 8860 12900 8888
rect 11793 8851 11851 8857
rect 12894 8848 12900 8860
rect 12952 8888 12958 8900
rect 13480 8891 13538 8897
rect 13480 8888 13492 8891
rect 12952 8860 13492 8888
rect 12952 8848 12958 8860
rect 13480 8857 13492 8860
rect 13526 8888 13538 8891
rect 14660 8888 14688 8987
rect 15838 8984 15844 8996
rect 15896 8984 15902 9036
rect 16117 8959 16175 8965
rect 16117 8925 16129 8959
rect 16163 8956 16175 8959
rect 16666 8956 16672 8968
rect 16163 8928 16672 8956
rect 16163 8925 16175 8928
rect 16117 8919 16175 8925
rect 16666 8916 16672 8928
rect 16724 8956 16730 8968
rect 16850 8956 16856 8968
rect 16724 8928 16856 8956
rect 16724 8916 16730 8928
rect 16850 8916 16856 8928
rect 16908 8916 16914 8968
rect 17144 8956 17172 9064
rect 18138 9024 18144 9036
rect 18099 8996 18144 9024
rect 18138 8984 18144 8996
rect 18196 8984 18202 9036
rect 17957 8959 18015 8965
rect 17957 8956 17969 8959
rect 17144 8928 17969 8956
rect 17957 8925 17969 8928
rect 18003 8956 18015 8959
rect 18417 8959 18475 8965
rect 18417 8956 18429 8959
rect 18003 8928 18429 8956
rect 18003 8925 18015 8928
rect 17957 8919 18015 8925
rect 18417 8925 18429 8928
rect 18463 8925 18475 8959
rect 18417 8919 18475 8925
rect 13526 8860 14688 8888
rect 13526 8857 13538 8860
rect 13480 8851 13538 8857
rect 14734 8848 14740 8900
rect 14792 8888 14798 8900
rect 15289 8891 15347 8897
rect 15289 8888 15301 8891
rect 14792 8860 15301 8888
rect 14792 8848 14798 8860
rect 15289 8857 15301 8860
rect 15335 8888 15347 8891
rect 16206 8888 16212 8900
rect 15335 8860 16212 8888
rect 15335 8857 15347 8860
rect 15289 8851 15347 8857
rect 16206 8848 16212 8860
rect 16264 8848 16270 8900
rect 16390 8897 16396 8900
rect 16384 8851 16396 8897
rect 16448 8888 16454 8900
rect 16448 8860 16484 8888
rect 16390 8848 16396 8851
rect 16448 8848 16454 8860
rect 9217 8823 9275 8829
rect 9217 8820 9229 8823
rect 6880 8792 9229 8820
rect 6880 8780 6886 8792
rect 9217 8789 9229 8792
rect 9263 8789 9275 8823
rect 9398 8820 9404 8832
rect 9359 8792 9404 8820
rect 9217 8783 9275 8789
rect 9398 8780 9404 8792
rect 9456 8780 9462 8832
rect 9582 8820 9588 8832
rect 9543 8792 9588 8820
rect 9582 8780 9588 8792
rect 9640 8780 9646 8832
rect 10502 8780 10508 8832
rect 10560 8820 10566 8832
rect 10781 8823 10839 8829
rect 10781 8820 10793 8823
rect 10560 8792 10793 8820
rect 10560 8780 10566 8792
rect 10781 8789 10793 8792
rect 10827 8789 10839 8823
rect 11238 8820 11244 8832
rect 11199 8792 11244 8820
rect 10781 8783 10839 8789
rect 11238 8780 11244 8792
rect 11296 8780 11302 8832
rect 11514 8780 11520 8832
rect 11572 8820 11578 8832
rect 11885 8823 11943 8829
rect 11885 8820 11897 8823
rect 11572 8792 11897 8820
rect 11572 8780 11578 8792
rect 11885 8789 11897 8792
rect 11931 8820 11943 8823
rect 12342 8820 12348 8832
rect 11931 8792 12348 8820
rect 11931 8789 11943 8792
rect 11885 8783 11943 8789
rect 12342 8780 12348 8792
rect 12400 8780 12406 8832
rect 13814 8820 13820 8832
rect 13775 8792 13820 8820
rect 13814 8780 13820 8792
rect 13872 8780 13878 8832
rect 14461 8823 14519 8829
rect 14461 8789 14473 8823
rect 14507 8820 14519 8823
rect 14642 8820 14648 8832
rect 14507 8792 14648 8820
rect 14507 8789 14519 8792
rect 14461 8783 14519 8789
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 14921 8823 14979 8829
rect 14921 8789 14933 8823
rect 14967 8820 14979 8823
rect 15102 8820 15108 8832
rect 14967 8792 15108 8820
rect 14967 8789 14979 8792
rect 14921 8783 14979 8789
rect 15102 8780 15108 8792
rect 15160 8780 15166 8832
rect 15381 8823 15439 8829
rect 15381 8789 15393 8823
rect 15427 8820 15439 8823
rect 15470 8820 15476 8832
rect 15427 8792 15476 8820
rect 15427 8789 15439 8792
rect 15381 8783 15439 8789
rect 15470 8780 15476 8792
rect 15528 8820 15534 8832
rect 15933 8823 15991 8829
rect 15933 8820 15945 8823
rect 15528 8792 15945 8820
rect 15528 8780 15534 8792
rect 15933 8789 15945 8792
rect 15979 8820 15991 8823
rect 16298 8820 16304 8832
rect 15979 8792 16304 8820
rect 15979 8789 15991 8792
rect 15933 8783 15991 8789
rect 16298 8780 16304 8792
rect 16356 8780 16362 8832
rect 17497 8823 17555 8829
rect 17497 8789 17509 8823
rect 17543 8820 17555 8823
rect 17586 8820 17592 8832
rect 17543 8792 17592 8820
rect 17543 8789 17555 8792
rect 17497 8783 17555 8789
rect 17586 8780 17592 8792
rect 17644 8780 17650 8832
rect 18046 8780 18052 8832
rect 18104 8820 18110 8832
rect 18104 8792 18149 8820
rect 18104 8780 18110 8792
rect 1104 8730 18860 8752
rect 1104 8678 5398 8730
rect 5450 8678 5462 8730
rect 5514 8678 5526 8730
rect 5578 8678 5590 8730
rect 5642 8678 5654 8730
rect 5706 8678 9846 8730
rect 9898 8678 9910 8730
rect 9962 8678 9974 8730
rect 10026 8678 10038 8730
rect 10090 8678 10102 8730
rect 10154 8678 14294 8730
rect 14346 8678 14358 8730
rect 14410 8678 14422 8730
rect 14474 8678 14486 8730
rect 14538 8678 14550 8730
rect 14602 8678 18860 8730
rect 1104 8656 18860 8678
rect 2222 8576 2228 8628
rect 2280 8616 2286 8628
rect 2961 8619 3019 8625
rect 2961 8616 2973 8619
rect 2280 8588 2973 8616
rect 2280 8576 2286 8588
rect 2961 8585 2973 8588
rect 3007 8585 3019 8619
rect 3418 8616 3424 8628
rect 3379 8588 3424 8616
rect 2961 8579 3019 8585
rect 3418 8576 3424 8588
rect 3476 8576 3482 8628
rect 4798 8616 4804 8628
rect 4711 8588 4804 8616
rect 4798 8576 4804 8588
rect 4856 8616 4862 8628
rect 5902 8616 5908 8628
rect 4856 8588 5908 8616
rect 4856 8576 4862 8588
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 6641 8619 6699 8625
rect 6641 8585 6653 8619
rect 6687 8616 6699 8619
rect 6914 8616 6920 8628
rect 6687 8588 6920 8616
rect 6687 8585 6699 8588
rect 6641 8579 6699 8585
rect 6914 8576 6920 8588
rect 6972 8576 6978 8628
rect 7098 8616 7104 8628
rect 7059 8588 7104 8616
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 8113 8619 8171 8625
rect 8113 8585 8125 8619
rect 8159 8616 8171 8619
rect 8570 8616 8576 8628
rect 8159 8588 8576 8616
rect 8159 8585 8171 8588
rect 8113 8579 8171 8585
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 10870 8616 10876 8628
rect 10831 8588 10876 8616
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 12894 8616 12900 8628
rect 12855 8588 12900 8616
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 13722 8616 13728 8628
rect 13683 8588 13728 8616
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 14093 8619 14151 8625
rect 14093 8585 14105 8619
rect 14139 8616 14151 8619
rect 14645 8619 14703 8625
rect 14645 8616 14657 8619
rect 14139 8588 14657 8616
rect 14139 8585 14151 8588
rect 14093 8579 14151 8585
rect 14645 8585 14657 8588
rect 14691 8585 14703 8619
rect 15102 8616 15108 8628
rect 15063 8588 15108 8616
rect 14645 8579 14703 8585
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 15473 8619 15531 8625
rect 15473 8585 15485 8619
rect 15519 8585 15531 8619
rect 15473 8579 15531 8585
rect 3050 8508 3056 8560
rect 3108 8548 3114 8560
rect 3329 8551 3387 8557
rect 3329 8548 3341 8551
rect 3108 8520 3341 8548
rect 3108 8508 3114 8520
rect 3329 8517 3341 8520
rect 3375 8517 3387 8551
rect 3329 8511 3387 8517
rect 4157 8551 4215 8557
rect 4157 8517 4169 8551
rect 4203 8548 4215 8551
rect 4246 8548 4252 8560
rect 4203 8520 4252 8548
rect 4203 8517 4215 8520
rect 4157 8511 4215 8517
rect 4246 8508 4252 8520
rect 4304 8508 4310 8560
rect 6730 8548 6736 8560
rect 4356 8520 6736 8548
rect 2521 8483 2579 8489
rect 2521 8449 2533 8483
rect 2567 8480 2579 8483
rect 4356 8480 4384 8520
rect 6730 8508 6736 8520
rect 6788 8508 6794 8560
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 9585 8551 9643 8557
rect 9585 8548 9597 8551
rect 8352 8520 9597 8548
rect 8352 8508 8358 8520
rect 9585 8517 9597 8520
rect 9631 8517 9643 8551
rect 9585 8511 9643 8517
rect 11330 8508 11336 8560
rect 11388 8548 11394 8560
rect 13265 8551 13323 8557
rect 13265 8548 13277 8551
rect 11388 8520 13277 8548
rect 11388 8508 11394 8520
rect 13265 8517 13277 8520
rect 13311 8548 13323 8551
rect 13446 8548 13452 8560
rect 13311 8520 13452 8548
rect 13311 8517 13323 8520
rect 13265 8511 13323 8517
rect 13446 8508 13452 8520
rect 13504 8508 13510 8560
rect 14185 8551 14243 8557
rect 14185 8517 14197 8551
rect 14231 8548 14243 8551
rect 15488 8548 15516 8579
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 15841 8619 15899 8625
rect 15841 8616 15853 8619
rect 15620 8588 15853 8616
rect 15620 8576 15626 8588
rect 15841 8585 15853 8588
rect 15887 8616 15899 8619
rect 16206 8616 16212 8628
rect 15887 8588 16212 8616
rect 15887 8585 15899 8588
rect 15841 8579 15899 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16393 8619 16451 8625
rect 16393 8585 16405 8619
rect 16439 8616 16451 8619
rect 16482 8616 16488 8628
rect 16439 8588 16488 8616
rect 16439 8585 16451 8588
rect 16393 8579 16451 8585
rect 16482 8576 16488 8588
rect 16540 8576 16546 8628
rect 16914 8551 16972 8557
rect 16914 8548 16926 8551
rect 14231 8520 15516 8548
rect 15580 8520 16926 8548
rect 14231 8517 14243 8520
rect 14185 8511 14243 8517
rect 2567 8452 3280 8480
rect 2567 8449 2579 8452
rect 2521 8443 2579 8449
rect 2774 8372 2780 8424
rect 2832 8412 2838 8424
rect 3252 8412 3280 8452
rect 4264 8452 4384 8480
rect 4264 8424 4292 8452
rect 4982 8440 4988 8492
rect 5040 8480 5046 8492
rect 5914 8483 5972 8489
rect 5914 8480 5926 8483
rect 5040 8452 5926 8480
rect 5040 8440 5046 8452
rect 5914 8449 5926 8452
rect 5960 8449 5972 8483
rect 6178 8480 6184 8492
rect 6139 8452 6184 8480
rect 5914 8443 5972 8449
rect 6178 8440 6184 8452
rect 6236 8440 6242 8492
rect 7006 8480 7012 8492
rect 6967 8452 7012 8480
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 8754 8480 8760 8492
rect 7576 8452 8760 8480
rect 3510 8412 3516 8424
rect 2832 8384 2877 8412
rect 3252 8384 3516 8412
rect 2832 8372 2838 8384
rect 3510 8372 3516 8384
rect 3568 8412 3574 8424
rect 3605 8415 3663 8421
rect 3605 8412 3617 8415
rect 3568 8384 3617 8412
rect 3568 8372 3574 8384
rect 3605 8381 3617 8384
rect 3651 8412 3663 8415
rect 4246 8412 4252 8424
rect 3651 8384 4108 8412
rect 4159 8384 4252 8412
rect 3651 8381 3663 8384
rect 3605 8375 3663 8381
rect 4080 8356 4108 8384
rect 4246 8372 4252 8384
rect 4304 8372 4310 8424
rect 4341 8415 4399 8421
rect 4341 8381 4353 8415
rect 4387 8381 4399 8415
rect 4341 8375 4399 8381
rect 1394 8344 1400 8356
rect 1355 8316 1400 8344
rect 1394 8304 1400 8316
rect 1452 8304 1458 8356
rect 4062 8304 4068 8356
rect 4120 8344 4126 8356
rect 4356 8344 4384 8375
rect 6362 8372 6368 8424
rect 6420 8372 6426 8424
rect 7285 8415 7343 8421
rect 7285 8381 7297 8415
rect 7331 8412 7343 8415
rect 7466 8412 7472 8424
rect 7331 8384 7472 8412
rect 7331 8381 7343 8384
rect 7285 8375 7343 8381
rect 7466 8372 7472 8384
rect 7524 8372 7530 8424
rect 4120 8316 4384 8344
rect 4120 8304 4126 8316
rect 6178 8304 6184 8356
rect 6236 8344 6242 8356
rect 6380 8344 6408 8372
rect 6457 8347 6515 8353
rect 6457 8344 6469 8347
rect 6236 8316 6469 8344
rect 6236 8304 6242 8316
rect 6457 8313 6469 8316
rect 6503 8313 6515 8347
rect 6457 8307 6515 8313
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 7576 8353 7604 8452
rect 8754 8440 8760 8452
rect 8812 8440 8818 8492
rect 9237 8483 9295 8489
rect 9237 8449 9249 8483
rect 9283 8480 9295 8483
rect 9858 8480 9864 8492
rect 9283 8452 9864 8480
rect 9283 8449 9295 8452
rect 9237 8443 9295 8449
rect 9858 8440 9864 8452
rect 9916 8480 9922 8492
rect 10226 8480 10232 8492
rect 9916 8452 10232 8480
rect 9916 8440 9922 8452
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 11784 8483 11842 8489
rect 11784 8449 11796 8483
rect 11830 8480 11842 8483
rect 12526 8480 12532 8492
rect 11830 8452 12532 8480
rect 11830 8449 11842 8452
rect 11784 8443 11842 8449
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 12986 8440 12992 8492
rect 13044 8480 13050 8492
rect 13357 8483 13415 8489
rect 13357 8480 13369 8483
rect 13044 8452 13369 8480
rect 13044 8440 13050 8452
rect 13357 8449 13369 8452
rect 13403 8480 13415 8483
rect 14826 8480 14832 8492
rect 13403 8452 14832 8480
rect 13403 8449 13415 8452
rect 13357 8443 13415 8449
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 15010 8480 15016 8492
rect 14971 8452 15016 8480
rect 15010 8440 15016 8452
rect 15068 8440 15074 8492
rect 15102 8440 15108 8492
rect 15160 8480 15166 8492
rect 15580 8480 15608 8520
rect 16914 8517 16926 8520
rect 16960 8517 16972 8551
rect 16914 8511 16972 8517
rect 15160 8452 15608 8480
rect 15933 8483 15991 8489
rect 15160 8440 15166 8452
rect 15933 8449 15945 8483
rect 15979 8480 15991 8483
rect 16666 8480 16672 8492
rect 15979 8452 16252 8480
rect 16627 8452 16672 8480
rect 15979 8449 15991 8452
rect 15933 8443 15991 8449
rect 7837 8415 7895 8421
rect 7837 8381 7849 8415
rect 7883 8412 7895 8415
rect 8110 8412 8116 8424
rect 7883 8384 8116 8412
rect 7883 8381 7895 8384
rect 7837 8375 7895 8381
rect 8110 8372 8116 8384
rect 8168 8372 8174 8424
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8412 9551 8415
rect 9766 8412 9772 8424
rect 9539 8384 9772 8412
rect 9539 8381 9551 8384
rect 9493 8375 9551 8381
rect 9766 8372 9772 8384
rect 9824 8412 9830 8424
rect 11330 8412 11336 8424
rect 9824 8384 11336 8412
rect 9824 8372 9830 8384
rect 11330 8372 11336 8384
rect 11388 8412 11394 8424
rect 11517 8415 11575 8421
rect 11517 8412 11529 8415
rect 11388 8384 11529 8412
rect 11388 8372 11394 8384
rect 11517 8381 11529 8384
rect 11563 8381 11575 8415
rect 11517 8375 11575 8381
rect 12894 8372 12900 8424
rect 12952 8412 12958 8424
rect 13081 8415 13139 8421
rect 13081 8412 13093 8415
rect 12952 8384 13093 8412
rect 12952 8372 12958 8384
rect 13081 8381 13093 8384
rect 13127 8381 13139 8415
rect 13081 8375 13139 8381
rect 14001 8415 14059 8421
rect 14001 8381 14013 8415
rect 14047 8412 14059 8415
rect 14918 8412 14924 8424
rect 14047 8384 14924 8412
rect 14047 8381 14059 8384
rect 14001 8375 14059 8381
rect 14918 8372 14924 8384
rect 14976 8372 14982 8424
rect 15289 8415 15347 8421
rect 15289 8381 15301 8415
rect 15335 8381 15347 8415
rect 16114 8412 16120 8424
rect 16075 8384 16120 8412
rect 15289 8375 15347 8381
rect 7561 8347 7619 8353
rect 7561 8344 7573 8347
rect 6972 8316 7573 8344
rect 6972 8304 6978 8316
rect 7561 8313 7573 8316
rect 7607 8313 7619 8347
rect 7561 8307 7619 8313
rect 8021 8347 8079 8353
rect 8021 8313 8033 8347
rect 8067 8344 8079 8347
rect 8478 8344 8484 8356
rect 8067 8316 8484 8344
rect 8067 8313 8079 8316
rect 8021 8307 8079 8313
rect 8478 8304 8484 8316
rect 8536 8304 8542 8356
rect 11146 8344 11152 8356
rect 9600 8316 11152 8344
rect 1762 8236 1768 8288
rect 1820 8276 1826 8288
rect 3789 8279 3847 8285
rect 3789 8276 3801 8279
rect 1820 8248 3801 8276
rect 1820 8236 1826 8248
rect 3789 8245 3801 8248
rect 3835 8245 3847 8279
rect 3789 8239 3847 8245
rect 4614 8236 4620 8288
rect 4672 8276 4678 8288
rect 4709 8279 4767 8285
rect 4709 8276 4721 8279
rect 4672 8248 4721 8276
rect 4672 8236 4678 8248
rect 4709 8245 4721 8248
rect 4755 8276 4767 8279
rect 5258 8276 5264 8288
rect 4755 8248 5264 8276
rect 4755 8245 4767 8248
rect 4709 8239 4767 8245
rect 5258 8236 5264 8248
rect 5316 8236 5322 8288
rect 6362 8236 6368 8288
rect 6420 8276 6426 8288
rect 8846 8276 8852 8288
rect 6420 8248 8852 8276
rect 6420 8236 6426 8248
rect 8846 8236 8852 8248
rect 8904 8276 8910 8288
rect 9600 8276 9628 8316
rect 11146 8304 11152 8316
rect 11204 8304 11210 8356
rect 14936 8344 14964 8372
rect 15102 8344 15108 8356
rect 14936 8316 15108 8344
rect 15102 8304 15108 8316
rect 15160 8304 15166 8356
rect 15304 8344 15332 8375
rect 16114 8372 16120 8384
rect 16172 8372 16178 8424
rect 16224 8412 16252 8452
rect 16666 8440 16672 8452
rect 16724 8440 16730 8492
rect 17770 8480 17776 8492
rect 16776 8452 17776 8480
rect 16298 8412 16304 8424
rect 16224 8384 16304 8412
rect 16298 8372 16304 8384
rect 16356 8412 16362 8424
rect 16776 8412 16804 8452
rect 17770 8440 17776 8452
rect 17828 8440 17834 8492
rect 17954 8440 17960 8492
rect 18012 8480 18018 8492
rect 18141 8483 18199 8489
rect 18141 8480 18153 8483
rect 18012 8452 18153 8480
rect 18012 8440 18018 8452
rect 18141 8449 18153 8452
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 16356 8384 16804 8412
rect 16356 8372 16362 8384
rect 15378 8344 15384 8356
rect 15291 8316 15384 8344
rect 15378 8304 15384 8316
rect 15436 8344 15442 8356
rect 16132 8344 16160 8372
rect 15436 8316 16160 8344
rect 15436 8304 15442 8316
rect 17954 8304 17960 8356
rect 18012 8344 18018 8356
rect 18049 8347 18107 8353
rect 18049 8344 18061 8347
rect 18012 8316 18061 8344
rect 18012 8304 18018 8316
rect 18049 8313 18061 8316
rect 18095 8313 18107 8347
rect 18322 8344 18328 8356
rect 18283 8316 18328 8344
rect 18049 8307 18107 8313
rect 18322 8304 18328 8316
rect 18380 8304 18386 8356
rect 14550 8276 14556 8288
rect 8904 8248 9628 8276
rect 14511 8248 14556 8276
rect 8904 8236 8910 8248
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 14826 8236 14832 8288
rect 14884 8276 14890 8288
rect 15286 8276 15292 8288
rect 14884 8248 15292 8276
rect 14884 8236 14890 8248
rect 15286 8236 15292 8248
rect 15344 8236 15350 8288
rect 1104 8186 18860 8208
rect 1104 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 3430 8186
rect 3482 8134 7622 8186
rect 7674 8134 7686 8186
rect 7738 8134 7750 8186
rect 7802 8134 7814 8186
rect 7866 8134 7878 8186
rect 7930 8134 12070 8186
rect 12122 8134 12134 8186
rect 12186 8134 12198 8186
rect 12250 8134 12262 8186
rect 12314 8134 12326 8186
rect 12378 8134 16518 8186
rect 16570 8134 16582 8186
rect 16634 8134 16646 8186
rect 16698 8134 16710 8186
rect 16762 8134 16774 8186
rect 16826 8134 18860 8186
rect 1104 8112 18860 8134
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 4154 8072 4160 8084
rect 1636 8044 2544 8072
rect 4115 8044 4160 8072
rect 1636 8032 1642 8044
rect 1949 8007 2007 8013
rect 1949 7973 1961 8007
rect 1995 7973 2007 8007
rect 1949 7967 2007 7973
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7868 1915 7871
rect 1964 7868 1992 7967
rect 2130 7896 2136 7948
rect 2188 7936 2194 7948
rect 2516 7945 2544 8044
rect 4154 8032 4160 8044
rect 4212 8032 4218 8084
rect 4890 8072 4896 8084
rect 4264 8044 4896 8072
rect 3694 7964 3700 8016
rect 3752 8004 3758 8016
rect 4264 8004 4292 8044
rect 4890 8032 4896 8044
rect 4948 8072 4954 8084
rect 6178 8072 6184 8084
rect 4948 8044 6184 8072
rect 4948 8032 4954 8044
rect 6178 8032 6184 8044
rect 6236 8072 6242 8084
rect 6236 8044 6408 8072
rect 6236 8032 6242 8044
rect 4982 8004 4988 8016
rect 3752 7976 4292 8004
rect 4943 7976 4988 8004
rect 3752 7964 3758 7976
rect 4982 7964 4988 7976
rect 5040 7964 5046 8016
rect 2409 7939 2467 7945
rect 2409 7936 2421 7939
rect 2188 7908 2421 7936
rect 2188 7896 2194 7908
rect 2409 7905 2421 7908
rect 2455 7905 2467 7939
rect 2409 7899 2467 7905
rect 2501 7939 2559 7945
rect 2501 7905 2513 7939
rect 2547 7905 2559 7939
rect 3510 7936 3516 7948
rect 3471 7908 3516 7936
rect 2501 7899 2559 7905
rect 3510 7896 3516 7908
rect 3568 7896 3574 7948
rect 4798 7936 4804 7948
rect 4759 7908 4804 7936
rect 4798 7896 4804 7908
rect 4856 7896 4862 7948
rect 5166 7936 5172 7948
rect 4908 7908 5172 7936
rect 1903 7840 1992 7868
rect 1903 7837 1915 7840
rect 1857 7831 1915 7837
rect 2038 7828 2044 7880
rect 2096 7868 2102 7880
rect 2317 7871 2375 7877
rect 2317 7868 2329 7871
rect 2096 7840 2329 7868
rect 2096 7828 2102 7840
rect 2317 7837 2329 7840
rect 2363 7837 2375 7871
rect 2317 7831 2375 7837
rect 4065 7871 4123 7877
rect 4065 7837 4077 7871
rect 4111 7868 4123 7871
rect 4430 7868 4436 7880
rect 4111 7840 4436 7868
rect 4111 7837 4123 7840
rect 4065 7831 4123 7837
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 4908 7868 4936 7908
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 6380 7936 6408 8044
rect 6454 8032 6460 8084
rect 6512 8072 6518 8084
rect 6914 8072 6920 8084
rect 6512 8044 6920 8072
rect 6512 8032 6518 8044
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 11057 8075 11115 8081
rect 11057 8072 11069 8075
rect 9324 8044 11069 8072
rect 9125 8007 9183 8013
rect 9125 7973 9137 8007
rect 9171 8004 9183 8007
rect 9214 8004 9220 8016
rect 9171 7976 9220 8004
rect 9171 7973 9183 7976
rect 9125 7967 9183 7973
rect 9214 7964 9220 7976
rect 9272 7964 9278 8016
rect 7742 7936 7748 7948
rect 6380 7908 6776 7936
rect 7703 7908 7748 7936
rect 4571 7840 4936 7868
rect 5000 7840 6224 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 1210 7760 1216 7812
rect 1268 7800 1274 7812
rect 1581 7803 1639 7809
rect 1581 7800 1593 7803
rect 1268 7772 1593 7800
rect 1268 7760 1274 7772
rect 1581 7769 1593 7772
rect 1627 7769 1639 7803
rect 1581 7763 1639 7769
rect 3237 7803 3295 7809
rect 3237 7769 3249 7803
rect 3283 7800 3295 7803
rect 5000 7800 5028 7840
rect 6086 7800 6092 7812
rect 6144 7809 6150 7812
rect 3283 7772 5028 7800
rect 6056 7772 6092 7800
rect 3283 7769 3295 7772
rect 3237 7763 3295 7769
rect 6086 7760 6092 7772
rect 6144 7763 6156 7809
rect 6196 7800 6224 7840
rect 6270 7828 6276 7880
rect 6328 7868 6334 7880
rect 6748 7877 6776 7908
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 8386 7936 8392 7948
rect 8347 7908 8392 7936
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 8570 7936 8576 7948
rect 8531 7908 8576 7936
rect 8570 7896 8576 7908
rect 8628 7896 8634 7948
rect 6365 7871 6423 7877
rect 6365 7868 6377 7871
rect 6328 7840 6377 7868
rect 6328 7828 6334 7840
rect 6365 7837 6377 7840
rect 6411 7837 6423 7871
rect 6365 7831 6423 7837
rect 6733 7871 6791 7877
rect 6733 7837 6745 7871
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7868 7527 7871
rect 9324 7868 9352 8044
rect 11057 8041 11069 8044
rect 11103 8041 11115 8075
rect 12526 8072 12532 8084
rect 12487 8044 12532 8072
rect 11057 8035 11115 8041
rect 12526 8032 12532 8044
rect 12584 8032 12590 8084
rect 12897 8075 12955 8081
rect 12897 8041 12909 8075
rect 12943 8072 12955 8075
rect 13170 8072 13176 8084
rect 12943 8044 13176 8072
rect 12943 8041 12955 8044
rect 12897 8035 12955 8041
rect 13170 8032 13176 8044
rect 13228 8032 13234 8084
rect 13446 8032 13452 8084
rect 13504 8072 13510 8084
rect 13504 8044 16804 8072
rect 13504 8032 13510 8044
rect 9858 8004 9864 8016
rect 9508 7976 9864 8004
rect 9508 7945 9536 7976
rect 9858 7964 9864 7976
rect 9916 7964 9922 8016
rect 10137 8007 10195 8013
rect 10137 7973 10149 8007
rect 10183 8004 10195 8007
rect 10183 7976 11560 8004
rect 10183 7973 10195 7976
rect 10137 7967 10195 7973
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7905 9551 7939
rect 9674 7936 9680 7948
rect 9635 7908 9680 7936
rect 9493 7899 9551 7905
rect 9674 7896 9680 7908
rect 9732 7896 9738 7948
rect 9876 7936 9904 7964
rect 10321 7939 10379 7945
rect 10321 7936 10333 7939
rect 9876 7908 10333 7936
rect 10321 7905 10333 7908
rect 10367 7905 10379 7939
rect 10962 7936 10968 7948
rect 10321 7899 10379 7905
rect 10428 7908 10968 7936
rect 7515 7840 9352 7868
rect 7515 7837 7527 7840
rect 7469 7831 7527 7837
rect 9398 7828 9404 7880
rect 9456 7868 9462 7880
rect 9769 7871 9827 7877
rect 9769 7868 9781 7871
rect 9456 7840 9781 7868
rect 9456 7828 9462 7840
rect 9769 7837 9781 7840
rect 9815 7868 9827 7871
rect 10428 7868 10456 7908
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 11532 7945 11560 7976
rect 12434 7964 12440 8016
rect 12492 8004 12498 8016
rect 12989 8007 13047 8013
rect 12989 8004 13001 8007
rect 12492 7976 13001 8004
rect 12492 7964 12498 7976
rect 12989 7973 13001 7976
rect 13035 7973 13047 8007
rect 15378 8004 15384 8016
rect 12989 7967 13047 7973
rect 13372 7976 15384 8004
rect 11517 7939 11575 7945
rect 11517 7905 11529 7939
rect 11563 7905 11575 7939
rect 11698 7936 11704 7948
rect 11659 7908 11704 7936
rect 11517 7899 11575 7905
rect 11698 7896 11704 7908
rect 11756 7896 11762 7948
rect 13372 7945 13400 7976
rect 15378 7964 15384 7976
rect 15436 7964 15442 8016
rect 15473 8007 15531 8013
rect 15473 7973 15485 8007
rect 15519 8004 15531 8007
rect 15930 8004 15936 8016
rect 15519 7976 15936 8004
rect 15519 7973 15531 7976
rect 15473 7967 15531 7973
rect 13357 7939 13415 7945
rect 13357 7905 13369 7939
rect 13403 7905 13415 7939
rect 13357 7899 13415 7905
rect 14277 7939 14335 7945
rect 14277 7905 14289 7939
rect 14323 7905 14335 7939
rect 14277 7899 14335 7905
rect 14369 7939 14427 7945
rect 14369 7905 14381 7939
rect 14415 7936 14427 7939
rect 14550 7936 14556 7948
rect 14415 7908 14556 7936
rect 14415 7905 14427 7908
rect 14369 7899 14427 7905
rect 9815 7840 10456 7868
rect 10597 7871 10655 7877
rect 9815 7837 9827 7840
rect 9769 7831 9827 7837
rect 10597 7837 10609 7871
rect 10643 7868 10655 7871
rect 11238 7868 11244 7880
rect 10643 7840 11244 7868
rect 10643 7837 10655 7840
rect 10597 7831 10655 7837
rect 11238 7828 11244 7840
rect 11296 7828 11302 7880
rect 11885 7871 11943 7877
rect 11885 7837 11897 7871
rect 11931 7837 11943 7871
rect 14292 7868 14320 7899
rect 14550 7896 14556 7908
rect 14608 7896 14614 7948
rect 14642 7896 14648 7948
rect 14700 7936 14706 7948
rect 15488 7936 15516 7967
rect 15930 7964 15936 7976
rect 15988 7964 15994 8016
rect 16776 8004 16804 8044
rect 16850 8032 16856 8084
rect 16908 8072 16914 8084
rect 16945 8075 17003 8081
rect 16945 8072 16957 8075
rect 16908 8044 16957 8072
rect 16908 8032 16914 8044
rect 16945 8041 16957 8044
rect 16991 8041 17003 8075
rect 16945 8035 17003 8041
rect 18046 8032 18052 8084
rect 18104 8072 18110 8084
rect 18233 8075 18291 8081
rect 18233 8072 18245 8075
rect 18104 8044 18245 8072
rect 18104 8032 18110 8044
rect 18233 8041 18245 8044
rect 18279 8041 18291 8075
rect 18233 8035 18291 8041
rect 17678 8004 17684 8016
rect 16776 7976 17684 8004
rect 17678 7964 17684 7976
rect 17736 8004 17742 8016
rect 17736 7976 17816 8004
rect 17736 7964 17742 7976
rect 14700 7908 15516 7936
rect 14700 7896 14706 7908
rect 16298 7896 16304 7948
rect 16356 7936 16362 7948
rect 16758 7936 16764 7948
rect 16356 7908 16764 7936
rect 16356 7896 16362 7908
rect 16758 7896 16764 7908
rect 16816 7896 16822 7948
rect 17218 7896 17224 7948
rect 17276 7936 17282 7948
rect 17402 7936 17408 7948
rect 17276 7908 17408 7936
rect 17276 7896 17282 7908
rect 17402 7896 17408 7908
rect 17460 7896 17466 7948
rect 17586 7936 17592 7948
rect 17547 7908 17592 7936
rect 17586 7896 17592 7908
rect 17644 7896 17650 7948
rect 17788 7945 17816 7976
rect 17773 7939 17831 7945
rect 17773 7905 17785 7939
rect 17819 7936 17831 7939
rect 18325 7939 18383 7945
rect 18325 7936 18337 7939
rect 17819 7908 18337 7936
rect 17819 7905 17831 7908
rect 17773 7899 17831 7905
rect 18325 7905 18337 7908
rect 18371 7905 18383 7939
rect 18325 7899 18383 7905
rect 17126 7868 17132 7880
rect 14292 7840 17132 7868
rect 11885 7831 11943 7837
rect 6825 7803 6883 7809
rect 6825 7800 6837 7803
rect 6196 7772 6837 7800
rect 6825 7769 6837 7772
rect 6871 7769 6883 7803
rect 6825 7763 6883 7769
rect 8297 7803 8355 7809
rect 8297 7769 8309 7803
rect 8343 7800 8355 7803
rect 9582 7800 9588 7812
rect 8343 7772 9588 7800
rect 8343 7769 8355 7772
rect 8297 7763 8355 7769
rect 6144 7760 6150 7763
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 11425 7803 11483 7809
rect 11425 7800 11437 7803
rect 10980 7772 11437 7800
rect 2130 7692 2136 7744
rect 2188 7732 2194 7744
rect 2869 7735 2927 7741
rect 2869 7732 2881 7735
rect 2188 7704 2881 7732
rect 2188 7692 2194 7704
rect 2869 7701 2881 7704
rect 2915 7701 2927 7735
rect 2869 7695 2927 7701
rect 3326 7692 3332 7744
rect 3384 7732 3390 7744
rect 3878 7732 3884 7744
rect 3384 7704 3429 7732
rect 3839 7704 3884 7732
rect 3384 7692 3390 7704
rect 3878 7692 3884 7704
rect 3936 7692 3942 7744
rect 4614 7692 4620 7744
rect 4672 7732 4678 7744
rect 4672 7704 4717 7732
rect 4672 7692 4678 7704
rect 5902 7692 5908 7744
rect 5960 7732 5966 7744
rect 6549 7735 6607 7741
rect 6549 7732 6561 7735
rect 5960 7704 6561 7732
rect 5960 7692 5966 7704
rect 6549 7701 6561 7704
rect 6595 7701 6607 7735
rect 7098 7732 7104 7744
rect 7059 7704 7104 7732
rect 6549 7695 6607 7701
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 7561 7735 7619 7741
rect 7561 7701 7573 7735
rect 7607 7732 7619 7735
rect 7929 7735 7987 7741
rect 7929 7732 7941 7735
rect 7607 7704 7941 7732
rect 7607 7701 7619 7704
rect 7561 7695 7619 7701
rect 7929 7701 7941 7704
rect 7975 7701 7987 7735
rect 7929 7695 7987 7701
rect 9309 7735 9367 7741
rect 9309 7701 9321 7735
rect 9355 7732 9367 7735
rect 9674 7732 9680 7744
rect 9355 7704 9680 7732
rect 9355 7701 9367 7704
rect 9309 7695 9367 7701
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 10502 7732 10508 7744
rect 10463 7704 10508 7732
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 10980 7741 11008 7772
rect 11425 7769 11437 7772
rect 11471 7769 11483 7803
rect 11425 7763 11483 7769
rect 11606 7760 11612 7812
rect 11664 7800 11670 7812
rect 11900 7800 11928 7831
rect 17126 7828 17132 7840
rect 17184 7868 17190 7880
rect 17954 7868 17960 7880
rect 17184 7840 17960 7868
rect 17184 7828 17190 7840
rect 17954 7828 17960 7840
rect 18012 7828 18018 7880
rect 11664 7772 11928 7800
rect 13541 7803 13599 7809
rect 11664 7760 11670 7772
rect 13541 7769 13553 7803
rect 13587 7800 13599 7803
rect 14921 7803 14979 7809
rect 14921 7800 14933 7803
rect 13587 7772 14933 7800
rect 13587 7769 13599 7772
rect 13541 7763 13599 7769
rect 14921 7769 14933 7772
rect 14967 7769 14979 7803
rect 14921 7763 14979 7769
rect 15657 7803 15715 7809
rect 15657 7769 15669 7803
rect 15703 7800 15715 7803
rect 16298 7800 16304 7812
rect 15703 7772 16304 7800
rect 15703 7769 15715 7772
rect 15657 7763 15715 7769
rect 16298 7760 16304 7772
rect 16356 7760 16362 7812
rect 17862 7800 17868 7812
rect 17823 7772 17868 7800
rect 17862 7760 17868 7772
rect 17920 7760 17926 7812
rect 10965 7735 11023 7741
rect 10965 7701 10977 7735
rect 11011 7701 11023 7735
rect 10965 7695 11023 7701
rect 12713 7735 12771 7741
rect 12713 7701 12725 7735
rect 12759 7732 12771 7735
rect 12894 7732 12900 7744
rect 12759 7704 12900 7732
rect 12759 7701 12771 7704
rect 12713 7695 12771 7701
rect 12894 7692 12900 7704
rect 12952 7692 12958 7744
rect 13446 7732 13452 7744
rect 13407 7704 13452 7732
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13906 7732 13912 7744
rect 13867 7704 13912 7732
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 14182 7692 14188 7744
rect 14240 7732 14246 7744
rect 14461 7735 14519 7741
rect 14461 7732 14473 7735
rect 14240 7704 14473 7732
rect 14240 7692 14246 7704
rect 14461 7701 14473 7704
rect 14507 7701 14519 7735
rect 14826 7732 14832 7744
rect 14787 7704 14832 7732
rect 14461 7695 14519 7701
rect 14826 7692 14832 7704
rect 14884 7692 14890 7744
rect 15286 7732 15292 7744
rect 15199 7704 15292 7732
rect 15286 7692 15292 7704
rect 15344 7732 15350 7744
rect 15562 7732 15568 7744
rect 15344 7704 15568 7732
rect 15344 7692 15350 7704
rect 15562 7692 15568 7704
rect 15620 7732 15626 7744
rect 17880 7732 17908 7760
rect 15620 7704 17908 7732
rect 15620 7692 15626 7704
rect 1104 7642 18860 7664
rect 1104 7590 5398 7642
rect 5450 7590 5462 7642
rect 5514 7590 5526 7642
rect 5578 7590 5590 7642
rect 5642 7590 5654 7642
rect 5706 7590 9846 7642
rect 9898 7590 9910 7642
rect 9962 7590 9974 7642
rect 10026 7590 10038 7642
rect 10090 7590 10102 7642
rect 10154 7590 14294 7642
rect 14346 7590 14358 7642
rect 14410 7590 14422 7642
rect 14474 7590 14486 7642
rect 14538 7590 14550 7642
rect 14602 7590 18860 7642
rect 1104 7568 18860 7590
rect 1486 7528 1492 7540
rect 1447 7500 1492 7528
rect 1486 7488 1492 7500
rect 1544 7488 1550 7540
rect 3050 7488 3056 7540
rect 3108 7528 3114 7540
rect 4985 7531 5043 7537
rect 4985 7528 4997 7531
rect 3108 7500 4997 7528
rect 3108 7488 3114 7500
rect 4985 7497 4997 7500
rect 5031 7497 5043 7531
rect 4985 7491 5043 7497
rect 5258 7488 5264 7540
rect 5316 7528 5322 7540
rect 5316 7500 6868 7528
rect 5316 7488 5322 7500
rect 2774 7420 2780 7472
rect 2832 7460 2838 7472
rect 4341 7463 4399 7469
rect 2832 7432 2877 7460
rect 2832 7420 2838 7432
rect 4341 7429 4353 7463
rect 4387 7460 4399 7463
rect 5074 7460 5080 7472
rect 4387 7432 5080 7460
rect 4387 7429 4399 7432
rect 4341 7423 4399 7429
rect 5074 7420 5080 7432
rect 5132 7420 5138 7472
rect 5166 7420 5172 7472
rect 5224 7460 5230 7472
rect 5534 7460 5540 7472
rect 5224 7432 5540 7460
rect 5224 7420 5230 7432
rect 5534 7420 5540 7432
rect 5592 7420 5598 7472
rect 5626 7420 5632 7472
rect 5684 7460 5690 7472
rect 5721 7463 5779 7469
rect 5721 7460 5733 7463
rect 5684 7432 5733 7460
rect 5684 7420 5690 7432
rect 5721 7429 5733 7432
rect 5767 7429 5779 7463
rect 5721 7423 5779 7429
rect 1670 7392 1676 7404
rect 1631 7364 1676 7392
rect 1670 7352 1676 7364
rect 1728 7352 1734 7404
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7392 2191 7395
rect 2314 7392 2320 7404
rect 2179 7364 2320 7392
rect 2179 7361 2191 7364
rect 2133 7355 2191 7361
rect 2314 7352 2320 7364
rect 2372 7352 2378 7404
rect 4246 7352 4252 7404
rect 4304 7392 4310 7404
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 4304 7364 4445 7392
rect 4304 7352 4310 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 6178 7392 6184 7404
rect 5859 7364 6184 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 6178 7352 6184 7364
rect 6236 7352 6242 7404
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7392 6699 7395
rect 6730 7392 6736 7404
rect 6687 7364 6736 7392
rect 6687 7361 6699 7364
rect 6641 7355 6699 7361
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 6840 7392 6868 7500
rect 6914 7488 6920 7540
rect 6972 7528 6978 7540
rect 8481 7531 8539 7537
rect 6972 7500 7017 7528
rect 6972 7488 6978 7500
rect 8481 7497 8493 7531
rect 8527 7497 8539 7531
rect 8481 7491 8539 7497
rect 11885 7531 11943 7537
rect 11885 7497 11897 7531
rect 11931 7528 11943 7531
rect 12345 7531 12403 7537
rect 12345 7528 12357 7531
rect 11931 7500 12357 7528
rect 11931 7497 11943 7500
rect 11885 7491 11943 7497
rect 12345 7497 12357 7500
rect 12391 7497 12403 7531
rect 12345 7491 12403 7497
rect 12805 7531 12863 7537
rect 12805 7497 12817 7531
rect 12851 7528 12863 7531
rect 13173 7531 13231 7537
rect 13173 7528 13185 7531
rect 12851 7500 13185 7528
rect 12851 7497 12863 7500
rect 12805 7491 12863 7497
rect 13173 7497 13185 7500
rect 13219 7497 13231 7531
rect 13630 7528 13636 7540
rect 13591 7500 13636 7528
rect 13173 7491 13231 7497
rect 7285 7395 7343 7401
rect 7285 7392 7297 7395
rect 6840 7364 7297 7392
rect 7285 7361 7297 7364
rect 7331 7361 7343 7395
rect 7742 7392 7748 7404
rect 7655 7364 7748 7392
rect 7285 7355 7343 7361
rect 7742 7352 7748 7364
rect 7800 7392 7806 7404
rect 8496 7392 8524 7491
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 14182 7488 14188 7540
rect 14240 7528 14246 7540
rect 14277 7531 14335 7537
rect 14277 7528 14289 7531
rect 14240 7500 14289 7528
rect 14240 7488 14246 7500
rect 14277 7497 14289 7500
rect 14323 7497 14335 7531
rect 14277 7491 14335 7497
rect 16390 7488 16396 7540
rect 16448 7528 16454 7540
rect 16761 7531 16819 7537
rect 16761 7528 16773 7531
rect 16448 7500 16773 7528
rect 16448 7488 16454 7500
rect 16761 7497 16773 7500
rect 16807 7497 16819 7531
rect 17494 7528 17500 7540
rect 17455 7500 17500 7528
rect 16761 7491 16819 7497
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 18414 7528 18420 7540
rect 18375 7500 18420 7528
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 8570 7420 8576 7472
rect 8628 7460 8634 7472
rect 9616 7463 9674 7469
rect 9616 7460 9628 7463
rect 8628 7432 9628 7460
rect 8628 7420 8634 7432
rect 9616 7429 9628 7432
rect 9662 7460 9674 7463
rect 11698 7460 11704 7472
rect 9662 7432 11704 7460
rect 9662 7429 9674 7432
rect 9616 7423 9674 7429
rect 11698 7420 11704 7432
rect 11756 7420 11762 7472
rect 12526 7420 12532 7472
rect 12584 7460 12590 7472
rect 13648 7460 13676 7488
rect 12584 7432 13676 7460
rect 12584 7420 12590 7432
rect 13906 7420 13912 7472
rect 13964 7460 13970 7472
rect 14645 7463 14703 7469
rect 14645 7460 14657 7463
rect 13964 7432 14657 7460
rect 13964 7420 13970 7432
rect 14645 7429 14657 7432
rect 14691 7429 14703 7463
rect 16850 7460 16856 7472
rect 14645 7423 14703 7429
rect 15120 7432 16856 7460
rect 7800 7364 8524 7392
rect 7800 7352 7806 7364
rect 9766 7352 9772 7404
rect 9824 7392 9830 7404
rect 9861 7395 9919 7401
rect 9861 7392 9873 7395
rect 9824 7364 9873 7392
rect 9824 7352 9830 7364
rect 9861 7361 9873 7364
rect 9907 7392 9919 7395
rect 9953 7395 10011 7401
rect 9953 7392 9965 7395
rect 9907 7364 9965 7392
rect 9907 7361 9919 7364
rect 9861 7355 9919 7361
rect 9953 7361 9965 7364
rect 9999 7361 10011 7395
rect 9953 7355 10011 7361
rect 10042 7352 10048 7404
rect 10100 7392 10106 7404
rect 10220 7395 10278 7401
rect 10220 7392 10232 7395
rect 10100 7364 10232 7392
rect 10100 7352 10106 7364
rect 10220 7361 10232 7364
rect 10266 7392 10278 7395
rect 12710 7392 12716 7404
rect 10266 7364 12434 7392
rect 12671 7364 12716 7392
rect 10266 7361 10278 7364
rect 10220 7355 10278 7361
rect 12406 7336 12434 7364
rect 12710 7352 12716 7364
rect 12768 7352 12774 7404
rect 13541 7395 13599 7401
rect 13541 7361 13553 7395
rect 13587 7392 13599 7395
rect 13814 7392 13820 7404
rect 13587 7364 13820 7392
rect 13587 7361 13599 7364
rect 13541 7355 13599 7361
rect 13814 7352 13820 7364
rect 13872 7392 13878 7404
rect 14090 7392 14096 7404
rect 13872 7364 14096 7392
rect 13872 7352 13878 7364
rect 14090 7352 14096 7364
rect 14148 7352 14154 7404
rect 15120 7401 15148 7432
rect 16850 7420 16856 7432
rect 16908 7420 16914 7472
rect 15105 7395 15163 7401
rect 15105 7361 15117 7395
rect 15151 7361 15163 7395
rect 15105 7355 15163 7361
rect 15372 7395 15430 7401
rect 15372 7361 15384 7395
rect 15418 7392 15430 7395
rect 16114 7392 16120 7404
rect 15418 7364 16120 7392
rect 15418 7361 15430 7364
rect 15372 7355 15430 7361
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 17126 7352 17132 7404
rect 17184 7392 17190 7404
rect 17405 7395 17463 7401
rect 17405 7392 17417 7395
rect 17184 7364 17417 7392
rect 17184 7352 17190 7364
rect 17405 7361 17417 7364
rect 17451 7361 17463 7395
rect 17405 7355 17463 7361
rect 17586 7352 17592 7404
rect 17644 7392 17650 7404
rect 18141 7395 18199 7401
rect 18141 7392 18153 7395
rect 17644 7364 18153 7392
rect 17644 7352 17650 7364
rect 18141 7361 18153 7364
rect 18187 7361 18199 7395
rect 18141 7355 18199 7361
rect 18233 7395 18291 7401
rect 18233 7361 18245 7395
rect 18279 7392 18291 7395
rect 18279 7364 18460 7392
rect 18279 7361 18291 7364
rect 18233 7355 18291 7361
rect 18432 7336 18460 7364
rect 1949 7327 2007 7333
rect 1949 7293 1961 7327
rect 1995 7293 2007 7327
rect 1949 7287 2007 7293
rect 2041 7327 2099 7333
rect 2041 7293 2053 7327
rect 2087 7324 2099 7327
rect 4706 7324 4712 7336
rect 2087 7296 4712 7324
rect 2087 7293 2099 7296
rect 2041 7287 2099 7293
rect 1964 7256 1992 7287
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7293 4859 7327
rect 4801 7287 4859 7293
rect 4893 7327 4951 7333
rect 4893 7293 4905 7327
rect 4939 7324 4951 7327
rect 5258 7324 5264 7336
rect 4939 7296 5264 7324
rect 4939 7293 4951 7296
rect 4893 7287 4951 7293
rect 3510 7256 3516 7268
rect 1964 7228 3516 7256
rect 3510 7216 3516 7228
rect 3568 7216 3574 7268
rect 4816 7256 4844 7287
rect 5258 7284 5264 7296
rect 5316 7284 5322 7336
rect 5629 7327 5687 7333
rect 5629 7293 5641 7327
rect 5675 7293 5687 7327
rect 5629 7287 5687 7293
rect 5644 7256 5672 7287
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7377 7327 7435 7333
rect 7377 7324 7389 7327
rect 6972 7296 7389 7324
rect 6972 7284 6978 7296
rect 7377 7293 7389 7296
rect 7423 7293 7435 7327
rect 7377 7287 7435 7293
rect 7466 7284 7472 7336
rect 7524 7324 7530 7336
rect 11606 7324 11612 7336
rect 7524 7296 7569 7324
rect 11348 7296 11612 7324
rect 7524 7284 7530 7296
rect 6086 7256 6092 7268
rect 4816 7228 6092 7256
rect 6086 7216 6092 7228
rect 6144 7256 6150 7268
rect 6270 7256 6276 7268
rect 6144 7228 6276 7256
rect 6144 7216 6150 7228
rect 6270 7216 6276 7228
rect 6328 7216 6334 7268
rect 11348 7265 11376 7296
rect 11606 7284 11612 7296
rect 11664 7284 11670 7336
rect 11790 7324 11796 7336
rect 11751 7296 11796 7324
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 12406 7296 12440 7336
rect 12434 7284 12440 7296
rect 12492 7324 12498 7336
rect 12897 7327 12955 7333
rect 12897 7324 12909 7327
rect 12492 7296 12909 7324
rect 12492 7284 12498 7296
rect 12897 7293 12909 7296
rect 12943 7293 12955 7327
rect 12897 7287 12955 7293
rect 13722 7284 13728 7336
rect 13780 7324 13786 7336
rect 14001 7327 14059 7333
rect 13780 7296 13825 7324
rect 13780 7284 13786 7296
rect 14001 7293 14013 7327
rect 14047 7293 14059 7327
rect 14734 7324 14740 7336
rect 14695 7296 14740 7324
rect 14001 7287 14059 7293
rect 11333 7259 11391 7265
rect 11333 7225 11345 7259
rect 11379 7225 11391 7259
rect 11333 7219 11391 7225
rect 13078 7216 13084 7268
rect 13136 7256 13142 7268
rect 14016 7256 14044 7287
rect 14734 7284 14740 7296
rect 14792 7284 14798 7336
rect 14918 7324 14924 7336
rect 14879 7296 14924 7324
rect 14918 7284 14924 7296
rect 14976 7284 14982 7336
rect 18414 7284 18420 7336
rect 18472 7284 18478 7336
rect 13136 7228 14044 7256
rect 13136 7216 13142 7228
rect 2498 7188 2504 7200
rect 2459 7160 2504 7188
rect 2498 7148 2504 7160
rect 2556 7148 2562 7200
rect 5166 7148 5172 7200
rect 5224 7188 5230 7200
rect 5353 7191 5411 7197
rect 5353 7188 5365 7191
rect 5224 7160 5365 7188
rect 5224 7148 5230 7160
rect 5353 7157 5365 7160
rect 5399 7157 5411 7191
rect 6178 7188 6184 7200
rect 6139 7160 6184 7188
rect 5353 7151 5411 7157
rect 6178 7148 6184 7160
rect 6236 7148 6242 7200
rect 6454 7188 6460 7200
rect 6415 7160 6460 7188
rect 6454 7148 6460 7160
rect 6512 7148 6518 7200
rect 6638 7148 6644 7200
rect 6696 7188 6702 7200
rect 6733 7191 6791 7197
rect 6733 7188 6745 7191
rect 6696 7160 6745 7188
rect 6696 7148 6702 7160
rect 6733 7157 6745 7160
rect 6779 7188 6791 7191
rect 6914 7188 6920 7200
rect 6779 7160 6920 7188
rect 6779 7157 6791 7160
rect 6733 7151 6791 7157
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 8386 7188 8392 7200
rect 8347 7160 8392 7188
rect 8386 7148 8392 7160
rect 8444 7148 8450 7200
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 12253 7191 12311 7197
rect 12253 7188 12265 7191
rect 12032 7160 12265 7188
rect 12032 7148 12038 7160
rect 12253 7157 12265 7160
rect 12299 7157 12311 7191
rect 14936 7188 14964 7284
rect 16485 7191 16543 7197
rect 16485 7188 16497 7191
rect 14936 7160 16497 7188
rect 12253 7151 12311 7157
rect 16485 7157 16497 7160
rect 16531 7157 16543 7191
rect 16485 7151 16543 7157
rect 17494 7148 17500 7200
rect 17552 7188 17558 7200
rect 17862 7188 17868 7200
rect 17552 7160 17868 7188
rect 17552 7148 17558 7160
rect 17862 7148 17868 7160
rect 17920 7148 17926 7200
rect 1104 7098 18860 7120
rect 1104 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 3430 7098
rect 3482 7046 7622 7098
rect 7674 7046 7686 7098
rect 7738 7046 7750 7098
rect 7802 7046 7814 7098
rect 7866 7046 7878 7098
rect 7930 7046 12070 7098
rect 12122 7046 12134 7098
rect 12186 7046 12198 7098
rect 12250 7046 12262 7098
rect 12314 7046 12326 7098
rect 12378 7046 16518 7098
rect 16570 7046 16582 7098
rect 16634 7046 16646 7098
rect 16698 7046 16710 7098
rect 16762 7046 16774 7098
rect 16826 7046 18860 7098
rect 1104 7024 18860 7046
rect 2314 6944 2320 6996
rect 2372 6984 2378 6996
rect 2372 6956 5580 6984
rect 2372 6944 2378 6956
rect 5552 6916 5580 6956
rect 5994 6944 6000 6996
rect 6052 6984 6058 6996
rect 6549 6987 6607 6993
rect 6549 6984 6561 6987
rect 6052 6956 6561 6984
rect 6052 6944 6058 6956
rect 6549 6953 6561 6956
rect 6595 6953 6607 6987
rect 9953 6987 10011 6993
rect 6549 6947 6607 6953
rect 7116 6956 9904 6984
rect 7116 6916 7144 6956
rect 7282 6916 7288 6928
rect 5552 6888 7144 6916
rect 7208 6888 7288 6916
rect 3142 6808 3148 6860
rect 3200 6848 3206 6860
rect 3200 6820 3556 6848
rect 3200 6808 3206 6820
rect 3528 6789 3556 6820
rect 4982 6808 4988 6860
rect 5040 6848 5046 6860
rect 6178 6848 6184 6860
rect 5040 6820 6040 6848
rect 6139 6820 6184 6848
rect 5040 6808 5046 6820
rect 1581 6783 1639 6789
rect 1581 6749 1593 6783
rect 1627 6780 1639 6783
rect 3513 6783 3571 6789
rect 1627 6752 3372 6780
rect 1627 6749 1639 6752
rect 1581 6743 1639 6749
rect 1394 6672 1400 6724
rect 1452 6712 1458 6724
rect 1826 6715 1884 6721
rect 1826 6712 1838 6715
rect 1452 6684 1838 6712
rect 1452 6672 1458 6684
rect 1826 6681 1838 6684
rect 1872 6681 1884 6715
rect 1826 6675 1884 6681
rect 2774 6672 2780 6724
rect 2832 6712 2838 6724
rect 3237 6715 3295 6721
rect 3237 6712 3249 6715
rect 2832 6684 3249 6712
rect 2832 6672 2838 6684
rect 3237 6681 3249 6684
rect 3283 6681 3295 6715
rect 3344 6712 3372 6752
rect 3513 6749 3525 6783
rect 3559 6749 3571 6783
rect 3513 6743 3571 6749
rect 3881 6783 3939 6789
rect 3881 6749 3893 6783
rect 3927 6780 3939 6783
rect 3970 6780 3976 6792
rect 3927 6752 3976 6780
rect 3927 6749 3939 6752
rect 3881 6743 3939 6749
rect 3896 6712 3924 6743
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 5626 6780 5632 6792
rect 5587 6752 5632 6780
rect 5626 6740 5632 6752
rect 5684 6740 5690 6792
rect 6012 6780 6040 6820
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 7208 6857 7236 6888
rect 7282 6876 7288 6888
rect 7340 6876 7346 6928
rect 8938 6876 8944 6928
rect 8996 6916 9002 6928
rect 9876 6916 9904 6956
rect 9953 6953 9965 6987
rect 9999 6984 10011 6987
rect 10042 6984 10048 6996
rect 9999 6956 10048 6984
rect 9999 6953 10011 6956
rect 9953 6947 10011 6953
rect 10042 6944 10048 6956
rect 10100 6944 10106 6996
rect 10410 6984 10416 6996
rect 10323 6956 10416 6984
rect 10410 6944 10416 6956
rect 10468 6984 10474 6996
rect 10962 6984 10968 6996
rect 10468 6956 10968 6984
rect 10468 6944 10474 6956
rect 10962 6944 10968 6956
rect 11020 6944 11026 6996
rect 11517 6987 11575 6993
rect 11517 6953 11529 6987
rect 11563 6984 11575 6987
rect 11790 6984 11796 6996
rect 11563 6956 11796 6984
rect 11563 6953 11575 6956
rect 11517 6947 11575 6953
rect 11790 6944 11796 6956
rect 11848 6944 11854 6996
rect 12710 6984 12716 6996
rect 12671 6956 12716 6984
rect 12710 6944 12716 6956
rect 12768 6944 12774 6996
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 16850 6984 16856 6996
rect 12952 6956 15056 6984
rect 16811 6956 16856 6984
rect 12952 6944 12958 6956
rect 10428 6916 10456 6944
rect 12434 6916 12440 6928
rect 8996 6888 9168 6916
rect 9876 6888 10456 6916
rect 12176 6888 12440 6916
rect 8996 6876 9002 6888
rect 6273 6851 6331 6857
rect 6273 6817 6285 6851
rect 6319 6817 6331 6851
rect 6273 6811 6331 6817
rect 7193 6851 7251 6857
rect 7193 6817 7205 6851
rect 7239 6817 7251 6851
rect 9030 6848 9036 6860
rect 8991 6820 9036 6848
rect 7193 6811 7251 6817
rect 6288 6780 6316 6811
rect 9030 6808 9036 6820
rect 9088 6808 9094 6860
rect 9140 6848 9168 6888
rect 9490 6848 9496 6860
rect 9140 6820 9496 6848
rect 9490 6808 9496 6820
rect 9548 6848 9554 6860
rect 9769 6851 9827 6857
rect 9769 6848 9781 6851
rect 9548 6820 9781 6848
rect 9548 6808 9554 6820
rect 9769 6817 9781 6820
rect 9815 6817 9827 6851
rect 11330 6848 11336 6860
rect 11291 6820 11336 6848
rect 9769 6811 9827 6817
rect 11330 6808 11336 6820
rect 11388 6808 11394 6860
rect 12176 6857 12204 6888
rect 12434 6876 12440 6888
rect 12492 6876 12498 6928
rect 12618 6876 12624 6928
rect 12676 6916 12682 6928
rect 13446 6916 13452 6928
rect 12676 6888 13452 6916
rect 12676 6876 12682 6888
rect 13446 6876 13452 6888
rect 13504 6876 13510 6928
rect 15028 6916 15056 6956
rect 16850 6944 16856 6956
rect 16908 6944 16914 6996
rect 17405 6987 17463 6993
rect 17405 6953 17417 6987
rect 17451 6984 17463 6987
rect 17494 6984 17500 6996
rect 17451 6956 17500 6984
rect 17451 6953 17463 6956
rect 17405 6947 17463 6953
rect 17494 6944 17500 6956
rect 17552 6944 17558 6996
rect 18230 6916 18236 6928
rect 15028 6888 18236 6916
rect 18230 6876 18236 6888
rect 18288 6876 18294 6928
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6817 12219 6851
rect 13354 6848 13360 6860
rect 13267 6820 13360 6848
rect 12161 6811 12219 6817
rect 13354 6808 13360 6820
rect 13412 6848 13418 6860
rect 13722 6848 13728 6860
rect 13412 6820 13728 6848
rect 13412 6808 13418 6820
rect 13722 6808 13728 6820
rect 13780 6848 13786 6860
rect 16114 6848 16120 6860
rect 13780 6820 14228 6848
rect 16075 6820 16120 6848
rect 13780 6808 13786 6820
rect 6012 6752 6316 6780
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 7009 6783 7067 6789
rect 7009 6780 7021 6783
rect 6972 6752 7021 6780
rect 6972 6740 6978 6752
rect 7009 6749 7021 6752
rect 7055 6749 7067 6783
rect 7009 6743 7067 6749
rect 7374 6740 7380 6792
rect 7432 6780 7438 6792
rect 8018 6780 8024 6792
rect 7432 6752 8024 6780
rect 7432 6740 7438 6752
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 8757 6783 8815 6789
rect 8757 6780 8769 6783
rect 8260 6752 8769 6780
rect 8260 6740 8266 6752
rect 8757 6749 8769 6752
rect 8803 6749 8815 6783
rect 11238 6780 11244 6792
rect 8757 6743 8815 6749
rect 9048 6752 11244 6780
rect 4154 6721 4160 6724
rect 4148 6712 4160 6721
rect 3344 6684 3924 6712
rect 4115 6684 4160 6712
rect 3237 6675 3295 6681
rect 4148 6675 4160 6684
rect 4154 6672 4160 6675
rect 4212 6672 4218 6724
rect 4264 6684 5488 6712
rect 1302 6604 1308 6656
rect 1360 6644 1366 6656
rect 1489 6647 1547 6653
rect 1489 6644 1501 6647
rect 1360 6616 1501 6644
rect 1360 6604 1366 6616
rect 1489 6613 1501 6616
rect 1535 6644 1547 6647
rect 2682 6644 2688 6656
rect 1535 6616 2688 6644
rect 1535 6613 1547 6616
rect 1489 6607 1547 6613
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 2958 6644 2964 6656
rect 2919 6616 2964 6644
rect 2958 6604 2964 6616
rect 3016 6644 3022 6656
rect 3510 6644 3516 6656
rect 3016 6616 3516 6644
rect 3016 6604 3022 6616
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 3878 6604 3884 6656
rect 3936 6644 3942 6656
rect 4264 6644 4292 6684
rect 3936 6616 4292 6644
rect 3936 6604 3942 6616
rect 4890 6604 4896 6656
rect 4948 6644 4954 6656
rect 5460 6653 5488 6684
rect 5534 6672 5540 6724
rect 5592 6712 5598 6724
rect 8512 6715 8570 6721
rect 5592 6684 5764 6712
rect 5592 6672 5598 6684
rect 5736 6653 5764 6684
rect 8512 6681 8524 6715
rect 8558 6712 8570 6715
rect 9048 6712 9076 6752
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 12437 6783 12495 6789
rect 12437 6749 12449 6783
rect 12483 6780 12495 6783
rect 12526 6780 12532 6792
rect 12483 6752 12532 6780
rect 12483 6749 12495 6752
rect 12437 6743 12495 6749
rect 12526 6740 12532 6752
rect 12584 6740 12590 6792
rect 13078 6780 13084 6792
rect 13039 6752 13084 6780
rect 13078 6740 13084 6752
rect 13136 6740 13142 6792
rect 13538 6780 13544 6792
rect 13499 6752 13544 6780
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 13814 6780 13820 6792
rect 13775 6752 13820 6780
rect 13814 6740 13820 6752
rect 13872 6740 13878 6792
rect 14090 6780 14096 6792
rect 14051 6752 14096 6780
rect 14090 6740 14096 6752
rect 14148 6740 14154 6792
rect 14200 6780 14228 6820
rect 16114 6808 16120 6820
rect 16172 6808 16178 6860
rect 16206 6808 16212 6860
rect 16264 6848 16270 6860
rect 16393 6851 16451 6857
rect 16393 6848 16405 6851
rect 16264 6820 16405 6848
rect 16264 6808 16270 6820
rect 16393 6817 16405 6820
rect 16439 6817 16451 6851
rect 17954 6848 17960 6860
rect 16393 6811 16451 6817
rect 16960 6820 17960 6848
rect 15930 6780 15936 6792
rect 14200 6752 14504 6780
rect 15891 6752 15936 6780
rect 8558 6684 9076 6712
rect 8558 6681 8570 6684
rect 8512 6675 8570 6681
rect 9122 6672 9128 6724
rect 9180 6712 9186 6724
rect 9309 6715 9367 6721
rect 9309 6712 9321 6715
rect 9180 6684 9321 6712
rect 9180 6672 9186 6684
rect 9309 6681 9321 6684
rect 9355 6681 9367 6715
rect 11088 6715 11146 6721
rect 9309 6675 9367 6681
rect 9692 6684 11008 6712
rect 5261 6647 5319 6653
rect 5261 6644 5273 6647
rect 4948 6616 5273 6644
rect 4948 6604 4954 6616
rect 5261 6613 5273 6616
rect 5307 6613 5319 6647
rect 5261 6607 5319 6613
rect 5445 6647 5503 6653
rect 5445 6613 5457 6647
rect 5491 6613 5503 6647
rect 5445 6607 5503 6613
rect 5721 6647 5779 6653
rect 5721 6613 5733 6647
rect 5767 6613 5779 6647
rect 6086 6644 6092 6656
rect 6047 6616 6092 6644
rect 5721 6607 5779 6613
rect 6086 6604 6092 6616
rect 6144 6604 6150 6656
rect 6178 6604 6184 6656
rect 6236 6644 6242 6656
rect 6914 6644 6920 6656
rect 6236 6616 6920 6644
rect 6236 6604 6242 6616
rect 6914 6604 6920 6616
rect 6972 6604 6978 6656
rect 7374 6644 7380 6656
rect 7335 6616 7380 6644
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 9214 6644 9220 6656
rect 9175 6616 9220 6644
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 9692 6653 9720 6684
rect 9677 6647 9735 6653
rect 9677 6613 9689 6647
rect 9723 6613 9735 6647
rect 10980 6644 11008 6684
rect 11088 6681 11100 6715
rect 11134 6712 11146 6715
rect 13354 6712 13360 6724
rect 11134 6684 13360 6712
rect 11134 6681 11146 6684
rect 11088 6675 11146 6681
rect 13354 6672 13360 6684
rect 13412 6672 13418 6724
rect 13630 6672 13636 6724
rect 13688 6712 13694 6724
rect 14338 6715 14396 6721
rect 14338 6712 14350 6715
rect 13688 6684 14350 6712
rect 13688 6672 13694 6684
rect 14338 6681 14350 6684
rect 14384 6681 14396 6715
rect 14338 6675 14396 6681
rect 11422 6644 11428 6656
rect 10980 6616 11428 6644
rect 9677 6607 9735 6613
rect 11422 6604 11428 6616
rect 11480 6604 11486 6656
rect 11882 6644 11888 6656
rect 11843 6616 11888 6644
rect 11882 6604 11888 6616
rect 11940 6604 11946 6656
rect 11977 6647 12035 6653
rect 11977 6613 11989 6647
rect 12023 6644 12035 6647
rect 12158 6644 12164 6656
rect 12023 6616 12164 6644
rect 12023 6613 12035 6616
rect 11977 6607 12035 6613
rect 12158 6604 12164 6616
rect 12216 6604 12222 6656
rect 13173 6647 13231 6653
rect 13173 6613 13185 6647
rect 13219 6644 13231 6647
rect 13262 6644 13268 6656
rect 13219 6616 13268 6644
rect 13219 6613 13231 6616
rect 13173 6607 13231 6613
rect 13262 6604 13268 6616
rect 13320 6604 13326 6656
rect 14476 6644 14504 6752
rect 15930 6740 15936 6752
rect 15988 6780 15994 6792
rect 16960 6789 16988 6820
rect 17954 6808 17960 6820
rect 18012 6848 18018 6860
rect 18012 6820 18276 6848
rect 18012 6808 18018 6820
rect 16945 6783 17003 6789
rect 16945 6780 16957 6783
rect 15988 6752 16957 6780
rect 15988 6740 15994 6752
rect 16945 6749 16957 6752
rect 16991 6749 17003 6783
rect 16945 6743 17003 6749
rect 17126 6740 17132 6792
rect 17184 6780 17190 6792
rect 17497 6783 17555 6789
rect 17497 6780 17509 6783
rect 17184 6752 17509 6780
rect 17184 6740 17190 6752
rect 17497 6749 17509 6752
rect 17543 6749 17555 6783
rect 17497 6743 17555 6749
rect 17586 6740 17592 6792
rect 17644 6780 17650 6792
rect 18248 6789 18276 6820
rect 17865 6783 17923 6789
rect 17865 6780 17877 6783
rect 17644 6752 17877 6780
rect 17644 6740 17650 6752
rect 17865 6749 17877 6752
rect 17911 6749 17923 6783
rect 17865 6743 17923 6749
rect 18233 6783 18291 6789
rect 18233 6749 18245 6783
rect 18279 6749 18291 6783
rect 18233 6743 18291 6749
rect 14734 6672 14740 6724
rect 14792 6712 14798 6724
rect 14792 6684 15608 6712
rect 14792 6672 14798 6684
rect 15580 6653 15608 6684
rect 16298 6672 16304 6724
rect 16356 6712 16362 6724
rect 16577 6715 16635 6721
rect 16577 6712 16589 6715
rect 16356 6684 16589 6712
rect 16356 6672 16362 6684
rect 16577 6681 16589 6684
rect 16623 6681 16635 6715
rect 16577 6675 16635 6681
rect 17770 6672 17776 6724
rect 17828 6712 17834 6724
rect 17828 6684 18460 6712
rect 17828 6672 17834 6684
rect 15473 6647 15531 6653
rect 15473 6644 15485 6647
rect 14476 6616 15485 6644
rect 15473 6613 15485 6616
rect 15519 6613 15531 6647
rect 15473 6607 15531 6613
rect 15565 6647 15623 6653
rect 15565 6613 15577 6647
rect 15611 6613 15623 6647
rect 15565 6607 15623 6613
rect 16025 6647 16083 6653
rect 16025 6613 16037 6647
rect 16071 6644 16083 6647
rect 16114 6644 16120 6656
rect 16071 6616 16120 6644
rect 16071 6613 16083 6616
rect 16025 6607 16083 6613
rect 16114 6604 16120 6616
rect 16172 6644 16178 6656
rect 17129 6647 17187 6653
rect 17129 6644 17141 6647
rect 16172 6616 17141 6644
rect 16172 6604 16178 6616
rect 17129 6613 17141 6616
rect 17175 6613 17187 6647
rect 17678 6644 17684 6656
rect 17639 6616 17684 6644
rect 17129 6607 17187 6613
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 18049 6647 18107 6653
rect 18049 6613 18061 6647
rect 18095 6644 18107 6647
rect 18138 6644 18144 6656
rect 18095 6616 18144 6644
rect 18095 6613 18107 6616
rect 18049 6607 18107 6613
rect 18138 6604 18144 6616
rect 18196 6604 18202 6656
rect 18432 6653 18460 6684
rect 18417 6647 18475 6653
rect 18417 6613 18429 6647
rect 18463 6613 18475 6647
rect 18417 6607 18475 6613
rect 1104 6554 18860 6576
rect 1104 6502 5398 6554
rect 5450 6502 5462 6554
rect 5514 6502 5526 6554
rect 5578 6502 5590 6554
rect 5642 6502 5654 6554
rect 5706 6502 9846 6554
rect 9898 6502 9910 6554
rect 9962 6502 9974 6554
rect 10026 6502 10038 6554
rect 10090 6502 10102 6554
rect 10154 6502 14294 6554
rect 14346 6502 14358 6554
rect 14410 6502 14422 6554
rect 14474 6502 14486 6554
rect 14538 6502 14550 6554
rect 14602 6502 18860 6554
rect 1104 6480 18860 6502
rect 2225 6443 2283 6449
rect 2225 6409 2237 6443
rect 2271 6440 2283 6443
rect 2682 6440 2688 6452
rect 2271 6412 2688 6440
rect 2271 6409 2283 6412
rect 2225 6403 2283 6409
rect 2682 6400 2688 6412
rect 2740 6400 2746 6452
rect 4614 6440 4620 6452
rect 3528 6412 4384 6440
rect 4575 6412 4620 6440
rect 2317 6375 2375 6381
rect 2317 6341 2329 6375
rect 2363 6372 2375 6375
rect 3528 6372 3556 6412
rect 2363 6344 3556 6372
rect 2363 6341 2375 6344
rect 2317 6335 2375 6341
rect 3602 6332 3608 6384
rect 3660 6372 3666 6384
rect 3890 6375 3948 6381
rect 3890 6372 3902 6375
rect 3660 6344 3902 6372
rect 3660 6332 3666 6344
rect 3890 6341 3902 6344
rect 3936 6341 3948 6375
rect 3890 6335 3948 6341
rect 1762 6264 1768 6316
rect 1820 6304 1826 6316
rect 1857 6307 1915 6313
rect 1857 6304 1869 6307
rect 1820 6276 1869 6304
rect 1820 6264 1826 6276
rect 1857 6273 1869 6276
rect 1903 6273 1915 6307
rect 4246 6304 4252 6316
rect 1857 6267 1915 6273
rect 2700 6276 4252 6304
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 1946 6236 1952 6248
rect 1719 6208 1952 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 1946 6196 1952 6208
rect 2004 6196 2010 6248
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6205 2191 6239
rect 2133 6199 2191 6205
rect 2148 6100 2176 6199
rect 2700 6177 2728 6276
rect 4246 6264 4252 6276
rect 4304 6264 4310 6316
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6205 4215 6239
rect 4157 6199 4215 6205
rect 2685 6171 2743 6177
rect 2685 6137 2697 6171
rect 2731 6137 2743 6171
rect 2685 6131 2743 6137
rect 3142 6128 3148 6180
rect 3200 6128 3206 6180
rect 2777 6103 2835 6109
rect 2777 6100 2789 6103
rect 2148 6072 2789 6100
rect 2777 6069 2789 6072
rect 2823 6100 2835 6103
rect 2958 6100 2964 6112
rect 2823 6072 2964 6100
rect 2823 6069 2835 6072
rect 2777 6063 2835 6069
rect 2958 6060 2964 6072
rect 3016 6060 3022 6112
rect 3160 6100 3188 6128
rect 3510 6100 3516 6112
rect 3160 6072 3516 6100
rect 3510 6060 3516 6072
rect 3568 6060 3574 6112
rect 3970 6060 3976 6112
rect 4028 6100 4034 6112
rect 4163 6100 4191 6199
rect 4356 6168 4384 6412
rect 4614 6400 4620 6412
rect 4672 6400 4678 6452
rect 4985 6443 5043 6449
rect 4985 6409 4997 6443
rect 5031 6440 5043 6443
rect 5445 6443 5503 6449
rect 5445 6440 5457 6443
rect 5031 6412 5457 6440
rect 5031 6409 5043 6412
rect 4985 6403 5043 6409
rect 5445 6409 5457 6412
rect 5491 6409 5503 6443
rect 5810 6440 5816 6452
rect 5771 6412 5816 6440
rect 5445 6403 5503 6409
rect 5810 6400 5816 6412
rect 5868 6400 5874 6452
rect 6086 6400 6092 6452
rect 6144 6440 6150 6452
rect 7837 6443 7895 6449
rect 7837 6440 7849 6443
rect 6144 6412 7849 6440
rect 6144 6400 6150 6412
rect 7837 6409 7849 6412
rect 7883 6409 7895 6443
rect 7837 6403 7895 6409
rect 8110 6400 8116 6452
rect 8168 6440 8174 6452
rect 8205 6443 8263 6449
rect 8205 6440 8217 6443
rect 8168 6412 8217 6440
rect 8168 6400 8174 6412
rect 8205 6409 8217 6412
rect 8251 6409 8263 6443
rect 8662 6440 8668 6452
rect 8623 6412 8668 6440
rect 8205 6403 8263 6409
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 9033 6443 9091 6449
rect 9033 6440 9045 6443
rect 8812 6412 9045 6440
rect 8812 6400 8818 6412
rect 9033 6409 9045 6412
rect 9079 6409 9091 6443
rect 9033 6403 9091 6409
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 11793 6443 11851 6449
rect 11793 6440 11805 6443
rect 11664 6412 11805 6440
rect 11664 6400 11670 6412
rect 11793 6409 11805 6412
rect 11839 6409 11851 6443
rect 11793 6403 11851 6409
rect 11882 6400 11888 6452
rect 11940 6440 11946 6452
rect 11977 6443 12035 6449
rect 11977 6440 11989 6443
rect 11940 6412 11989 6440
rect 11940 6400 11946 6412
rect 11977 6409 11989 6412
rect 12023 6409 12035 6443
rect 11977 6403 12035 6409
rect 12158 6400 12164 6452
rect 12216 6440 12222 6452
rect 12805 6443 12863 6449
rect 12805 6440 12817 6443
rect 12216 6412 12817 6440
rect 12216 6400 12222 6412
rect 12805 6409 12817 6412
rect 12851 6409 12863 6443
rect 12805 6403 12863 6409
rect 13265 6443 13323 6449
rect 13265 6409 13277 6443
rect 13311 6440 13323 6443
rect 14461 6443 14519 6449
rect 14461 6440 14473 6443
rect 13311 6412 14473 6440
rect 13311 6409 13323 6412
rect 13265 6403 13323 6409
rect 14461 6409 14473 6412
rect 14507 6409 14519 6443
rect 14461 6403 14519 6409
rect 14921 6443 14979 6449
rect 14921 6409 14933 6443
rect 14967 6440 14979 6443
rect 15470 6440 15476 6452
rect 14967 6412 15476 6440
rect 14967 6409 14979 6412
rect 14921 6403 14979 6409
rect 15470 6400 15476 6412
rect 15528 6440 15534 6452
rect 15528 6412 16160 6440
rect 15528 6400 15534 6412
rect 5077 6375 5135 6381
rect 5077 6341 5089 6375
rect 5123 6372 5135 6375
rect 5166 6372 5172 6384
rect 5123 6344 5172 6372
rect 5123 6341 5135 6344
rect 5077 6335 5135 6341
rect 5166 6332 5172 6344
rect 5224 6332 5230 6384
rect 6914 6372 6920 6384
rect 6380 6344 6920 6372
rect 4522 6304 4528 6316
rect 4483 6276 4528 6304
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 4706 6264 4712 6316
rect 4764 6304 4770 6316
rect 6380 6313 6408 6344
rect 6914 6332 6920 6344
rect 6972 6332 6978 6384
rect 7926 6332 7932 6384
rect 7984 6372 7990 6384
rect 8570 6372 8576 6384
rect 7984 6344 8576 6372
rect 7984 6332 7990 6344
rect 8570 6332 8576 6344
rect 8628 6372 8634 6384
rect 11517 6375 11575 6381
rect 11517 6372 11529 6375
rect 8628 6344 9674 6372
rect 8628 6332 8634 6344
rect 6638 6313 6644 6316
rect 5905 6307 5963 6313
rect 5905 6304 5917 6307
rect 4764 6276 5917 6304
rect 4764 6264 4770 6276
rect 5905 6273 5917 6276
rect 5951 6273 5963 6307
rect 5905 6267 5963 6273
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6632 6267 6644 6313
rect 6696 6304 6702 6316
rect 6696 6276 6732 6304
rect 6638 6264 6644 6267
rect 6696 6264 6702 6276
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7432 6276 8432 6304
rect 7432 6264 7438 6276
rect 4982 6196 4988 6248
rect 5040 6236 5046 6248
rect 5169 6239 5227 6245
rect 5169 6236 5181 6239
rect 5040 6208 5181 6236
rect 5040 6196 5046 6208
rect 5169 6205 5181 6208
rect 5215 6205 5227 6239
rect 5169 6199 5227 6205
rect 6089 6239 6147 6245
rect 6089 6205 6101 6239
rect 6135 6236 6147 6239
rect 6270 6236 6276 6248
rect 6135 6208 6276 6236
rect 6135 6205 6147 6208
rect 6089 6199 6147 6205
rect 6270 6196 6276 6208
rect 6328 6236 6334 6248
rect 6328 6208 6408 6236
rect 6328 6196 6334 6208
rect 6178 6168 6184 6180
rect 4356 6140 6184 6168
rect 6178 6128 6184 6140
rect 6236 6128 6242 6180
rect 4028 6072 4191 6100
rect 4341 6103 4399 6109
rect 4028 6060 4034 6072
rect 4341 6069 4353 6103
rect 4387 6100 4399 6103
rect 4522 6100 4528 6112
rect 4387 6072 4528 6100
rect 4387 6069 4399 6072
rect 4341 6063 4399 6069
rect 4522 6060 4528 6072
rect 4580 6060 4586 6112
rect 6380 6100 6408 6208
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 8110 6236 8116 6248
rect 7524 6208 8116 6236
rect 7524 6196 7530 6208
rect 8110 6196 8116 6208
rect 8168 6236 8174 6248
rect 8404 6245 8432 6276
rect 8297 6239 8355 6245
rect 8297 6236 8309 6239
rect 8168 6208 8309 6236
rect 8168 6196 8174 6208
rect 8297 6205 8309 6208
rect 8343 6205 8355 6239
rect 8297 6199 8355 6205
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6205 8447 6239
rect 8389 6199 8447 6205
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 9125 6239 9183 6245
rect 9125 6236 9137 6239
rect 8996 6208 9137 6236
rect 8996 6196 9002 6208
rect 9125 6205 9137 6208
rect 9171 6205 9183 6239
rect 9306 6236 9312 6248
rect 9267 6208 9312 6236
rect 9125 6199 9183 6205
rect 9306 6196 9312 6208
rect 9364 6196 9370 6248
rect 7926 6168 7932 6180
rect 7760 6140 7932 6168
rect 7374 6100 7380 6112
rect 6380 6072 7380 6100
rect 7374 6060 7380 6072
rect 7432 6060 7438 6112
rect 7760 6109 7788 6140
rect 7926 6128 7932 6140
rect 7984 6128 7990 6180
rect 9646 6168 9674 6344
rect 9784 6344 11529 6372
rect 9784 6313 9812 6344
rect 11517 6341 11529 6344
rect 11563 6372 11575 6375
rect 12526 6372 12532 6384
rect 11563 6344 12532 6372
rect 11563 6341 11575 6344
rect 11517 6335 11575 6341
rect 12526 6332 12532 6344
rect 12584 6332 12590 6384
rect 13814 6332 13820 6384
rect 13872 6372 13878 6384
rect 14093 6375 14151 6381
rect 14093 6372 14105 6375
rect 13872 6344 14105 6372
rect 13872 6332 13878 6344
rect 14093 6341 14105 6344
rect 14139 6372 14151 6375
rect 15838 6372 15844 6384
rect 14139 6344 15844 6372
rect 14139 6341 14151 6344
rect 14093 6335 14151 6341
rect 15838 6332 15844 6344
rect 15896 6372 15902 6384
rect 16025 6375 16083 6381
rect 16025 6372 16037 6375
rect 15896 6344 16037 6372
rect 15896 6332 15902 6344
rect 16025 6341 16037 6344
rect 16071 6341 16083 6375
rect 16132 6372 16160 6412
rect 16206 6400 16212 6452
rect 16264 6440 16270 6452
rect 17037 6443 17095 6449
rect 17037 6440 17049 6443
rect 16264 6412 17049 6440
rect 16264 6400 16270 6412
rect 17037 6409 17049 6412
rect 17083 6440 17095 6443
rect 17678 6440 17684 6452
rect 17083 6412 17684 6440
rect 17083 6409 17095 6412
rect 17037 6403 17095 6409
rect 17678 6400 17684 6412
rect 17736 6400 17742 6452
rect 17862 6400 17868 6452
rect 17920 6440 17926 6452
rect 18417 6443 18475 6449
rect 18417 6440 18429 6443
rect 17920 6412 18429 6440
rect 17920 6400 17926 6412
rect 18417 6409 18429 6412
rect 18463 6409 18475 6443
rect 18417 6403 18475 6409
rect 16850 6372 16856 6384
rect 16132 6344 16344 6372
rect 16811 6344 16856 6372
rect 16025 6335 16083 6341
rect 9769 6307 9827 6313
rect 9769 6273 9781 6307
rect 9815 6273 9827 6307
rect 9769 6267 9827 6273
rect 10985 6307 11043 6313
rect 10985 6273 10997 6307
rect 11031 6304 11043 6307
rect 11146 6304 11152 6316
rect 11031 6276 11152 6304
rect 11031 6273 11043 6276
rect 10985 6267 11043 6273
rect 11146 6264 11152 6276
rect 11204 6264 11210 6316
rect 11241 6307 11299 6313
rect 11241 6273 11253 6307
rect 11287 6304 11299 6307
rect 11330 6304 11336 6316
rect 11287 6276 11336 6304
rect 11287 6273 11299 6276
rect 11241 6267 11299 6273
rect 11330 6264 11336 6276
rect 11388 6264 11394 6316
rect 11606 6264 11612 6316
rect 11664 6304 11670 6316
rect 12342 6304 12348 6316
rect 11664 6276 12348 6304
rect 11664 6264 11670 6276
rect 12342 6264 12348 6276
rect 12400 6264 12406 6316
rect 13170 6304 13176 6316
rect 13131 6276 13176 6304
rect 13170 6264 13176 6276
rect 13228 6264 13234 6316
rect 14001 6307 14059 6313
rect 14001 6273 14013 6307
rect 14047 6304 14059 6307
rect 14047 6276 14596 6304
rect 14047 6273 14059 6276
rect 14001 6267 14059 6273
rect 12437 6239 12495 6245
rect 12437 6205 12449 6239
rect 12483 6205 12495 6239
rect 12437 6199 12495 6205
rect 12621 6239 12679 6245
rect 12621 6205 12633 6239
rect 12667 6236 12679 6239
rect 13354 6236 13360 6248
rect 12667 6208 13360 6236
rect 12667 6205 12679 6208
rect 12621 6199 12679 6205
rect 12452 6168 12480 6199
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 13814 6196 13820 6248
rect 13872 6236 13878 6248
rect 14016 6236 14044 6267
rect 13872 6208 14044 6236
rect 14185 6239 14243 6245
rect 13872 6196 13878 6208
rect 14185 6205 14197 6239
rect 14231 6205 14243 6239
rect 14568 6236 14596 6276
rect 14642 6264 14648 6316
rect 14700 6304 14706 6316
rect 14829 6307 14887 6313
rect 14829 6304 14841 6307
rect 14700 6276 14841 6304
rect 14700 6264 14706 6276
rect 14829 6273 14841 6276
rect 14875 6273 14887 6307
rect 15194 6304 15200 6316
rect 14829 6267 14887 6273
rect 14936 6276 15200 6304
rect 14936 6236 14964 6276
rect 15194 6264 15200 6276
rect 15252 6264 15258 6316
rect 15289 6307 15347 6313
rect 15289 6273 15301 6307
rect 15335 6273 15347 6307
rect 15930 6304 15936 6316
rect 15891 6276 15936 6304
rect 15289 6267 15347 6273
rect 14568 6208 14964 6236
rect 15013 6239 15071 6245
rect 14185 6199 14243 6205
rect 15013 6205 15025 6239
rect 15059 6205 15071 6239
rect 15013 6199 15071 6205
rect 13633 6171 13691 6177
rect 13633 6168 13645 6171
rect 9646 6140 10364 6168
rect 12452 6140 13645 6168
rect 7745 6103 7803 6109
rect 7745 6069 7757 6103
rect 7791 6069 7803 6103
rect 9582 6100 9588 6112
rect 9543 6072 9588 6100
rect 7745 6063 7803 6069
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 9861 6103 9919 6109
rect 9861 6069 9873 6103
rect 9907 6100 9919 6103
rect 10226 6100 10232 6112
rect 9907 6072 10232 6100
rect 9907 6069 9919 6072
rect 9861 6063 9919 6069
rect 10226 6060 10232 6072
rect 10284 6060 10290 6112
rect 10336 6100 10364 6140
rect 13633 6137 13645 6140
rect 13679 6137 13691 6171
rect 13633 6131 13691 6137
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 14200 6168 14228 6199
rect 15028 6168 15056 6199
rect 13780 6140 15056 6168
rect 13780 6128 13786 6140
rect 15304 6100 15332 6267
rect 15930 6264 15936 6276
rect 15988 6264 15994 6316
rect 16316 6245 16344 6344
rect 16850 6332 16856 6344
rect 16908 6332 16914 6384
rect 16868 6304 16896 6332
rect 16592 6276 16896 6304
rect 16301 6239 16359 6245
rect 16301 6205 16313 6239
rect 16347 6236 16359 6239
rect 16390 6236 16396 6248
rect 16347 6208 16396 6236
rect 16347 6205 16359 6208
rect 16301 6199 16359 6205
rect 16390 6196 16396 6208
rect 16448 6196 16454 6248
rect 15378 6128 15384 6180
rect 15436 6168 15442 6180
rect 16485 6171 16543 6177
rect 16485 6168 16497 6171
rect 15436 6140 16497 6168
rect 15436 6128 15442 6140
rect 16485 6137 16497 6140
rect 16531 6137 16543 6171
rect 16485 6131 16543 6137
rect 10336 6072 15332 6100
rect 15930 6060 15936 6112
rect 15988 6100 15994 6112
rect 16592 6100 16620 6276
rect 17034 6264 17040 6316
rect 17092 6304 17098 6316
rect 17497 6307 17555 6313
rect 17497 6304 17509 6307
rect 17092 6276 17509 6304
rect 17092 6264 17098 6276
rect 17497 6273 17509 6276
rect 17543 6304 17555 6307
rect 17586 6304 17592 6316
rect 17543 6276 17592 6304
rect 17543 6273 17555 6276
rect 17497 6267 17555 6273
rect 17586 6264 17592 6276
rect 17644 6264 17650 6316
rect 17862 6304 17868 6316
rect 17823 6276 17868 6304
rect 17862 6264 17868 6276
rect 17920 6264 17926 6316
rect 18138 6264 18144 6316
rect 18196 6304 18202 6316
rect 18233 6307 18291 6313
rect 18233 6304 18245 6307
rect 18196 6276 18245 6304
rect 18196 6264 18202 6276
rect 18233 6273 18245 6276
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 16761 6239 16819 6245
rect 16761 6205 16773 6239
rect 16807 6236 16819 6239
rect 16850 6236 16856 6248
rect 16807 6208 16856 6236
rect 16807 6205 16819 6208
rect 16761 6199 16819 6205
rect 16850 6196 16856 6208
rect 16908 6196 16914 6248
rect 17773 6239 17831 6245
rect 17773 6205 17785 6239
rect 17819 6236 17831 6239
rect 18414 6236 18420 6248
rect 17819 6208 18420 6236
rect 17819 6205 17831 6208
rect 17773 6199 17831 6205
rect 18414 6196 18420 6208
rect 18472 6196 18478 6248
rect 18046 6168 18052 6180
rect 18007 6140 18052 6168
rect 18046 6128 18052 6140
rect 18104 6128 18110 6180
rect 15988 6072 16620 6100
rect 15988 6060 15994 6072
rect 17126 6060 17132 6112
rect 17184 6100 17190 6112
rect 17313 6103 17371 6109
rect 17313 6100 17325 6103
rect 17184 6072 17325 6100
rect 17184 6060 17190 6072
rect 17313 6069 17325 6072
rect 17359 6069 17371 6103
rect 17313 6063 17371 6069
rect 1104 6010 18860 6032
rect 1104 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 3430 6010
rect 3482 5958 7622 6010
rect 7674 5958 7686 6010
rect 7738 5958 7750 6010
rect 7802 5958 7814 6010
rect 7866 5958 7878 6010
rect 7930 5958 12070 6010
rect 12122 5958 12134 6010
rect 12186 5958 12198 6010
rect 12250 5958 12262 6010
rect 12314 5958 12326 6010
rect 12378 5958 16518 6010
rect 16570 5958 16582 6010
rect 16634 5958 16646 6010
rect 16698 5958 16710 6010
rect 16762 5958 16774 6010
rect 16826 5958 18860 6010
rect 1104 5936 18860 5958
rect 1581 5899 1639 5905
rect 1581 5865 1593 5899
rect 1627 5896 1639 5899
rect 1854 5896 1860 5908
rect 1627 5868 1860 5896
rect 1627 5865 1639 5868
rect 1581 5859 1639 5865
rect 1854 5856 1860 5868
rect 1912 5896 1918 5908
rect 2314 5896 2320 5908
rect 1912 5868 2320 5896
rect 1912 5856 1918 5868
rect 2314 5856 2320 5868
rect 2372 5856 2378 5908
rect 2590 5856 2596 5908
rect 2648 5896 2654 5908
rect 6086 5896 6092 5908
rect 2648 5868 6092 5896
rect 2648 5856 2654 5868
rect 6086 5856 6092 5868
rect 6144 5856 6150 5908
rect 6733 5899 6791 5905
rect 6733 5865 6745 5899
rect 6779 5896 6791 5899
rect 6914 5896 6920 5908
rect 6779 5868 6920 5896
rect 6779 5865 6791 5868
rect 6733 5859 6791 5865
rect 6914 5856 6920 5868
rect 6972 5896 6978 5908
rect 7374 5896 7380 5908
rect 6972 5868 7380 5896
rect 6972 5856 6978 5868
rect 7374 5856 7380 5868
rect 7432 5896 7438 5908
rect 8202 5896 8208 5908
rect 7432 5868 8208 5896
rect 7432 5856 7438 5868
rect 8202 5856 8208 5868
rect 8260 5896 8266 5908
rect 8260 5868 8524 5896
rect 8260 5856 8266 5868
rect 4890 5828 4896 5840
rect 2976 5800 4896 5828
rect 2976 5760 3004 5800
rect 4890 5788 4896 5800
rect 4948 5788 4954 5840
rect 5169 5831 5227 5837
rect 5169 5797 5181 5831
rect 5215 5828 5227 5831
rect 7466 5828 7472 5840
rect 5215 5800 7472 5828
rect 5215 5797 5227 5800
rect 5169 5791 5227 5797
rect 7466 5788 7472 5800
rect 7524 5788 7530 5840
rect 2884 5732 3004 5760
rect 2705 5695 2763 5701
rect 2705 5661 2717 5695
rect 2751 5692 2763 5695
rect 2884 5692 2912 5732
rect 3050 5720 3056 5772
rect 3108 5760 3114 5772
rect 8496 5769 8524 5868
rect 8846 5856 8852 5908
rect 8904 5896 8910 5908
rect 10873 5899 10931 5905
rect 8904 5868 10824 5896
rect 8904 5856 8910 5868
rect 10796 5828 10824 5868
rect 10873 5865 10885 5899
rect 10919 5896 10931 5899
rect 11330 5896 11336 5908
rect 10919 5868 11336 5896
rect 10919 5865 10931 5868
rect 10873 5859 10931 5865
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 12618 5896 12624 5908
rect 11440 5868 12624 5896
rect 11440 5828 11468 5868
rect 12618 5856 12624 5868
rect 12676 5856 12682 5908
rect 16393 5899 16451 5905
rect 16393 5896 16405 5899
rect 14200 5868 16405 5896
rect 14090 5828 14096 5840
rect 10796 5800 11468 5828
rect 13280 5800 14096 5828
rect 4525 5763 4583 5769
rect 4525 5760 4537 5763
rect 3108 5732 4537 5760
rect 3108 5720 3114 5732
rect 4525 5729 4537 5732
rect 4571 5760 4583 5763
rect 8481 5763 8539 5769
rect 4571 5732 5488 5760
rect 4571 5729 4583 5732
rect 4525 5723 4583 5729
rect 2751 5664 2912 5692
rect 2961 5695 3019 5701
rect 2751 5661 2763 5664
rect 2705 5655 2763 5661
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 3513 5695 3571 5701
rect 3007 5664 3372 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 3050 5584 3056 5636
rect 3108 5624 3114 5636
rect 3237 5627 3295 5633
rect 3237 5624 3249 5627
rect 3108 5596 3249 5624
rect 3108 5584 3114 5596
rect 3237 5593 3249 5596
rect 3283 5593 3295 5627
rect 3344 5624 3372 5664
rect 3513 5661 3525 5695
rect 3559 5692 3571 5695
rect 3694 5692 3700 5704
rect 3559 5664 3700 5692
rect 3559 5661 3571 5664
rect 3513 5655 3571 5661
rect 3694 5652 3700 5664
rect 3752 5652 3758 5704
rect 4341 5695 4399 5701
rect 4341 5661 4353 5695
rect 4387 5692 4399 5695
rect 4430 5692 4436 5704
rect 4387 5664 4436 5692
rect 4387 5661 4399 5664
rect 4341 5655 4399 5661
rect 4430 5652 4436 5664
rect 4488 5652 4494 5704
rect 4801 5695 4859 5701
rect 4801 5661 4813 5695
rect 4847 5692 4859 5695
rect 4982 5692 4988 5704
rect 4847 5664 4988 5692
rect 4847 5661 4859 5664
rect 4801 5655 4859 5661
rect 4982 5652 4988 5664
rect 5040 5652 5046 5704
rect 5074 5652 5080 5704
rect 5132 5692 5138 5704
rect 5261 5695 5319 5701
rect 5261 5692 5273 5695
rect 5132 5664 5273 5692
rect 5132 5652 5138 5664
rect 5261 5661 5273 5664
rect 5307 5661 5319 5695
rect 5460 5692 5488 5732
rect 8481 5729 8493 5763
rect 8527 5760 8539 5763
rect 8941 5763 8999 5769
rect 8941 5760 8953 5763
rect 8527 5732 8953 5760
rect 8527 5729 8539 5732
rect 8481 5723 8539 5729
rect 8941 5729 8953 5732
rect 8987 5729 8999 5763
rect 8941 5723 8999 5729
rect 5460 5664 8340 5692
rect 5261 5655 5319 5661
rect 3970 5624 3976 5636
rect 3344 5596 3976 5624
rect 3237 5587 3295 5593
rect 3970 5584 3976 5596
rect 4028 5584 4034 5636
rect 4062 5584 4068 5636
rect 4120 5624 4126 5636
rect 8214 5627 8272 5633
rect 4120 5596 4165 5624
rect 4120 5584 4126 5596
rect 8214 5593 8226 5627
rect 8260 5593 8272 5627
rect 8312 5624 8340 5664
rect 8386 5652 8392 5704
rect 8444 5692 8450 5704
rect 9197 5695 9255 5701
rect 9197 5692 9209 5695
rect 8444 5664 9209 5692
rect 8444 5652 8450 5664
rect 9197 5661 9209 5664
rect 9243 5661 9255 5695
rect 9197 5655 9255 5661
rect 11054 5652 11060 5704
rect 11112 5692 11118 5704
rect 12161 5695 12219 5701
rect 12161 5692 12173 5695
rect 11112 5664 12173 5692
rect 11112 5652 11118 5664
rect 12161 5661 12173 5664
rect 12207 5661 12219 5695
rect 12161 5655 12219 5661
rect 12253 5695 12311 5701
rect 12253 5661 12265 5695
rect 12299 5692 12311 5695
rect 13280 5692 13308 5800
rect 14090 5788 14096 5800
rect 14148 5788 14154 5840
rect 14200 5760 14228 5868
rect 16393 5865 16405 5868
rect 16439 5865 16451 5899
rect 17310 5896 17316 5908
rect 17271 5868 17316 5896
rect 16393 5859 16451 5865
rect 17310 5856 17316 5868
rect 17368 5856 17374 5908
rect 17773 5899 17831 5905
rect 17773 5865 17785 5899
rect 17819 5896 17831 5899
rect 17954 5896 17960 5908
rect 17819 5868 17960 5896
rect 17819 5865 17831 5868
rect 17773 5859 17831 5865
rect 17954 5856 17960 5868
rect 18012 5856 18018 5908
rect 14921 5831 14979 5837
rect 14921 5828 14933 5831
rect 12299 5664 13308 5692
rect 13464 5732 14228 5760
rect 14476 5800 14933 5828
rect 12299 5661 12311 5664
rect 12253 5655 12311 5661
rect 9030 5624 9036 5636
rect 8312 5596 9036 5624
rect 8214 5587 8272 5593
rect 1489 5559 1547 5565
rect 1489 5525 1501 5559
rect 1535 5556 1547 5559
rect 2590 5556 2596 5568
rect 1535 5528 2596 5556
rect 1535 5525 1547 5528
rect 1489 5519 1547 5525
rect 2590 5516 2596 5528
rect 2648 5516 2654 5568
rect 4706 5516 4712 5568
rect 4764 5556 4770 5568
rect 4764 5528 4809 5556
rect 4764 5516 4770 5528
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 7101 5559 7159 5565
rect 7101 5556 7113 5559
rect 6604 5528 7113 5556
rect 6604 5516 6610 5528
rect 7101 5525 7113 5528
rect 7147 5556 7159 5559
rect 7466 5556 7472 5568
rect 7147 5528 7472 5556
rect 7147 5525 7159 5528
rect 7101 5519 7159 5525
rect 7466 5516 7472 5528
rect 7524 5516 7530 5568
rect 8229 5556 8257 5587
rect 9030 5584 9036 5596
rect 9088 5584 9094 5636
rect 11330 5624 11336 5636
rect 10244 5596 11336 5624
rect 8570 5556 8576 5568
rect 8229 5528 8576 5556
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 8754 5556 8760 5568
rect 8715 5528 8760 5556
rect 8754 5516 8760 5528
rect 8812 5516 8818 5568
rect 8938 5516 8944 5568
rect 8996 5556 9002 5568
rect 10244 5556 10272 5596
rect 11330 5584 11336 5596
rect 11388 5584 11394 5636
rect 8996 5528 10272 5556
rect 10321 5559 10379 5565
rect 8996 5516 9002 5528
rect 10321 5525 10333 5559
rect 10367 5556 10379 5559
rect 10962 5556 10968 5568
rect 10367 5528 10968 5556
rect 10367 5525 10379 5528
rect 10321 5519 10379 5525
rect 10962 5516 10968 5528
rect 11020 5516 11026 5568
rect 12176 5556 12204 5655
rect 12520 5627 12578 5633
rect 12520 5593 12532 5627
rect 12566 5624 12578 5627
rect 13464 5624 13492 5732
rect 13538 5652 13544 5704
rect 13596 5692 13602 5704
rect 14366 5692 14372 5704
rect 13596 5664 14372 5692
rect 13596 5652 13602 5664
rect 14366 5652 14372 5664
rect 14424 5652 14430 5704
rect 14476 5701 14504 5800
rect 14921 5797 14933 5800
rect 14967 5797 14979 5831
rect 16850 5828 16856 5840
rect 14921 5791 14979 5797
rect 15120 5800 16856 5828
rect 14642 5760 14648 5772
rect 14603 5732 14648 5760
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 14734 5720 14740 5772
rect 14792 5760 14798 5772
rect 15120 5760 15148 5800
rect 16850 5788 16856 5800
rect 16908 5788 16914 5840
rect 14792 5732 15148 5760
rect 14792 5720 14798 5732
rect 15194 5720 15200 5772
rect 15252 5760 15258 5772
rect 15473 5763 15531 5769
rect 15473 5760 15485 5763
rect 15252 5732 15485 5760
rect 15252 5720 15258 5732
rect 15473 5729 15485 5732
rect 15519 5729 15531 5763
rect 15473 5723 15531 5729
rect 14461 5695 14519 5701
rect 14461 5661 14473 5695
rect 14507 5661 14519 5695
rect 14461 5655 14519 5661
rect 14550 5652 14556 5704
rect 14608 5692 14614 5704
rect 15749 5695 15807 5701
rect 15749 5692 15761 5695
rect 14608 5664 15761 5692
rect 14608 5652 14614 5664
rect 15749 5661 15761 5664
rect 15795 5661 15807 5695
rect 15749 5655 15807 5661
rect 17310 5652 17316 5704
rect 17368 5692 17374 5704
rect 17865 5695 17923 5701
rect 17865 5692 17877 5695
rect 17368 5664 17877 5692
rect 17368 5652 17374 5664
rect 17865 5661 17877 5664
rect 17911 5661 17923 5695
rect 18230 5692 18236 5704
rect 18191 5664 18236 5692
rect 17865 5655 17923 5661
rect 18230 5652 18236 5664
rect 18288 5652 18294 5704
rect 13817 5627 13875 5633
rect 13817 5624 13829 5627
rect 12566 5596 13492 5624
rect 13556 5596 13829 5624
rect 12566 5593 12578 5596
rect 12520 5587 12578 5593
rect 13556 5556 13584 5596
rect 13817 5593 13829 5596
rect 13863 5624 13875 5627
rect 14734 5624 14740 5636
rect 13863 5596 14740 5624
rect 13863 5593 13875 5596
rect 13817 5587 13875 5593
rect 14734 5584 14740 5596
rect 14792 5624 14798 5636
rect 16298 5624 16304 5636
rect 14792 5596 16304 5624
rect 14792 5584 14798 5596
rect 16298 5584 16304 5596
rect 16356 5584 16362 5636
rect 12176 5528 13584 5556
rect 13630 5516 13636 5568
rect 13688 5556 13694 5568
rect 13688 5528 13733 5556
rect 13688 5516 13694 5528
rect 13906 5516 13912 5568
rect 13964 5556 13970 5568
rect 14093 5559 14151 5565
rect 14093 5556 14105 5559
rect 13964 5528 14105 5556
rect 13964 5516 13970 5528
rect 14093 5525 14105 5528
rect 14139 5525 14151 5559
rect 14093 5519 14151 5525
rect 14553 5559 14611 5565
rect 14553 5525 14565 5559
rect 14599 5556 14611 5559
rect 14918 5556 14924 5568
rect 14599 5528 14924 5556
rect 14599 5525 14611 5528
rect 14553 5519 14611 5525
rect 14918 5516 14924 5528
rect 14976 5516 14982 5568
rect 15286 5556 15292 5568
rect 15247 5528 15292 5556
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 15378 5516 15384 5568
rect 15436 5556 15442 5568
rect 16485 5559 16543 5565
rect 16485 5556 16497 5559
rect 15436 5528 16497 5556
rect 15436 5516 15442 5528
rect 16485 5525 16497 5528
rect 16531 5556 16543 5559
rect 16666 5556 16672 5568
rect 16531 5528 16672 5556
rect 16531 5525 16543 5528
rect 16485 5519 16543 5525
rect 16666 5516 16672 5528
rect 16724 5516 16730 5568
rect 17034 5516 17040 5568
rect 17092 5556 17098 5568
rect 17497 5559 17555 5565
rect 17497 5556 17509 5559
rect 17092 5528 17509 5556
rect 17092 5516 17098 5528
rect 17497 5525 17509 5528
rect 17543 5556 17555 5559
rect 17862 5556 17868 5568
rect 17543 5528 17868 5556
rect 17543 5525 17555 5528
rect 17497 5519 17555 5525
rect 17862 5516 17868 5528
rect 17920 5516 17926 5568
rect 18046 5556 18052 5568
rect 18007 5528 18052 5556
rect 18046 5516 18052 5528
rect 18104 5516 18110 5568
rect 18414 5556 18420 5568
rect 18375 5528 18420 5556
rect 18414 5516 18420 5528
rect 18472 5516 18478 5568
rect 106 5448 112 5500
rect 164 5488 170 5500
rect 934 5488 940 5500
rect 164 5460 940 5488
rect 164 5448 170 5460
rect 934 5448 940 5460
rect 992 5448 998 5500
rect 1104 5466 18860 5488
rect 1104 5414 5398 5466
rect 5450 5414 5462 5466
rect 5514 5414 5526 5466
rect 5578 5414 5590 5466
rect 5642 5414 5654 5466
rect 5706 5414 9846 5466
rect 9898 5414 9910 5466
rect 9962 5414 9974 5466
rect 10026 5414 10038 5466
rect 10090 5414 10102 5466
rect 10154 5414 14294 5466
rect 14346 5414 14358 5466
rect 14410 5414 14422 5466
rect 14474 5414 14486 5466
rect 14538 5414 14550 5466
rect 14602 5414 18860 5466
rect 1104 5392 18860 5414
rect 2222 5352 2228 5364
rect 2183 5324 2228 5352
rect 2222 5312 2228 5324
rect 2280 5312 2286 5364
rect 4338 5352 4344 5364
rect 2424 5324 4344 5352
rect 2424 5284 2452 5324
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 4798 5312 4804 5364
rect 4856 5312 4862 5364
rect 4985 5355 5043 5361
rect 4985 5321 4997 5355
rect 5031 5352 5043 5355
rect 5353 5355 5411 5361
rect 5031 5324 5304 5352
rect 5031 5321 5043 5324
rect 4985 5315 5043 5321
rect 2590 5284 2596 5296
rect 1688 5256 2452 5284
rect 2503 5256 2596 5284
rect 1688 5225 1716 5256
rect 2590 5244 2596 5256
rect 2648 5284 2654 5296
rect 3878 5284 3884 5296
rect 2648 5256 3884 5284
rect 2648 5244 2654 5256
rect 3878 5244 3884 5256
rect 3936 5244 3942 5296
rect 4525 5287 4583 5293
rect 4525 5253 4537 5287
rect 4571 5284 4583 5287
rect 4816 5284 4844 5312
rect 4571 5256 4844 5284
rect 4571 5253 4583 5256
rect 4525 5247 4583 5253
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 1673 5179 1731 5185
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5216 2191 5219
rect 2498 5216 2504 5228
rect 2179 5188 2504 5216
rect 2179 5185 2191 5188
rect 2133 5179 2191 5185
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 4816 5216 4844 5256
rect 5276 5216 5304 5324
rect 5353 5321 5365 5355
rect 5399 5352 5411 5355
rect 5905 5355 5963 5361
rect 5905 5352 5917 5355
rect 5399 5324 5917 5352
rect 5399 5321 5411 5324
rect 5353 5315 5411 5321
rect 5905 5321 5917 5324
rect 5951 5321 5963 5355
rect 5905 5315 5963 5321
rect 7009 5355 7067 5361
rect 7009 5321 7021 5355
rect 7055 5321 7067 5355
rect 7009 5315 7067 5321
rect 7469 5355 7527 5361
rect 7469 5321 7481 5355
rect 7515 5352 7527 5355
rect 8662 5352 8668 5364
rect 7515 5324 8668 5352
rect 7515 5321 7527 5324
rect 7469 5315 7527 5321
rect 5813 5287 5871 5293
rect 5813 5253 5825 5287
rect 5859 5284 5871 5287
rect 7024 5284 7052 5315
rect 8662 5312 8668 5324
rect 8720 5312 8726 5364
rect 9033 5355 9091 5361
rect 9033 5321 9045 5355
rect 9079 5352 9091 5355
rect 9585 5355 9643 5361
rect 9585 5352 9597 5355
rect 9079 5324 9597 5352
rect 9079 5321 9091 5324
rect 9033 5315 9091 5321
rect 9585 5321 9597 5324
rect 9631 5321 9643 5355
rect 9585 5315 9643 5321
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 9953 5355 10011 5361
rect 9953 5352 9965 5355
rect 9732 5324 9965 5352
rect 9732 5312 9738 5324
rect 9953 5321 9965 5324
rect 9999 5321 10011 5355
rect 9953 5315 10011 5321
rect 10045 5355 10103 5361
rect 10045 5321 10057 5355
rect 10091 5352 10103 5355
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 10091 5324 10425 5352
rect 10091 5321 10103 5324
rect 10045 5315 10103 5321
rect 10413 5321 10425 5324
rect 10459 5321 10471 5355
rect 10413 5315 10471 5321
rect 10686 5312 10692 5364
rect 10744 5352 10750 5364
rect 10873 5355 10931 5361
rect 10873 5352 10885 5355
rect 10744 5324 10885 5352
rect 10744 5312 10750 5324
rect 10873 5321 10885 5324
rect 10919 5321 10931 5355
rect 10873 5315 10931 5321
rect 12989 5355 13047 5361
rect 12989 5321 13001 5355
rect 13035 5352 13047 5355
rect 13170 5352 13176 5364
rect 13035 5324 13176 5352
rect 13035 5321 13047 5324
rect 12989 5315 13047 5321
rect 13170 5312 13176 5324
rect 13228 5312 13234 5364
rect 13262 5312 13268 5364
rect 13320 5352 13326 5364
rect 13817 5355 13875 5361
rect 13817 5352 13829 5355
rect 13320 5324 13829 5352
rect 13320 5312 13326 5324
rect 13817 5321 13829 5324
rect 13863 5321 13875 5355
rect 15010 5352 15016 5364
rect 13817 5315 13875 5321
rect 14200 5324 15016 5352
rect 5859 5256 7052 5284
rect 7377 5287 7435 5293
rect 5859 5253 5871 5256
rect 5813 5247 5871 5253
rect 7377 5253 7389 5287
rect 7423 5284 7435 5287
rect 8386 5284 8392 5296
rect 7423 5256 8392 5284
rect 7423 5253 7435 5256
rect 7377 5247 7435 5253
rect 8386 5244 8392 5256
rect 8444 5244 8450 5296
rect 10594 5284 10600 5296
rect 8496 5256 10600 5284
rect 5350 5216 5356 5228
rect 4816 5188 5028 5216
rect 5276 5188 5356 5216
rect 1578 5108 1584 5160
rect 1636 5148 1642 5160
rect 2317 5151 2375 5157
rect 2317 5148 2329 5151
rect 1636 5120 2329 5148
rect 1636 5108 1642 5120
rect 2317 5117 2329 5120
rect 2363 5117 2375 5151
rect 2317 5111 2375 5117
rect 4709 5151 4767 5157
rect 4709 5117 4721 5151
rect 4755 5117 4767 5151
rect 4890 5148 4896 5160
rect 4851 5120 4896 5148
rect 4709 5111 4767 5117
rect 1489 5083 1547 5089
rect 1489 5049 1501 5083
rect 1535 5080 1547 5083
rect 2866 5080 2872 5092
rect 1535 5052 2872 5080
rect 1535 5049 1547 5052
rect 1489 5043 1547 5049
rect 2866 5040 2872 5052
rect 2924 5040 2930 5092
rect 1765 5015 1823 5021
rect 1765 4981 1777 5015
rect 1811 5012 1823 5015
rect 2038 5012 2044 5024
rect 1811 4984 2044 5012
rect 1811 4981 1823 4984
rect 1765 4975 1823 4981
rect 2038 4972 2044 4984
rect 2096 4972 2102 5024
rect 3881 5015 3939 5021
rect 3881 4981 3893 5015
rect 3927 5012 3939 5015
rect 3970 5012 3976 5024
rect 3927 4984 3976 5012
rect 3927 4981 3939 4984
rect 3881 4975 3939 4981
rect 3970 4972 3976 4984
rect 4028 4972 4034 5024
rect 4724 5012 4752 5111
rect 4890 5108 4896 5120
rect 4948 5108 4954 5160
rect 5000 5148 5028 5188
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 6917 5219 6975 5225
rect 6917 5185 6929 5219
rect 6963 5216 6975 5219
rect 7190 5216 7196 5228
rect 6963 5188 7196 5216
rect 6963 5185 6975 5188
rect 6917 5179 6975 5185
rect 7190 5176 7196 5188
rect 7248 5176 7254 5228
rect 8205 5219 8263 5225
rect 8205 5185 8217 5219
rect 8251 5216 8263 5219
rect 8496 5216 8524 5256
rect 10594 5244 10600 5256
rect 10652 5284 10658 5296
rect 10781 5287 10839 5293
rect 10781 5284 10793 5287
rect 10652 5256 10793 5284
rect 10652 5244 10658 5256
rect 10781 5253 10793 5256
rect 10827 5284 10839 5287
rect 11241 5287 11299 5293
rect 11241 5284 11253 5287
rect 10827 5256 11253 5284
rect 10827 5253 10839 5256
rect 10781 5247 10839 5253
rect 11241 5253 11253 5256
rect 11287 5253 11299 5287
rect 11241 5247 11299 5253
rect 11784 5287 11842 5293
rect 11784 5253 11796 5287
rect 11830 5284 11842 5287
rect 13722 5284 13728 5296
rect 11830 5256 13728 5284
rect 11830 5253 11842 5256
rect 11784 5247 11842 5253
rect 13722 5244 13728 5256
rect 13780 5244 13786 5296
rect 8251 5188 8524 5216
rect 9125 5219 9183 5225
rect 8251 5185 8263 5188
rect 8205 5179 8263 5185
rect 9125 5185 9137 5219
rect 9171 5216 9183 5219
rect 9766 5216 9772 5228
rect 9171 5188 9772 5216
rect 9171 5185 9183 5188
rect 9125 5179 9183 5185
rect 5994 5148 6000 5160
rect 5000 5120 5856 5148
rect 5955 5120 6000 5148
rect 5166 5040 5172 5092
rect 5224 5080 5230 5092
rect 5445 5083 5503 5089
rect 5445 5080 5457 5083
rect 5224 5052 5457 5080
rect 5224 5040 5230 5052
rect 5445 5049 5457 5052
rect 5491 5049 5503 5083
rect 5828 5080 5856 5120
rect 5994 5108 6000 5120
rect 6052 5108 6058 5160
rect 6733 5151 6791 5157
rect 6733 5117 6745 5151
rect 6779 5148 6791 5151
rect 7006 5148 7012 5160
rect 6779 5120 7012 5148
rect 6779 5117 6791 5120
rect 6733 5111 6791 5117
rect 7006 5108 7012 5120
rect 7064 5108 7070 5160
rect 7466 5108 7472 5160
rect 7524 5148 7530 5160
rect 7561 5151 7619 5157
rect 7561 5148 7573 5151
rect 7524 5120 7573 5148
rect 7524 5108 7530 5120
rect 7561 5117 7573 5120
rect 7607 5117 7619 5151
rect 8220 5148 8248 5179
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 13354 5216 13360 5228
rect 13315 5188 13360 5216
rect 13354 5176 13360 5188
rect 13412 5176 13418 5228
rect 13446 5176 13452 5228
rect 13504 5216 13510 5228
rect 14200 5216 14228 5324
rect 15010 5312 15016 5324
rect 15068 5312 15074 5364
rect 15286 5312 15292 5364
rect 15344 5352 15350 5364
rect 15565 5355 15623 5361
rect 15565 5352 15577 5355
rect 15344 5324 15577 5352
rect 15344 5312 15350 5324
rect 15565 5321 15577 5324
rect 15611 5321 15623 5355
rect 16022 5352 16028 5364
rect 15983 5324 16028 5352
rect 15565 5315 15623 5321
rect 16022 5312 16028 5324
rect 16080 5312 16086 5364
rect 16298 5352 16304 5364
rect 16259 5324 16304 5352
rect 16298 5312 16304 5324
rect 16356 5312 16362 5364
rect 16482 5352 16488 5364
rect 16443 5324 16488 5352
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 16666 5352 16672 5364
rect 16627 5324 16672 5352
rect 16666 5312 16672 5324
rect 16724 5312 16730 5364
rect 16850 5352 16856 5364
rect 16811 5324 16856 5352
rect 16850 5312 16856 5324
rect 16908 5312 16914 5364
rect 17678 5352 17684 5364
rect 17639 5324 17684 5352
rect 17678 5312 17684 5324
rect 17736 5312 17742 5364
rect 18230 5312 18236 5364
rect 18288 5352 18294 5364
rect 18417 5355 18475 5361
rect 18417 5352 18429 5355
rect 18288 5324 18429 5352
rect 18288 5312 18294 5324
rect 18417 5321 18429 5324
rect 18463 5321 18475 5355
rect 18417 5315 18475 5321
rect 14642 5244 14648 5296
rect 14700 5284 14706 5296
rect 15930 5284 15936 5296
rect 14700 5256 15240 5284
rect 15891 5256 15936 5284
rect 14700 5244 14706 5256
rect 14366 5225 14372 5228
rect 13504 5188 14228 5216
rect 13504 5176 13510 5188
rect 14360 5179 14372 5225
rect 14424 5216 14430 5228
rect 14424 5188 14460 5216
rect 14366 5176 14372 5179
rect 14424 5176 14430 5188
rect 7561 5111 7619 5117
rect 7668 5120 8248 5148
rect 8297 5151 8355 5157
rect 7668 5080 7696 5120
rect 8297 5117 8309 5151
rect 8343 5117 8355 5151
rect 8478 5148 8484 5160
rect 8439 5120 8484 5148
rect 8297 5111 8355 5117
rect 5828 5052 7696 5080
rect 5445 5043 5503 5049
rect 8110 5040 8116 5092
rect 8168 5080 8174 5092
rect 8312 5080 8340 5111
rect 8478 5108 8484 5120
rect 8536 5108 8542 5160
rect 8941 5151 8999 5157
rect 8941 5117 8953 5151
rect 8987 5148 8999 5151
rect 9674 5148 9680 5160
rect 8987 5120 9680 5148
rect 8987 5117 8999 5120
rect 8941 5111 8999 5117
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 10226 5148 10232 5160
rect 10187 5120 10232 5148
rect 10226 5108 10232 5120
rect 10284 5108 10290 5160
rect 10962 5108 10968 5160
rect 11020 5148 11026 5160
rect 11514 5148 11520 5160
rect 11020 5120 11065 5148
rect 11475 5120 11520 5148
rect 11020 5108 11026 5120
rect 11514 5108 11520 5120
rect 11572 5108 11578 5160
rect 13630 5148 13636 5160
rect 13591 5120 13636 5148
rect 13630 5108 13636 5120
rect 13688 5108 13694 5160
rect 14090 5148 14096 5160
rect 14051 5120 14096 5148
rect 14090 5108 14096 5120
rect 14148 5108 14154 5160
rect 10686 5080 10692 5092
rect 8168 5052 10692 5080
rect 8168 5040 8174 5052
rect 10686 5040 10692 5052
rect 10744 5040 10750 5092
rect 12897 5083 12955 5089
rect 12897 5049 12909 5083
rect 12943 5080 12955 5083
rect 13078 5080 13084 5092
rect 12943 5052 13084 5080
rect 12943 5049 12955 5052
rect 12897 5043 12955 5049
rect 13078 5040 13084 5052
rect 13136 5080 13142 5092
rect 13538 5080 13544 5092
rect 13136 5052 13544 5080
rect 13136 5040 13142 5052
rect 13538 5040 13544 5052
rect 13596 5040 13602 5092
rect 15212 5080 15240 5256
rect 15930 5244 15936 5256
rect 15988 5244 15994 5296
rect 16040 5284 16068 5312
rect 16206 5284 16212 5296
rect 16040 5256 16212 5284
rect 16206 5244 16212 5256
rect 16264 5244 16270 5296
rect 16500 5284 16528 5312
rect 17310 5284 17316 5296
rect 16500 5256 17316 5284
rect 17310 5244 17316 5256
rect 17368 5244 17374 5296
rect 17696 5216 17724 5312
rect 17865 5219 17923 5225
rect 17865 5216 17877 5219
rect 17696 5188 17877 5216
rect 17865 5185 17877 5188
rect 17911 5185 17923 5219
rect 17865 5179 17923 5185
rect 18138 5176 18144 5228
rect 18196 5216 18202 5228
rect 18233 5219 18291 5225
rect 18233 5216 18245 5219
rect 18196 5188 18245 5216
rect 18196 5176 18202 5188
rect 18233 5185 18245 5188
rect 18279 5185 18291 5219
rect 18233 5179 18291 5185
rect 15473 5083 15531 5089
rect 15473 5080 15485 5083
rect 15212 5052 15485 5080
rect 15473 5049 15485 5052
rect 15519 5049 15531 5083
rect 15473 5043 15531 5049
rect 4798 5012 4804 5024
rect 4724 4984 4804 5012
rect 4798 4972 4804 4984
rect 4856 4972 4862 5024
rect 5258 4972 5264 5024
rect 5316 5012 5322 5024
rect 7837 5015 7895 5021
rect 7837 5012 7849 5015
rect 5316 4984 7849 5012
rect 5316 4972 5322 4984
rect 7837 4981 7849 4984
rect 7883 4981 7895 5015
rect 7837 4975 7895 4981
rect 9398 4972 9404 5024
rect 9456 5012 9462 5024
rect 9493 5015 9551 5021
rect 9493 5012 9505 5015
rect 9456 4984 9505 5012
rect 9456 4972 9462 4984
rect 9493 4981 9505 4984
rect 9539 4981 9551 5015
rect 10704 5012 10732 5040
rect 11238 5012 11244 5024
rect 10704 4984 11244 5012
rect 9493 4975 9551 4981
rect 11238 4972 11244 4984
rect 11296 5012 11302 5024
rect 11882 5012 11888 5024
rect 11296 4984 11888 5012
rect 11296 4972 11302 4984
rect 11882 4972 11888 4984
rect 11940 5012 11946 5024
rect 15378 5012 15384 5024
rect 11940 4984 15384 5012
rect 11940 4972 11946 4984
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 18046 5012 18052 5024
rect 18007 4984 18052 5012
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 1104 4922 18860 4944
rect 1104 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 3430 4922
rect 3482 4870 7622 4922
rect 7674 4870 7686 4922
rect 7738 4870 7750 4922
rect 7802 4870 7814 4922
rect 7866 4870 7878 4922
rect 7930 4870 12070 4922
rect 12122 4870 12134 4922
rect 12186 4870 12198 4922
rect 12250 4870 12262 4922
rect 12314 4870 12326 4922
rect 12378 4870 16518 4922
rect 16570 4870 16582 4922
rect 16634 4870 16646 4922
rect 16698 4870 16710 4922
rect 16762 4870 16774 4922
rect 16826 4870 18860 4922
rect 1104 4848 18860 4870
rect 3878 4808 3884 4820
rect 3839 4780 3884 4808
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 10686 4808 10692 4820
rect 7248 4780 10692 4808
rect 7248 4768 7254 4780
rect 10686 4768 10692 4780
rect 10744 4768 10750 4820
rect 11146 4768 11152 4820
rect 11204 4808 11210 4820
rect 13909 4811 13967 4817
rect 13909 4808 13921 4811
rect 11204 4780 13921 4808
rect 11204 4768 11210 4780
rect 13909 4777 13921 4780
rect 13955 4777 13967 4811
rect 13909 4771 13967 4777
rect 15378 4768 15384 4820
rect 15436 4808 15442 4820
rect 16298 4808 16304 4820
rect 15436 4780 16304 4808
rect 15436 4768 15442 4780
rect 16298 4768 16304 4780
rect 16356 4808 16362 4820
rect 16669 4811 16727 4817
rect 16669 4808 16681 4811
rect 16356 4780 16681 4808
rect 16356 4768 16362 4780
rect 16669 4777 16681 4780
rect 16715 4777 16727 4811
rect 16669 4771 16727 4777
rect 16942 4768 16948 4820
rect 17000 4808 17006 4820
rect 17681 4811 17739 4817
rect 17681 4808 17693 4811
rect 17000 4780 17693 4808
rect 17000 4768 17006 4780
rect 17681 4777 17693 4780
rect 17727 4777 17739 4811
rect 17681 4771 17739 4777
rect 10962 4700 10968 4752
rect 11020 4740 11026 4752
rect 14918 4740 14924 4752
rect 11020 4712 12434 4740
rect 14879 4712 14924 4740
rect 11020 4700 11026 4712
rect 1578 4672 1584 4684
rect 1539 4644 1584 4672
rect 1578 4632 1584 4644
rect 1636 4632 1642 4684
rect 1670 4632 1676 4684
rect 1728 4672 1734 4684
rect 2130 4672 2136 4684
rect 1728 4644 1773 4672
rect 2056 4644 2136 4672
rect 1728 4632 1734 4644
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 2056 4604 2084 4644
rect 2130 4632 2136 4644
rect 2188 4632 2194 4684
rect 6825 4675 6883 4681
rect 6825 4641 6837 4675
rect 6871 4672 6883 4675
rect 7374 4672 7380 4684
rect 6871 4644 7380 4672
rect 6871 4641 6883 4644
rect 6825 4635 6883 4641
rect 7374 4632 7380 4644
rect 7432 4632 7438 4684
rect 11609 4675 11667 4681
rect 11609 4672 11621 4675
rect 10888 4644 11621 4672
rect 10888 4616 10916 4644
rect 11609 4641 11621 4644
rect 11655 4641 11667 4675
rect 11609 4635 11667 4641
rect 11882 4632 11888 4684
rect 11940 4672 11946 4684
rect 12161 4675 12219 4681
rect 12161 4672 12173 4675
rect 11940 4644 12173 4672
rect 11940 4632 11946 4644
rect 12161 4641 12173 4644
rect 12207 4641 12219 4675
rect 12161 4635 12219 4641
rect 1811 4576 2084 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 2222 4564 2228 4616
rect 2280 4604 2286 4616
rect 3970 4604 3976 4616
rect 2280 4576 3976 4604
rect 2280 4564 2286 4576
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 6546 4604 6552 4616
rect 6604 4613 6610 4616
rect 4856 4576 6552 4604
rect 4856 4564 4862 4576
rect 6546 4564 6552 4576
rect 6604 4567 6616 4613
rect 6604 4564 6610 4567
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 6788 4576 7205 4604
rect 6788 4564 6794 4576
rect 7193 4573 7205 4576
rect 7239 4604 7251 4607
rect 8018 4604 8024 4616
rect 7239 4576 8024 4604
rect 7239 4573 7251 4576
rect 7193 4567 7251 4573
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 9030 4604 9036 4616
rect 8991 4576 9036 4604
rect 9030 4564 9036 4576
rect 9088 4564 9094 4616
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 9640 4564 9674 4604
rect 10226 4564 10232 4616
rect 10284 4604 10290 4616
rect 10698 4607 10756 4613
rect 10698 4604 10710 4607
rect 10284 4576 10710 4604
rect 10284 4564 10290 4576
rect 10698 4573 10710 4576
rect 10744 4604 10756 4607
rect 10870 4604 10876 4616
rect 10744 4576 10876 4604
rect 10744 4573 10756 4576
rect 10698 4567 10756 4573
rect 10870 4564 10876 4576
rect 10928 4564 10934 4616
rect 10965 4607 11023 4613
rect 10965 4573 10977 4607
rect 11011 4604 11023 4607
rect 11514 4604 11520 4616
rect 11011 4576 11520 4604
rect 11011 4573 11023 4576
rect 10965 4567 11023 4573
rect 11514 4564 11520 4576
rect 11572 4564 11578 4616
rect 12406 4604 12434 4712
rect 14918 4700 14924 4712
rect 14976 4700 14982 4752
rect 15010 4700 15016 4752
rect 15068 4740 15074 4752
rect 15068 4712 15608 4740
rect 15068 4700 15074 4712
rect 13078 4672 13084 4684
rect 13039 4644 13084 4672
rect 13078 4632 13084 4644
rect 13136 4632 13142 4684
rect 14642 4672 14648 4684
rect 14603 4644 14648 4672
rect 14642 4632 14648 4644
rect 14700 4632 14706 4684
rect 15194 4632 15200 4684
rect 15252 4672 15258 4684
rect 15473 4675 15531 4681
rect 15473 4672 15485 4675
rect 15252 4644 15485 4672
rect 15252 4632 15258 4644
rect 15473 4641 15485 4644
rect 15519 4641 15531 4675
rect 15580 4672 15608 4712
rect 15654 4700 15660 4752
rect 15712 4740 15718 4752
rect 17221 4743 17279 4749
rect 17221 4740 17233 4743
rect 15712 4712 17233 4740
rect 15712 4700 15718 4712
rect 17221 4709 17233 4712
rect 17267 4709 17279 4743
rect 17221 4703 17279 4709
rect 17497 4675 17555 4681
rect 17497 4672 17509 4675
rect 15580 4644 17509 4672
rect 15473 4635 15531 4641
rect 17497 4641 17509 4644
rect 17543 4641 17555 4675
rect 17497 4635 17555 4641
rect 13265 4607 13323 4613
rect 13265 4604 13277 4607
rect 12406 4576 13277 4604
rect 13265 4573 13277 4576
rect 13311 4573 13323 4607
rect 13265 4567 13323 4573
rect 13814 4564 13820 4616
rect 13872 4604 13878 4616
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 13872 4576 15761 4604
rect 13872 4564 13878 4576
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 15930 4564 15936 4616
rect 15988 4604 15994 4616
rect 16390 4604 16396 4616
rect 15988 4576 16396 4604
rect 15988 4564 15994 4576
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 17696 4604 17724 4771
rect 17865 4607 17923 4613
rect 17865 4604 17877 4607
rect 17696 4576 17877 4604
rect 17865 4573 17877 4576
rect 17911 4573 17923 4607
rect 17865 4567 17923 4573
rect 2498 4545 2504 4548
rect 2492 4536 2504 4545
rect 2459 4508 2504 4536
rect 2492 4499 2504 4508
rect 2498 4496 2504 4499
rect 2556 4496 2562 4548
rect 4240 4539 4298 4545
rect 4240 4505 4252 4539
rect 4286 4536 4298 4539
rect 4338 4536 4344 4548
rect 4286 4508 4344 4536
rect 4286 4505 4298 4508
rect 4240 4499 4298 4505
rect 4338 4496 4344 4508
rect 4396 4496 4402 4548
rect 7622 4539 7680 4545
rect 7622 4536 7634 4539
rect 7392 4508 7634 4536
rect 2130 4468 2136 4480
rect 2091 4440 2136 4468
rect 2130 4428 2136 4440
rect 2188 4428 2194 4480
rect 3418 4428 3424 4480
rect 3476 4468 3482 4480
rect 3605 4471 3663 4477
rect 3605 4468 3617 4471
rect 3476 4440 3617 4468
rect 3476 4428 3482 4440
rect 3605 4437 3617 4440
rect 3651 4437 3663 4471
rect 3605 4431 3663 4437
rect 5074 4428 5080 4480
rect 5132 4468 5138 4480
rect 5353 4471 5411 4477
rect 5353 4468 5365 4471
rect 5132 4440 5365 4468
rect 5132 4428 5138 4440
rect 5353 4437 5365 4440
rect 5399 4437 5411 4471
rect 5353 4431 5411 4437
rect 5445 4471 5503 4477
rect 5445 4437 5457 4471
rect 5491 4468 5503 4471
rect 5994 4468 6000 4480
rect 5491 4440 6000 4468
rect 5491 4437 5503 4440
rect 5445 4431 5503 4437
rect 5994 4428 6000 4440
rect 6052 4428 6058 4480
rect 6822 4428 6828 4480
rect 6880 4468 6886 4480
rect 7009 4471 7067 4477
rect 7009 4468 7021 4471
rect 6880 4440 7021 4468
rect 6880 4428 6886 4440
rect 7009 4437 7021 4440
rect 7055 4437 7067 4471
rect 7009 4431 7067 4437
rect 7190 4428 7196 4480
rect 7248 4468 7254 4480
rect 7392 4468 7420 4508
rect 7622 4505 7634 4508
rect 7668 4505 7680 4539
rect 9306 4536 9312 4548
rect 9267 4508 9312 4536
rect 7622 4499 7680 4505
rect 9306 4496 9312 4508
rect 9364 4496 9370 4548
rect 9646 4536 9674 4564
rect 11146 4536 11152 4548
rect 9646 4508 11152 4536
rect 11146 4496 11152 4508
rect 11204 4496 11210 4548
rect 11425 4539 11483 4545
rect 11425 4505 11437 4539
rect 11471 4536 11483 4539
rect 11885 4539 11943 4545
rect 11885 4536 11897 4539
rect 11471 4508 11897 4536
rect 11471 4505 11483 4508
rect 11425 4499 11483 4505
rect 11885 4505 11897 4508
rect 11931 4505 11943 4539
rect 11885 4499 11943 4505
rect 12897 4539 12955 4545
rect 12897 4505 12909 4539
rect 12943 4536 12955 4539
rect 14461 4539 14519 4545
rect 12943 4508 14136 4536
rect 12943 4505 12955 4508
rect 12897 4499 12955 4505
rect 7248 4440 7420 4468
rect 7248 4428 7254 4440
rect 7466 4428 7472 4480
rect 7524 4468 7530 4480
rect 8110 4468 8116 4480
rect 7524 4440 8116 4468
rect 7524 4428 7530 4440
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 8662 4428 8668 4480
rect 8720 4468 8726 4480
rect 8757 4471 8815 4477
rect 8757 4468 8769 4471
rect 8720 4440 8769 4468
rect 8720 4428 8726 4440
rect 8757 4437 8769 4440
rect 8803 4437 8815 4471
rect 8757 4431 8815 4437
rect 9585 4471 9643 4477
rect 9585 4437 9597 4471
rect 9631 4468 9643 4471
rect 9674 4468 9680 4480
rect 9631 4440 9680 4468
rect 9631 4437 9643 4440
rect 9585 4431 9643 4437
rect 9674 4428 9680 4440
rect 9732 4468 9738 4480
rect 10318 4468 10324 4480
rect 9732 4440 10324 4468
rect 9732 4428 9738 4440
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 11054 4468 11060 4480
rect 11015 4440 11060 4468
rect 11054 4428 11060 4440
rect 11112 4428 11118 4480
rect 11517 4471 11575 4477
rect 11517 4437 11529 4471
rect 11563 4468 11575 4471
rect 11974 4468 11980 4480
rect 11563 4440 11980 4468
rect 11563 4437 11575 4440
rect 11517 4431 11575 4437
rect 11974 4428 11980 4440
rect 12032 4428 12038 4480
rect 12342 4428 12348 4480
rect 12400 4468 12406 4480
rect 12437 4471 12495 4477
rect 12437 4468 12449 4471
rect 12400 4440 12449 4468
rect 12400 4428 12406 4440
rect 12437 4437 12449 4440
rect 12483 4437 12495 4471
rect 12437 4431 12495 4437
rect 12805 4471 12863 4477
rect 12805 4437 12817 4471
rect 12851 4468 12863 4471
rect 13906 4468 13912 4480
rect 12851 4440 13912 4468
rect 12851 4437 12863 4440
rect 12805 4431 12863 4437
rect 13906 4428 13912 4440
rect 13964 4428 13970 4480
rect 14108 4477 14136 4508
rect 14461 4505 14473 4539
rect 14507 4536 14519 4539
rect 14642 4536 14648 4548
rect 14507 4508 14648 4536
rect 14507 4505 14519 4508
rect 14461 4499 14519 4505
rect 14642 4496 14648 4508
rect 14700 4496 14706 4548
rect 15289 4539 15347 4545
rect 15289 4536 15301 4539
rect 15212 4508 15301 4536
rect 14093 4471 14151 4477
rect 14093 4437 14105 4471
rect 14139 4437 14151 4471
rect 14093 4431 14151 4437
rect 14553 4471 14611 4477
rect 14553 4437 14565 4471
rect 14599 4468 14611 4471
rect 14826 4468 14832 4480
rect 14599 4440 14832 4468
rect 14599 4437 14611 4440
rect 14553 4431 14611 4437
rect 14826 4428 14832 4440
rect 14884 4428 14890 4480
rect 15102 4428 15108 4480
rect 15160 4468 15166 4480
rect 15212 4468 15240 4508
rect 15289 4505 15301 4508
rect 15335 4536 15347 4539
rect 16485 4539 16543 4545
rect 16485 4536 16497 4539
rect 15335 4508 16497 4536
rect 15335 4505 15347 4508
rect 15289 4499 15347 4505
rect 16485 4505 16497 4508
rect 16531 4536 16543 4539
rect 17126 4536 17132 4548
rect 16531 4508 17132 4536
rect 16531 4505 16543 4508
rect 16485 4499 16543 4505
rect 17126 4496 17132 4508
rect 17184 4496 17190 4548
rect 17954 4496 17960 4548
rect 18012 4536 18018 4548
rect 18417 4539 18475 4545
rect 18417 4536 18429 4539
rect 18012 4508 18429 4536
rect 18012 4496 18018 4508
rect 18417 4505 18429 4508
rect 18463 4505 18475 4539
rect 18417 4499 18475 4505
rect 15378 4468 15384 4480
rect 15160 4440 15240 4468
rect 15339 4440 15384 4468
rect 15160 4428 15166 4440
rect 15378 4428 15384 4440
rect 15436 4428 15442 4480
rect 15470 4428 15476 4480
rect 15528 4468 15534 4480
rect 16393 4471 16451 4477
rect 16393 4468 16405 4471
rect 15528 4440 16405 4468
rect 15528 4428 15534 4440
rect 16393 4437 16405 4440
rect 16439 4437 16451 4471
rect 16850 4468 16856 4480
rect 16811 4440 16856 4468
rect 16393 4431 16451 4437
rect 16850 4428 16856 4440
rect 16908 4428 16914 4480
rect 17034 4468 17040 4480
rect 16995 4440 17040 4468
rect 17034 4428 17040 4440
rect 17092 4428 17098 4480
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 18049 4471 18107 4477
rect 18049 4468 18061 4471
rect 17920 4440 18061 4468
rect 17920 4428 17926 4440
rect 18049 4437 18061 4440
rect 18095 4437 18107 4471
rect 18322 4468 18328 4480
rect 18283 4440 18328 4468
rect 18049 4431 18107 4437
rect 18322 4428 18328 4440
rect 18380 4428 18386 4480
rect 1104 4378 18860 4400
rect 1104 4326 5398 4378
rect 5450 4326 5462 4378
rect 5514 4326 5526 4378
rect 5578 4326 5590 4378
rect 5642 4326 5654 4378
rect 5706 4326 9846 4378
rect 9898 4326 9910 4378
rect 9962 4326 9974 4378
rect 10026 4326 10038 4378
rect 10090 4326 10102 4378
rect 10154 4326 14294 4378
rect 14346 4326 14358 4378
rect 14410 4326 14422 4378
rect 14474 4326 14486 4378
rect 14538 4326 14550 4378
rect 14602 4326 18860 4378
rect 1104 4304 18860 4326
rect 2130 4264 2136 4276
rect 2091 4236 2136 4264
rect 2130 4224 2136 4236
rect 2188 4224 2194 4276
rect 2593 4267 2651 4273
rect 2593 4233 2605 4267
rect 2639 4264 2651 4267
rect 4338 4264 4344 4276
rect 2639 4236 4344 4264
rect 2639 4233 2651 4236
rect 2593 4227 2651 4233
rect 4338 4224 4344 4236
rect 4396 4224 4402 4276
rect 4890 4224 4896 4276
rect 4948 4264 4954 4276
rect 5353 4267 5411 4273
rect 5353 4264 5365 4267
rect 4948 4236 5365 4264
rect 4948 4224 4954 4236
rect 5353 4233 5365 4236
rect 5399 4233 5411 4267
rect 8021 4267 8079 4273
rect 8021 4264 8033 4267
rect 5353 4227 5411 4233
rect 5460 4236 8033 4264
rect 2038 4156 2044 4208
rect 2096 4196 2102 4208
rect 2225 4199 2283 4205
rect 2225 4196 2237 4199
rect 2096 4168 2237 4196
rect 2096 4156 2102 4168
rect 2225 4165 2237 4168
rect 2271 4165 2283 4199
rect 2225 4159 2283 4165
rect 3418 4156 3424 4208
rect 3476 4196 3482 4208
rect 3694 4196 3700 4208
rect 3752 4205 3758 4208
rect 3476 4168 3700 4196
rect 3476 4156 3482 4168
rect 3694 4156 3700 4168
rect 3752 4159 3764 4205
rect 3752 4156 3758 4159
rect 3878 4156 3884 4208
rect 3936 4196 3942 4208
rect 5460 4196 5488 4236
rect 8021 4233 8033 4236
rect 8067 4233 8079 4267
rect 8386 4264 8392 4276
rect 8347 4236 8392 4264
rect 8021 4227 8079 4233
rect 8386 4224 8392 4236
rect 8444 4224 8450 4276
rect 8754 4264 8760 4276
rect 8715 4236 8760 4264
rect 8754 4224 8760 4236
rect 8812 4224 8818 4276
rect 10045 4267 10103 4273
rect 10045 4233 10057 4267
rect 10091 4264 10103 4267
rect 11054 4264 11060 4276
rect 10091 4236 11060 4264
rect 10091 4233 10103 4236
rect 10045 4227 10103 4233
rect 11054 4224 11060 4236
rect 11112 4224 11118 4276
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 13446 4264 13452 4276
rect 11204 4236 13452 4264
rect 11204 4224 11210 4236
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 14826 4224 14832 4276
rect 14884 4264 14890 4276
rect 15105 4267 15163 4273
rect 15105 4264 15117 4267
rect 14884 4236 15117 4264
rect 14884 4224 14890 4236
rect 15105 4233 15117 4236
rect 15151 4233 15163 4267
rect 15105 4227 15163 4233
rect 15473 4267 15531 4273
rect 15473 4233 15485 4267
rect 15519 4264 15531 4267
rect 15654 4264 15660 4276
rect 15519 4236 15660 4264
rect 15519 4233 15531 4236
rect 15473 4227 15531 4233
rect 15654 4224 15660 4236
rect 15712 4264 15718 4276
rect 16301 4267 16359 4273
rect 16301 4264 16313 4267
rect 15712 4236 16313 4264
rect 15712 4224 15718 4236
rect 16301 4233 16313 4236
rect 16347 4233 16359 4267
rect 16942 4264 16948 4276
rect 16903 4236 16948 4264
rect 16301 4227 16359 4233
rect 3936 4168 5488 4196
rect 5813 4199 5871 4205
rect 3936 4156 3942 4168
rect 5813 4165 5825 4199
rect 5859 4196 5871 4199
rect 6362 4196 6368 4208
rect 5859 4168 6368 4196
rect 5859 4165 5871 4168
rect 5813 4159 5871 4165
rect 6362 4156 6368 4168
rect 6420 4156 6426 4208
rect 7374 4156 7380 4208
rect 7432 4196 7438 4208
rect 10318 4196 10324 4208
rect 7432 4168 7880 4196
rect 10231 4168 10324 4196
rect 7432 4156 7438 4168
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4128 1731 4131
rect 2130 4128 2136 4140
rect 1719 4100 2136 4128
rect 1719 4097 1731 4100
rect 1673 4091 1731 4097
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 4249 4131 4307 4137
rect 4249 4097 4261 4131
rect 4295 4128 4307 4131
rect 4295 4100 4384 4128
rect 4295 4097 4307 4100
rect 4249 4091 4307 4097
rect 2409 4063 2467 4069
rect 2409 4029 2421 4063
rect 2455 4060 2467 4063
rect 3970 4060 3976 4072
rect 2455 4032 2774 4060
rect 3931 4032 3976 4060
rect 2455 4029 2467 4032
rect 2409 4023 2467 4029
rect 1486 3992 1492 4004
rect 1447 3964 1492 3992
rect 1486 3952 1492 3964
rect 1544 3952 1550 4004
rect 1762 3992 1768 4004
rect 1723 3964 1768 3992
rect 1762 3952 1768 3964
rect 1820 3952 1826 4004
rect 2746 3924 2774 4032
rect 3970 4020 3976 4032
rect 4028 4020 4034 4072
rect 3602 3924 3608 3936
rect 2746 3896 3608 3924
rect 3602 3884 3608 3896
rect 3660 3884 3666 3936
rect 4356 3924 4384 4100
rect 4430 4088 4436 4140
rect 4488 4128 4494 4140
rect 4525 4131 4583 4137
rect 4525 4128 4537 4131
rect 4488 4100 4537 4128
rect 4488 4088 4494 4100
rect 4525 4097 4537 4100
rect 4571 4097 4583 4131
rect 4890 4128 4896 4140
rect 4851 4100 4896 4128
rect 4525 4091 4583 4097
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 4985 4131 5043 4137
rect 4985 4097 4997 4131
rect 5031 4128 5043 4131
rect 5442 4128 5448 4140
rect 5031 4100 5448 4128
rect 5031 4097 5043 4100
rect 4985 4091 5043 4097
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 7852 4137 7880 4168
rect 10318 4156 10324 4168
rect 10376 4196 10382 4208
rect 10376 4168 11008 4196
rect 10376 4156 10382 4168
rect 7581 4131 7639 4137
rect 7581 4097 7593 4131
rect 7627 4128 7639 4131
rect 7837 4131 7895 4137
rect 7627 4100 7788 4128
rect 7627 4097 7639 4100
rect 7581 4091 7639 4097
rect 4709 4063 4767 4069
rect 4709 4029 4721 4063
rect 4755 4060 4767 4063
rect 5902 4060 5908 4072
rect 4755 4032 4844 4060
rect 4755 4029 4767 4032
rect 4709 4023 4767 4029
rect 4816 3992 4844 4032
rect 5000 4032 5764 4060
rect 5863 4032 5908 4060
rect 5000 3992 5028 4032
rect 4816 3964 5028 3992
rect 5258 3952 5264 4004
rect 5316 3992 5322 4004
rect 5445 3995 5503 4001
rect 5445 3992 5457 3995
rect 5316 3964 5457 3992
rect 5316 3952 5322 3964
rect 5445 3961 5457 3964
rect 5491 3961 5503 3995
rect 5736 3992 5764 4032
rect 5902 4020 5908 4032
rect 5960 4020 5966 4072
rect 5997 4063 6055 4069
rect 5997 4029 6009 4063
rect 6043 4060 6055 4063
rect 6546 4060 6552 4072
rect 6043 4032 6552 4060
rect 6043 4029 6055 4032
rect 5997 4023 6055 4029
rect 6012 3992 6040 4023
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 7760 4060 7788 4100
rect 7837 4097 7849 4131
rect 7883 4097 7895 4131
rect 8202 4128 8208 4140
rect 8163 4100 8208 4128
rect 7837 4091 7895 4097
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 9490 4128 9496 4140
rect 9451 4100 9496 4128
rect 9490 4088 9496 4100
rect 9548 4088 9554 4140
rect 8110 4060 8116 4072
rect 7760 4032 8116 4060
rect 8110 4020 8116 4032
rect 8168 4020 8174 4072
rect 8570 4020 8576 4072
rect 8628 4060 8634 4072
rect 10336 4069 10364 4156
rect 10778 4088 10784 4140
rect 10836 4128 10842 4140
rect 10873 4131 10931 4137
rect 10873 4128 10885 4131
rect 10836 4100 10885 4128
rect 10836 4088 10842 4100
rect 10873 4097 10885 4100
rect 10919 4097 10931 4131
rect 10980 4128 11008 4168
rect 11974 4156 11980 4208
rect 12032 4196 12038 4208
rect 14090 4196 14096 4208
rect 12032 4168 13308 4196
rect 12032 4156 12038 4168
rect 13280 4140 13308 4168
rect 13832 4168 14096 4196
rect 11773 4131 11831 4137
rect 11773 4128 11785 4131
rect 10980 4100 11785 4128
rect 10873 4091 10931 4097
rect 11773 4097 11785 4100
rect 11819 4097 11831 4131
rect 13262 4128 13268 4140
rect 13223 4100 13268 4128
rect 11773 4091 11831 4097
rect 13262 4088 13268 4100
rect 13320 4088 13326 4140
rect 13446 4088 13452 4140
rect 13504 4128 13510 4140
rect 13633 4131 13691 4137
rect 13633 4128 13645 4131
rect 13504 4100 13645 4128
rect 13504 4088 13510 4100
rect 13633 4097 13645 4100
rect 13679 4128 13691 4131
rect 13832 4128 13860 4168
rect 14090 4156 14096 4168
rect 14148 4156 14154 4208
rect 16316 4196 16344 4227
rect 16942 4224 16948 4236
rect 17000 4224 17006 4276
rect 17310 4264 17316 4276
rect 17271 4236 17316 4264
rect 17310 4224 17316 4236
rect 17368 4224 17374 4276
rect 17034 4196 17040 4208
rect 16316 4168 17040 4196
rect 17034 4156 17040 4168
rect 17092 4196 17098 4208
rect 17957 4199 18015 4205
rect 17957 4196 17969 4199
rect 17092 4168 17969 4196
rect 17092 4156 17098 4168
rect 17957 4165 17969 4168
rect 18003 4165 18015 4199
rect 17957 4159 18015 4165
rect 13679 4100 13860 4128
rect 13900 4131 13958 4137
rect 13679 4097 13691 4100
rect 13633 4091 13691 4097
rect 13900 4097 13912 4131
rect 13946 4128 13958 4131
rect 15378 4128 15384 4140
rect 13946 4100 15384 4128
rect 13946 4097 13958 4100
rect 13900 4091 13958 4097
rect 15378 4088 15384 4100
rect 15436 4088 15442 4140
rect 16114 4128 16120 4140
rect 16075 4100 16120 4128
rect 16114 4088 16120 4100
rect 16172 4088 16178 4140
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 18325 4131 18383 4137
rect 18325 4128 18337 4131
rect 16356 4100 18337 4128
rect 16356 4088 16362 4100
rect 18325 4097 18337 4100
rect 18371 4097 18383 4131
rect 18325 4091 18383 4097
rect 8849 4063 8907 4069
rect 8849 4060 8861 4063
rect 8628 4032 8861 4060
rect 8628 4020 8634 4032
rect 8849 4029 8861 4032
rect 8895 4029 8907 4063
rect 8849 4023 8907 4029
rect 8941 4063 8999 4069
rect 8941 4029 8953 4063
rect 8987 4029 8999 4063
rect 8941 4023 8999 4029
rect 10137 4063 10195 4069
rect 10137 4029 10149 4063
rect 10183 4029 10195 4063
rect 10137 4023 10195 4029
rect 10321 4063 10379 4069
rect 10321 4029 10333 4063
rect 10367 4029 10379 4063
rect 10962 4060 10968 4072
rect 10923 4032 10968 4060
rect 10321 4023 10379 4029
rect 6730 3992 6736 4004
rect 5736 3964 6040 3992
rect 6380 3964 6736 3992
rect 5445 3955 5503 3961
rect 6380 3924 6408 3964
rect 6730 3952 6736 3964
rect 6788 3952 6794 4004
rect 8386 3952 8392 4004
rect 8444 3992 8450 4004
rect 8662 3992 8668 4004
rect 8444 3964 8668 3992
rect 8444 3952 8450 3964
rect 8662 3952 8668 3964
rect 8720 3992 8726 4004
rect 8956 3992 8984 4023
rect 8720 3964 8984 3992
rect 8720 3952 8726 3964
rect 9214 3952 9220 4004
rect 9272 3992 9278 4004
rect 9309 3995 9367 4001
rect 9309 3992 9321 3995
rect 9272 3964 9321 3992
rect 9272 3952 9278 3964
rect 9309 3961 9321 3964
rect 9355 3961 9367 3995
rect 10152 3992 10180 4023
rect 10962 4020 10968 4032
rect 11020 4020 11026 4072
rect 11057 4063 11115 4069
rect 11057 4029 11069 4063
rect 11103 4029 11115 4063
rect 11514 4060 11520 4072
rect 11475 4032 11520 4060
rect 11057 4023 11115 4029
rect 10505 3995 10563 4001
rect 10505 3992 10517 3995
rect 10152 3964 10517 3992
rect 9309 3955 9367 3961
rect 10505 3961 10517 3964
rect 10551 3961 10563 3995
rect 10505 3955 10563 3961
rect 10870 3952 10876 4004
rect 10928 3992 10934 4004
rect 11072 3992 11100 4023
rect 11514 4020 11520 4032
rect 11572 4020 11578 4072
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4060 13139 4063
rect 13538 4060 13544 4072
rect 13127 4032 13544 4060
rect 13127 4029 13139 4032
rect 13081 4023 13139 4029
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 15562 4060 15568 4072
rect 15523 4032 15568 4060
rect 15562 4020 15568 4032
rect 15620 4020 15626 4072
rect 15657 4063 15715 4069
rect 15657 4029 15669 4063
rect 15703 4029 15715 4063
rect 15930 4060 15936 4072
rect 15891 4032 15936 4060
rect 15657 4023 15715 4029
rect 15194 3992 15200 4004
rect 10928 3964 11100 3992
rect 15028 3964 15200 3992
rect 10928 3952 10934 3964
rect 4356 3896 6408 3924
rect 6457 3927 6515 3933
rect 6457 3893 6469 3927
rect 6503 3924 6515 3927
rect 7190 3924 7196 3936
rect 6503 3896 7196 3924
rect 6503 3893 6515 3896
rect 6457 3887 6515 3893
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 9674 3924 9680 3936
rect 9635 3896 9680 3924
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 10318 3884 10324 3936
rect 10376 3924 10382 3936
rect 12897 3927 12955 3933
rect 12897 3924 12909 3927
rect 10376 3896 12909 3924
rect 10376 3884 10382 3896
rect 12897 3893 12909 3896
rect 12943 3924 12955 3927
rect 13814 3924 13820 3936
rect 12943 3896 13820 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 14274 3884 14280 3936
rect 14332 3924 14338 3936
rect 15028 3933 15056 3964
rect 15194 3952 15200 3964
rect 15252 3992 15258 4004
rect 15672 3992 15700 4023
rect 15930 4020 15936 4032
rect 15988 4020 15994 4072
rect 16761 4063 16819 4069
rect 16761 4029 16773 4063
rect 16807 4060 16819 4063
rect 16850 4060 16856 4072
rect 16807 4032 16856 4060
rect 16807 4029 16819 4032
rect 16761 4023 16819 4029
rect 16850 4020 16856 4032
rect 16908 4020 16914 4072
rect 16942 4020 16948 4072
rect 17000 4060 17006 4072
rect 17773 4063 17831 4069
rect 17773 4060 17785 4063
rect 17000 4032 17785 4060
rect 17000 4020 17006 4032
rect 17773 4029 17785 4032
rect 17819 4029 17831 4063
rect 17773 4023 17831 4029
rect 15252 3964 15700 3992
rect 15252 3952 15258 3964
rect 16022 3952 16028 4004
rect 16080 3992 16086 4004
rect 17589 3995 17647 4001
rect 17589 3992 17601 3995
rect 16080 3964 17601 3992
rect 16080 3952 16086 3964
rect 17589 3961 17601 3964
rect 17635 3961 17647 3995
rect 17589 3955 17647 3961
rect 15013 3927 15071 3933
rect 15013 3924 15025 3927
rect 14332 3896 15025 3924
rect 14332 3884 14338 3896
rect 15013 3893 15025 3896
rect 15059 3893 15071 3927
rect 15013 3887 15071 3893
rect 17129 3927 17187 3933
rect 17129 3893 17141 3927
rect 17175 3924 17187 3927
rect 17494 3924 17500 3936
rect 17175 3896 17500 3924
rect 17175 3893 17187 3896
rect 17129 3887 17187 3893
rect 17494 3884 17500 3896
rect 17552 3884 17558 3936
rect 18230 3924 18236 3936
rect 18191 3896 18236 3924
rect 18230 3884 18236 3896
rect 18288 3884 18294 3936
rect 1104 3834 18860 3856
rect 1104 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 3430 3834
rect 3482 3782 7622 3834
rect 7674 3782 7686 3834
rect 7738 3782 7750 3834
rect 7802 3782 7814 3834
rect 7866 3782 7878 3834
rect 7930 3782 12070 3834
rect 12122 3782 12134 3834
rect 12186 3782 12198 3834
rect 12250 3782 12262 3834
rect 12314 3782 12326 3834
rect 12378 3782 16518 3834
rect 16570 3782 16582 3834
rect 16634 3782 16646 3834
rect 16698 3782 16710 3834
rect 16762 3782 16774 3834
rect 16826 3782 18860 3834
rect 1104 3760 18860 3782
rect 3605 3723 3663 3729
rect 3605 3689 3617 3723
rect 3651 3720 3663 3723
rect 4154 3720 4160 3732
rect 3651 3692 4160 3720
rect 3651 3689 3663 3692
rect 3605 3683 3663 3689
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 4614 3720 4620 3732
rect 4575 3692 4620 3720
rect 4614 3680 4620 3692
rect 4672 3680 4678 3732
rect 5000 3692 5212 3720
rect 2498 3612 2504 3664
rect 2556 3652 2562 3664
rect 2869 3655 2927 3661
rect 2869 3652 2881 3655
rect 2556 3624 2881 3652
rect 2556 3612 2562 3624
rect 2869 3621 2881 3624
rect 2915 3652 2927 3655
rect 4430 3652 4436 3664
rect 2915 3624 4436 3652
rect 2915 3621 2927 3624
rect 2869 3615 2927 3621
rect 4430 3612 4436 3624
rect 4488 3612 4494 3664
rect 4525 3655 4583 3661
rect 4525 3621 4537 3655
rect 4571 3652 4583 3655
rect 4706 3652 4712 3664
rect 4571 3624 4712 3652
rect 4571 3621 4583 3624
rect 4525 3615 4583 3621
rect 4706 3612 4712 3624
rect 4764 3612 4770 3664
rect 3970 3584 3976 3596
rect 3931 3556 3976 3584
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 4065 3587 4123 3593
rect 4065 3553 4077 3587
rect 4111 3584 4123 3587
rect 4246 3584 4252 3596
rect 4111 3556 4252 3584
rect 4111 3553 4123 3556
rect 4065 3547 4123 3553
rect 4246 3544 4252 3556
rect 4304 3544 4310 3596
rect 5000 3584 5028 3692
rect 5184 3652 5212 3692
rect 5442 3680 5448 3732
rect 5500 3720 5506 3732
rect 7929 3723 7987 3729
rect 7929 3720 7941 3723
rect 5500 3692 7941 3720
rect 5500 3680 5506 3692
rect 7929 3689 7941 3692
rect 7975 3689 7987 3723
rect 7929 3683 7987 3689
rect 8941 3723 8999 3729
rect 8941 3689 8953 3723
rect 8987 3720 8999 3723
rect 9030 3720 9036 3732
rect 8987 3692 9036 3720
rect 8987 3689 8999 3692
rect 8941 3683 8999 3689
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 9769 3723 9827 3729
rect 9769 3720 9781 3723
rect 9640 3692 9781 3720
rect 9640 3680 9646 3692
rect 9769 3689 9781 3692
rect 9815 3689 9827 3723
rect 9769 3683 9827 3689
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 10045 3723 10103 3729
rect 10045 3720 10057 3723
rect 9916 3692 10057 3720
rect 9916 3680 9922 3692
rect 10045 3689 10057 3692
rect 10091 3689 10103 3723
rect 10045 3683 10103 3689
rect 10686 3680 10692 3732
rect 10744 3720 10750 3732
rect 10873 3723 10931 3729
rect 10873 3720 10885 3723
rect 10744 3692 10885 3720
rect 10744 3680 10750 3692
rect 10873 3689 10885 3692
rect 10919 3689 10931 3723
rect 10873 3683 10931 3689
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 13538 3720 13544 3732
rect 11020 3692 13544 3720
rect 11020 3680 11026 3692
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 13906 3720 13912 3732
rect 13867 3692 13912 3720
rect 13906 3680 13912 3692
rect 13964 3680 13970 3732
rect 14642 3680 14648 3732
rect 14700 3720 14706 3732
rect 14829 3723 14887 3729
rect 14829 3720 14841 3723
rect 14700 3692 14841 3720
rect 14700 3680 14706 3692
rect 14829 3689 14841 3692
rect 14875 3689 14887 3723
rect 14829 3683 14887 3689
rect 15378 3680 15384 3732
rect 15436 3720 15442 3732
rect 15565 3723 15623 3729
rect 15565 3720 15577 3723
rect 15436 3692 15577 3720
rect 15436 3680 15442 3692
rect 15565 3689 15577 3692
rect 15611 3689 15623 3723
rect 15565 3683 15623 3689
rect 15654 3680 15660 3732
rect 15712 3720 15718 3732
rect 15838 3720 15844 3732
rect 15712 3692 15757 3720
rect 15799 3692 15844 3720
rect 15712 3680 15718 3692
rect 15838 3680 15844 3692
rect 15896 3720 15902 3732
rect 16298 3720 16304 3732
rect 15896 3692 16304 3720
rect 15896 3680 15902 3692
rect 16298 3680 16304 3692
rect 16356 3680 16362 3732
rect 16853 3723 16911 3729
rect 16853 3689 16865 3723
rect 16899 3720 16911 3723
rect 17034 3720 17040 3732
rect 16899 3692 17040 3720
rect 16899 3689 16911 3692
rect 16853 3683 16911 3689
rect 17034 3680 17040 3692
rect 17092 3720 17098 3732
rect 17310 3720 17316 3732
rect 17092 3692 17316 3720
rect 17092 3680 17098 3692
rect 17310 3680 17316 3692
rect 17368 3680 17374 3732
rect 6638 3652 6644 3664
rect 5184 3624 6644 3652
rect 6638 3612 6644 3624
rect 6696 3612 6702 3664
rect 11793 3655 11851 3661
rect 9232 3624 10548 3652
rect 5077 3587 5135 3593
rect 5077 3584 5089 3587
rect 5000 3556 5089 3584
rect 5077 3553 5089 3556
rect 5123 3553 5135 3587
rect 5077 3547 5135 3553
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 5316 3556 5361 3584
rect 5316 3544 5322 3556
rect 7282 3544 7288 3596
rect 7340 3584 7346 3596
rect 8481 3587 8539 3593
rect 8481 3584 8493 3587
rect 7340 3556 8493 3584
rect 7340 3544 7346 3556
rect 8481 3553 8493 3556
rect 8527 3553 8539 3587
rect 8481 3547 8539 3553
rect 1489 3519 1547 3525
rect 1489 3485 1501 3519
rect 1535 3516 1547 3519
rect 2222 3516 2228 3528
rect 1535 3488 2228 3516
rect 1535 3485 1547 3488
rect 1489 3479 1547 3485
rect 2222 3476 2228 3488
rect 2280 3476 2286 3528
rect 2958 3516 2964 3528
rect 2919 3488 2964 3516
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3516 5043 3519
rect 5718 3516 5724 3528
rect 5031 3488 5724 3516
rect 5031 3485 5043 3488
rect 4985 3479 5043 3485
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3516 7895 3519
rect 9232 3516 9260 3624
rect 9398 3584 9404 3596
rect 9359 3556 9404 3584
rect 9398 3544 9404 3556
rect 9456 3544 9462 3596
rect 9585 3587 9643 3593
rect 9585 3553 9597 3587
rect 9631 3584 9643 3587
rect 10318 3584 10324 3596
rect 9631 3556 10324 3584
rect 9631 3553 9643 3556
rect 9585 3547 9643 3553
rect 10318 3544 10324 3556
rect 10376 3544 10382 3596
rect 7883 3488 9260 3516
rect 9309 3519 9367 3525
rect 7883 3485 7895 3488
rect 7837 3479 7895 3485
rect 9309 3485 9321 3519
rect 9355 3516 9367 3519
rect 9674 3516 9680 3528
rect 9355 3488 9680 3516
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9674 3476 9680 3488
rect 9732 3476 9738 3528
rect 10410 3516 10416 3528
rect 10371 3488 10416 3516
rect 10410 3476 10416 3488
rect 10468 3476 10474 3528
rect 10520 3525 10548 3624
rect 11793 3621 11805 3655
rect 11839 3652 11851 3655
rect 11882 3652 11888 3664
rect 11839 3624 11888 3652
rect 11839 3621 11851 3624
rect 11793 3615 11851 3621
rect 11882 3612 11888 3624
rect 11940 3612 11946 3664
rect 16206 3652 16212 3664
rect 14384 3624 16212 3652
rect 10689 3587 10747 3593
rect 10689 3553 10701 3587
rect 10735 3584 10747 3587
rect 10870 3584 10876 3596
rect 10735 3556 10876 3584
rect 10735 3553 10747 3556
rect 10689 3547 10747 3553
rect 10870 3544 10876 3556
rect 10928 3544 10934 3596
rect 11054 3544 11060 3596
rect 11112 3584 11118 3596
rect 11425 3587 11483 3593
rect 11425 3584 11437 3587
rect 11112 3556 11437 3584
rect 11112 3544 11118 3556
rect 11425 3553 11437 3556
rect 11471 3553 11483 3587
rect 11425 3547 11483 3553
rect 11514 3544 11520 3596
rect 11572 3584 11578 3596
rect 11572 3556 12204 3584
rect 11572 3544 11578 3556
rect 10505 3519 10563 3525
rect 10505 3485 10517 3519
rect 10551 3516 10563 3519
rect 11606 3516 11612 3528
rect 10551 3488 11612 3516
rect 10551 3485 10563 3488
rect 10505 3479 10563 3485
rect 11606 3476 11612 3488
rect 11664 3476 11670 3528
rect 11977 3519 12035 3525
rect 11977 3485 11989 3519
rect 12023 3516 12035 3519
rect 12066 3516 12072 3528
rect 12023 3488 12072 3516
rect 12023 3485 12035 3488
rect 11977 3479 12035 3485
rect 12066 3476 12072 3488
rect 12124 3476 12130 3528
rect 12176 3525 12204 3556
rect 13354 3544 13360 3596
rect 13412 3584 13418 3596
rect 14274 3584 14280 3596
rect 13412 3556 13768 3584
rect 14235 3556 14280 3584
rect 13412 3544 13418 3556
rect 13740 3528 13768 3556
rect 14274 3544 14280 3556
rect 14332 3544 14338 3596
rect 14384 3593 14412 3624
rect 16206 3612 16212 3624
rect 16264 3612 16270 3664
rect 17681 3655 17739 3661
rect 17681 3621 17693 3655
rect 17727 3652 17739 3655
rect 18138 3652 18144 3664
rect 17727 3624 18144 3652
rect 17727 3621 17739 3624
rect 17681 3615 17739 3621
rect 18138 3612 18144 3624
rect 18196 3612 18202 3664
rect 18414 3652 18420 3664
rect 18375 3624 18420 3652
rect 18414 3612 18420 3624
rect 18472 3612 18478 3664
rect 14369 3587 14427 3593
rect 14369 3553 14381 3587
rect 14415 3553 14427 3587
rect 16022 3584 16028 3596
rect 15983 3556 16028 3584
rect 14369 3547 14427 3553
rect 16022 3544 16028 3556
rect 16080 3544 16086 3596
rect 16942 3584 16948 3596
rect 16408 3556 16948 3584
rect 12161 3519 12219 3525
rect 12161 3485 12173 3519
rect 12207 3516 12219 3519
rect 13446 3516 13452 3528
rect 12207 3488 13452 3516
rect 12207 3485 12219 3488
rect 12161 3479 12219 3485
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 13722 3516 13728 3528
rect 13683 3488 13728 3516
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 13906 3476 13912 3528
rect 13964 3516 13970 3528
rect 14090 3516 14096 3528
rect 13964 3488 14096 3516
rect 13964 3476 13970 3488
rect 14090 3476 14096 3488
rect 14148 3516 14154 3528
rect 14921 3519 14979 3525
rect 14921 3516 14933 3519
rect 14148 3488 14933 3516
rect 14148 3476 14154 3488
rect 14921 3485 14933 3488
rect 14967 3485 14979 3519
rect 14921 3479 14979 3485
rect 1756 3451 1814 3457
rect 1756 3417 1768 3451
rect 1802 3448 1814 3451
rect 1854 3448 1860 3460
rect 1802 3420 1860 3448
rect 1802 3417 1814 3420
rect 1756 3411 1814 3417
rect 1854 3408 1860 3420
rect 1912 3408 1918 3460
rect 3694 3408 3700 3460
rect 3752 3448 3758 3460
rect 3752 3420 4292 3448
rect 3752 3408 3758 3420
rect 4154 3380 4160 3392
rect 4115 3352 4160 3380
rect 4154 3340 4160 3352
rect 4212 3340 4218 3392
rect 4264 3380 4292 3420
rect 4430 3408 4436 3460
rect 4488 3448 4494 3460
rect 5445 3451 5503 3457
rect 5445 3448 5457 3451
rect 4488 3420 5457 3448
rect 4488 3408 4494 3420
rect 5445 3417 5457 3420
rect 5491 3417 5503 3451
rect 7374 3448 7380 3460
rect 5445 3411 5503 3417
rect 6012 3420 7380 3448
rect 6012 3380 6040 3420
rect 7374 3408 7380 3420
rect 7432 3408 7438 3460
rect 7469 3451 7527 3457
rect 7469 3417 7481 3451
rect 7515 3448 7527 3451
rect 11054 3448 11060 3460
rect 7515 3420 11060 3448
rect 7515 3417 7527 3420
rect 7469 3411 7527 3417
rect 11054 3408 11060 3420
rect 11112 3408 11118 3460
rect 11241 3451 11299 3457
rect 11241 3417 11253 3451
rect 11287 3448 11299 3451
rect 11422 3448 11428 3460
rect 11287 3420 11428 3448
rect 11287 3417 11299 3420
rect 11241 3411 11299 3417
rect 11422 3408 11428 3420
rect 11480 3408 11486 3460
rect 11514 3408 11520 3460
rect 11572 3448 11578 3460
rect 11698 3448 11704 3460
rect 11572 3420 11704 3448
rect 11572 3408 11578 3420
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 12428 3451 12486 3457
rect 12428 3417 12440 3451
rect 12474 3448 12486 3451
rect 15470 3448 15476 3460
rect 12474 3420 15476 3448
rect 12474 3417 12486 3420
rect 12428 3411 12486 3417
rect 15470 3408 15476 3420
rect 15528 3408 15534 3460
rect 16408 3457 16436 3556
rect 16942 3544 16948 3556
rect 17000 3584 17006 3596
rect 17000 3556 17908 3584
rect 17000 3544 17006 3556
rect 17129 3519 17187 3525
rect 17129 3516 17141 3519
rect 16500 3488 17141 3516
rect 16393 3451 16451 3457
rect 16393 3448 16405 3451
rect 15580 3420 16405 3448
rect 6178 3380 6184 3392
rect 4264 3352 6040 3380
rect 6139 3352 6184 3380
rect 6178 3340 6184 3352
rect 6236 3340 6242 3392
rect 7190 3340 7196 3392
rect 7248 3380 7254 3392
rect 7653 3383 7711 3389
rect 7653 3380 7665 3383
rect 7248 3352 7665 3380
rect 7248 3340 7254 3352
rect 7653 3349 7665 3352
rect 7699 3349 7711 3383
rect 7653 3343 7711 3349
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 8297 3383 8355 3389
rect 8297 3380 8309 3383
rect 8076 3352 8309 3380
rect 8076 3340 8082 3352
rect 8297 3349 8309 3352
rect 8343 3349 8355 3383
rect 8297 3343 8355 3349
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 11330 3380 11336 3392
rect 8444 3352 8489 3380
rect 11291 3352 11336 3380
rect 8444 3340 8450 3352
rect 11330 3340 11336 3352
rect 11388 3340 11394 3392
rect 13541 3383 13599 3389
rect 13541 3349 13553 3383
rect 13587 3380 13599 3383
rect 13906 3380 13912 3392
rect 13587 3352 13912 3380
rect 13587 3349 13599 3352
rect 13541 3343 13599 3349
rect 13906 3340 13912 3352
rect 13964 3340 13970 3392
rect 13998 3340 14004 3392
rect 14056 3380 14062 3392
rect 14461 3383 14519 3389
rect 14461 3380 14473 3383
rect 14056 3352 14473 3380
rect 14056 3340 14062 3352
rect 14461 3349 14473 3352
rect 14507 3380 14519 3383
rect 15580 3380 15608 3420
rect 16393 3417 16405 3420
rect 16439 3417 16451 3451
rect 16393 3411 16451 3417
rect 14507 3352 15608 3380
rect 14507 3349 14519 3352
rect 14461 3343 14519 3349
rect 16206 3340 16212 3392
rect 16264 3380 16270 3392
rect 16500 3380 16528 3488
rect 17129 3485 17141 3488
rect 17175 3516 17187 3519
rect 17313 3519 17371 3525
rect 17313 3516 17325 3519
rect 17175 3488 17325 3516
rect 17175 3485 17187 3488
rect 17129 3479 17187 3485
rect 17313 3485 17325 3488
rect 17359 3485 17371 3519
rect 17494 3516 17500 3528
rect 17455 3488 17500 3516
rect 17313 3479 17371 3485
rect 17494 3476 17500 3488
rect 17552 3476 17558 3528
rect 17880 3525 17908 3556
rect 17865 3519 17923 3525
rect 17865 3485 17877 3519
rect 17911 3485 17923 3519
rect 18230 3516 18236 3528
rect 18191 3488 18236 3516
rect 17865 3479 17923 3485
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 16574 3408 16580 3460
rect 16632 3448 16638 3460
rect 16942 3448 16948 3460
rect 16632 3420 16677 3448
rect 16903 3420 16948 3448
rect 16632 3408 16638 3420
rect 16942 3408 16948 3420
rect 17000 3448 17006 3460
rect 19426 3448 19432 3460
rect 17000 3420 19432 3448
rect 17000 3408 17006 3420
rect 19426 3408 19432 3420
rect 19484 3408 19490 3460
rect 18046 3380 18052 3392
rect 16264 3352 16528 3380
rect 18007 3352 18052 3380
rect 16264 3340 16270 3352
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 1104 3290 18860 3312
rect 1104 3238 5398 3290
rect 5450 3238 5462 3290
rect 5514 3238 5526 3290
rect 5578 3238 5590 3290
rect 5642 3238 5654 3290
rect 5706 3238 9846 3290
rect 9898 3238 9910 3290
rect 9962 3238 9974 3290
rect 10026 3238 10038 3290
rect 10090 3238 10102 3290
rect 10154 3238 14294 3290
rect 14346 3238 14358 3290
rect 14410 3238 14422 3290
rect 14474 3238 14486 3290
rect 14538 3238 14550 3290
rect 14602 3238 18860 3290
rect 1104 3216 18860 3238
rect 1394 3136 1400 3188
rect 1452 3176 1458 3188
rect 1489 3179 1547 3185
rect 1489 3176 1501 3179
rect 1452 3148 1501 3176
rect 1452 3136 1458 3148
rect 1489 3145 1501 3148
rect 1535 3145 1547 3179
rect 1489 3139 1547 3145
rect 2130 3136 2136 3188
rect 2188 3176 2194 3188
rect 2958 3176 2964 3188
rect 2188 3148 2964 3176
rect 2188 3136 2194 3148
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 3053 3179 3111 3185
rect 3053 3145 3065 3179
rect 3099 3176 3111 3179
rect 3510 3176 3516 3188
rect 3099 3148 3516 3176
rect 3099 3145 3111 3148
rect 3053 3139 3111 3145
rect 3510 3136 3516 3148
rect 3568 3136 3574 3188
rect 4525 3179 4583 3185
rect 4525 3176 4537 3179
rect 3620 3148 4537 3176
rect 1872 3080 2774 3108
rect 1670 3040 1676 3052
rect 1631 3012 1676 3040
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 1872 2981 1900 3080
rect 2130 3040 2136 3052
rect 2091 3012 2136 3040
rect 2130 3000 2136 3012
rect 2188 3000 2194 3052
rect 2746 3040 2774 3080
rect 2866 3068 2872 3120
rect 2924 3108 2930 3120
rect 3620 3108 3648 3148
rect 4525 3145 4537 3148
rect 4571 3145 4583 3179
rect 4525 3139 4583 3145
rect 4614 3136 4620 3188
rect 4672 3176 4678 3188
rect 5074 3176 5080 3188
rect 4672 3148 5080 3176
rect 4672 3136 4678 3148
rect 5074 3136 5080 3148
rect 5132 3136 5138 3188
rect 5902 3136 5908 3188
rect 5960 3176 5966 3188
rect 7009 3179 7067 3185
rect 7009 3176 7021 3179
rect 5960 3148 7021 3176
rect 5960 3136 5966 3148
rect 7009 3145 7021 3148
rect 7055 3145 7067 3179
rect 7009 3139 7067 3145
rect 7374 3136 7380 3188
rect 7432 3176 7438 3188
rect 10137 3179 10195 3185
rect 7432 3148 7972 3176
rect 7432 3136 7438 3148
rect 2924 3080 3648 3108
rect 4341 3111 4399 3117
rect 2924 3068 2930 3080
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 6178 3108 6184 3120
rect 4387 3080 6184 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 6178 3068 6184 3080
rect 6236 3108 6242 3120
rect 7837 3111 7895 3117
rect 7837 3108 7849 3111
rect 6236 3080 7849 3108
rect 6236 3068 6242 3080
rect 7837 3077 7849 3080
rect 7883 3077 7895 3111
rect 7837 3071 7895 3077
rect 4614 3040 4620 3052
rect 2746 3012 4620 3040
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3009 4767 3043
rect 4709 3003 4767 3009
rect 1857 2975 1915 2981
rect 1857 2941 1869 2975
rect 1903 2941 1915 2975
rect 1857 2935 1915 2941
rect 2041 2975 2099 2981
rect 2041 2941 2053 2975
rect 2087 2972 2099 2975
rect 3786 2972 3792 2984
rect 2087 2944 3792 2972
rect 2087 2941 2099 2944
rect 2041 2935 2099 2941
rect 3786 2932 3792 2944
rect 3844 2932 3850 2984
rect 4614 2904 4620 2916
rect 2746 2876 4620 2904
rect 2501 2839 2559 2845
rect 2501 2805 2513 2839
rect 2547 2836 2559 2839
rect 2746 2836 2774 2876
rect 4614 2864 4620 2876
rect 4672 2864 4678 2916
rect 2547 2808 2774 2836
rect 2547 2805 2559 2808
rect 2501 2799 2559 2805
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 4430 2836 4436 2848
rect 3568 2808 4436 2836
rect 3568 2796 3574 2808
rect 4430 2796 4436 2808
rect 4488 2796 4494 2848
rect 4724 2836 4752 3003
rect 4798 3000 4804 3052
rect 4856 3040 4862 3052
rect 5074 3049 5080 3052
rect 5068 3040 5080 3049
rect 4856 3012 4901 3040
rect 5035 3012 5080 3040
rect 4856 3000 4862 3012
rect 5068 3003 5080 3012
rect 5074 3000 5080 3003
rect 5132 3000 5138 3052
rect 5534 3000 5540 3052
rect 5592 3040 5598 3052
rect 6454 3040 6460 3052
rect 5592 3012 6460 3040
rect 5592 3000 5598 3012
rect 6454 3000 6460 3012
rect 6512 3000 6518 3052
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3040 6975 3043
rect 7098 3040 7104 3052
rect 6963 3012 7104 3040
rect 6963 3009 6975 3012
rect 6917 3003 6975 3009
rect 7098 3000 7104 3012
rect 7156 3000 7162 3052
rect 7374 3040 7380 3052
rect 7335 3012 7380 3040
rect 7374 3000 7380 3012
rect 7432 3000 7438 3052
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3040 7527 3043
rect 7650 3040 7656 3052
rect 7515 3012 7656 3040
rect 7515 3009 7527 3012
rect 7469 3003 7527 3009
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 6733 2975 6791 2981
rect 6733 2941 6745 2975
rect 6779 2941 6791 2975
rect 6733 2935 6791 2941
rect 6748 2904 6776 2935
rect 7558 2932 7564 2984
rect 7616 2972 7622 2984
rect 7944 2972 7972 3148
rect 10137 3145 10149 3179
rect 10183 3176 10195 3179
rect 10502 3176 10508 3188
rect 10183 3148 10508 3176
rect 10183 3145 10195 3148
rect 10137 3139 10195 3145
rect 10502 3136 10508 3148
rect 10560 3136 10566 3188
rect 10594 3136 10600 3188
rect 10652 3176 10658 3188
rect 10873 3179 10931 3185
rect 10873 3176 10885 3179
rect 10652 3148 10885 3176
rect 10652 3136 10658 3148
rect 10873 3145 10885 3148
rect 10919 3145 10931 3179
rect 10873 3139 10931 3145
rect 11241 3179 11299 3185
rect 11241 3145 11253 3179
rect 11287 3176 11299 3179
rect 11977 3179 12035 3185
rect 11977 3176 11989 3179
rect 11287 3148 11989 3176
rect 11287 3145 11299 3148
rect 11241 3139 11299 3145
rect 11977 3145 11989 3148
rect 12023 3145 12035 3179
rect 11977 3139 12035 3145
rect 12066 3136 12072 3188
rect 12124 3176 12130 3188
rect 13446 3176 13452 3188
rect 12124 3148 13308 3176
rect 13407 3148 13452 3176
rect 12124 3136 12130 3148
rect 10318 3068 10324 3120
rect 10376 3108 10382 3120
rect 12621 3111 12679 3117
rect 12621 3108 12633 3111
rect 10376 3080 12633 3108
rect 10376 3068 10382 3080
rect 12621 3077 12633 3080
rect 12667 3077 12679 3111
rect 12621 3071 12679 3077
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 9732 3012 10057 3040
rect 9732 3000 9738 3012
rect 10045 3009 10057 3012
rect 10091 3040 10103 3043
rect 10410 3040 10416 3052
rect 10091 3012 10416 3040
rect 10091 3009 10103 3012
rect 10045 3003 10103 3009
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 10781 3043 10839 3049
rect 10781 3009 10793 3043
rect 10827 3040 10839 3043
rect 10962 3040 10968 3052
rect 10827 3012 10968 3040
rect 10827 3009 10839 3012
rect 10781 3003 10839 3009
rect 10962 3000 10968 3012
rect 11020 3000 11026 3052
rect 11514 3040 11520 3052
rect 11164 3012 11520 3040
rect 10229 2975 10287 2981
rect 7616 2944 7661 2972
rect 7944 2944 10088 2972
rect 7616 2932 7622 2944
rect 8478 2904 8484 2916
rect 6748 2876 8484 2904
rect 8478 2864 8484 2876
rect 8536 2864 8542 2916
rect 10060 2904 10088 2944
rect 10229 2941 10241 2975
rect 10275 2972 10287 2975
rect 10597 2975 10655 2981
rect 10597 2972 10609 2975
rect 10275 2944 10609 2972
rect 10275 2941 10287 2944
rect 10229 2935 10287 2941
rect 10597 2941 10609 2944
rect 10643 2941 10655 2975
rect 10597 2935 10655 2941
rect 10244 2904 10272 2935
rect 10060 2876 10272 2904
rect 10612 2904 10640 2935
rect 11164 2904 11192 3012
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 11882 3040 11888 3052
rect 11843 3012 11888 3040
rect 11882 3000 11888 3012
rect 11940 3000 11946 3052
rect 12342 3040 12348 3052
rect 12303 3012 12348 3040
rect 12342 3000 12348 3012
rect 12400 3000 12406 3052
rect 13280 3040 13308 3148
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 13906 3136 13912 3188
rect 13964 3176 13970 3188
rect 13964 3148 16252 3176
rect 13964 3136 13970 3148
rect 13998 3068 14004 3120
rect 14056 3108 14062 3120
rect 14182 3108 14188 3120
rect 14056 3080 14188 3108
rect 14056 3068 14062 3080
rect 14182 3068 14188 3080
rect 14240 3068 14246 3120
rect 15654 3108 15660 3120
rect 14292 3080 15660 3108
rect 14292 3040 14320 3080
rect 15654 3068 15660 3080
rect 15712 3108 15718 3120
rect 16114 3108 16120 3120
rect 15712 3080 16120 3108
rect 15712 3068 15718 3080
rect 16114 3068 16120 3080
rect 16172 3068 16178 3120
rect 16224 3117 16252 3148
rect 16209 3111 16267 3117
rect 16209 3077 16221 3111
rect 16255 3077 16267 3111
rect 16209 3071 16267 3077
rect 16298 3068 16304 3120
rect 16356 3108 16362 3120
rect 16356 3080 17908 3108
rect 16356 3068 16362 3080
rect 13280 3012 14320 3040
rect 14737 3043 14795 3049
rect 14737 3009 14749 3043
rect 14783 3009 14795 3043
rect 14737 3003 14795 3009
rect 11330 2932 11336 2984
rect 11388 2972 11394 2984
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 11388 2944 12081 2972
rect 11388 2932 11394 2944
rect 12069 2941 12081 2944
rect 12115 2941 12127 2975
rect 12069 2935 12127 2941
rect 14752 2916 14780 3003
rect 14826 3000 14832 3052
rect 14884 3040 14890 3052
rect 14884 3012 14929 3040
rect 14884 3000 14890 3012
rect 15286 3000 15292 3052
rect 15344 3040 15350 3052
rect 15381 3043 15439 3049
rect 15381 3040 15393 3043
rect 15344 3012 15393 3040
rect 15344 3000 15350 3012
rect 15381 3009 15393 3012
rect 15427 3009 15439 3043
rect 15381 3003 15439 3009
rect 15746 3000 15752 3052
rect 15804 3040 15810 3052
rect 15933 3043 15991 3049
rect 15933 3040 15945 3043
rect 15804 3012 15945 3040
rect 15804 3000 15810 3012
rect 15933 3009 15945 3012
rect 15979 3009 15991 3043
rect 15933 3003 15991 3009
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3040 17003 3043
rect 17034 3040 17040 3052
rect 16991 3012 17040 3040
rect 16991 3009 17003 3012
rect 16945 3003 17003 3009
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 17129 3043 17187 3049
rect 17129 3009 17141 3043
rect 17175 3009 17187 3043
rect 17129 3003 17187 3009
rect 15105 2975 15163 2981
rect 15105 2941 15117 2975
rect 15151 2972 15163 2975
rect 15194 2972 15200 2984
rect 15151 2944 15200 2972
rect 15151 2941 15163 2944
rect 15105 2935 15163 2941
rect 15194 2932 15200 2944
rect 15252 2932 15258 2984
rect 15565 2975 15623 2981
rect 15565 2941 15577 2975
rect 15611 2941 15623 2975
rect 15565 2935 15623 2941
rect 10612 2876 11192 2904
rect 14734 2864 14740 2916
rect 14792 2864 14798 2916
rect 14826 2864 14832 2916
rect 14884 2904 14890 2916
rect 15580 2904 15608 2935
rect 16022 2932 16028 2984
rect 16080 2972 16086 2984
rect 17144 2972 17172 3003
rect 17310 3000 17316 3052
rect 17368 3040 17374 3052
rect 17880 3049 17908 3080
rect 17497 3043 17555 3049
rect 17497 3040 17509 3043
rect 17368 3012 17509 3040
rect 17368 3000 17374 3012
rect 17497 3009 17509 3012
rect 17543 3009 17555 3043
rect 17497 3003 17555 3009
rect 17865 3043 17923 3049
rect 17865 3009 17877 3043
rect 17911 3009 17923 3043
rect 17865 3003 17923 3009
rect 18233 3043 18291 3049
rect 18233 3009 18245 3043
rect 18279 3040 18291 3043
rect 18322 3040 18328 3052
rect 18279 3012 18328 3040
rect 18279 3009 18291 3012
rect 18233 3003 18291 3009
rect 18322 3000 18328 3012
rect 18380 3000 18386 3052
rect 16080 2944 17172 2972
rect 16080 2932 16086 2944
rect 16298 2904 16304 2916
rect 14884 2876 15608 2904
rect 15672 2876 16304 2904
rect 14884 2864 14890 2876
rect 5534 2836 5540 2848
rect 4724 2808 5540 2836
rect 5534 2796 5540 2808
rect 5592 2796 5598 2848
rect 6178 2836 6184 2848
rect 6139 2808 6184 2836
rect 6178 2796 6184 2808
rect 6236 2796 6242 2848
rect 6362 2796 6368 2848
rect 6420 2836 6426 2848
rect 6914 2836 6920 2848
rect 6420 2808 6920 2836
rect 6420 2796 6426 2808
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7098 2796 7104 2848
rect 7156 2836 7162 2848
rect 7282 2836 7288 2848
rect 7156 2808 7288 2836
rect 7156 2796 7162 2808
rect 7282 2796 7288 2808
rect 7340 2796 7346 2848
rect 8754 2796 8760 2848
rect 8812 2836 8818 2848
rect 9125 2839 9183 2845
rect 9125 2836 9137 2839
rect 8812 2808 9137 2836
rect 8812 2796 8818 2808
rect 9125 2805 9137 2808
rect 9171 2805 9183 2839
rect 9125 2799 9183 2805
rect 9214 2796 9220 2848
rect 9272 2836 9278 2848
rect 9677 2839 9735 2845
rect 9677 2836 9689 2839
rect 9272 2808 9689 2836
rect 9272 2796 9278 2808
rect 9677 2805 9689 2808
rect 9723 2805 9735 2839
rect 9677 2799 9735 2805
rect 11054 2796 11060 2848
rect 11112 2836 11118 2848
rect 11517 2839 11575 2845
rect 11517 2836 11529 2839
rect 11112 2808 11529 2836
rect 11112 2796 11118 2808
rect 11517 2805 11529 2808
rect 11563 2805 11575 2839
rect 11517 2799 11575 2805
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 13722 2836 13728 2848
rect 12492 2808 13728 2836
rect 12492 2796 12498 2808
rect 13722 2796 13728 2808
rect 13780 2836 13786 2848
rect 15672 2836 15700 2876
rect 16298 2864 16304 2876
rect 16356 2904 16362 2916
rect 16574 2904 16580 2916
rect 16356 2876 16580 2904
rect 16356 2864 16362 2876
rect 16574 2864 16580 2876
rect 16632 2864 16638 2916
rect 16758 2904 16764 2916
rect 16719 2876 16764 2904
rect 16758 2864 16764 2876
rect 16816 2864 16822 2916
rect 18690 2904 18696 2916
rect 16868 2876 18696 2904
rect 13780 2808 15700 2836
rect 13780 2796 13786 2808
rect 15746 2796 15752 2848
rect 15804 2836 15810 2848
rect 16868 2836 16896 2876
rect 18690 2864 18696 2876
rect 18748 2864 18754 2916
rect 17310 2836 17316 2848
rect 15804 2808 16896 2836
rect 17271 2808 17316 2836
rect 15804 2796 15810 2808
rect 17310 2796 17316 2808
rect 17368 2796 17374 2848
rect 17678 2836 17684 2848
rect 17639 2808 17684 2836
rect 17678 2796 17684 2808
rect 17736 2796 17742 2848
rect 18046 2836 18052 2848
rect 18007 2808 18052 2836
rect 18046 2796 18052 2808
rect 18104 2796 18110 2848
rect 18417 2839 18475 2845
rect 18417 2805 18429 2839
rect 18463 2836 18475 2839
rect 18874 2836 18880 2848
rect 18463 2808 18880 2836
rect 18463 2805 18475 2808
rect 18417 2799 18475 2805
rect 18874 2796 18880 2808
rect 18932 2796 18938 2848
rect 1104 2746 18860 2768
rect 1104 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 3430 2746
rect 3482 2694 7622 2746
rect 7674 2694 7686 2746
rect 7738 2694 7750 2746
rect 7802 2694 7814 2746
rect 7866 2694 7878 2746
rect 7930 2694 12070 2746
rect 12122 2694 12134 2746
rect 12186 2694 12198 2746
rect 12250 2694 12262 2746
rect 12314 2694 12326 2746
rect 12378 2694 16518 2746
rect 16570 2694 16582 2746
rect 16634 2694 16646 2746
rect 16698 2694 16710 2746
rect 16762 2694 16774 2746
rect 16826 2694 18860 2746
rect 1104 2672 18860 2694
rect 2130 2592 2136 2644
rect 2188 2632 2194 2644
rect 2869 2635 2927 2641
rect 2869 2632 2881 2635
rect 2188 2604 2881 2632
rect 2188 2592 2194 2604
rect 2869 2601 2881 2604
rect 2915 2601 2927 2635
rect 2869 2595 2927 2601
rect 3786 2592 3792 2644
rect 3844 2632 3850 2644
rect 4982 2632 4988 2644
rect 3844 2604 4988 2632
rect 3844 2592 3850 2604
rect 4982 2592 4988 2604
rect 5040 2592 5046 2644
rect 5077 2635 5135 2641
rect 5077 2601 5089 2635
rect 5123 2632 5135 2635
rect 6181 2635 6239 2641
rect 6181 2632 6193 2635
rect 5123 2604 6193 2632
rect 5123 2601 5135 2604
rect 5077 2595 5135 2601
rect 6181 2601 6193 2604
rect 6227 2632 6239 2635
rect 6270 2632 6276 2644
rect 6227 2604 6276 2632
rect 6227 2601 6239 2604
rect 6181 2595 6239 2601
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 9048 2604 9996 2632
rect 2148 2536 3924 2564
rect 2148 2505 2176 2536
rect 3896 2508 3924 2536
rect 4890 2524 4896 2576
rect 4948 2564 4954 2576
rect 6549 2567 6607 2573
rect 6549 2564 6561 2567
rect 4948 2536 6561 2564
rect 4948 2524 4954 2536
rect 6549 2533 6561 2536
rect 6595 2533 6607 2567
rect 9048 2564 9076 2604
rect 6549 2527 6607 2533
rect 6647 2536 9076 2564
rect 2133 2499 2191 2505
rect 2133 2465 2145 2499
rect 2179 2465 2191 2499
rect 2314 2496 2320 2508
rect 2275 2468 2320 2496
rect 2133 2459 2191 2465
rect 2314 2456 2320 2468
rect 2372 2456 2378 2508
rect 2958 2456 2964 2508
rect 3016 2496 3022 2508
rect 3329 2499 3387 2505
rect 3329 2496 3341 2499
rect 3016 2468 3341 2496
rect 3016 2456 3022 2468
rect 3329 2465 3341 2468
rect 3375 2465 3387 2499
rect 3329 2459 3387 2465
rect 3513 2499 3571 2505
rect 3513 2465 3525 2499
rect 3559 2465 3571 2499
rect 3513 2459 3571 2465
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2428 2007 2431
rect 2222 2428 2228 2440
rect 1995 2400 2228 2428
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 2222 2388 2228 2400
rect 2280 2388 2286 2440
rect 2406 2428 2412 2440
rect 2367 2400 2412 2428
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 3528 2428 3556 2459
rect 3878 2456 3884 2508
rect 3936 2496 3942 2508
rect 4157 2499 4215 2505
rect 4157 2496 4169 2499
rect 3936 2468 4169 2496
rect 3936 2456 3942 2468
rect 4157 2465 4169 2468
rect 4203 2465 4215 2499
rect 4157 2459 4215 2465
rect 4338 2456 4344 2508
rect 4396 2496 4402 2508
rect 5813 2499 5871 2505
rect 5813 2496 5825 2499
rect 4396 2468 4441 2496
rect 4816 2468 5825 2496
rect 4396 2456 4402 2468
rect 4246 2428 4252 2440
rect 3528 2400 4252 2428
rect 4246 2388 4252 2400
rect 4304 2428 4310 2440
rect 4816 2428 4844 2468
rect 5813 2465 5825 2468
rect 5859 2496 5871 2499
rect 6647 2496 6675 2536
rect 7098 2496 7104 2508
rect 5859 2468 6675 2496
rect 7059 2468 7104 2496
rect 5859 2465 5871 2468
rect 5813 2459 5871 2465
rect 7098 2456 7104 2468
rect 7156 2496 7162 2508
rect 7466 2496 7472 2508
rect 7156 2468 7472 2496
rect 7156 2456 7162 2468
rect 7466 2456 7472 2468
rect 7524 2456 7530 2508
rect 8205 2499 8263 2505
rect 8205 2465 8217 2499
rect 8251 2496 8263 2499
rect 8294 2496 8300 2508
rect 8251 2468 8300 2496
rect 8251 2465 8263 2468
rect 8205 2459 8263 2465
rect 8294 2456 8300 2468
rect 8352 2456 8358 2508
rect 9048 2505 9076 2536
rect 9677 2567 9735 2573
rect 9677 2533 9689 2567
rect 9723 2564 9735 2567
rect 9968 2564 9996 2604
rect 10226 2592 10232 2644
rect 10284 2632 10290 2644
rect 10597 2635 10655 2641
rect 10597 2632 10609 2635
rect 10284 2604 10609 2632
rect 10284 2592 10290 2604
rect 10597 2601 10609 2604
rect 10643 2601 10655 2635
rect 11330 2632 11336 2644
rect 10597 2595 10655 2601
rect 10704 2604 11336 2632
rect 10704 2564 10732 2604
rect 11330 2592 11336 2604
rect 11388 2592 11394 2644
rect 11517 2635 11575 2641
rect 11517 2601 11529 2635
rect 11563 2632 11575 2635
rect 11882 2632 11888 2644
rect 11563 2604 11888 2632
rect 11563 2601 11575 2604
rect 11517 2595 11575 2601
rect 11882 2592 11888 2604
rect 11940 2592 11946 2644
rect 11974 2592 11980 2644
rect 12032 2632 12038 2644
rect 13909 2635 13967 2641
rect 12032 2604 13124 2632
rect 12032 2592 12038 2604
rect 12986 2564 12992 2576
rect 9723 2536 9904 2564
rect 9968 2536 10732 2564
rect 11164 2536 12434 2564
rect 12947 2536 12992 2564
rect 9723 2533 9735 2536
rect 9677 2527 9735 2533
rect 9033 2499 9091 2505
rect 8404 2468 8892 2496
rect 4304 2400 4844 2428
rect 5537 2431 5595 2437
rect 4304 2388 4310 2400
rect 5537 2397 5549 2431
rect 5583 2428 5595 2431
rect 5718 2428 5724 2440
rect 5583 2400 5724 2428
rect 5583 2397 5595 2400
rect 5537 2391 5595 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 6457 2431 6515 2437
rect 6457 2397 6469 2431
rect 6503 2428 6515 2431
rect 6914 2428 6920 2440
rect 6503 2400 6776 2428
rect 6875 2400 6920 2428
rect 6503 2397 6515 2400
rect 6457 2391 6515 2397
rect 1673 2363 1731 2369
rect 1673 2329 1685 2363
rect 1719 2360 1731 2363
rect 3973 2363 4031 2369
rect 1719 2332 3924 2360
rect 1719 2329 1731 2332
rect 1673 2323 1731 2329
rect 2777 2295 2835 2301
rect 2777 2261 2789 2295
rect 2823 2292 2835 2295
rect 2866 2292 2872 2304
rect 2823 2264 2872 2292
rect 2823 2261 2835 2264
rect 2777 2255 2835 2261
rect 2866 2252 2872 2264
rect 2924 2252 2930 2304
rect 3237 2295 3295 2301
rect 3237 2261 3249 2295
rect 3283 2292 3295 2295
rect 3510 2292 3516 2304
rect 3283 2264 3516 2292
rect 3283 2261 3295 2264
rect 3237 2255 3295 2261
rect 3510 2252 3516 2264
rect 3568 2252 3574 2304
rect 3896 2292 3924 2332
rect 3973 2329 3985 2363
rect 4019 2360 4031 2363
rect 4433 2363 4491 2369
rect 4433 2360 4445 2363
rect 4019 2332 4445 2360
rect 4019 2329 4031 2332
rect 3973 2323 4031 2329
rect 4433 2329 4445 2332
rect 4479 2329 4491 2363
rect 6748 2360 6776 2400
rect 6914 2388 6920 2400
rect 6972 2388 6978 2440
rect 7653 2431 7711 2437
rect 7653 2428 7665 2431
rect 7024 2400 7665 2428
rect 7024 2360 7052 2400
rect 7653 2397 7665 2400
rect 7699 2428 7711 2431
rect 8404 2428 8432 2468
rect 8754 2428 8760 2440
rect 7699 2400 8432 2428
rect 8715 2400 8760 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 8864 2428 8892 2468
rect 9033 2465 9045 2499
rect 9079 2465 9091 2499
rect 9214 2496 9220 2508
rect 9175 2468 9220 2496
rect 9033 2459 9091 2465
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 9674 2428 9680 2440
rect 8864 2400 9680 2428
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 6748 2332 7052 2360
rect 9876 2360 9904 2536
rect 11164 2508 11192 2536
rect 9950 2456 9956 2508
rect 10008 2496 10014 2508
rect 11054 2496 11060 2508
rect 10008 2468 10053 2496
rect 10336 2468 11060 2496
rect 10008 2456 10014 2468
rect 10045 2431 10103 2437
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10336 2428 10364 2468
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 11146 2456 11152 2508
rect 11204 2496 11210 2508
rect 11204 2468 11249 2496
rect 11204 2456 11210 2468
rect 11514 2456 11520 2508
rect 11572 2496 11578 2508
rect 12069 2499 12127 2505
rect 12069 2496 12081 2499
rect 11572 2468 12081 2496
rect 11572 2456 11578 2468
rect 12069 2465 12081 2468
rect 12115 2465 12127 2499
rect 12406 2496 12434 2536
rect 12986 2524 12992 2536
rect 13044 2524 13050 2576
rect 13096 2564 13124 2604
rect 13909 2601 13921 2635
rect 13955 2632 13967 2635
rect 13998 2632 14004 2644
rect 13955 2604 14004 2632
rect 13955 2601 13967 2604
rect 13909 2595 13967 2601
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 14734 2592 14740 2644
rect 14792 2632 14798 2644
rect 16209 2635 16267 2641
rect 16209 2632 16221 2635
rect 14792 2604 16221 2632
rect 14792 2592 14798 2604
rect 16209 2601 16221 2604
rect 16255 2601 16267 2635
rect 16209 2595 16267 2601
rect 16298 2592 16304 2644
rect 16356 2632 16362 2644
rect 16393 2635 16451 2641
rect 16393 2632 16405 2635
rect 16356 2604 16405 2632
rect 16356 2592 16362 2604
rect 16393 2601 16405 2604
rect 16439 2601 16451 2635
rect 16393 2595 16451 2601
rect 16945 2635 17003 2641
rect 16945 2601 16957 2635
rect 16991 2632 17003 2635
rect 17218 2632 17224 2644
rect 16991 2604 17224 2632
rect 16991 2601 17003 2604
rect 16945 2595 17003 2601
rect 17218 2592 17224 2604
rect 17276 2592 17282 2644
rect 14918 2564 14924 2576
rect 13096 2536 14924 2564
rect 14918 2524 14924 2536
rect 14976 2524 14982 2576
rect 15010 2524 15016 2576
rect 15068 2564 15074 2576
rect 15068 2536 15240 2564
rect 15068 2524 15074 2536
rect 12406 2468 13124 2496
rect 12069 2459 12127 2465
rect 11422 2428 11428 2440
rect 10091 2400 10364 2428
rect 10428 2400 11428 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 10137 2363 10195 2369
rect 10137 2360 10149 2363
rect 9876 2332 10149 2360
rect 4433 2323 4491 2329
rect 10137 2329 10149 2332
rect 10183 2329 10195 2363
rect 10137 2323 10195 2329
rect 4706 2292 4712 2304
rect 3896 2264 4712 2292
rect 4706 2252 4712 2264
rect 4764 2252 4770 2304
rect 4798 2252 4804 2304
rect 4856 2292 4862 2304
rect 4856 2264 4901 2292
rect 4856 2252 4862 2264
rect 4982 2252 4988 2304
rect 5040 2292 5046 2304
rect 5169 2295 5227 2301
rect 5169 2292 5181 2295
rect 5040 2264 5181 2292
rect 5040 2252 5046 2264
rect 5169 2261 5181 2264
rect 5215 2261 5227 2295
rect 5169 2255 5227 2261
rect 5629 2295 5687 2301
rect 5629 2261 5641 2295
rect 5675 2292 5687 2295
rect 5902 2292 5908 2304
rect 5675 2264 5908 2292
rect 5675 2261 5687 2264
rect 5629 2255 5687 2261
rect 5902 2252 5908 2264
rect 5960 2252 5966 2304
rect 6914 2252 6920 2304
rect 6972 2292 6978 2304
rect 7009 2295 7067 2301
rect 7009 2292 7021 2295
rect 6972 2264 7021 2292
rect 6972 2252 6978 2264
rect 7009 2261 7021 2264
rect 7055 2261 7067 2295
rect 7466 2292 7472 2304
rect 7427 2264 7472 2292
rect 7009 2255 7067 2261
rect 7466 2252 7472 2264
rect 7524 2252 7530 2304
rect 9309 2295 9367 2301
rect 9309 2261 9321 2295
rect 9355 2292 9367 2295
rect 10428 2292 10456 2400
rect 11422 2388 11428 2400
rect 11480 2388 11486 2440
rect 12342 2428 12348 2440
rect 12303 2400 12348 2428
rect 12342 2388 12348 2400
rect 12400 2388 12406 2440
rect 13096 2437 13124 2468
rect 14090 2456 14096 2508
rect 14148 2496 14154 2508
rect 15212 2505 15240 2536
rect 16666 2524 16672 2576
rect 16724 2564 16730 2576
rect 18230 2564 18236 2576
rect 16724 2536 18236 2564
rect 16724 2524 16730 2536
rect 18230 2524 18236 2536
rect 18288 2524 18294 2576
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 14148 2468 14197 2496
rect 14148 2456 14154 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 15197 2499 15255 2505
rect 14185 2459 14243 2465
rect 14292 2468 15148 2496
rect 13081 2431 13139 2437
rect 13081 2397 13093 2431
rect 13127 2397 13139 2431
rect 14292 2428 14320 2468
rect 15120 2440 15148 2468
rect 15197 2465 15209 2499
rect 15243 2465 15255 2499
rect 16025 2499 16083 2505
rect 16025 2496 16037 2499
rect 15197 2459 15255 2465
rect 15304 2468 16037 2496
rect 13081 2391 13139 2397
rect 14016 2400 14320 2428
rect 14369 2431 14427 2437
rect 11057 2363 11115 2369
rect 11057 2360 11069 2363
rect 10520 2332 11069 2360
rect 10520 2301 10548 2332
rect 11057 2329 11069 2332
rect 11103 2329 11115 2363
rect 11057 2323 11115 2329
rect 11977 2363 12035 2369
rect 11977 2329 11989 2363
rect 12023 2360 12035 2363
rect 14016 2360 14044 2400
rect 14369 2397 14381 2431
rect 14415 2428 14427 2431
rect 14642 2428 14648 2440
rect 14415 2400 14648 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 14642 2388 14648 2400
rect 14700 2388 14706 2440
rect 14918 2388 14924 2440
rect 14976 2428 14982 2440
rect 14976 2400 15021 2428
rect 14976 2388 14982 2400
rect 15102 2388 15108 2440
rect 15160 2428 15166 2440
rect 15304 2428 15332 2468
rect 16025 2465 16037 2468
rect 16071 2465 16083 2499
rect 16025 2459 16083 2465
rect 15470 2428 15476 2440
rect 15160 2400 15332 2428
rect 15431 2400 15476 2428
rect 15160 2388 15166 2400
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 16040 2428 16068 2459
rect 17681 2431 17739 2437
rect 17681 2428 17693 2431
rect 16040 2400 17693 2428
rect 17681 2397 17693 2400
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 17954 2388 17960 2440
rect 18012 2428 18018 2440
rect 18049 2431 18107 2437
rect 18049 2428 18061 2431
rect 18012 2400 18061 2428
rect 18012 2388 18018 2400
rect 18049 2397 18061 2400
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 12023 2332 14044 2360
rect 12023 2329 12035 2332
rect 11977 2323 12035 2329
rect 14090 2320 14096 2372
rect 14148 2360 14154 2372
rect 15749 2363 15807 2369
rect 15749 2360 15761 2363
rect 14148 2332 15761 2360
rect 14148 2320 14154 2332
rect 15749 2329 15761 2332
rect 15795 2329 15807 2363
rect 17405 2363 17463 2369
rect 17405 2360 17417 2363
rect 15749 2323 15807 2329
rect 16132 2332 17417 2360
rect 16132 2304 16160 2332
rect 17405 2329 17417 2332
rect 17451 2360 17463 2363
rect 18417 2363 18475 2369
rect 18417 2360 18429 2363
rect 17451 2332 18429 2360
rect 17451 2329 17463 2332
rect 17405 2323 17463 2329
rect 18417 2329 18429 2332
rect 18463 2329 18475 2363
rect 18417 2323 18475 2329
rect 9355 2264 10456 2292
rect 10505 2295 10563 2301
rect 9355 2261 9367 2264
rect 9309 2255 9367 2261
rect 10505 2261 10517 2295
rect 10551 2261 10563 2295
rect 10962 2292 10968 2304
rect 10923 2264 10968 2292
rect 10505 2255 10563 2261
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11885 2295 11943 2301
rect 11885 2292 11897 2295
rect 11664 2264 11897 2292
rect 11664 2252 11670 2264
rect 11885 2261 11897 2264
rect 11931 2292 11943 2295
rect 12434 2292 12440 2304
rect 11931 2264 12440 2292
rect 11931 2261 11943 2264
rect 11885 2255 11943 2261
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 13722 2292 13728 2304
rect 13683 2264 13728 2292
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 14461 2295 14519 2301
rect 14461 2261 14473 2295
rect 14507 2292 14519 2295
rect 14734 2292 14740 2304
rect 14507 2264 14740 2292
rect 14507 2261 14519 2264
rect 14461 2255 14519 2261
rect 14734 2252 14740 2264
rect 14792 2252 14798 2304
rect 14829 2295 14887 2301
rect 14829 2261 14841 2295
rect 14875 2292 14887 2295
rect 15562 2292 15568 2304
rect 14875 2264 15568 2292
rect 14875 2261 14887 2264
rect 14829 2255 14887 2261
rect 15562 2252 15568 2264
rect 15620 2252 15626 2304
rect 16114 2252 16120 2304
rect 16172 2252 16178 2304
rect 16666 2292 16672 2304
rect 16627 2264 16672 2292
rect 16666 2252 16672 2264
rect 16724 2252 16730 2304
rect 17034 2292 17040 2304
rect 16995 2264 17040 2292
rect 17034 2252 17040 2264
rect 17092 2252 17098 2304
rect 17218 2292 17224 2304
rect 17179 2264 17224 2292
rect 17218 2252 17224 2264
rect 17276 2252 17282 2304
rect 17862 2292 17868 2304
rect 17823 2264 17868 2292
rect 17862 2252 17868 2264
rect 17920 2252 17926 2304
rect 18230 2292 18236 2304
rect 18191 2264 18236 2292
rect 18230 2252 18236 2264
rect 18288 2252 18294 2304
rect 1104 2202 18860 2224
rect 1104 2150 5398 2202
rect 5450 2150 5462 2202
rect 5514 2150 5526 2202
rect 5578 2150 5590 2202
rect 5642 2150 5654 2202
rect 5706 2150 9846 2202
rect 9898 2150 9910 2202
rect 9962 2150 9974 2202
rect 10026 2150 10038 2202
rect 10090 2150 10102 2202
rect 10154 2150 14294 2202
rect 14346 2150 14358 2202
rect 14410 2150 14422 2202
rect 14474 2150 14486 2202
rect 14538 2150 14550 2202
rect 14602 2150 18860 2202
rect 1104 2128 18860 2150
rect 4798 2048 4804 2100
rect 4856 2088 4862 2100
rect 9122 2088 9128 2100
rect 4856 2060 9128 2088
rect 4856 2048 4862 2060
rect 9122 2048 9128 2060
rect 9180 2048 9186 2100
rect 11146 2088 11152 2100
rect 10244 2060 11152 2088
rect 6178 1980 6184 2032
rect 6236 2020 6242 2032
rect 10244 2020 10272 2060
rect 11146 2048 11152 2060
rect 11204 2048 11210 2100
rect 11330 2048 11336 2100
rect 11388 2088 11394 2100
rect 13722 2088 13728 2100
rect 11388 2060 13728 2088
rect 11388 2048 11394 2060
rect 13722 2048 13728 2060
rect 13780 2048 13786 2100
rect 14734 2048 14740 2100
rect 14792 2088 14798 2100
rect 16114 2088 16120 2100
rect 14792 2060 16120 2088
rect 14792 2048 14798 2060
rect 16114 2048 16120 2060
rect 16172 2048 16178 2100
rect 6236 1992 10272 2020
rect 6236 1980 6242 1992
rect 10410 1980 10416 2032
rect 10468 2020 10474 2032
rect 13630 2020 13636 2032
rect 10468 1992 13636 2020
rect 10468 1980 10474 1992
rect 13630 1980 13636 1992
rect 13688 2020 13694 2032
rect 17218 2020 17224 2032
rect 13688 1992 17224 2020
rect 13688 1980 13694 1992
rect 17218 1980 17224 1992
rect 17276 1980 17282 2032
rect 5994 1912 6000 1964
rect 6052 1952 6058 1964
rect 12342 1952 12348 1964
rect 6052 1924 12348 1952
rect 6052 1912 6058 1924
rect 12342 1912 12348 1924
rect 12400 1912 12406 1964
rect 14642 1912 14648 1964
rect 14700 1952 14706 1964
rect 17034 1952 17040 1964
rect 14700 1924 17040 1952
rect 14700 1912 14706 1924
rect 17034 1912 17040 1924
rect 17092 1952 17098 1964
rect 17494 1952 17500 1964
rect 17092 1924 17500 1952
rect 17092 1912 17098 1924
rect 17494 1912 17500 1924
rect 17552 1912 17558 1964
rect 4062 1844 4068 1896
rect 4120 1884 4126 1896
rect 6822 1884 6828 1896
rect 4120 1856 6828 1884
rect 4120 1844 4126 1856
rect 6822 1844 6828 1856
rect 6880 1844 6886 1896
rect 8110 1844 8116 1896
rect 8168 1884 8174 1896
rect 11330 1884 11336 1896
rect 8168 1856 11336 1884
rect 8168 1844 8174 1856
rect 11330 1844 11336 1856
rect 11388 1844 11394 1896
rect 12158 1844 12164 1896
rect 12216 1884 12222 1896
rect 14090 1884 14096 1896
rect 12216 1856 14096 1884
rect 12216 1844 12222 1856
rect 14090 1844 14096 1856
rect 14148 1844 14154 1896
rect 5718 1776 5724 1828
rect 5776 1816 5782 1828
rect 10594 1816 10600 1828
rect 5776 1788 10600 1816
rect 5776 1776 5782 1788
rect 10594 1776 10600 1788
rect 10652 1776 10658 1828
rect 11422 1776 11428 1828
rect 11480 1816 11486 1828
rect 16666 1816 16672 1828
rect 11480 1788 16672 1816
rect 11480 1776 11486 1788
rect 16666 1776 16672 1788
rect 16724 1776 16730 1828
rect 5074 1708 5080 1760
rect 5132 1748 5138 1760
rect 9766 1748 9772 1760
rect 5132 1720 9772 1748
rect 5132 1708 5138 1720
rect 9766 1708 9772 1720
rect 9824 1708 9830 1760
rect 3878 1640 3884 1692
rect 3936 1680 3942 1692
rect 7466 1680 7472 1692
rect 3936 1652 7472 1680
rect 3936 1640 3942 1652
rect 7466 1640 7472 1652
rect 7524 1640 7530 1692
rect 13078 1504 13084 1556
rect 13136 1544 13142 1556
rect 15194 1544 15200 1556
rect 13136 1516 15200 1544
rect 13136 1504 13142 1516
rect 15194 1504 15200 1516
rect 15252 1504 15258 1556
rect 3326 1436 3332 1488
rect 3384 1476 3390 1488
rect 7190 1476 7196 1488
rect 3384 1448 7196 1476
rect 3384 1436 3390 1448
rect 7190 1436 7196 1448
rect 7248 1436 7254 1488
rect 3694 1232 3700 1284
rect 3752 1272 3758 1284
rect 5810 1272 5816 1284
rect 3752 1244 5816 1272
rect 3752 1232 3758 1244
rect 5810 1232 5816 1244
rect 5868 1232 5874 1284
rect 11238 1164 11244 1216
rect 11296 1204 11302 1216
rect 15010 1204 15016 1216
rect 11296 1176 15016 1204
rect 11296 1164 11302 1176
rect 15010 1164 15016 1176
rect 15068 1164 15074 1216
rect 4062 1028 4068 1080
rect 4120 1068 4126 1080
rect 11790 1068 11796 1080
rect 4120 1040 11796 1068
rect 4120 1028 4126 1040
rect 11790 1028 11796 1040
rect 11848 1028 11854 1080
<< via1 >>
rect 3700 15376 3752 15428
rect 7472 15376 7524 15428
rect 13176 15308 13228 15360
rect 18052 15308 18104 15360
rect 3516 15172 3568 15224
rect 9220 15172 9272 15224
rect 13268 15172 13320 15224
rect 15200 15172 15252 15224
rect 3174 14662 3226 14714
rect 3238 14662 3290 14714
rect 3302 14662 3354 14714
rect 3366 14662 3418 14714
rect 3430 14662 3482 14714
rect 7622 14662 7674 14714
rect 7686 14662 7738 14714
rect 7750 14662 7802 14714
rect 7814 14662 7866 14714
rect 7878 14662 7930 14714
rect 12070 14662 12122 14714
rect 12134 14662 12186 14714
rect 12198 14662 12250 14714
rect 12262 14662 12314 14714
rect 12326 14662 12378 14714
rect 16518 14662 16570 14714
rect 16582 14662 16634 14714
rect 16646 14662 16698 14714
rect 16710 14662 16762 14714
rect 16774 14662 16826 14714
rect 3792 14424 3844 14476
rect 10508 14424 10560 14476
rect 10600 14424 10652 14476
rect 15292 14424 15344 14476
rect 1124 14356 1176 14408
rect 13084 14356 13136 14408
rect 5540 14288 5592 14340
rect 18052 14288 18104 14340
rect 4068 14220 4120 14272
rect 7196 14220 7248 14272
rect 7564 14220 7616 14272
rect 15660 14220 15712 14272
rect 5398 14118 5450 14170
rect 5462 14118 5514 14170
rect 5526 14118 5578 14170
rect 5590 14118 5642 14170
rect 5654 14118 5706 14170
rect 9846 14118 9898 14170
rect 9910 14118 9962 14170
rect 9974 14118 10026 14170
rect 10038 14118 10090 14170
rect 10102 14118 10154 14170
rect 14294 14118 14346 14170
rect 14358 14118 14410 14170
rect 14422 14118 14474 14170
rect 14486 14118 14538 14170
rect 14550 14118 14602 14170
rect 3884 14016 3936 14068
rect 2136 13948 2188 14000
rect 4988 13948 5040 14000
rect 4896 13923 4948 13932
rect 4896 13889 4905 13923
rect 4905 13889 4939 13923
rect 4939 13889 4948 13923
rect 4896 13880 4948 13889
rect 10968 14016 11020 14068
rect 5172 13948 5224 14000
rect 7564 13948 7616 14000
rect 15200 14016 15252 14068
rect 18052 14059 18104 14068
rect 13084 13991 13136 14000
rect 13084 13957 13093 13991
rect 13093 13957 13127 13991
rect 13127 13957 13136 13991
rect 13084 13948 13136 13957
rect 14188 13948 14240 14000
rect 15108 13948 15160 14000
rect 16948 13948 17000 14000
rect 18052 14025 18061 14059
rect 18061 14025 18095 14059
rect 18095 14025 18104 14059
rect 18052 14016 18104 14025
rect 18512 14016 18564 14068
rect 18788 13948 18840 14000
rect 13636 13923 13688 13932
rect 13636 13889 13645 13923
rect 13645 13889 13679 13923
rect 13679 13889 13688 13923
rect 13636 13880 13688 13889
rect 17868 13923 17920 13932
rect 4804 13855 4856 13864
rect 4804 13821 4813 13855
rect 4813 13821 4847 13855
rect 4847 13821 4856 13855
rect 4804 13812 4856 13821
rect 6920 13855 6972 13864
rect 6920 13821 6929 13855
rect 6929 13821 6963 13855
rect 6963 13821 6972 13855
rect 6920 13812 6972 13821
rect 13452 13812 13504 13864
rect 13544 13812 13596 13864
rect 17868 13889 17877 13923
rect 17877 13889 17911 13923
rect 17911 13889 17920 13923
rect 17868 13880 17920 13889
rect 18052 13880 18104 13932
rect 5172 13744 5224 13796
rect 4436 13676 4488 13728
rect 5816 13676 5868 13728
rect 6092 13676 6144 13728
rect 15568 13744 15620 13796
rect 16856 13812 16908 13864
rect 17040 13855 17092 13864
rect 17040 13821 17049 13855
rect 17049 13821 17083 13855
rect 17083 13821 17092 13855
rect 17040 13812 17092 13821
rect 17132 13744 17184 13796
rect 9404 13676 9456 13728
rect 10600 13676 10652 13728
rect 14740 13719 14792 13728
rect 14740 13685 14749 13719
rect 14749 13685 14783 13719
rect 14783 13685 14792 13719
rect 14740 13676 14792 13685
rect 3174 13574 3226 13626
rect 3238 13574 3290 13626
rect 3302 13574 3354 13626
rect 3366 13574 3418 13626
rect 3430 13574 3482 13626
rect 7622 13574 7674 13626
rect 7686 13574 7738 13626
rect 7750 13574 7802 13626
rect 7814 13574 7866 13626
rect 7878 13574 7930 13626
rect 12070 13574 12122 13626
rect 12134 13574 12186 13626
rect 12198 13574 12250 13626
rect 12262 13574 12314 13626
rect 12326 13574 12378 13626
rect 16518 13574 16570 13626
rect 16582 13574 16634 13626
rect 16646 13574 16698 13626
rect 16710 13574 16762 13626
rect 16774 13574 16826 13626
rect 3884 13515 3936 13524
rect 3884 13481 3893 13515
rect 3893 13481 3927 13515
rect 3927 13481 3936 13515
rect 3884 13472 3936 13481
rect 4896 13472 4948 13524
rect 3976 13404 4028 13456
rect 5264 13404 5316 13456
rect 4160 13268 4212 13320
rect 4620 13336 4672 13388
rect 8484 13472 8536 13524
rect 10232 13472 10284 13524
rect 13636 13472 13688 13524
rect 16856 13472 16908 13524
rect 10508 13447 10560 13456
rect 10508 13413 10517 13447
rect 10517 13413 10551 13447
rect 10551 13413 10560 13447
rect 10508 13404 10560 13413
rect 16948 13404 17000 13456
rect 5724 13379 5776 13388
rect 5724 13345 5733 13379
rect 5733 13345 5767 13379
rect 5767 13345 5776 13379
rect 5724 13336 5776 13345
rect 6552 13379 6604 13388
rect 6552 13345 6561 13379
rect 6561 13345 6595 13379
rect 6595 13345 6604 13379
rect 6552 13336 6604 13345
rect 8484 13336 8536 13388
rect 9404 13379 9456 13388
rect 9404 13345 9413 13379
rect 9413 13345 9447 13379
rect 9447 13345 9456 13379
rect 9404 13336 9456 13345
rect 9680 13336 9732 13388
rect 11888 13336 11940 13388
rect 15108 13336 15160 13388
rect 6920 13268 6972 13320
rect 7840 13268 7892 13320
rect 9036 13268 9088 13320
rect 10968 13268 11020 13320
rect 12164 13268 12216 13320
rect 15200 13311 15252 13320
rect 15200 13277 15209 13311
rect 15209 13277 15243 13311
rect 15243 13277 15252 13311
rect 15200 13268 15252 13277
rect 18052 13311 18104 13320
rect 18052 13277 18061 13311
rect 18061 13277 18095 13311
rect 18095 13277 18104 13311
rect 18052 13268 18104 13277
rect 1952 13132 2004 13184
rect 3884 13132 3936 13184
rect 4896 13132 4948 13184
rect 5264 13200 5316 13252
rect 5816 13132 5868 13184
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 6920 13175 6972 13184
rect 6920 13141 6929 13175
rect 6929 13141 6963 13175
rect 6963 13141 6972 13175
rect 6920 13132 6972 13141
rect 7012 13175 7064 13184
rect 7012 13141 7021 13175
rect 7021 13141 7055 13175
rect 7055 13141 7064 13175
rect 8024 13200 8076 13252
rect 8944 13175 8996 13184
rect 7012 13132 7064 13141
rect 8944 13141 8953 13175
rect 8953 13141 8987 13175
rect 8987 13141 8996 13175
rect 8944 13132 8996 13141
rect 9312 13175 9364 13184
rect 9312 13141 9321 13175
rect 9321 13141 9355 13175
rect 9355 13141 9364 13175
rect 9312 13132 9364 13141
rect 10416 13175 10468 13184
rect 10416 13141 10425 13175
rect 10425 13141 10459 13175
rect 10459 13141 10468 13175
rect 10416 13132 10468 13141
rect 14740 13200 14792 13252
rect 17132 13200 17184 13252
rect 18696 13200 18748 13252
rect 14004 13132 14056 13184
rect 15292 13132 15344 13184
rect 17224 13132 17276 13184
rect 17868 13132 17920 13184
rect 5398 13030 5450 13082
rect 5462 13030 5514 13082
rect 5526 13030 5578 13082
rect 5590 13030 5642 13082
rect 5654 13030 5706 13082
rect 9846 13030 9898 13082
rect 9910 13030 9962 13082
rect 9974 13030 10026 13082
rect 10038 13030 10090 13082
rect 10102 13030 10154 13082
rect 14294 13030 14346 13082
rect 14358 13030 14410 13082
rect 14422 13030 14474 13082
rect 14486 13030 14538 13082
rect 14550 13030 14602 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 3884 12860 3936 12912
rect 4436 12928 4488 12980
rect 4804 12928 4856 12980
rect 5816 12928 5868 12980
rect 8944 12928 8996 12980
rect 4712 12860 4764 12912
rect 7380 12860 7432 12912
rect 5816 12835 5868 12844
rect 2780 12767 2832 12776
rect 2780 12733 2789 12767
rect 2789 12733 2823 12767
rect 2823 12733 2832 12767
rect 2780 12724 2832 12733
rect 4620 12724 4672 12776
rect 5080 12767 5132 12776
rect 5080 12733 5089 12767
rect 5089 12733 5123 12767
rect 5123 12733 5132 12767
rect 5080 12724 5132 12733
rect 1952 12631 2004 12640
rect 1952 12597 1961 12631
rect 1961 12597 1995 12631
rect 1995 12597 2004 12631
rect 1952 12588 2004 12597
rect 2136 12631 2188 12640
rect 2136 12597 2145 12631
rect 2145 12597 2179 12631
rect 2179 12597 2188 12631
rect 2136 12588 2188 12597
rect 5816 12801 5825 12835
rect 5825 12801 5859 12835
rect 5859 12801 5868 12835
rect 5816 12792 5868 12801
rect 6092 12792 6144 12844
rect 7012 12792 7064 12844
rect 8116 12860 8168 12912
rect 13084 12928 13136 12980
rect 13544 12971 13596 12980
rect 13544 12937 13553 12971
rect 13553 12937 13587 12971
rect 13587 12937 13596 12971
rect 13544 12928 13596 12937
rect 9680 12860 9732 12912
rect 7840 12835 7892 12844
rect 7840 12801 7849 12835
rect 7849 12801 7883 12835
rect 7883 12801 7892 12835
rect 7840 12792 7892 12801
rect 10968 12860 11020 12912
rect 18144 12928 18196 12980
rect 13820 12860 13872 12912
rect 14832 12903 14884 12912
rect 14832 12869 14850 12903
rect 14850 12869 14884 12903
rect 14832 12860 14884 12869
rect 5908 12767 5960 12776
rect 5908 12733 5917 12767
rect 5917 12733 5951 12767
rect 5951 12733 5960 12767
rect 5908 12724 5960 12733
rect 4160 12631 4212 12640
rect 4160 12597 4169 12631
rect 4169 12597 4203 12631
rect 4203 12597 4212 12631
rect 5724 12656 5776 12708
rect 6552 12656 6604 12708
rect 4160 12588 4212 12597
rect 4528 12631 4580 12640
rect 4528 12597 4537 12631
rect 4537 12597 4571 12631
rect 4571 12597 4580 12631
rect 4528 12588 4580 12597
rect 5816 12588 5868 12640
rect 7104 12588 7156 12640
rect 10232 12792 10284 12844
rect 8392 12767 8444 12776
rect 8392 12733 8401 12767
rect 8401 12733 8435 12767
rect 8435 12733 8444 12767
rect 8392 12724 8444 12733
rect 12164 12767 12216 12776
rect 12164 12733 12173 12767
rect 12173 12733 12207 12767
rect 12207 12733 12216 12767
rect 12164 12724 12216 12733
rect 13820 12724 13872 12776
rect 14556 12792 14608 12844
rect 15016 12792 15068 12844
rect 9036 12656 9088 12708
rect 17500 12792 17552 12844
rect 18328 12792 18380 12844
rect 15844 12767 15896 12776
rect 15844 12733 15853 12767
rect 15853 12733 15887 12767
rect 15887 12733 15896 12767
rect 15844 12724 15896 12733
rect 18144 12767 18196 12776
rect 18144 12733 18153 12767
rect 18153 12733 18187 12767
rect 18187 12733 18196 12767
rect 18144 12724 18196 12733
rect 8852 12631 8904 12640
rect 8852 12597 8861 12631
rect 8861 12597 8895 12631
rect 8895 12597 8904 12631
rect 8852 12588 8904 12597
rect 9588 12588 9640 12640
rect 11060 12631 11112 12640
rect 11060 12597 11069 12631
rect 11069 12597 11103 12631
rect 11103 12597 11112 12631
rect 11060 12588 11112 12597
rect 11796 12588 11848 12640
rect 15108 12588 15160 12640
rect 15384 12631 15436 12640
rect 15384 12597 15393 12631
rect 15393 12597 15427 12631
rect 15427 12597 15436 12631
rect 15384 12588 15436 12597
rect 17040 12588 17092 12640
rect 17776 12656 17828 12708
rect 17592 12631 17644 12640
rect 17592 12597 17601 12631
rect 17601 12597 17635 12631
rect 17635 12597 17644 12631
rect 17592 12588 17644 12597
rect 3174 12486 3226 12538
rect 3238 12486 3290 12538
rect 3302 12486 3354 12538
rect 3366 12486 3418 12538
rect 3430 12486 3482 12538
rect 7622 12486 7674 12538
rect 7686 12486 7738 12538
rect 7750 12486 7802 12538
rect 7814 12486 7866 12538
rect 7878 12486 7930 12538
rect 12070 12486 12122 12538
rect 12134 12486 12186 12538
rect 12198 12486 12250 12538
rect 12262 12486 12314 12538
rect 12326 12486 12378 12538
rect 16518 12486 16570 12538
rect 16582 12486 16634 12538
rect 16646 12486 16698 12538
rect 16710 12486 16762 12538
rect 16774 12486 16826 12538
rect 4804 12384 4856 12436
rect 5080 12384 5132 12436
rect 5908 12384 5960 12436
rect 8760 12427 8812 12436
rect 8760 12393 8769 12427
rect 8769 12393 8803 12427
rect 8803 12393 8812 12427
rect 8760 12384 8812 12393
rect 10232 12384 10284 12436
rect 5172 12359 5224 12368
rect 5172 12325 5181 12359
rect 5181 12325 5215 12359
rect 5215 12325 5224 12359
rect 5172 12316 5224 12325
rect 2320 12180 2372 12232
rect 2964 12223 3016 12232
rect 2964 12189 2973 12223
rect 2973 12189 3007 12223
rect 3007 12189 3016 12223
rect 2964 12180 3016 12189
rect 3792 12223 3844 12232
rect 3792 12189 3801 12223
rect 3801 12189 3835 12223
rect 3835 12189 3844 12223
rect 3792 12180 3844 12189
rect 5724 12248 5776 12300
rect 7196 12316 7248 12368
rect 9680 12316 9732 12368
rect 7012 12248 7064 12300
rect 7380 12291 7432 12300
rect 7380 12257 7389 12291
rect 7389 12257 7423 12291
rect 7423 12257 7432 12291
rect 7380 12248 7432 12257
rect 9312 12248 9364 12300
rect 9588 12248 9640 12300
rect 14740 12384 14792 12436
rect 14556 12316 14608 12368
rect 7104 12180 7156 12232
rect 10416 12180 10468 12232
rect 10508 12223 10560 12232
rect 10508 12189 10517 12223
rect 10517 12189 10551 12223
rect 10551 12189 10560 12223
rect 10508 12180 10560 12189
rect 11336 12180 11388 12232
rect 12440 12180 12492 12232
rect 12992 12180 13044 12232
rect 13452 12223 13504 12232
rect 13452 12189 13461 12223
rect 13461 12189 13495 12223
rect 13495 12189 13504 12223
rect 13452 12180 13504 12189
rect 15384 12291 15436 12300
rect 15384 12257 15393 12291
rect 15393 12257 15427 12291
rect 15427 12257 15436 12291
rect 15384 12248 15436 12257
rect 15936 12316 15988 12368
rect 18144 12248 18196 12300
rect 14924 12180 14976 12232
rect 17408 12223 17460 12232
rect 17408 12189 17417 12223
rect 17417 12189 17451 12223
rect 17451 12189 17460 12223
rect 17408 12180 17460 12189
rect 17776 12180 17828 12232
rect 2044 12112 2096 12164
rect 2596 12155 2648 12164
rect 2596 12121 2605 12155
rect 2605 12121 2639 12155
rect 2639 12121 2648 12155
rect 2596 12112 2648 12121
rect 1492 12087 1544 12096
rect 1492 12053 1501 12087
rect 1501 12053 1535 12087
rect 1535 12053 1544 12087
rect 1492 12044 1544 12053
rect 1768 12087 1820 12096
rect 1768 12053 1777 12087
rect 1777 12053 1811 12087
rect 1811 12053 1820 12087
rect 1768 12044 1820 12053
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 3608 12087 3660 12096
rect 3608 12053 3617 12087
rect 3617 12053 3651 12087
rect 3651 12053 3660 12087
rect 3608 12044 3660 12053
rect 4160 12112 4212 12164
rect 4252 12112 4304 12164
rect 4528 12112 4580 12164
rect 6736 12112 6788 12164
rect 9496 12112 9548 12164
rect 5264 12044 5316 12096
rect 5724 12087 5776 12096
rect 5724 12053 5733 12087
rect 5733 12053 5767 12087
rect 5767 12053 5776 12087
rect 5724 12044 5776 12053
rect 6552 12044 6604 12096
rect 6828 12044 6880 12096
rect 8944 12044 8996 12096
rect 9772 12087 9824 12096
rect 9772 12053 9781 12087
rect 9781 12053 9815 12087
rect 9815 12053 9824 12087
rect 9772 12044 9824 12053
rect 10600 12087 10652 12096
rect 10600 12053 10609 12087
rect 10609 12053 10643 12087
rect 10643 12053 10652 12087
rect 10600 12044 10652 12053
rect 10784 12044 10836 12096
rect 11520 12044 11572 12096
rect 11704 12044 11756 12096
rect 14188 12112 14240 12164
rect 14096 12087 14148 12096
rect 14096 12053 14105 12087
rect 14105 12053 14139 12087
rect 14139 12053 14148 12087
rect 14096 12044 14148 12053
rect 17316 12112 17368 12164
rect 14648 12044 14700 12096
rect 15200 12044 15252 12096
rect 16488 12044 16540 12096
rect 18420 12112 18472 12164
rect 17868 12044 17920 12096
rect 5398 11942 5450 11994
rect 5462 11942 5514 11994
rect 5526 11942 5578 11994
rect 5590 11942 5642 11994
rect 5654 11942 5706 11994
rect 9846 11942 9898 11994
rect 9910 11942 9962 11994
rect 9974 11942 10026 11994
rect 10038 11942 10090 11994
rect 10102 11942 10154 11994
rect 14294 11942 14346 11994
rect 14358 11942 14410 11994
rect 14422 11942 14474 11994
rect 14486 11942 14538 11994
rect 14550 11942 14602 11994
rect 2688 11840 2740 11892
rect 4252 11840 4304 11892
rect 5724 11840 5776 11892
rect 6552 11840 6604 11892
rect 7656 11840 7708 11892
rect 1676 11772 1728 11824
rect 1952 11772 2004 11824
rect 3516 11815 3568 11824
rect 3516 11781 3525 11815
rect 3525 11781 3559 11815
rect 3559 11781 3568 11815
rect 3516 11772 3568 11781
rect 4068 11772 4120 11824
rect 1584 11704 1636 11756
rect 3700 11704 3752 11756
rect 4712 11704 4764 11756
rect 2228 11636 2280 11688
rect 3516 11636 3568 11688
rect 3792 11636 3844 11688
rect 4068 11679 4120 11688
rect 4068 11645 4077 11679
rect 4077 11645 4111 11679
rect 4111 11645 4120 11679
rect 4068 11636 4120 11645
rect 5172 11704 5224 11756
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 6828 11679 6880 11688
rect 6828 11645 6837 11679
rect 6837 11645 6871 11679
rect 6871 11645 6880 11679
rect 6828 11636 6880 11645
rect 6736 11568 6788 11620
rect 8208 11704 8260 11756
rect 7012 11679 7064 11688
rect 7012 11645 7021 11679
rect 7021 11645 7055 11679
rect 7055 11645 7064 11679
rect 7012 11636 7064 11645
rect 7196 11636 7248 11688
rect 7656 11679 7708 11688
rect 7656 11645 7665 11679
rect 7665 11645 7699 11679
rect 7699 11645 7708 11679
rect 7656 11636 7708 11645
rect 2044 11500 2096 11552
rect 2504 11500 2556 11552
rect 3792 11543 3844 11552
rect 3792 11509 3801 11543
rect 3801 11509 3835 11543
rect 3835 11509 3844 11543
rect 3792 11500 3844 11509
rect 5448 11543 5500 11552
rect 5448 11509 5457 11543
rect 5457 11509 5491 11543
rect 5491 11509 5500 11543
rect 5448 11500 5500 11509
rect 7196 11500 7248 11552
rect 8852 11840 8904 11892
rect 9404 11883 9456 11892
rect 9404 11849 9413 11883
rect 9413 11849 9447 11883
rect 9447 11849 9456 11883
rect 9404 11840 9456 11849
rect 9772 11883 9824 11892
rect 9772 11849 9781 11883
rect 9781 11849 9815 11883
rect 9815 11849 9824 11883
rect 9772 11840 9824 11849
rect 10784 11840 10836 11892
rect 11888 11883 11940 11892
rect 11888 11849 11897 11883
rect 11897 11849 11931 11883
rect 11931 11849 11940 11883
rect 12532 11883 12584 11892
rect 11888 11840 11940 11849
rect 12532 11849 12541 11883
rect 12541 11849 12575 11883
rect 12575 11849 12584 11883
rect 12532 11840 12584 11849
rect 14096 11840 14148 11892
rect 14188 11883 14240 11892
rect 14188 11849 14197 11883
rect 14197 11849 14231 11883
rect 14231 11849 14240 11883
rect 15200 11883 15252 11892
rect 14188 11840 14240 11849
rect 15200 11849 15209 11883
rect 15209 11849 15243 11883
rect 15243 11849 15252 11883
rect 15200 11840 15252 11849
rect 15568 11883 15620 11892
rect 15568 11849 15577 11883
rect 15577 11849 15611 11883
rect 15611 11849 15620 11883
rect 15568 11840 15620 11849
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 17500 11840 17552 11849
rect 8944 11772 8996 11824
rect 14648 11772 14700 11824
rect 15476 11772 15528 11824
rect 16120 11772 16172 11824
rect 17132 11815 17184 11824
rect 17132 11781 17141 11815
rect 17141 11781 17175 11815
rect 17175 11781 17184 11815
rect 17132 11772 17184 11781
rect 8760 11679 8812 11688
rect 8760 11645 8769 11679
rect 8769 11645 8803 11679
rect 8803 11645 8812 11679
rect 8760 11636 8812 11645
rect 9036 11704 9088 11756
rect 9220 11704 9272 11756
rect 9496 11704 9548 11756
rect 10508 11704 10560 11756
rect 10784 11704 10836 11756
rect 8392 11568 8444 11620
rect 9680 11636 9732 11688
rect 10416 11636 10468 11688
rect 10876 11636 10928 11688
rect 10140 11568 10192 11620
rect 10232 11568 10284 11620
rect 11704 11636 11756 11688
rect 11520 11611 11572 11620
rect 11520 11577 11529 11611
rect 11529 11577 11563 11611
rect 11563 11577 11572 11611
rect 11520 11568 11572 11577
rect 13084 11704 13136 11756
rect 13544 11679 13596 11688
rect 13544 11645 13553 11679
rect 13553 11645 13587 11679
rect 13587 11645 13596 11679
rect 13544 11636 13596 11645
rect 14004 11704 14056 11756
rect 15568 11704 15620 11756
rect 16856 11704 16908 11756
rect 14464 11568 14516 11620
rect 14740 11679 14792 11688
rect 14740 11645 14749 11679
rect 14749 11645 14783 11679
rect 14783 11645 14792 11679
rect 14740 11636 14792 11645
rect 16212 11636 16264 11688
rect 17776 11704 17828 11756
rect 17316 11679 17368 11688
rect 17316 11645 17325 11679
rect 17325 11645 17359 11679
rect 17359 11645 17368 11679
rect 17316 11636 17368 11645
rect 15476 11568 15528 11620
rect 16120 11568 16172 11620
rect 17132 11568 17184 11620
rect 13084 11500 13136 11552
rect 13268 11543 13320 11552
rect 13268 11509 13277 11543
rect 13277 11509 13311 11543
rect 13311 11509 13320 11543
rect 13268 11500 13320 11509
rect 14096 11543 14148 11552
rect 14096 11509 14105 11543
rect 14105 11509 14139 11543
rect 14139 11509 14148 11543
rect 14096 11500 14148 11509
rect 16396 11500 16448 11552
rect 3174 11398 3226 11450
rect 3238 11398 3290 11450
rect 3302 11398 3354 11450
rect 3366 11398 3418 11450
rect 3430 11398 3482 11450
rect 7622 11398 7674 11450
rect 7686 11398 7738 11450
rect 7750 11398 7802 11450
rect 7814 11398 7866 11450
rect 7878 11398 7930 11450
rect 12070 11398 12122 11450
rect 12134 11398 12186 11450
rect 12198 11398 12250 11450
rect 12262 11398 12314 11450
rect 12326 11398 12378 11450
rect 16518 11398 16570 11450
rect 16582 11398 16634 11450
rect 16646 11398 16698 11450
rect 16710 11398 16762 11450
rect 16774 11398 16826 11450
rect 2044 11296 2096 11348
rect 6828 11296 6880 11348
rect 7472 11296 7524 11348
rect 8852 11296 8904 11348
rect 9404 11339 9456 11348
rect 9404 11305 9413 11339
rect 9413 11305 9447 11339
rect 9447 11305 9456 11339
rect 9404 11296 9456 11305
rect 10232 11296 10284 11348
rect 10600 11296 10652 11348
rect 11704 11296 11756 11348
rect 4160 11271 4212 11280
rect 4160 11237 4169 11271
rect 4169 11237 4203 11271
rect 4203 11237 4212 11271
rect 4160 11228 4212 11237
rect 4344 11228 4396 11280
rect 6276 11228 6328 11280
rect 3700 11160 3752 11212
rect 3884 11160 3936 11212
rect 1952 11024 2004 11076
rect 2780 11092 2832 11144
rect 4068 11092 4120 11144
rect 6368 11160 6420 11212
rect 6644 11228 6696 11280
rect 7932 11228 7984 11280
rect 9220 11228 9272 11280
rect 6736 11160 6788 11212
rect 2964 11024 3016 11076
rect 3516 11024 3568 11076
rect 2504 10956 2556 11008
rect 4988 11024 5040 11076
rect 5448 11067 5500 11076
rect 5448 11033 5466 11067
rect 5466 11033 5500 11067
rect 5448 11024 5500 11033
rect 6828 11092 6880 11144
rect 6092 11024 6144 11076
rect 6460 11067 6512 11076
rect 6460 11033 6469 11067
rect 6469 11033 6503 11067
rect 6503 11033 6512 11067
rect 6460 11024 6512 11033
rect 7012 11067 7064 11076
rect 7012 11033 7021 11067
rect 7021 11033 7055 11067
rect 7055 11033 7064 11067
rect 7012 11024 7064 11033
rect 8116 11203 8168 11212
rect 8116 11169 8125 11203
rect 8125 11169 8159 11203
rect 8159 11169 8168 11203
rect 8116 11160 8168 11169
rect 8208 11160 8260 11212
rect 9956 11160 10008 11212
rect 11244 11160 11296 11212
rect 14464 11296 14516 11348
rect 12624 11228 12676 11280
rect 8576 11092 8628 11144
rect 11520 11092 11572 11144
rect 11612 11135 11664 11144
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 17316 11296 17368 11348
rect 17776 11296 17828 11348
rect 16396 11228 16448 11280
rect 12900 11203 12952 11212
rect 12900 11169 12909 11203
rect 12909 11169 12943 11203
rect 12943 11169 12952 11203
rect 12900 11160 12952 11169
rect 13268 11160 13320 11212
rect 13728 11203 13780 11212
rect 13728 11169 13737 11203
rect 13737 11169 13771 11203
rect 13771 11169 13780 11203
rect 14924 11203 14976 11212
rect 13728 11160 13780 11169
rect 14924 11169 14933 11203
rect 14933 11169 14967 11203
rect 14967 11169 14976 11203
rect 14924 11160 14976 11169
rect 11612 11092 11664 11101
rect 14096 11092 14148 11144
rect 7932 11067 7984 11076
rect 7932 11033 7941 11067
rect 7941 11033 7975 11067
rect 7975 11033 7984 11067
rect 7932 11024 7984 11033
rect 4620 10956 4672 11008
rect 5080 10956 5132 11008
rect 6552 10999 6604 11008
rect 6552 10965 6561 10999
rect 6561 10965 6595 10999
rect 6595 10965 6604 10999
rect 6552 10956 6604 10965
rect 6920 10999 6972 11008
rect 6920 10965 6929 10999
rect 6929 10965 6963 10999
rect 6963 10965 6972 10999
rect 6920 10956 6972 10965
rect 8208 11024 8260 11076
rect 9220 11067 9272 11076
rect 9220 11033 9229 11067
rect 9229 11033 9263 11067
rect 9263 11033 9272 11067
rect 9220 11024 9272 11033
rect 10692 11067 10744 11076
rect 10692 11033 10710 11067
rect 10710 11033 10744 11067
rect 10692 11024 10744 11033
rect 12256 11067 12308 11076
rect 8300 10956 8352 11008
rect 8852 10956 8904 11008
rect 9036 10999 9088 11008
rect 9036 10965 9045 10999
rect 9045 10965 9079 10999
rect 9079 10965 9088 10999
rect 9036 10956 9088 10965
rect 12256 11033 12265 11067
rect 12265 11033 12299 11067
rect 12299 11033 12308 11067
rect 12256 11024 12308 11033
rect 17408 11092 17460 11144
rect 18144 11092 18196 11144
rect 15292 11024 15344 11076
rect 11888 10956 11940 11008
rect 12808 10999 12860 11008
rect 12808 10965 12817 10999
rect 12817 10965 12851 10999
rect 12851 10965 12860 10999
rect 12808 10956 12860 10965
rect 14832 10999 14884 11008
rect 14832 10965 14841 10999
rect 14841 10965 14875 10999
rect 14875 10965 14884 10999
rect 14832 10956 14884 10965
rect 16672 10999 16724 11008
rect 16672 10965 16681 10999
rect 16681 10965 16715 10999
rect 16715 10965 16724 10999
rect 16672 10956 16724 10965
rect 16856 10956 16908 11008
rect 17684 10956 17736 11008
rect 5398 10854 5450 10906
rect 5462 10854 5514 10906
rect 5526 10854 5578 10906
rect 5590 10854 5642 10906
rect 5654 10854 5706 10906
rect 9846 10854 9898 10906
rect 9910 10854 9962 10906
rect 9974 10854 10026 10906
rect 10038 10854 10090 10906
rect 10102 10854 10154 10906
rect 14294 10854 14346 10906
rect 14358 10854 14410 10906
rect 14422 10854 14474 10906
rect 14486 10854 14538 10906
rect 14550 10854 14602 10906
rect 4160 10752 4212 10804
rect 4804 10752 4856 10804
rect 6368 10752 6420 10804
rect 6644 10795 6696 10804
rect 6644 10761 6653 10795
rect 6653 10761 6687 10795
rect 6687 10761 6696 10795
rect 6644 10752 6696 10761
rect 6920 10752 6972 10804
rect 2504 10727 2556 10736
rect 2504 10693 2522 10727
rect 2522 10693 2556 10727
rect 2504 10684 2556 10693
rect 4620 10684 4672 10736
rect 4896 10684 4948 10736
rect 6460 10684 6512 10736
rect 8300 10752 8352 10804
rect 8576 10795 8628 10804
rect 8576 10761 8585 10795
rect 8585 10761 8619 10795
rect 8619 10761 8628 10795
rect 8576 10752 8628 10761
rect 7380 10684 7432 10736
rect 4160 10616 4212 10668
rect 4344 10616 4396 10668
rect 5908 10616 5960 10668
rect 6644 10616 6696 10668
rect 2780 10591 2832 10600
rect 2780 10557 2789 10591
rect 2789 10557 2823 10591
rect 2823 10557 2832 10591
rect 2780 10548 2832 10557
rect 3056 10548 3108 10600
rect 3516 10591 3568 10600
rect 3516 10557 3525 10591
rect 3525 10557 3559 10591
rect 3559 10557 3568 10591
rect 3516 10548 3568 10557
rect 6828 10616 6880 10668
rect 7472 10659 7524 10668
rect 7472 10625 7506 10659
rect 7506 10625 7524 10659
rect 10692 10752 10744 10804
rect 11152 10752 11204 10804
rect 7472 10616 7524 10625
rect 3792 10523 3844 10532
rect 3792 10489 3801 10523
rect 3801 10489 3835 10523
rect 3835 10489 3844 10523
rect 3792 10480 3844 10489
rect 4804 10480 4856 10532
rect 4988 10480 5040 10532
rect 1584 10412 1636 10464
rect 2504 10412 2556 10464
rect 3884 10455 3936 10464
rect 3884 10421 3893 10455
rect 3893 10421 3927 10455
rect 3927 10421 3936 10455
rect 3884 10412 3936 10421
rect 5724 10412 5776 10464
rect 7104 10548 7156 10600
rect 10876 10616 10928 10668
rect 11060 10548 11112 10600
rect 15384 10752 15436 10804
rect 15844 10752 15896 10804
rect 17868 10752 17920 10804
rect 18328 10795 18380 10804
rect 18328 10761 18337 10795
rect 18337 10761 18371 10795
rect 18371 10761 18380 10795
rect 18328 10752 18380 10761
rect 12716 10684 12768 10736
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 12992 10659 13044 10668
rect 12992 10625 13001 10659
rect 13001 10625 13035 10659
rect 13035 10625 13044 10659
rect 12992 10616 13044 10625
rect 7472 10412 7524 10464
rect 8300 10412 8352 10464
rect 10048 10455 10100 10464
rect 10048 10421 10057 10455
rect 10057 10421 10091 10455
rect 10091 10421 10100 10455
rect 10048 10412 10100 10421
rect 12532 10548 12584 10600
rect 12900 10548 12952 10600
rect 14924 10684 14976 10736
rect 15292 10616 15344 10668
rect 16304 10684 16356 10736
rect 16856 10616 16908 10668
rect 16672 10548 16724 10600
rect 16948 10548 17000 10600
rect 17316 10616 17368 10668
rect 17592 10616 17644 10668
rect 12532 10412 12584 10464
rect 13728 10412 13780 10464
rect 14096 10412 14148 10464
rect 15200 10412 15252 10464
rect 15476 10412 15528 10464
rect 15660 10412 15712 10464
rect 16304 10412 16356 10464
rect 17500 10455 17552 10464
rect 17500 10421 17509 10455
rect 17509 10421 17543 10455
rect 17543 10421 17552 10455
rect 17500 10412 17552 10421
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 3430 10310 3482 10362
rect 7622 10310 7674 10362
rect 7686 10310 7738 10362
rect 7750 10310 7802 10362
rect 7814 10310 7866 10362
rect 7878 10310 7930 10362
rect 12070 10310 12122 10362
rect 12134 10310 12186 10362
rect 12198 10310 12250 10362
rect 12262 10310 12314 10362
rect 12326 10310 12378 10362
rect 16518 10310 16570 10362
rect 16582 10310 16634 10362
rect 16646 10310 16698 10362
rect 16710 10310 16762 10362
rect 16774 10310 16826 10362
rect 112 10140 164 10192
rect 3056 10208 3108 10260
rect 6644 10208 6696 10260
rect 6828 10208 6880 10260
rect 7104 10208 7156 10260
rect 9404 10251 9456 10260
rect 9404 10217 9413 10251
rect 9413 10217 9447 10251
rect 9447 10217 9456 10251
rect 9404 10208 9456 10217
rect 10968 10208 11020 10260
rect 12716 10208 12768 10260
rect 12808 10208 12860 10260
rect 2596 10115 2648 10124
rect 2596 10081 2605 10115
rect 2605 10081 2639 10115
rect 2639 10081 2648 10115
rect 2596 10072 2648 10081
rect 4344 10140 4396 10192
rect 7564 10183 7616 10192
rect 7564 10149 7573 10183
rect 7573 10149 7607 10183
rect 7607 10149 7616 10183
rect 7564 10140 7616 10149
rect 7748 10140 7800 10192
rect 9312 10183 9364 10192
rect 9312 10149 9321 10183
rect 9321 10149 9355 10183
rect 9355 10149 9364 10183
rect 9312 10140 9364 10149
rect 11796 10140 11848 10192
rect 3516 10115 3568 10124
rect 3516 10081 3525 10115
rect 3525 10081 3559 10115
rect 3559 10081 3568 10115
rect 3516 10072 3568 10081
rect 4160 10072 4212 10124
rect 4620 10072 4672 10124
rect 4988 10115 5040 10124
rect 4988 10081 4997 10115
rect 4997 10081 5031 10115
rect 5031 10081 5040 10115
rect 4988 10072 5040 10081
rect 6736 10072 6788 10124
rect 8024 10072 8076 10124
rect 8116 10072 8168 10124
rect 10048 10072 10100 10124
rect 10784 10072 10836 10124
rect 11520 10072 11572 10124
rect 11980 10072 12032 10124
rect 12992 10140 13044 10192
rect 14096 10140 14148 10192
rect 15844 10140 15896 10192
rect 16856 10140 16908 10192
rect 13728 10115 13780 10124
rect 13728 10081 13737 10115
rect 13737 10081 13771 10115
rect 13771 10081 13780 10115
rect 13728 10072 13780 10081
rect 15200 10072 15252 10124
rect 16948 10115 17000 10124
rect 16948 10081 16957 10115
rect 16957 10081 16991 10115
rect 16991 10081 17000 10115
rect 16948 10072 17000 10081
rect 18144 10072 18196 10124
rect 3884 10004 3936 10056
rect 4068 10004 4120 10056
rect 4896 10047 4948 10056
rect 4896 10013 4905 10047
rect 4905 10013 4939 10047
rect 4939 10013 4948 10047
rect 4896 10004 4948 10013
rect 5264 10047 5316 10056
rect 5264 10013 5273 10047
rect 5273 10013 5307 10047
rect 5307 10013 5316 10047
rect 5264 10004 5316 10013
rect 10876 10004 10928 10056
rect 12624 10047 12676 10056
rect 12624 10013 12633 10047
rect 12633 10013 12667 10047
rect 12667 10013 12676 10047
rect 12624 10004 12676 10013
rect 14924 10004 14976 10056
rect 17500 10004 17552 10056
rect 17960 10004 18012 10056
rect 2688 9936 2740 9988
rect 2136 9868 2188 9920
rect 3332 9868 3384 9920
rect 6000 9936 6052 9988
rect 8208 9936 8260 9988
rect 9404 9936 9456 9988
rect 4896 9868 4948 9920
rect 7748 9868 7800 9920
rect 8668 9868 8720 9920
rect 8852 9868 8904 9920
rect 9036 9911 9088 9920
rect 9036 9877 9045 9911
rect 9045 9877 9079 9911
rect 9079 9877 9088 9911
rect 9036 9868 9088 9877
rect 9588 9911 9640 9920
rect 9588 9877 9597 9911
rect 9597 9877 9631 9911
rect 9631 9877 9640 9911
rect 9588 9868 9640 9877
rect 10232 9936 10284 9988
rect 14188 9936 14240 9988
rect 14832 9936 14884 9988
rect 12348 9868 12400 9920
rect 12992 9911 13044 9920
rect 12992 9877 13001 9911
rect 13001 9877 13035 9911
rect 13035 9877 13044 9911
rect 12992 9868 13044 9877
rect 13084 9868 13136 9920
rect 13360 9868 13412 9920
rect 13544 9911 13596 9920
rect 13544 9877 13553 9911
rect 13553 9877 13587 9911
rect 13587 9877 13596 9911
rect 13544 9868 13596 9877
rect 15476 9868 15528 9920
rect 15752 9868 15804 9920
rect 17132 9868 17184 9920
rect 18604 9936 18656 9988
rect 5398 9766 5450 9818
rect 5462 9766 5514 9818
rect 5526 9766 5578 9818
rect 5590 9766 5642 9818
rect 5654 9766 5706 9818
rect 9846 9766 9898 9818
rect 9910 9766 9962 9818
rect 9974 9766 10026 9818
rect 10038 9766 10090 9818
rect 10102 9766 10154 9818
rect 14294 9766 14346 9818
rect 14358 9766 14410 9818
rect 14422 9766 14474 9818
rect 14486 9766 14538 9818
rect 14550 9766 14602 9818
rect 1676 9664 1728 9716
rect 2780 9596 2832 9648
rect 2964 9596 3016 9648
rect 6000 9664 6052 9716
rect 5080 9596 5132 9648
rect 7380 9664 7432 9716
rect 7472 9664 7524 9716
rect 9588 9664 9640 9716
rect 10232 9664 10284 9716
rect 14648 9664 14700 9716
rect 14924 9664 14976 9716
rect 2228 9571 2280 9580
rect 2228 9537 2262 9571
rect 2262 9537 2280 9571
rect 2228 9528 2280 9537
rect 4896 9528 4948 9580
rect 5172 9528 5224 9580
rect 6184 9528 6236 9580
rect 6828 9596 6880 9648
rect 7288 9596 7340 9648
rect 8944 9596 8996 9648
rect 1308 9324 1360 9376
rect 1492 9324 1544 9376
rect 1676 9367 1728 9376
rect 1676 9333 1685 9367
rect 1685 9333 1719 9367
rect 1719 9333 1728 9367
rect 1676 9324 1728 9333
rect 1952 9324 2004 9376
rect 6000 9460 6052 9512
rect 6920 9528 6972 9580
rect 8116 9528 8168 9580
rect 8484 9503 8536 9512
rect 8484 9469 8493 9503
rect 8493 9469 8527 9503
rect 8527 9469 8536 9503
rect 8484 9460 8536 9469
rect 9312 9528 9364 9580
rect 10784 9571 10836 9580
rect 10784 9537 10802 9571
rect 10802 9537 10836 9571
rect 10784 9528 10836 9537
rect 9128 9503 9180 9512
rect 9128 9469 9137 9503
rect 9137 9469 9171 9503
rect 9171 9469 9180 9503
rect 9128 9460 9180 9469
rect 12532 9596 12584 9648
rect 12716 9596 12768 9648
rect 12072 9503 12124 9512
rect 12072 9469 12081 9503
rect 12081 9469 12115 9503
rect 12115 9469 12124 9503
rect 12072 9460 12124 9469
rect 4068 9324 4120 9376
rect 5172 9367 5224 9376
rect 5172 9333 5181 9367
rect 5181 9333 5215 9367
rect 5215 9333 5224 9367
rect 5172 9324 5224 9333
rect 7104 9324 7156 9376
rect 7380 9324 7432 9376
rect 8392 9324 8444 9376
rect 8852 9324 8904 9376
rect 9128 9324 9180 9376
rect 9588 9367 9640 9376
rect 9588 9333 9597 9367
rect 9597 9333 9631 9367
rect 9631 9333 9640 9367
rect 9588 9324 9640 9333
rect 11980 9392 12032 9444
rect 12348 9392 12400 9444
rect 12808 9528 12860 9580
rect 13728 9596 13780 9648
rect 13084 9503 13136 9512
rect 13084 9469 13093 9503
rect 13093 9469 13127 9503
rect 13127 9469 13136 9503
rect 13084 9460 13136 9469
rect 14096 9528 14148 9580
rect 13728 9460 13780 9512
rect 18144 9664 18196 9716
rect 17960 9596 18012 9648
rect 15844 9571 15896 9580
rect 15844 9537 15853 9571
rect 15853 9537 15887 9571
rect 15887 9537 15896 9571
rect 15844 9528 15896 9537
rect 17500 9528 17552 9580
rect 16856 9503 16908 9512
rect 16856 9469 16865 9503
rect 16865 9469 16899 9503
rect 16899 9469 16908 9503
rect 16856 9460 16908 9469
rect 13452 9435 13504 9444
rect 13452 9401 13461 9435
rect 13461 9401 13495 9435
rect 13495 9401 13504 9435
rect 13452 9392 13504 9401
rect 10140 9324 10192 9376
rect 10876 9324 10928 9376
rect 15384 9324 15436 9376
rect 16212 9324 16264 9376
rect 16764 9392 16816 9444
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 3430 9222 3482 9274
rect 7622 9222 7674 9274
rect 7686 9222 7738 9274
rect 7750 9222 7802 9274
rect 7814 9222 7866 9274
rect 7878 9222 7930 9274
rect 12070 9222 12122 9274
rect 12134 9222 12186 9274
rect 12198 9222 12250 9274
rect 12262 9222 12314 9274
rect 12326 9222 12378 9274
rect 16518 9222 16570 9274
rect 16582 9222 16634 9274
rect 16646 9222 16698 9274
rect 16710 9222 16762 9274
rect 16774 9222 16826 9274
rect 4160 9120 4212 9172
rect 4344 9163 4396 9172
rect 4344 9129 4353 9163
rect 4353 9129 4387 9163
rect 4387 9129 4396 9163
rect 4344 9120 4396 9129
rect 7288 9120 7340 9172
rect 2780 9052 2832 9104
rect 2504 9027 2556 9036
rect 2504 8993 2513 9027
rect 2513 8993 2547 9027
rect 2547 8993 2556 9027
rect 2504 8984 2556 8993
rect 2596 9027 2648 9036
rect 2596 8993 2605 9027
rect 2605 8993 2639 9027
rect 2639 8993 2648 9027
rect 2964 9027 3016 9036
rect 2596 8984 2648 8993
rect 2964 8993 2973 9027
rect 2973 8993 3007 9027
rect 3007 8993 3016 9027
rect 2964 8984 3016 8993
rect 3516 8984 3568 9036
rect 4988 9027 5040 9036
rect 4988 8993 4997 9027
rect 4997 8993 5031 9027
rect 5031 8993 5040 9027
rect 4988 8984 5040 8993
rect 6920 9052 6972 9104
rect 2412 8959 2464 8968
rect 2412 8925 2421 8959
rect 2421 8925 2455 8959
rect 2455 8925 2464 8959
rect 2412 8916 2464 8925
rect 3700 8916 3752 8968
rect 3976 8916 4028 8968
rect 5724 8916 5776 8968
rect 6184 8916 6236 8968
rect 8484 9120 8536 9172
rect 13084 9120 13136 9172
rect 14096 9163 14148 9172
rect 14096 9129 14105 9163
rect 14105 9129 14139 9163
rect 14139 9129 14148 9163
rect 14096 9120 14148 9129
rect 8944 9052 8996 9104
rect 9404 9052 9456 9104
rect 10508 9052 10560 9104
rect 12716 9052 12768 9104
rect 9588 8984 9640 9036
rect 10232 9027 10284 9036
rect 10232 8993 10241 9027
rect 10241 8993 10275 9027
rect 10275 8993 10284 9027
rect 10232 8984 10284 8993
rect 10784 8984 10836 9036
rect 9956 8959 10008 8968
rect 9956 8925 9965 8959
rect 9965 8925 9999 8959
rect 9999 8925 10008 8959
rect 9956 8916 10008 8925
rect 2596 8848 2648 8900
rect 5080 8848 5132 8900
rect 6920 8848 6972 8900
rect 7380 8848 7432 8900
rect 2044 8823 2096 8832
rect 2044 8789 2053 8823
rect 2053 8789 2087 8823
rect 2087 8789 2096 8823
rect 2044 8780 2096 8789
rect 3424 8780 3476 8832
rect 3792 8780 3844 8832
rect 3976 8780 4028 8832
rect 6828 8780 6880 8832
rect 11336 8848 11388 8900
rect 11704 8848 11756 8900
rect 14188 8984 14240 9036
rect 15660 9052 15712 9104
rect 17132 9120 17184 9172
rect 11980 8916 12032 8968
rect 12900 8848 12952 8900
rect 15844 8984 15896 9036
rect 16672 8916 16724 8968
rect 16856 8916 16908 8968
rect 18144 9027 18196 9036
rect 18144 8993 18153 9027
rect 18153 8993 18187 9027
rect 18187 8993 18196 9027
rect 18144 8984 18196 8993
rect 14740 8848 14792 8900
rect 16212 8848 16264 8900
rect 16396 8891 16448 8900
rect 16396 8857 16430 8891
rect 16430 8857 16448 8891
rect 16396 8848 16448 8857
rect 9404 8823 9456 8832
rect 9404 8789 9413 8823
rect 9413 8789 9447 8823
rect 9447 8789 9456 8823
rect 9404 8780 9456 8789
rect 9588 8823 9640 8832
rect 9588 8789 9597 8823
rect 9597 8789 9631 8823
rect 9631 8789 9640 8823
rect 9588 8780 9640 8789
rect 10508 8780 10560 8832
rect 11244 8823 11296 8832
rect 11244 8789 11253 8823
rect 11253 8789 11287 8823
rect 11287 8789 11296 8823
rect 11244 8780 11296 8789
rect 11520 8780 11572 8832
rect 12348 8780 12400 8832
rect 13820 8823 13872 8832
rect 13820 8789 13829 8823
rect 13829 8789 13863 8823
rect 13863 8789 13872 8823
rect 13820 8780 13872 8789
rect 14648 8780 14700 8832
rect 15108 8780 15160 8832
rect 15476 8780 15528 8832
rect 16304 8780 16356 8832
rect 17592 8780 17644 8832
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 5398 8678 5450 8730
rect 5462 8678 5514 8730
rect 5526 8678 5578 8730
rect 5590 8678 5642 8730
rect 5654 8678 5706 8730
rect 9846 8678 9898 8730
rect 9910 8678 9962 8730
rect 9974 8678 10026 8730
rect 10038 8678 10090 8730
rect 10102 8678 10154 8730
rect 14294 8678 14346 8730
rect 14358 8678 14410 8730
rect 14422 8678 14474 8730
rect 14486 8678 14538 8730
rect 14550 8678 14602 8730
rect 2228 8576 2280 8628
rect 3424 8619 3476 8628
rect 3424 8585 3433 8619
rect 3433 8585 3467 8619
rect 3467 8585 3476 8619
rect 3424 8576 3476 8585
rect 4804 8619 4856 8628
rect 4804 8585 4813 8619
rect 4813 8585 4847 8619
rect 4847 8585 4856 8619
rect 4804 8576 4856 8585
rect 5908 8576 5960 8628
rect 6920 8576 6972 8628
rect 7104 8619 7156 8628
rect 7104 8585 7113 8619
rect 7113 8585 7147 8619
rect 7147 8585 7156 8619
rect 7104 8576 7156 8585
rect 8576 8576 8628 8628
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 12900 8619 12952 8628
rect 12900 8585 12909 8619
rect 12909 8585 12943 8619
rect 12943 8585 12952 8619
rect 12900 8576 12952 8585
rect 13728 8619 13780 8628
rect 13728 8585 13737 8619
rect 13737 8585 13771 8619
rect 13771 8585 13780 8619
rect 13728 8576 13780 8585
rect 15108 8619 15160 8628
rect 15108 8585 15117 8619
rect 15117 8585 15151 8619
rect 15151 8585 15160 8619
rect 15108 8576 15160 8585
rect 3056 8508 3108 8560
rect 4252 8508 4304 8560
rect 6736 8508 6788 8560
rect 8300 8508 8352 8560
rect 11336 8508 11388 8560
rect 13452 8508 13504 8560
rect 15568 8576 15620 8628
rect 16212 8576 16264 8628
rect 16488 8576 16540 8628
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 4988 8440 5040 8492
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 2780 8372 2832 8381
rect 3516 8372 3568 8424
rect 4252 8415 4304 8424
rect 4252 8381 4261 8415
rect 4261 8381 4295 8415
rect 4295 8381 4304 8415
rect 4252 8372 4304 8381
rect 1400 8347 1452 8356
rect 1400 8313 1409 8347
rect 1409 8313 1443 8347
rect 1443 8313 1452 8347
rect 1400 8304 1452 8313
rect 4068 8304 4120 8356
rect 6368 8372 6420 8424
rect 7472 8372 7524 8424
rect 6184 8304 6236 8356
rect 6920 8304 6972 8356
rect 8760 8440 8812 8492
rect 9864 8440 9916 8492
rect 10232 8440 10284 8492
rect 12532 8440 12584 8492
rect 12992 8440 13044 8492
rect 14832 8440 14884 8492
rect 15016 8483 15068 8492
rect 15016 8449 15025 8483
rect 15025 8449 15059 8483
rect 15059 8449 15068 8483
rect 15016 8440 15068 8449
rect 15108 8440 15160 8492
rect 16672 8483 16724 8492
rect 8116 8372 8168 8424
rect 9772 8372 9824 8424
rect 11336 8372 11388 8424
rect 12900 8372 12952 8424
rect 14924 8372 14976 8424
rect 16120 8415 16172 8424
rect 8484 8304 8536 8356
rect 1768 8236 1820 8288
rect 4620 8236 4672 8288
rect 5264 8236 5316 8288
rect 6368 8236 6420 8288
rect 8852 8236 8904 8288
rect 11152 8304 11204 8356
rect 15108 8304 15160 8356
rect 16120 8381 16129 8415
rect 16129 8381 16163 8415
rect 16163 8381 16172 8415
rect 16120 8372 16172 8381
rect 16672 8449 16681 8483
rect 16681 8449 16715 8483
rect 16715 8449 16724 8483
rect 16672 8440 16724 8449
rect 16304 8372 16356 8424
rect 17776 8440 17828 8492
rect 17960 8440 18012 8492
rect 15384 8304 15436 8356
rect 17960 8304 18012 8356
rect 18328 8347 18380 8356
rect 18328 8313 18337 8347
rect 18337 8313 18371 8347
rect 18371 8313 18380 8347
rect 18328 8304 18380 8313
rect 14556 8279 14608 8288
rect 14556 8245 14565 8279
rect 14565 8245 14599 8279
rect 14599 8245 14608 8279
rect 14556 8236 14608 8245
rect 14832 8236 14884 8288
rect 15292 8236 15344 8288
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 3430 8134 3482 8186
rect 7622 8134 7674 8186
rect 7686 8134 7738 8186
rect 7750 8134 7802 8186
rect 7814 8134 7866 8186
rect 7878 8134 7930 8186
rect 12070 8134 12122 8186
rect 12134 8134 12186 8186
rect 12198 8134 12250 8186
rect 12262 8134 12314 8186
rect 12326 8134 12378 8186
rect 16518 8134 16570 8186
rect 16582 8134 16634 8186
rect 16646 8134 16698 8186
rect 16710 8134 16762 8186
rect 16774 8134 16826 8186
rect 1584 8032 1636 8084
rect 4160 8075 4212 8084
rect 2136 7896 2188 7948
rect 4160 8041 4169 8075
rect 4169 8041 4203 8075
rect 4203 8041 4212 8075
rect 4160 8032 4212 8041
rect 3700 7964 3752 8016
rect 4896 8032 4948 8084
rect 6184 8032 6236 8084
rect 4988 8007 5040 8016
rect 4988 7973 4997 8007
rect 4997 7973 5031 8007
rect 5031 7973 5040 8007
rect 4988 7964 5040 7973
rect 3516 7939 3568 7948
rect 3516 7905 3525 7939
rect 3525 7905 3559 7939
rect 3559 7905 3568 7939
rect 3516 7896 3568 7905
rect 4804 7939 4856 7948
rect 4804 7905 4813 7939
rect 4813 7905 4847 7939
rect 4847 7905 4856 7939
rect 4804 7896 4856 7905
rect 2044 7828 2096 7880
rect 4436 7828 4488 7880
rect 5172 7896 5224 7948
rect 6460 8032 6512 8084
rect 6920 8032 6972 8084
rect 9220 7964 9272 8016
rect 7748 7939 7800 7948
rect 1216 7760 1268 7812
rect 6092 7803 6144 7812
rect 6092 7769 6110 7803
rect 6110 7769 6144 7803
rect 6092 7760 6144 7769
rect 6276 7828 6328 7880
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 8392 7939 8444 7948
rect 8392 7905 8401 7939
rect 8401 7905 8435 7939
rect 8435 7905 8444 7939
rect 8392 7896 8444 7905
rect 8576 7939 8628 7948
rect 8576 7905 8585 7939
rect 8585 7905 8619 7939
rect 8619 7905 8628 7939
rect 8576 7896 8628 7905
rect 12532 8075 12584 8084
rect 12532 8041 12541 8075
rect 12541 8041 12575 8075
rect 12575 8041 12584 8075
rect 12532 8032 12584 8041
rect 13176 8032 13228 8084
rect 13452 8032 13504 8084
rect 9864 7964 9916 8016
rect 9680 7939 9732 7948
rect 9680 7905 9689 7939
rect 9689 7905 9723 7939
rect 9723 7905 9732 7939
rect 9680 7896 9732 7905
rect 9404 7828 9456 7880
rect 10968 7896 11020 7948
rect 12440 7964 12492 8016
rect 11704 7939 11756 7948
rect 11704 7905 11713 7939
rect 11713 7905 11747 7939
rect 11747 7905 11756 7939
rect 11704 7896 11756 7905
rect 15384 7964 15436 8016
rect 11244 7828 11296 7880
rect 14556 7896 14608 7948
rect 14648 7896 14700 7948
rect 15936 7964 15988 8016
rect 16856 8032 16908 8084
rect 18052 8032 18104 8084
rect 17684 7964 17736 8016
rect 16304 7896 16356 7948
rect 16764 7896 16816 7948
rect 17224 7896 17276 7948
rect 17408 7896 17460 7948
rect 17592 7939 17644 7948
rect 17592 7905 17601 7939
rect 17601 7905 17635 7939
rect 17635 7905 17644 7939
rect 17592 7896 17644 7905
rect 9588 7760 9640 7812
rect 2136 7692 2188 7744
rect 3332 7735 3384 7744
rect 3332 7701 3341 7735
rect 3341 7701 3375 7735
rect 3375 7701 3384 7735
rect 3884 7735 3936 7744
rect 3332 7692 3384 7701
rect 3884 7701 3893 7735
rect 3893 7701 3927 7735
rect 3927 7701 3936 7735
rect 3884 7692 3936 7701
rect 4620 7735 4672 7744
rect 4620 7701 4629 7735
rect 4629 7701 4663 7735
rect 4663 7701 4672 7735
rect 4620 7692 4672 7701
rect 5908 7692 5960 7744
rect 7104 7735 7156 7744
rect 7104 7701 7113 7735
rect 7113 7701 7147 7735
rect 7147 7701 7156 7735
rect 7104 7692 7156 7701
rect 9680 7692 9732 7744
rect 10508 7735 10560 7744
rect 10508 7701 10517 7735
rect 10517 7701 10551 7735
rect 10551 7701 10560 7735
rect 10508 7692 10560 7701
rect 11612 7760 11664 7812
rect 17132 7828 17184 7880
rect 17960 7828 18012 7880
rect 16304 7760 16356 7812
rect 17868 7803 17920 7812
rect 17868 7769 17877 7803
rect 17877 7769 17911 7803
rect 17911 7769 17920 7803
rect 17868 7760 17920 7769
rect 12900 7692 12952 7744
rect 13452 7735 13504 7744
rect 13452 7701 13461 7735
rect 13461 7701 13495 7735
rect 13495 7701 13504 7735
rect 13452 7692 13504 7701
rect 13912 7735 13964 7744
rect 13912 7701 13921 7735
rect 13921 7701 13955 7735
rect 13955 7701 13964 7735
rect 13912 7692 13964 7701
rect 14188 7692 14240 7744
rect 14832 7735 14884 7744
rect 14832 7701 14841 7735
rect 14841 7701 14875 7735
rect 14875 7701 14884 7735
rect 14832 7692 14884 7701
rect 15292 7735 15344 7744
rect 15292 7701 15301 7735
rect 15301 7701 15335 7735
rect 15335 7701 15344 7735
rect 15292 7692 15344 7701
rect 15568 7692 15620 7744
rect 5398 7590 5450 7642
rect 5462 7590 5514 7642
rect 5526 7590 5578 7642
rect 5590 7590 5642 7642
rect 5654 7590 5706 7642
rect 9846 7590 9898 7642
rect 9910 7590 9962 7642
rect 9974 7590 10026 7642
rect 10038 7590 10090 7642
rect 10102 7590 10154 7642
rect 14294 7590 14346 7642
rect 14358 7590 14410 7642
rect 14422 7590 14474 7642
rect 14486 7590 14538 7642
rect 14550 7590 14602 7642
rect 1492 7531 1544 7540
rect 1492 7497 1501 7531
rect 1501 7497 1535 7531
rect 1535 7497 1544 7531
rect 1492 7488 1544 7497
rect 3056 7488 3108 7540
rect 5264 7488 5316 7540
rect 2780 7463 2832 7472
rect 2780 7429 2789 7463
rect 2789 7429 2823 7463
rect 2823 7429 2832 7463
rect 2780 7420 2832 7429
rect 5080 7420 5132 7472
rect 5172 7420 5224 7472
rect 5540 7420 5592 7472
rect 5632 7420 5684 7472
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 2320 7352 2372 7404
rect 4252 7352 4304 7404
rect 6184 7352 6236 7404
rect 6736 7352 6788 7404
rect 6920 7531 6972 7540
rect 6920 7497 6929 7531
rect 6929 7497 6963 7531
rect 6963 7497 6972 7531
rect 6920 7488 6972 7497
rect 13636 7531 13688 7540
rect 7748 7395 7800 7404
rect 7748 7361 7757 7395
rect 7757 7361 7791 7395
rect 7791 7361 7800 7395
rect 13636 7497 13645 7531
rect 13645 7497 13679 7531
rect 13679 7497 13688 7531
rect 13636 7488 13688 7497
rect 14188 7488 14240 7540
rect 16396 7488 16448 7540
rect 17500 7531 17552 7540
rect 17500 7497 17509 7531
rect 17509 7497 17543 7531
rect 17543 7497 17552 7531
rect 17500 7488 17552 7497
rect 18420 7531 18472 7540
rect 18420 7497 18429 7531
rect 18429 7497 18463 7531
rect 18463 7497 18472 7531
rect 18420 7488 18472 7497
rect 8576 7420 8628 7472
rect 11704 7420 11756 7472
rect 12532 7420 12584 7472
rect 13912 7420 13964 7472
rect 7748 7352 7800 7361
rect 9772 7352 9824 7404
rect 10048 7352 10100 7404
rect 12716 7395 12768 7404
rect 12716 7361 12725 7395
rect 12725 7361 12759 7395
rect 12759 7361 12768 7395
rect 12716 7352 12768 7361
rect 13820 7352 13872 7404
rect 14096 7352 14148 7404
rect 16856 7420 16908 7472
rect 16120 7352 16172 7404
rect 17132 7352 17184 7404
rect 17592 7352 17644 7404
rect 4712 7284 4764 7336
rect 3516 7216 3568 7268
rect 5264 7284 5316 7336
rect 6920 7284 6972 7336
rect 7472 7327 7524 7336
rect 7472 7293 7481 7327
rect 7481 7293 7515 7327
rect 7515 7293 7524 7327
rect 11612 7327 11664 7336
rect 7472 7284 7524 7293
rect 6092 7216 6144 7268
rect 6276 7216 6328 7268
rect 11612 7293 11621 7327
rect 11621 7293 11655 7327
rect 11655 7293 11664 7327
rect 11612 7284 11664 7293
rect 11796 7327 11848 7336
rect 11796 7293 11805 7327
rect 11805 7293 11839 7327
rect 11839 7293 11848 7327
rect 11796 7284 11848 7293
rect 12440 7284 12492 7336
rect 13728 7327 13780 7336
rect 13728 7293 13737 7327
rect 13737 7293 13771 7327
rect 13771 7293 13780 7327
rect 13728 7284 13780 7293
rect 14740 7327 14792 7336
rect 13084 7216 13136 7268
rect 14740 7293 14749 7327
rect 14749 7293 14783 7327
rect 14783 7293 14792 7327
rect 14740 7284 14792 7293
rect 14924 7327 14976 7336
rect 14924 7293 14933 7327
rect 14933 7293 14967 7327
rect 14967 7293 14976 7327
rect 14924 7284 14976 7293
rect 18420 7284 18472 7336
rect 2504 7191 2556 7200
rect 2504 7157 2513 7191
rect 2513 7157 2547 7191
rect 2547 7157 2556 7191
rect 2504 7148 2556 7157
rect 5172 7148 5224 7200
rect 6184 7191 6236 7200
rect 6184 7157 6193 7191
rect 6193 7157 6227 7191
rect 6227 7157 6236 7191
rect 6184 7148 6236 7157
rect 6460 7191 6512 7200
rect 6460 7157 6469 7191
rect 6469 7157 6503 7191
rect 6503 7157 6512 7191
rect 6460 7148 6512 7157
rect 6644 7148 6696 7200
rect 6920 7148 6972 7200
rect 8392 7191 8444 7200
rect 8392 7157 8401 7191
rect 8401 7157 8435 7191
rect 8435 7157 8444 7191
rect 8392 7148 8444 7157
rect 11980 7148 12032 7200
rect 17500 7148 17552 7200
rect 17868 7148 17920 7200
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 3430 7046 3482 7098
rect 7622 7046 7674 7098
rect 7686 7046 7738 7098
rect 7750 7046 7802 7098
rect 7814 7046 7866 7098
rect 7878 7046 7930 7098
rect 12070 7046 12122 7098
rect 12134 7046 12186 7098
rect 12198 7046 12250 7098
rect 12262 7046 12314 7098
rect 12326 7046 12378 7098
rect 16518 7046 16570 7098
rect 16582 7046 16634 7098
rect 16646 7046 16698 7098
rect 16710 7046 16762 7098
rect 16774 7046 16826 7098
rect 2320 6944 2372 6996
rect 6000 6944 6052 6996
rect 3148 6808 3200 6860
rect 4988 6808 5040 6860
rect 6184 6851 6236 6860
rect 1400 6672 1452 6724
rect 2780 6672 2832 6724
rect 3976 6740 4028 6792
rect 5632 6783 5684 6792
rect 5632 6749 5641 6783
rect 5641 6749 5675 6783
rect 5675 6749 5684 6783
rect 5632 6740 5684 6749
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 7288 6876 7340 6928
rect 8944 6876 8996 6928
rect 10048 6944 10100 6996
rect 10416 6944 10468 6996
rect 10968 6944 11020 6996
rect 11796 6944 11848 6996
rect 12716 6987 12768 6996
rect 12716 6953 12725 6987
rect 12725 6953 12759 6987
rect 12759 6953 12768 6987
rect 12716 6944 12768 6953
rect 12900 6944 12952 6996
rect 16856 6987 16908 6996
rect 9036 6851 9088 6860
rect 9036 6817 9045 6851
rect 9045 6817 9079 6851
rect 9079 6817 9088 6851
rect 9036 6808 9088 6817
rect 9496 6808 9548 6860
rect 11336 6851 11388 6860
rect 11336 6817 11345 6851
rect 11345 6817 11379 6851
rect 11379 6817 11388 6851
rect 11336 6808 11388 6817
rect 12440 6876 12492 6928
rect 12624 6919 12676 6928
rect 12624 6885 12633 6919
rect 12633 6885 12667 6919
rect 12667 6885 12676 6919
rect 12624 6876 12676 6885
rect 13452 6876 13504 6928
rect 16856 6953 16865 6987
rect 16865 6953 16899 6987
rect 16899 6953 16908 6987
rect 16856 6944 16908 6953
rect 17500 6944 17552 6996
rect 18236 6876 18288 6928
rect 13360 6851 13412 6860
rect 13360 6817 13369 6851
rect 13369 6817 13403 6851
rect 13403 6817 13412 6851
rect 13360 6808 13412 6817
rect 13728 6808 13780 6860
rect 16120 6851 16172 6860
rect 6920 6740 6972 6792
rect 7380 6740 7432 6792
rect 8024 6740 8076 6792
rect 8208 6740 8260 6792
rect 4160 6715 4212 6724
rect 4160 6681 4194 6715
rect 4194 6681 4212 6715
rect 4160 6672 4212 6681
rect 1308 6604 1360 6656
rect 2688 6604 2740 6656
rect 2964 6647 3016 6656
rect 2964 6613 2973 6647
rect 2973 6613 3007 6647
rect 3007 6613 3016 6647
rect 2964 6604 3016 6613
rect 3516 6604 3568 6656
rect 3884 6604 3936 6656
rect 4896 6604 4948 6656
rect 5540 6672 5592 6724
rect 11244 6740 11296 6792
rect 12532 6740 12584 6792
rect 13084 6783 13136 6792
rect 13084 6749 13093 6783
rect 13093 6749 13127 6783
rect 13127 6749 13136 6783
rect 13084 6740 13136 6749
rect 13544 6783 13596 6792
rect 13544 6749 13553 6783
rect 13553 6749 13587 6783
rect 13587 6749 13596 6783
rect 13544 6740 13596 6749
rect 13820 6783 13872 6792
rect 13820 6749 13829 6783
rect 13829 6749 13863 6783
rect 13863 6749 13872 6783
rect 13820 6740 13872 6749
rect 14096 6783 14148 6792
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 16120 6817 16129 6851
rect 16129 6817 16163 6851
rect 16163 6817 16172 6851
rect 16120 6808 16172 6817
rect 16212 6808 16264 6860
rect 15936 6783 15988 6792
rect 9128 6672 9180 6724
rect 6092 6647 6144 6656
rect 6092 6613 6101 6647
rect 6101 6613 6135 6647
rect 6135 6613 6144 6647
rect 6092 6604 6144 6613
rect 6184 6604 6236 6656
rect 6920 6647 6972 6656
rect 6920 6613 6929 6647
rect 6929 6613 6963 6647
rect 6963 6613 6972 6647
rect 6920 6604 6972 6613
rect 7380 6647 7432 6656
rect 7380 6613 7389 6647
rect 7389 6613 7423 6647
rect 7423 6613 7432 6647
rect 7380 6604 7432 6613
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 13360 6672 13412 6724
rect 13636 6672 13688 6724
rect 11428 6604 11480 6656
rect 11888 6647 11940 6656
rect 11888 6613 11897 6647
rect 11897 6613 11931 6647
rect 11931 6613 11940 6647
rect 11888 6604 11940 6613
rect 12164 6604 12216 6656
rect 13268 6604 13320 6656
rect 15936 6749 15945 6783
rect 15945 6749 15979 6783
rect 15979 6749 15988 6783
rect 17960 6808 18012 6860
rect 15936 6740 15988 6749
rect 17132 6740 17184 6792
rect 17592 6740 17644 6792
rect 14740 6672 14792 6724
rect 16304 6672 16356 6724
rect 17776 6672 17828 6724
rect 16120 6604 16172 6656
rect 17684 6647 17736 6656
rect 17684 6613 17693 6647
rect 17693 6613 17727 6647
rect 17727 6613 17736 6647
rect 17684 6604 17736 6613
rect 18144 6604 18196 6656
rect 5398 6502 5450 6554
rect 5462 6502 5514 6554
rect 5526 6502 5578 6554
rect 5590 6502 5642 6554
rect 5654 6502 5706 6554
rect 9846 6502 9898 6554
rect 9910 6502 9962 6554
rect 9974 6502 10026 6554
rect 10038 6502 10090 6554
rect 10102 6502 10154 6554
rect 14294 6502 14346 6554
rect 14358 6502 14410 6554
rect 14422 6502 14474 6554
rect 14486 6502 14538 6554
rect 14550 6502 14602 6554
rect 2688 6400 2740 6452
rect 4620 6443 4672 6452
rect 3608 6332 3660 6384
rect 1768 6264 1820 6316
rect 1952 6196 2004 6248
rect 4252 6264 4304 6316
rect 3148 6128 3200 6180
rect 2964 6060 3016 6112
rect 3516 6060 3568 6112
rect 3976 6060 4028 6112
rect 4620 6409 4629 6443
rect 4629 6409 4663 6443
rect 4663 6409 4672 6443
rect 4620 6400 4672 6409
rect 5816 6443 5868 6452
rect 5816 6409 5825 6443
rect 5825 6409 5859 6443
rect 5859 6409 5868 6443
rect 5816 6400 5868 6409
rect 6092 6400 6144 6452
rect 8116 6400 8168 6452
rect 8668 6443 8720 6452
rect 8668 6409 8677 6443
rect 8677 6409 8711 6443
rect 8711 6409 8720 6443
rect 8668 6400 8720 6409
rect 8760 6400 8812 6452
rect 11612 6400 11664 6452
rect 11888 6400 11940 6452
rect 12164 6400 12216 6452
rect 15476 6400 15528 6452
rect 5172 6332 5224 6384
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 4712 6264 4764 6316
rect 6920 6332 6972 6384
rect 7932 6332 7984 6384
rect 8576 6332 8628 6384
rect 6644 6307 6696 6316
rect 6644 6273 6678 6307
rect 6678 6273 6696 6307
rect 6644 6264 6696 6273
rect 7380 6264 7432 6316
rect 4988 6196 5040 6248
rect 6276 6196 6328 6248
rect 6184 6128 6236 6180
rect 4528 6060 4580 6112
rect 7472 6196 7524 6248
rect 8116 6196 8168 6248
rect 8944 6196 8996 6248
rect 9312 6239 9364 6248
rect 9312 6205 9321 6239
rect 9321 6205 9355 6239
rect 9355 6205 9364 6239
rect 9312 6196 9364 6205
rect 7380 6060 7432 6112
rect 7932 6128 7984 6180
rect 12532 6332 12584 6384
rect 13820 6332 13872 6384
rect 15844 6332 15896 6384
rect 16212 6400 16264 6452
rect 17684 6400 17736 6452
rect 17868 6400 17920 6452
rect 16856 6375 16908 6384
rect 11152 6264 11204 6316
rect 11336 6264 11388 6316
rect 11612 6264 11664 6316
rect 12348 6307 12400 6316
rect 12348 6273 12357 6307
rect 12357 6273 12391 6307
rect 12391 6273 12400 6307
rect 12348 6264 12400 6273
rect 13176 6307 13228 6316
rect 13176 6273 13185 6307
rect 13185 6273 13219 6307
rect 13219 6273 13228 6307
rect 13176 6264 13228 6273
rect 13360 6239 13412 6248
rect 13360 6205 13369 6239
rect 13369 6205 13403 6239
rect 13403 6205 13412 6239
rect 13360 6196 13412 6205
rect 13820 6196 13872 6248
rect 14648 6264 14700 6316
rect 15200 6264 15252 6316
rect 15936 6307 15988 6316
rect 9588 6103 9640 6112
rect 9588 6069 9597 6103
rect 9597 6069 9631 6103
rect 9631 6069 9640 6103
rect 9588 6060 9640 6069
rect 10232 6060 10284 6112
rect 13728 6128 13780 6180
rect 15936 6273 15945 6307
rect 15945 6273 15979 6307
rect 15979 6273 15988 6307
rect 15936 6264 15988 6273
rect 16856 6341 16865 6375
rect 16865 6341 16899 6375
rect 16899 6341 16908 6375
rect 16856 6332 16908 6341
rect 16396 6196 16448 6248
rect 15384 6128 15436 6180
rect 15936 6060 15988 6112
rect 17040 6264 17092 6316
rect 17592 6264 17644 6316
rect 17868 6307 17920 6316
rect 17868 6273 17877 6307
rect 17877 6273 17911 6307
rect 17911 6273 17920 6307
rect 17868 6264 17920 6273
rect 18144 6264 18196 6316
rect 16856 6196 16908 6248
rect 18420 6196 18472 6248
rect 18052 6171 18104 6180
rect 18052 6137 18061 6171
rect 18061 6137 18095 6171
rect 18095 6137 18104 6171
rect 18052 6128 18104 6137
rect 17132 6060 17184 6112
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 3430 5958 3482 6010
rect 7622 5958 7674 6010
rect 7686 5958 7738 6010
rect 7750 5958 7802 6010
rect 7814 5958 7866 6010
rect 7878 5958 7930 6010
rect 12070 5958 12122 6010
rect 12134 5958 12186 6010
rect 12198 5958 12250 6010
rect 12262 5958 12314 6010
rect 12326 5958 12378 6010
rect 16518 5958 16570 6010
rect 16582 5958 16634 6010
rect 16646 5958 16698 6010
rect 16710 5958 16762 6010
rect 16774 5958 16826 6010
rect 1860 5856 1912 5908
rect 2320 5856 2372 5908
rect 2596 5856 2648 5908
rect 6092 5856 6144 5908
rect 6920 5856 6972 5908
rect 7380 5856 7432 5908
rect 8208 5856 8260 5908
rect 4896 5788 4948 5840
rect 7472 5788 7524 5840
rect 3056 5720 3108 5772
rect 8852 5856 8904 5908
rect 11336 5856 11388 5908
rect 12624 5856 12676 5908
rect 3056 5584 3108 5636
rect 3700 5652 3752 5704
rect 4436 5652 4488 5704
rect 4988 5652 5040 5704
rect 5080 5652 5132 5704
rect 3976 5584 4028 5636
rect 4068 5627 4120 5636
rect 4068 5593 4077 5627
rect 4077 5593 4111 5627
rect 4111 5593 4120 5627
rect 4068 5584 4120 5593
rect 8392 5652 8444 5704
rect 11060 5652 11112 5704
rect 14096 5788 14148 5840
rect 17316 5899 17368 5908
rect 17316 5865 17325 5899
rect 17325 5865 17359 5899
rect 17359 5865 17368 5899
rect 17316 5856 17368 5865
rect 17960 5856 18012 5908
rect 2596 5516 2648 5568
rect 4712 5559 4764 5568
rect 4712 5525 4721 5559
rect 4721 5525 4755 5559
rect 4755 5525 4764 5559
rect 4712 5516 4764 5525
rect 6552 5516 6604 5568
rect 7472 5516 7524 5568
rect 9036 5584 9088 5636
rect 8576 5516 8628 5568
rect 8760 5559 8812 5568
rect 8760 5525 8769 5559
rect 8769 5525 8803 5559
rect 8803 5525 8812 5559
rect 8760 5516 8812 5525
rect 8944 5516 8996 5568
rect 11336 5584 11388 5636
rect 10968 5516 11020 5568
rect 13544 5652 13596 5704
rect 14372 5652 14424 5704
rect 14648 5763 14700 5772
rect 14648 5729 14657 5763
rect 14657 5729 14691 5763
rect 14691 5729 14700 5763
rect 14648 5720 14700 5729
rect 14740 5720 14792 5772
rect 16856 5788 16908 5840
rect 15200 5720 15252 5772
rect 14556 5652 14608 5704
rect 17316 5652 17368 5704
rect 18236 5695 18288 5704
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 14740 5584 14792 5636
rect 16304 5584 16356 5636
rect 13636 5559 13688 5568
rect 13636 5525 13645 5559
rect 13645 5525 13679 5559
rect 13679 5525 13688 5559
rect 13636 5516 13688 5525
rect 13912 5516 13964 5568
rect 14924 5516 14976 5568
rect 15292 5559 15344 5568
rect 15292 5525 15301 5559
rect 15301 5525 15335 5559
rect 15335 5525 15344 5559
rect 15292 5516 15344 5525
rect 15384 5559 15436 5568
rect 15384 5525 15393 5559
rect 15393 5525 15427 5559
rect 15427 5525 15436 5559
rect 15384 5516 15436 5525
rect 16672 5516 16724 5568
rect 17040 5516 17092 5568
rect 17868 5516 17920 5568
rect 18052 5559 18104 5568
rect 18052 5525 18061 5559
rect 18061 5525 18095 5559
rect 18095 5525 18104 5559
rect 18052 5516 18104 5525
rect 18420 5559 18472 5568
rect 18420 5525 18429 5559
rect 18429 5525 18463 5559
rect 18463 5525 18472 5559
rect 18420 5516 18472 5525
rect 112 5448 164 5500
rect 940 5448 992 5500
rect 5398 5414 5450 5466
rect 5462 5414 5514 5466
rect 5526 5414 5578 5466
rect 5590 5414 5642 5466
rect 5654 5414 5706 5466
rect 9846 5414 9898 5466
rect 9910 5414 9962 5466
rect 9974 5414 10026 5466
rect 10038 5414 10090 5466
rect 10102 5414 10154 5466
rect 14294 5414 14346 5466
rect 14358 5414 14410 5466
rect 14422 5414 14474 5466
rect 14486 5414 14538 5466
rect 14550 5414 14602 5466
rect 2228 5355 2280 5364
rect 2228 5321 2237 5355
rect 2237 5321 2271 5355
rect 2271 5321 2280 5355
rect 2228 5312 2280 5321
rect 4344 5312 4396 5364
rect 4804 5312 4856 5364
rect 2596 5287 2648 5296
rect 2596 5253 2605 5287
rect 2605 5253 2639 5287
rect 2639 5253 2648 5287
rect 2596 5244 2648 5253
rect 3884 5244 3936 5296
rect 2504 5176 2556 5228
rect 8668 5312 8720 5364
rect 9680 5312 9732 5364
rect 10692 5312 10744 5364
rect 13176 5312 13228 5364
rect 13268 5312 13320 5364
rect 8392 5244 8444 5296
rect 1584 5108 1636 5160
rect 4896 5151 4948 5160
rect 2872 5040 2924 5092
rect 2044 4972 2096 5024
rect 3976 4972 4028 5024
rect 4896 5117 4905 5151
rect 4905 5117 4939 5151
rect 4939 5117 4948 5151
rect 4896 5108 4948 5117
rect 5356 5176 5408 5228
rect 7196 5176 7248 5228
rect 10600 5244 10652 5296
rect 13728 5244 13780 5296
rect 6000 5151 6052 5160
rect 5172 5040 5224 5092
rect 6000 5117 6009 5151
rect 6009 5117 6043 5151
rect 6043 5117 6052 5151
rect 6000 5108 6052 5117
rect 7012 5108 7064 5160
rect 7472 5108 7524 5160
rect 9772 5176 9824 5228
rect 13360 5219 13412 5228
rect 13360 5185 13369 5219
rect 13369 5185 13403 5219
rect 13403 5185 13412 5219
rect 13360 5176 13412 5185
rect 13452 5219 13504 5228
rect 13452 5185 13461 5219
rect 13461 5185 13495 5219
rect 13495 5185 13504 5219
rect 15016 5312 15068 5364
rect 15292 5312 15344 5364
rect 16028 5355 16080 5364
rect 16028 5321 16037 5355
rect 16037 5321 16071 5355
rect 16071 5321 16080 5355
rect 16028 5312 16080 5321
rect 16304 5355 16356 5364
rect 16304 5321 16313 5355
rect 16313 5321 16347 5355
rect 16347 5321 16356 5355
rect 16304 5312 16356 5321
rect 16488 5355 16540 5364
rect 16488 5321 16497 5355
rect 16497 5321 16531 5355
rect 16531 5321 16540 5355
rect 16488 5312 16540 5321
rect 16672 5355 16724 5364
rect 16672 5321 16681 5355
rect 16681 5321 16715 5355
rect 16715 5321 16724 5355
rect 16672 5312 16724 5321
rect 16856 5355 16908 5364
rect 16856 5321 16865 5355
rect 16865 5321 16899 5355
rect 16899 5321 16908 5355
rect 16856 5312 16908 5321
rect 17684 5355 17736 5364
rect 17684 5321 17693 5355
rect 17693 5321 17727 5355
rect 17727 5321 17736 5355
rect 17684 5312 17736 5321
rect 18236 5312 18288 5364
rect 14648 5244 14700 5296
rect 15936 5287 15988 5296
rect 13452 5176 13504 5185
rect 14372 5219 14424 5228
rect 14372 5185 14406 5219
rect 14406 5185 14424 5219
rect 14372 5176 14424 5185
rect 8484 5151 8536 5160
rect 8116 5040 8168 5092
rect 8484 5117 8493 5151
rect 8493 5117 8527 5151
rect 8527 5117 8536 5151
rect 8484 5108 8536 5117
rect 9680 5108 9732 5160
rect 10232 5151 10284 5160
rect 10232 5117 10241 5151
rect 10241 5117 10275 5151
rect 10275 5117 10284 5151
rect 10232 5108 10284 5117
rect 10968 5151 11020 5160
rect 10968 5117 10977 5151
rect 10977 5117 11011 5151
rect 11011 5117 11020 5151
rect 11520 5151 11572 5160
rect 10968 5108 11020 5117
rect 11520 5117 11529 5151
rect 11529 5117 11563 5151
rect 11563 5117 11572 5151
rect 11520 5108 11572 5117
rect 13636 5151 13688 5160
rect 13636 5117 13645 5151
rect 13645 5117 13679 5151
rect 13679 5117 13688 5151
rect 13636 5108 13688 5117
rect 14096 5151 14148 5160
rect 14096 5117 14105 5151
rect 14105 5117 14139 5151
rect 14139 5117 14148 5151
rect 14096 5108 14148 5117
rect 10692 5040 10744 5092
rect 13084 5040 13136 5092
rect 13544 5040 13596 5092
rect 15936 5253 15945 5287
rect 15945 5253 15979 5287
rect 15979 5253 15988 5287
rect 15936 5244 15988 5253
rect 16212 5244 16264 5296
rect 17316 5244 17368 5296
rect 18144 5176 18196 5228
rect 4804 4972 4856 5024
rect 5264 4972 5316 5024
rect 9404 4972 9456 5024
rect 11244 4972 11296 5024
rect 11888 4972 11940 5024
rect 15384 4972 15436 5024
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 3430 4870 3482 4922
rect 7622 4870 7674 4922
rect 7686 4870 7738 4922
rect 7750 4870 7802 4922
rect 7814 4870 7866 4922
rect 7878 4870 7930 4922
rect 12070 4870 12122 4922
rect 12134 4870 12186 4922
rect 12198 4870 12250 4922
rect 12262 4870 12314 4922
rect 12326 4870 12378 4922
rect 16518 4870 16570 4922
rect 16582 4870 16634 4922
rect 16646 4870 16698 4922
rect 16710 4870 16762 4922
rect 16774 4870 16826 4922
rect 3884 4811 3936 4820
rect 3884 4777 3893 4811
rect 3893 4777 3927 4811
rect 3927 4777 3936 4811
rect 3884 4768 3936 4777
rect 7196 4768 7248 4820
rect 10692 4768 10744 4820
rect 11152 4768 11204 4820
rect 15384 4768 15436 4820
rect 16304 4768 16356 4820
rect 16948 4768 17000 4820
rect 10968 4700 11020 4752
rect 14924 4743 14976 4752
rect 1584 4675 1636 4684
rect 1584 4641 1593 4675
rect 1593 4641 1627 4675
rect 1627 4641 1636 4675
rect 1584 4632 1636 4641
rect 1676 4675 1728 4684
rect 1676 4641 1685 4675
rect 1685 4641 1719 4675
rect 1719 4641 1728 4675
rect 1676 4632 1728 4641
rect 2136 4632 2188 4684
rect 7380 4675 7432 4684
rect 7380 4641 7389 4675
rect 7389 4641 7423 4675
rect 7423 4641 7432 4675
rect 7380 4632 7432 4641
rect 11888 4632 11940 4684
rect 2228 4607 2280 4616
rect 2228 4573 2237 4607
rect 2237 4573 2271 4607
rect 2271 4573 2280 4607
rect 3976 4607 4028 4616
rect 2228 4564 2280 4573
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 4804 4564 4856 4616
rect 6552 4607 6604 4616
rect 6552 4573 6570 4607
rect 6570 4573 6604 4607
rect 6552 4564 6604 4573
rect 6736 4564 6788 4616
rect 8024 4564 8076 4616
rect 9036 4607 9088 4616
rect 9036 4573 9045 4607
rect 9045 4573 9079 4607
rect 9079 4573 9088 4607
rect 9036 4564 9088 4573
rect 9588 4564 9640 4616
rect 10232 4564 10284 4616
rect 10876 4564 10928 4616
rect 11520 4564 11572 4616
rect 14924 4709 14933 4743
rect 14933 4709 14967 4743
rect 14967 4709 14976 4743
rect 14924 4700 14976 4709
rect 15016 4700 15068 4752
rect 13084 4675 13136 4684
rect 13084 4641 13093 4675
rect 13093 4641 13127 4675
rect 13127 4641 13136 4675
rect 13084 4632 13136 4641
rect 14648 4675 14700 4684
rect 14648 4641 14657 4675
rect 14657 4641 14691 4675
rect 14691 4641 14700 4675
rect 14648 4632 14700 4641
rect 15200 4632 15252 4684
rect 15660 4700 15712 4752
rect 13820 4564 13872 4616
rect 15936 4564 15988 4616
rect 16396 4564 16448 4616
rect 2504 4539 2556 4548
rect 2504 4505 2538 4539
rect 2538 4505 2556 4539
rect 2504 4496 2556 4505
rect 4344 4496 4396 4548
rect 2136 4471 2188 4480
rect 2136 4437 2145 4471
rect 2145 4437 2179 4471
rect 2179 4437 2188 4471
rect 2136 4428 2188 4437
rect 3424 4428 3476 4480
rect 5080 4428 5132 4480
rect 6000 4428 6052 4480
rect 6828 4428 6880 4480
rect 7196 4428 7248 4480
rect 9312 4539 9364 4548
rect 9312 4505 9321 4539
rect 9321 4505 9355 4539
rect 9355 4505 9364 4539
rect 9312 4496 9364 4505
rect 11152 4496 11204 4548
rect 7472 4428 7524 4480
rect 8116 4428 8168 4480
rect 8668 4428 8720 4480
rect 9680 4428 9732 4480
rect 10324 4428 10376 4480
rect 11060 4471 11112 4480
rect 11060 4437 11069 4471
rect 11069 4437 11103 4471
rect 11103 4437 11112 4471
rect 11060 4428 11112 4437
rect 11980 4428 12032 4480
rect 12348 4428 12400 4480
rect 13912 4428 13964 4480
rect 14648 4496 14700 4548
rect 14832 4428 14884 4480
rect 15108 4428 15160 4480
rect 17132 4496 17184 4548
rect 17960 4496 18012 4548
rect 15384 4471 15436 4480
rect 15384 4437 15393 4471
rect 15393 4437 15427 4471
rect 15427 4437 15436 4471
rect 15384 4428 15436 4437
rect 15476 4428 15528 4480
rect 16856 4471 16908 4480
rect 16856 4437 16865 4471
rect 16865 4437 16899 4471
rect 16899 4437 16908 4471
rect 16856 4428 16908 4437
rect 17040 4471 17092 4480
rect 17040 4437 17049 4471
rect 17049 4437 17083 4471
rect 17083 4437 17092 4471
rect 17040 4428 17092 4437
rect 17868 4428 17920 4480
rect 18328 4471 18380 4480
rect 18328 4437 18337 4471
rect 18337 4437 18371 4471
rect 18371 4437 18380 4471
rect 18328 4428 18380 4437
rect 5398 4326 5450 4378
rect 5462 4326 5514 4378
rect 5526 4326 5578 4378
rect 5590 4326 5642 4378
rect 5654 4326 5706 4378
rect 9846 4326 9898 4378
rect 9910 4326 9962 4378
rect 9974 4326 10026 4378
rect 10038 4326 10090 4378
rect 10102 4326 10154 4378
rect 14294 4326 14346 4378
rect 14358 4326 14410 4378
rect 14422 4326 14474 4378
rect 14486 4326 14538 4378
rect 14550 4326 14602 4378
rect 2136 4267 2188 4276
rect 2136 4233 2145 4267
rect 2145 4233 2179 4267
rect 2179 4233 2188 4267
rect 2136 4224 2188 4233
rect 4344 4224 4396 4276
rect 4896 4224 4948 4276
rect 2044 4156 2096 4208
rect 3424 4156 3476 4208
rect 3700 4199 3752 4208
rect 3700 4165 3718 4199
rect 3718 4165 3752 4199
rect 3700 4156 3752 4165
rect 3884 4156 3936 4208
rect 8392 4267 8444 4276
rect 8392 4233 8401 4267
rect 8401 4233 8435 4267
rect 8435 4233 8444 4267
rect 8392 4224 8444 4233
rect 8760 4267 8812 4276
rect 8760 4233 8769 4267
rect 8769 4233 8803 4267
rect 8803 4233 8812 4267
rect 8760 4224 8812 4233
rect 11060 4224 11112 4276
rect 11152 4224 11204 4276
rect 13452 4267 13504 4276
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 14832 4224 14884 4276
rect 15660 4224 15712 4276
rect 16948 4267 17000 4276
rect 6368 4156 6420 4208
rect 7380 4156 7432 4208
rect 2136 4088 2188 4140
rect 3976 4063 4028 4072
rect 1492 3995 1544 4004
rect 1492 3961 1501 3995
rect 1501 3961 1535 3995
rect 1535 3961 1544 3995
rect 1492 3952 1544 3961
rect 1768 3995 1820 4004
rect 1768 3961 1777 3995
rect 1777 3961 1811 3995
rect 1811 3961 1820 3995
rect 1768 3952 1820 3961
rect 3976 4029 3985 4063
rect 3985 4029 4019 4063
rect 4019 4029 4028 4063
rect 3976 4020 4028 4029
rect 3608 3884 3660 3936
rect 4436 4088 4488 4140
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 4896 4088 4948 4097
rect 5448 4088 5500 4140
rect 10324 4156 10376 4208
rect 5908 4063 5960 4072
rect 5264 3952 5316 4004
rect 5908 4029 5917 4063
rect 5917 4029 5951 4063
rect 5951 4029 5960 4063
rect 5908 4020 5960 4029
rect 6552 4020 6604 4072
rect 8208 4131 8260 4140
rect 8208 4097 8217 4131
rect 8217 4097 8251 4131
rect 8251 4097 8260 4131
rect 8208 4088 8260 4097
rect 9496 4131 9548 4140
rect 9496 4097 9505 4131
rect 9505 4097 9539 4131
rect 9539 4097 9548 4131
rect 9496 4088 9548 4097
rect 8116 4020 8168 4072
rect 8576 4020 8628 4072
rect 10784 4088 10836 4140
rect 11980 4156 12032 4208
rect 13268 4131 13320 4140
rect 13268 4097 13277 4131
rect 13277 4097 13311 4131
rect 13311 4097 13320 4131
rect 13268 4088 13320 4097
rect 13452 4088 13504 4140
rect 14096 4156 14148 4208
rect 16948 4233 16957 4267
rect 16957 4233 16991 4267
rect 16991 4233 17000 4267
rect 16948 4224 17000 4233
rect 17316 4267 17368 4276
rect 17316 4233 17325 4267
rect 17325 4233 17359 4267
rect 17359 4233 17368 4267
rect 17316 4224 17368 4233
rect 17040 4156 17092 4208
rect 15384 4088 15436 4140
rect 16120 4131 16172 4140
rect 16120 4097 16129 4131
rect 16129 4097 16163 4131
rect 16163 4097 16172 4131
rect 16120 4088 16172 4097
rect 16304 4088 16356 4140
rect 10968 4063 11020 4072
rect 6736 3952 6788 4004
rect 8392 3952 8444 4004
rect 8668 3952 8720 4004
rect 9220 3952 9272 4004
rect 10968 4029 10977 4063
rect 10977 4029 11011 4063
rect 11011 4029 11020 4063
rect 10968 4020 11020 4029
rect 11520 4063 11572 4072
rect 10876 3952 10928 4004
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 13544 4020 13596 4072
rect 15568 4063 15620 4072
rect 15568 4029 15577 4063
rect 15577 4029 15611 4063
rect 15611 4029 15620 4063
rect 15568 4020 15620 4029
rect 15936 4063 15988 4072
rect 7196 3884 7248 3936
rect 9680 3927 9732 3936
rect 9680 3893 9689 3927
rect 9689 3893 9723 3927
rect 9723 3893 9732 3927
rect 9680 3884 9732 3893
rect 10324 3884 10376 3936
rect 13820 3884 13872 3936
rect 14280 3884 14332 3936
rect 15200 3952 15252 4004
rect 15936 4029 15945 4063
rect 15945 4029 15979 4063
rect 15979 4029 15988 4063
rect 15936 4020 15988 4029
rect 16856 4020 16908 4072
rect 16948 4020 17000 4072
rect 16028 3952 16080 4004
rect 17500 3927 17552 3936
rect 17500 3893 17509 3927
rect 17509 3893 17543 3927
rect 17543 3893 17552 3927
rect 17500 3884 17552 3893
rect 18236 3927 18288 3936
rect 18236 3893 18245 3927
rect 18245 3893 18279 3927
rect 18279 3893 18288 3927
rect 18236 3884 18288 3893
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 3430 3782 3482 3834
rect 7622 3782 7674 3834
rect 7686 3782 7738 3834
rect 7750 3782 7802 3834
rect 7814 3782 7866 3834
rect 7878 3782 7930 3834
rect 12070 3782 12122 3834
rect 12134 3782 12186 3834
rect 12198 3782 12250 3834
rect 12262 3782 12314 3834
rect 12326 3782 12378 3834
rect 16518 3782 16570 3834
rect 16582 3782 16634 3834
rect 16646 3782 16698 3834
rect 16710 3782 16762 3834
rect 16774 3782 16826 3834
rect 4160 3680 4212 3732
rect 4620 3723 4672 3732
rect 4620 3689 4629 3723
rect 4629 3689 4663 3723
rect 4663 3689 4672 3723
rect 4620 3680 4672 3689
rect 2504 3612 2556 3664
rect 4436 3612 4488 3664
rect 4712 3612 4764 3664
rect 3976 3587 4028 3596
rect 3976 3553 3985 3587
rect 3985 3553 4019 3587
rect 4019 3553 4028 3587
rect 3976 3544 4028 3553
rect 4252 3544 4304 3596
rect 5448 3680 5500 3732
rect 9036 3680 9088 3732
rect 9588 3680 9640 3732
rect 9864 3680 9916 3732
rect 10692 3680 10744 3732
rect 10968 3680 11020 3732
rect 13544 3680 13596 3732
rect 13912 3723 13964 3732
rect 13912 3689 13921 3723
rect 13921 3689 13955 3723
rect 13955 3689 13964 3723
rect 13912 3680 13964 3689
rect 14648 3680 14700 3732
rect 15384 3680 15436 3732
rect 15660 3723 15712 3732
rect 15660 3689 15669 3723
rect 15669 3689 15703 3723
rect 15703 3689 15712 3723
rect 15844 3723 15896 3732
rect 15660 3680 15712 3689
rect 15844 3689 15853 3723
rect 15853 3689 15887 3723
rect 15887 3689 15896 3723
rect 15844 3680 15896 3689
rect 16304 3680 16356 3732
rect 17040 3680 17092 3732
rect 17316 3680 17368 3732
rect 6644 3612 6696 3664
rect 5264 3587 5316 3596
rect 5264 3553 5273 3587
rect 5273 3553 5307 3587
rect 5307 3553 5316 3587
rect 5264 3544 5316 3553
rect 7288 3544 7340 3596
rect 2228 3476 2280 3528
rect 2964 3519 3016 3528
rect 2964 3485 2973 3519
rect 2973 3485 3007 3519
rect 3007 3485 3016 3519
rect 2964 3476 3016 3485
rect 5724 3476 5776 3528
rect 9404 3587 9456 3596
rect 9404 3553 9413 3587
rect 9413 3553 9447 3587
rect 9447 3553 9456 3587
rect 9404 3544 9456 3553
rect 10324 3544 10376 3596
rect 9680 3476 9732 3528
rect 10416 3519 10468 3528
rect 10416 3485 10425 3519
rect 10425 3485 10459 3519
rect 10459 3485 10468 3519
rect 10416 3476 10468 3485
rect 11888 3612 11940 3664
rect 16212 3655 16264 3664
rect 10876 3544 10928 3596
rect 11060 3544 11112 3596
rect 11520 3544 11572 3596
rect 11612 3476 11664 3528
rect 12072 3476 12124 3528
rect 13360 3544 13412 3596
rect 14280 3587 14332 3596
rect 14280 3553 14289 3587
rect 14289 3553 14323 3587
rect 14323 3553 14332 3587
rect 14280 3544 14332 3553
rect 16212 3621 16221 3655
rect 16221 3621 16255 3655
rect 16255 3621 16264 3655
rect 16212 3612 16264 3621
rect 18144 3612 18196 3664
rect 18420 3655 18472 3664
rect 18420 3621 18429 3655
rect 18429 3621 18463 3655
rect 18463 3621 18472 3655
rect 18420 3612 18472 3621
rect 16028 3587 16080 3596
rect 16028 3553 16037 3587
rect 16037 3553 16071 3587
rect 16071 3553 16080 3587
rect 16028 3544 16080 3553
rect 13452 3476 13504 3528
rect 13728 3519 13780 3528
rect 13728 3485 13737 3519
rect 13737 3485 13771 3519
rect 13771 3485 13780 3519
rect 13728 3476 13780 3485
rect 13912 3476 13964 3528
rect 14096 3476 14148 3528
rect 1860 3408 1912 3460
rect 3700 3408 3752 3460
rect 4160 3383 4212 3392
rect 4160 3349 4169 3383
rect 4169 3349 4203 3383
rect 4203 3349 4212 3383
rect 4160 3340 4212 3349
rect 4436 3408 4488 3460
rect 7380 3408 7432 3460
rect 11060 3408 11112 3460
rect 11428 3408 11480 3460
rect 11520 3408 11572 3460
rect 11704 3408 11756 3460
rect 15476 3408 15528 3460
rect 16948 3544 17000 3596
rect 6184 3383 6236 3392
rect 6184 3349 6193 3383
rect 6193 3349 6227 3383
rect 6227 3349 6236 3383
rect 6184 3340 6236 3349
rect 7196 3340 7248 3392
rect 8024 3340 8076 3392
rect 8392 3383 8444 3392
rect 8392 3349 8401 3383
rect 8401 3349 8435 3383
rect 8435 3349 8444 3383
rect 11336 3383 11388 3392
rect 8392 3340 8444 3349
rect 11336 3349 11345 3383
rect 11345 3349 11379 3383
rect 11379 3349 11388 3383
rect 11336 3340 11388 3349
rect 13912 3340 13964 3392
rect 14004 3340 14056 3392
rect 16212 3340 16264 3392
rect 17500 3519 17552 3528
rect 17500 3485 17509 3519
rect 17509 3485 17543 3519
rect 17543 3485 17552 3519
rect 17500 3476 17552 3485
rect 18236 3519 18288 3528
rect 18236 3485 18245 3519
rect 18245 3485 18279 3519
rect 18279 3485 18288 3519
rect 18236 3476 18288 3485
rect 16580 3451 16632 3460
rect 16580 3417 16589 3451
rect 16589 3417 16623 3451
rect 16623 3417 16632 3451
rect 16948 3451 17000 3460
rect 16580 3408 16632 3417
rect 16948 3417 16957 3451
rect 16957 3417 16991 3451
rect 16991 3417 17000 3451
rect 16948 3408 17000 3417
rect 19432 3408 19484 3460
rect 18052 3383 18104 3392
rect 18052 3349 18061 3383
rect 18061 3349 18095 3383
rect 18095 3349 18104 3383
rect 18052 3340 18104 3349
rect 5398 3238 5450 3290
rect 5462 3238 5514 3290
rect 5526 3238 5578 3290
rect 5590 3238 5642 3290
rect 5654 3238 5706 3290
rect 9846 3238 9898 3290
rect 9910 3238 9962 3290
rect 9974 3238 10026 3290
rect 10038 3238 10090 3290
rect 10102 3238 10154 3290
rect 14294 3238 14346 3290
rect 14358 3238 14410 3290
rect 14422 3238 14474 3290
rect 14486 3238 14538 3290
rect 14550 3238 14602 3290
rect 1400 3136 1452 3188
rect 2136 3136 2188 3188
rect 2964 3136 3016 3188
rect 3516 3136 3568 3188
rect 1676 3043 1728 3052
rect 1676 3009 1685 3043
rect 1685 3009 1719 3043
rect 1719 3009 1728 3043
rect 1676 3000 1728 3009
rect 2136 3043 2188 3052
rect 2136 3009 2145 3043
rect 2145 3009 2179 3043
rect 2179 3009 2188 3043
rect 2136 3000 2188 3009
rect 2872 3068 2924 3120
rect 4620 3136 4672 3188
rect 5080 3136 5132 3188
rect 5908 3136 5960 3188
rect 7380 3136 7432 3188
rect 6184 3068 6236 3120
rect 4620 3000 4672 3052
rect 3792 2932 3844 2984
rect 4620 2864 4672 2916
rect 3516 2796 3568 2848
rect 4436 2796 4488 2848
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 5080 3043 5132 3052
rect 4804 3000 4856 3009
rect 5080 3009 5114 3043
rect 5114 3009 5132 3043
rect 5080 3000 5132 3009
rect 5540 3000 5592 3052
rect 6460 3000 6512 3052
rect 7104 3000 7156 3052
rect 7380 3043 7432 3052
rect 7380 3009 7389 3043
rect 7389 3009 7423 3043
rect 7423 3009 7432 3043
rect 7380 3000 7432 3009
rect 7656 3000 7708 3052
rect 7564 2975 7616 2984
rect 7564 2941 7573 2975
rect 7573 2941 7607 2975
rect 7607 2941 7616 2975
rect 10508 3136 10560 3188
rect 10600 3136 10652 3188
rect 12072 3136 12124 3188
rect 13452 3179 13504 3188
rect 10324 3068 10376 3120
rect 9680 3000 9732 3052
rect 10416 3000 10468 3052
rect 10968 3000 11020 3052
rect 7564 2932 7616 2941
rect 8484 2864 8536 2916
rect 11520 3000 11572 3052
rect 11888 3043 11940 3052
rect 11888 3009 11897 3043
rect 11897 3009 11931 3043
rect 11931 3009 11940 3043
rect 11888 3000 11940 3009
rect 12348 3043 12400 3052
rect 12348 3009 12357 3043
rect 12357 3009 12391 3043
rect 12391 3009 12400 3043
rect 12348 3000 12400 3009
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 13912 3136 13964 3188
rect 14004 3068 14056 3120
rect 14188 3068 14240 3120
rect 15660 3068 15712 3120
rect 16120 3068 16172 3120
rect 16304 3068 16356 3120
rect 11336 2932 11388 2984
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 15292 3000 15344 3052
rect 15752 3000 15804 3052
rect 17040 3000 17092 3052
rect 15200 2932 15252 2984
rect 14740 2864 14792 2916
rect 14832 2864 14884 2916
rect 16028 2932 16080 2984
rect 17316 3000 17368 3052
rect 18328 3000 18380 3052
rect 5540 2796 5592 2848
rect 6184 2839 6236 2848
rect 6184 2805 6193 2839
rect 6193 2805 6227 2839
rect 6227 2805 6236 2839
rect 6184 2796 6236 2805
rect 6368 2796 6420 2848
rect 6920 2796 6972 2848
rect 7104 2796 7156 2848
rect 7288 2796 7340 2848
rect 8760 2796 8812 2848
rect 9220 2796 9272 2848
rect 11060 2796 11112 2848
rect 12440 2796 12492 2848
rect 13728 2796 13780 2848
rect 16304 2864 16356 2916
rect 16580 2864 16632 2916
rect 16764 2907 16816 2916
rect 16764 2873 16773 2907
rect 16773 2873 16807 2907
rect 16807 2873 16816 2907
rect 16764 2864 16816 2873
rect 15752 2796 15804 2848
rect 18696 2864 18748 2916
rect 17316 2839 17368 2848
rect 17316 2805 17325 2839
rect 17325 2805 17359 2839
rect 17359 2805 17368 2839
rect 17316 2796 17368 2805
rect 17684 2839 17736 2848
rect 17684 2805 17693 2839
rect 17693 2805 17727 2839
rect 17727 2805 17736 2839
rect 17684 2796 17736 2805
rect 18052 2839 18104 2848
rect 18052 2805 18061 2839
rect 18061 2805 18095 2839
rect 18095 2805 18104 2839
rect 18052 2796 18104 2805
rect 18880 2796 18932 2848
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 3430 2694 3482 2746
rect 7622 2694 7674 2746
rect 7686 2694 7738 2746
rect 7750 2694 7802 2746
rect 7814 2694 7866 2746
rect 7878 2694 7930 2746
rect 12070 2694 12122 2746
rect 12134 2694 12186 2746
rect 12198 2694 12250 2746
rect 12262 2694 12314 2746
rect 12326 2694 12378 2746
rect 16518 2694 16570 2746
rect 16582 2694 16634 2746
rect 16646 2694 16698 2746
rect 16710 2694 16762 2746
rect 16774 2694 16826 2746
rect 2136 2592 2188 2644
rect 3792 2592 3844 2644
rect 4988 2592 5040 2644
rect 6276 2592 6328 2644
rect 4896 2524 4948 2576
rect 2320 2499 2372 2508
rect 2320 2465 2329 2499
rect 2329 2465 2363 2499
rect 2363 2465 2372 2499
rect 2320 2456 2372 2465
rect 2964 2456 3016 2508
rect 2228 2388 2280 2440
rect 2412 2431 2464 2440
rect 2412 2397 2421 2431
rect 2421 2397 2455 2431
rect 2455 2397 2464 2431
rect 2412 2388 2464 2397
rect 3884 2456 3936 2508
rect 4344 2499 4396 2508
rect 4344 2465 4353 2499
rect 4353 2465 4387 2499
rect 4387 2465 4396 2499
rect 4344 2456 4396 2465
rect 4252 2388 4304 2440
rect 7104 2499 7156 2508
rect 7104 2465 7113 2499
rect 7113 2465 7147 2499
rect 7147 2465 7156 2499
rect 7104 2456 7156 2465
rect 7472 2456 7524 2508
rect 8300 2456 8352 2508
rect 10232 2592 10284 2644
rect 11336 2592 11388 2644
rect 11888 2592 11940 2644
rect 11980 2592 12032 2644
rect 12992 2567 13044 2576
rect 5724 2388 5776 2440
rect 6920 2431 6972 2440
rect 2872 2252 2924 2304
rect 3516 2252 3568 2304
rect 6920 2397 6929 2431
rect 6929 2397 6963 2431
rect 6963 2397 6972 2431
rect 6920 2388 6972 2397
rect 8760 2431 8812 2440
rect 8760 2397 8769 2431
rect 8769 2397 8803 2431
rect 8803 2397 8812 2431
rect 8760 2388 8812 2397
rect 9220 2499 9272 2508
rect 9220 2465 9229 2499
rect 9229 2465 9263 2499
rect 9263 2465 9272 2499
rect 9220 2456 9272 2465
rect 9680 2388 9732 2440
rect 9956 2499 10008 2508
rect 9956 2465 9965 2499
rect 9965 2465 9999 2499
rect 9999 2465 10008 2499
rect 9956 2456 10008 2465
rect 11060 2456 11112 2508
rect 11152 2499 11204 2508
rect 11152 2465 11161 2499
rect 11161 2465 11195 2499
rect 11195 2465 11204 2499
rect 11152 2456 11204 2465
rect 11520 2456 11572 2508
rect 12992 2533 13001 2567
rect 13001 2533 13035 2567
rect 13035 2533 13044 2567
rect 12992 2524 13044 2533
rect 14004 2592 14056 2644
rect 14740 2592 14792 2644
rect 16304 2592 16356 2644
rect 17224 2592 17276 2644
rect 14924 2524 14976 2576
rect 15016 2524 15068 2576
rect 4712 2252 4764 2304
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 4988 2252 5040 2304
rect 5908 2252 5960 2304
rect 6920 2252 6972 2304
rect 7472 2295 7524 2304
rect 7472 2261 7481 2295
rect 7481 2261 7515 2295
rect 7515 2261 7524 2295
rect 7472 2252 7524 2261
rect 11428 2388 11480 2440
rect 12348 2431 12400 2440
rect 12348 2397 12357 2431
rect 12357 2397 12391 2431
rect 12391 2397 12400 2431
rect 12348 2388 12400 2397
rect 14096 2456 14148 2508
rect 16672 2524 16724 2576
rect 18236 2524 18288 2576
rect 14648 2388 14700 2440
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 15108 2388 15160 2440
rect 15476 2431 15528 2440
rect 15476 2397 15485 2431
rect 15485 2397 15519 2431
rect 15519 2397 15528 2431
rect 15476 2388 15528 2397
rect 17960 2388 18012 2440
rect 14096 2320 14148 2372
rect 10968 2295 11020 2304
rect 10968 2261 10977 2295
rect 10977 2261 11011 2295
rect 11011 2261 11020 2295
rect 10968 2252 11020 2261
rect 11612 2252 11664 2304
rect 12440 2252 12492 2304
rect 13728 2295 13780 2304
rect 13728 2261 13737 2295
rect 13737 2261 13771 2295
rect 13771 2261 13780 2295
rect 13728 2252 13780 2261
rect 14740 2252 14792 2304
rect 15568 2252 15620 2304
rect 16120 2252 16172 2304
rect 16672 2295 16724 2304
rect 16672 2261 16681 2295
rect 16681 2261 16715 2295
rect 16715 2261 16724 2295
rect 16672 2252 16724 2261
rect 17040 2295 17092 2304
rect 17040 2261 17049 2295
rect 17049 2261 17083 2295
rect 17083 2261 17092 2295
rect 17040 2252 17092 2261
rect 17224 2295 17276 2304
rect 17224 2261 17233 2295
rect 17233 2261 17267 2295
rect 17267 2261 17276 2295
rect 17224 2252 17276 2261
rect 17868 2295 17920 2304
rect 17868 2261 17877 2295
rect 17877 2261 17911 2295
rect 17911 2261 17920 2295
rect 17868 2252 17920 2261
rect 18236 2295 18288 2304
rect 18236 2261 18245 2295
rect 18245 2261 18279 2295
rect 18279 2261 18288 2295
rect 18236 2252 18288 2261
rect 5398 2150 5450 2202
rect 5462 2150 5514 2202
rect 5526 2150 5578 2202
rect 5590 2150 5642 2202
rect 5654 2150 5706 2202
rect 9846 2150 9898 2202
rect 9910 2150 9962 2202
rect 9974 2150 10026 2202
rect 10038 2150 10090 2202
rect 10102 2150 10154 2202
rect 14294 2150 14346 2202
rect 14358 2150 14410 2202
rect 14422 2150 14474 2202
rect 14486 2150 14538 2202
rect 14550 2150 14602 2202
rect 4804 2048 4856 2100
rect 9128 2048 9180 2100
rect 6184 1980 6236 2032
rect 11152 2048 11204 2100
rect 11336 2048 11388 2100
rect 13728 2048 13780 2100
rect 14740 2048 14792 2100
rect 16120 2048 16172 2100
rect 10416 1980 10468 2032
rect 13636 1980 13688 2032
rect 17224 1980 17276 2032
rect 6000 1912 6052 1964
rect 12348 1912 12400 1964
rect 14648 1912 14700 1964
rect 17040 1912 17092 1964
rect 17500 1912 17552 1964
rect 4068 1844 4120 1896
rect 6828 1844 6880 1896
rect 8116 1844 8168 1896
rect 11336 1844 11388 1896
rect 12164 1844 12216 1896
rect 14096 1844 14148 1896
rect 5724 1776 5776 1828
rect 10600 1776 10652 1828
rect 11428 1776 11480 1828
rect 16672 1776 16724 1828
rect 5080 1708 5132 1760
rect 9772 1708 9824 1760
rect 3884 1640 3936 1692
rect 7472 1640 7524 1692
rect 13084 1504 13136 1556
rect 15200 1504 15252 1556
rect 3332 1436 3384 1488
rect 7196 1436 7248 1488
rect 3700 1232 3752 1284
rect 5816 1232 5868 1284
rect 11244 1164 11296 1216
rect 15016 1164 15068 1216
rect 4068 1028 4120 1080
rect 11796 1028 11848 1080
<< metal2 >>
rect 1122 16400 1178 17200
rect 3330 16538 3386 17200
rect 3698 16824 3754 16833
rect 3698 16759 3754 16768
rect 3330 16510 3648 16538
rect 3330 16400 3386 16510
rect 3514 16416 3570 16425
rect 1136 14414 1164 16400
rect 3514 16351 3570 16360
rect 3528 15230 3556 16351
rect 3516 15224 3568 15230
rect 1582 15192 1638 15201
rect 3516 15166 3568 15172
rect 1582 15127 1638 15136
rect 1124 14408 1176 14414
rect 1124 14350 1176 14356
rect 1596 12986 1624 15127
rect 2778 14784 2834 14793
rect 2778 14719 2834 14728
rect 2136 14000 2188 14006
rect 2136 13942 2188 13948
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1596 12481 1624 12922
rect 1964 12646 1992 13126
rect 2148 12646 2176 13942
rect 2792 12866 2820 14719
rect 3174 14716 3482 14736
rect 3174 14714 3180 14716
rect 3236 14714 3260 14716
rect 3316 14714 3340 14716
rect 3396 14714 3420 14716
rect 3476 14714 3482 14716
rect 3236 14662 3238 14714
rect 3418 14662 3420 14714
rect 3174 14660 3180 14662
rect 3236 14660 3260 14662
rect 3316 14660 3340 14662
rect 3396 14660 3420 14662
rect 3476 14660 3482 14662
rect 3174 14640 3482 14660
rect 3174 13628 3482 13648
rect 3174 13626 3180 13628
rect 3236 13626 3260 13628
rect 3316 13626 3340 13628
rect 3396 13626 3420 13628
rect 3476 13626 3482 13628
rect 3236 13574 3238 13626
rect 3418 13574 3420 13626
rect 3174 13572 3180 13574
rect 3236 13572 3260 13574
rect 3316 13572 3340 13574
rect 3396 13572 3420 13574
rect 3476 13572 3482 13574
rect 3174 13552 3482 13572
rect 3620 13297 3648 16510
rect 3712 15434 3740 16759
rect 5538 16400 5594 17200
rect 7746 16538 7802 17200
rect 9954 16538 10010 17200
rect 7746 16510 8064 16538
rect 7746 16400 7802 16510
rect 4066 16008 4122 16017
rect 4122 15966 4200 15994
rect 4066 15943 4122 15952
rect 3974 15600 4030 15609
rect 3974 15535 4030 15544
rect 3700 15428 3752 15434
rect 3700 15370 3752 15376
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3804 13977 3832 14418
rect 3884 14068 3936 14074
rect 3884 14010 3936 14016
rect 3790 13968 3846 13977
rect 3790 13903 3846 13912
rect 3896 13530 3924 14010
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3606 13288 3662 13297
rect 3606 13223 3662 13232
rect 3896 13190 3924 13466
rect 3988 13462 4016 15535
rect 4172 14634 4200 15966
rect 4172 14606 4384 14634
rect 4066 14376 4122 14385
rect 4066 14311 4122 14320
rect 4080 14278 4108 14311
rect 4068 14272 4120 14278
rect 4068 14214 4120 14220
rect 3976 13456 4028 13462
rect 3976 13398 4028 13404
rect 4066 13424 4122 13433
rect 4122 13382 4292 13410
rect 4066 13359 4122 13368
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 2700 12838 2820 12866
rect 3884 12912 3936 12918
rect 3884 12854 3936 12860
rect 1952 12640 2004 12646
rect 1872 12588 1952 12594
rect 2136 12640 2188 12646
rect 1872 12582 2004 12588
rect 2134 12608 2136 12617
rect 2188 12608 2190 12617
rect 1872 12566 1992 12582
rect 1582 12472 1638 12481
rect 1582 12407 1638 12416
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 112 10192 164 10198
rect 112 10134 164 10140
rect 124 5506 152 10134
rect 1504 9382 1532 12038
rect 1676 11824 1728 11830
rect 1676 11766 1728 11772
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1596 10470 1624 11698
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1308 9376 1360 9382
rect 1306 9344 1308 9353
rect 1492 9376 1544 9382
rect 1360 9344 1362 9353
rect 1492 9318 1544 9324
rect 1306 9279 1362 9288
rect 1216 7812 1268 7818
rect 1216 7754 1268 7760
rect 112 5500 164 5506
rect 112 5442 164 5448
rect 940 5500 992 5506
rect 940 5442 992 5448
rect 952 5137 980 5442
rect 938 5128 994 5137
rect 938 5063 994 5072
rect 938 2952 994 2961
rect 768 2910 938 2938
rect 400 870 520 898
rect 400 800 428 870
rect 386 0 442 800
rect 492 762 520 870
rect 768 762 796 2910
rect 938 2887 994 2896
rect 1228 800 1256 7754
rect 1320 6662 1348 9279
rect 1490 8528 1546 8537
rect 1490 8463 1546 8472
rect 1400 8356 1452 8362
rect 1400 8298 1452 8304
rect 1412 6730 1440 8298
rect 1504 7546 1532 8463
rect 1596 8090 1624 10406
rect 1688 9722 1716 11766
rect 1780 10849 1808 12038
rect 1766 10840 1822 10849
rect 1766 10775 1822 10784
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1676 9376 1728 9382
rect 1676 9318 1728 9324
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1688 7721 1716 9318
rect 1768 8288 1820 8294
rect 1768 8230 1820 8236
rect 1674 7712 1730 7721
rect 1674 7647 1730 7656
rect 1492 7540 1544 7546
rect 1492 7482 1544 7488
rect 1674 7440 1730 7449
rect 1674 7375 1676 7384
rect 1728 7375 1730 7384
rect 1676 7346 1728 7352
rect 1400 6724 1452 6730
rect 1400 6666 1452 6672
rect 1308 6656 1360 6662
rect 1308 6598 1360 6604
rect 1412 6610 1440 6666
rect 1412 6582 1624 6610
rect 1490 6488 1546 6497
rect 1490 6423 1546 6432
rect 1398 6080 1454 6089
rect 1398 6015 1454 6024
rect 1412 3194 1440 6015
rect 1504 4010 1532 6423
rect 1596 5166 1624 6582
rect 1780 6440 1808 8230
rect 1872 7721 1900 12566
rect 2134 12543 2190 12552
rect 2320 12232 2372 12238
rect 2320 12174 2372 12180
rect 2044 12164 2096 12170
rect 2044 12106 2096 12112
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1964 11830 1992 12038
rect 1952 11824 2004 11830
rect 1952 11766 2004 11772
rect 2056 11558 2084 12106
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 2056 11354 2084 11494
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 1952 11076 2004 11082
rect 1952 11018 2004 11024
rect 1964 9382 1992 11018
rect 2056 9761 2084 11290
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 2042 9752 2098 9761
rect 2042 9687 2098 9696
rect 1952 9376 2004 9382
rect 1952 9318 2004 9324
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 2056 7886 2084 8774
rect 2148 7954 2176 9862
rect 2240 9586 2268 11630
rect 2332 11393 2360 12174
rect 2596 12164 2648 12170
rect 2596 12106 2648 12112
rect 2504 11552 2556 11558
rect 2504 11494 2556 11500
rect 2318 11384 2374 11393
rect 2318 11319 2374 11328
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2136 7744 2188 7750
rect 1858 7712 1914 7721
rect 2136 7686 2188 7692
rect 1858 7647 1914 7656
rect 1688 6412 1808 6440
rect 1584 5160 1636 5166
rect 1584 5102 1636 5108
rect 1596 4690 1624 5102
rect 1688 4690 1716 6412
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1584 4684 1636 4690
rect 1584 4626 1636 4632
rect 1676 4684 1728 4690
rect 1676 4626 1728 4632
rect 1674 4040 1730 4049
rect 1492 4004 1544 4010
rect 1780 4010 1808 6258
rect 1952 6248 2004 6254
rect 1952 6190 2004 6196
rect 1860 5908 1912 5914
rect 1860 5850 1912 5856
rect 1674 3975 1730 3984
rect 1768 4004 1820 4010
rect 1492 3946 1544 3952
rect 1400 3188 1452 3194
rect 1400 3130 1452 3136
rect 1688 3058 1716 3975
rect 1768 3946 1820 3952
rect 1872 3466 1900 5850
rect 1860 3460 1912 3466
rect 1860 3402 1912 3408
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1964 2394 1992 6190
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 2056 4214 2084 4966
rect 2148 4690 2176 7686
rect 2240 5370 2268 8570
rect 2332 7410 2360 11319
rect 2516 11098 2544 11494
rect 2608 11370 2636 12106
rect 2700 11898 2728 12838
rect 2780 12776 2832 12782
rect 2780 12718 2832 12724
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2608 11342 2728 11370
rect 2424 11070 2544 11098
rect 2424 8974 2452 11070
rect 2504 11008 2556 11014
rect 2504 10950 2556 10956
rect 2516 10742 2544 10950
rect 2504 10736 2556 10742
rect 2504 10678 2556 10684
rect 2516 10554 2544 10678
rect 2516 10526 2636 10554
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 9042 2544 10406
rect 2608 10130 2636 10526
rect 2596 10124 2648 10130
rect 2596 10066 2648 10072
rect 2608 9042 2636 10066
rect 2700 9994 2728 11342
rect 2792 11150 2820 12718
rect 3174 12540 3482 12560
rect 3174 12538 3180 12540
rect 3236 12538 3260 12540
rect 3316 12538 3340 12540
rect 3396 12538 3420 12540
rect 3476 12538 3482 12540
rect 3236 12486 3238 12538
rect 3418 12486 3420 12538
rect 3174 12484 3180 12486
rect 3236 12484 3260 12486
rect 3316 12484 3340 12486
rect 3396 12484 3420 12486
rect 3476 12484 3482 12486
rect 3174 12464 3482 12484
rect 3896 12434 3924 12854
rect 4172 12646 4200 13262
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 3896 12406 4016 12434
rect 2964 12232 3016 12238
rect 2884 12192 2964 12220
rect 2780 11144 2832 11150
rect 2780 11086 2832 11092
rect 2792 10606 2820 11086
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2688 9988 2740 9994
rect 2688 9930 2740 9936
rect 2792 9654 2820 10542
rect 2780 9648 2832 9654
rect 2780 9590 2832 9596
rect 2792 9110 2820 9590
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2504 9036 2556 9042
rect 2504 8978 2556 8984
rect 2596 9036 2648 9042
rect 2596 8978 2648 8984
rect 2412 8968 2464 8974
rect 2412 8910 2464 8916
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2332 7002 2360 7346
rect 2504 7200 2556 7206
rect 2504 7142 2556 7148
rect 2320 6996 2372 7002
rect 2320 6938 2372 6944
rect 2410 6488 2466 6497
rect 2410 6423 2466 6432
rect 2318 6216 2374 6225
rect 2318 6151 2374 6160
rect 2332 5914 2360 6151
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 2136 4480 2188 4486
rect 2136 4422 2188 4428
rect 2148 4282 2176 4422
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 2044 4208 2096 4214
rect 2044 4150 2096 4156
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2148 4049 2176 4082
rect 2134 4040 2190 4049
rect 2134 3975 2190 3984
rect 2148 3194 2176 3975
rect 2240 3534 2268 4558
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2226 3360 2282 3369
rect 2226 3295 2282 3304
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 2148 2650 2176 2994
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 2240 2446 2268 3295
rect 2318 2680 2374 2689
rect 2318 2615 2374 2624
rect 2332 2514 2360 2615
rect 2320 2508 2372 2514
rect 2320 2450 2372 2456
rect 2424 2446 2452 6423
rect 2516 5234 2544 7142
rect 2608 5914 2636 8842
rect 2792 8430 2820 9046
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2792 7478 2820 8366
rect 2884 8242 2912 12192
rect 2964 12174 3016 12180
rect 3792 12232 3844 12238
rect 3792 12174 3844 12180
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3516 11824 3568 11830
rect 3514 11792 3516 11801
rect 3568 11792 3570 11801
rect 3514 11727 3570 11736
rect 3516 11688 3568 11694
rect 3516 11630 3568 11636
rect 3174 11452 3482 11472
rect 3174 11450 3180 11452
rect 3236 11450 3260 11452
rect 3316 11450 3340 11452
rect 3396 11450 3420 11452
rect 3476 11450 3482 11452
rect 3236 11398 3238 11450
rect 3418 11398 3420 11450
rect 3174 11396 3180 11398
rect 3236 11396 3260 11398
rect 3316 11396 3340 11398
rect 3396 11396 3420 11398
rect 3476 11396 3482 11398
rect 3174 11376 3482 11396
rect 3528 11082 3556 11630
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 2976 9654 3004 11018
rect 3528 10606 3556 11018
rect 3056 10600 3108 10606
rect 3056 10542 3108 10548
rect 3516 10600 3568 10606
rect 3516 10542 3568 10548
rect 3068 10266 3096 10542
rect 3174 10364 3482 10384
rect 3174 10362 3180 10364
rect 3236 10362 3260 10364
rect 3316 10362 3340 10364
rect 3396 10362 3420 10364
rect 3476 10362 3482 10364
rect 3236 10310 3238 10362
rect 3418 10310 3420 10362
rect 3174 10308 3180 10310
rect 3236 10308 3260 10310
rect 3316 10308 3340 10310
rect 3396 10308 3420 10310
rect 3476 10308 3482 10310
rect 3174 10288 3482 10308
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3528 10130 3556 10542
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3054 9752 3110 9761
rect 3054 9687 3110 9696
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2976 9042 3004 9590
rect 2964 9036 3016 9042
rect 2964 8978 3016 8984
rect 3068 8566 3096 9687
rect 3344 9466 3372 9862
rect 3344 9438 3556 9466
rect 3174 9276 3482 9296
rect 3174 9274 3180 9276
rect 3236 9274 3260 9276
rect 3316 9274 3340 9276
rect 3396 9274 3420 9276
rect 3476 9274 3482 9276
rect 3236 9222 3238 9274
rect 3418 9222 3420 9274
rect 3174 9220 3180 9222
rect 3236 9220 3260 9222
rect 3316 9220 3340 9222
rect 3396 9220 3420 9222
rect 3476 9220 3482 9222
rect 3174 9200 3482 9220
rect 3528 9042 3556 9438
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3528 8945 3556 8978
rect 3514 8936 3570 8945
rect 3514 8871 3570 8880
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 3436 8634 3464 8774
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2884 8214 3004 8242
rect 2870 8120 2926 8129
rect 2870 8055 2926 8064
rect 2780 7472 2832 7478
rect 2780 7414 2832 7420
rect 2686 6760 2742 6769
rect 2686 6695 2742 6704
rect 2780 6724 2832 6730
rect 2700 6662 2728 6695
rect 2780 6666 2832 6672
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 6458 2728 6598
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2596 5908 2648 5914
rect 2596 5850 2648 5856
rect 2596 5568 2648 5574
rect 2596 5510 2648 5516
rect 2608 5302 2636 5510
rect 2596 5296 2648 5302
rect 2596 5238 2648 5244
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 2504 4548 2556 4554
rect 2504 4490 2556 4496
rect 2516 3670 2544 4490
rect 2504 3664 2556 3670
rect 2504 3606 2556 3612
rect 2228 2440 2280 2446
rect 1964 2366 2176 2394
rect 2228 2382 2280 2388
rect 2412 2440 2464 2446
rect 2412 2382 2464 2388
rect 2148 800 2176 2366
rect 492 734 796 762
rect 1214 0 1270 800
rect 2134 0 2190 800
rect 2792 241 2820 6666
rect 2884 5098 2912 8055
rect 2976 6662 3004 8214
rect 3068 7546 3096 8502
rect 3516 8424 3568 8430
rect 3516 8366 3568 8372
rect 3174 8188 3482 8208
rect 3174 8186 3180 8188
rect 3236 8186 3260 8188
rect 3316 8186 3340 8188
rect 3396 8186 3420 8188
rect 3476 8186 3482 8188
rect 3236 8134 3238 8186
rect 3418 8134 3420 8186
rect 3174 8132 3180 8134
rect 3236 8132 3260 8134
rect 3316 8132 3340 8134
rect 3396 8132 3420 8134
rect 3476 8132 3482 8134
rect 3174 8112 3482 8132
rect 3528 7954 3556 8366
rect 3516 7948 3568 7954
rect 3516 7890 3568 7896
rect 3332 7744 3384 7750
rect 3330 7712 3332 7721
rect 3384 7712 3386 7721
rect 3330 7647 3386 7656
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3528 7274 3556 7890
rect 3516 7268 3568 7274
rect 3516 7210 3568 7216
rect 3174 7100 3482 7120
rect 3174 7098 3180 7100
rect 3236 7098 3260 7100
rect 3316 7098 3340 7100
rect 3396 7098 3420 7100
rect 3476 7098 3482 7100
rect 3236 7046 3238 7098
rect 3418 7046 3420 7098
rect 3174 7044 3180 7046
rect 3236 7044 3260 7046
rect 3316 7044 3340 7046
rect 3396 7044 3420 7046
rect 3476 7044 3482 7046
rect 3174 7024 3482 7044
rect 3148 6860 3200 6866
rect 3148 6802 3200 6808
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 3054 6216 3110 6225
rect 3160 6186 3188 6802
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3528 6202 3556 6598
rect 3620 6390 3648 12038
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3712 11218 3740 11698
rect 3804 11694 3832 12174
rect 3882 11928 3938 11937
rect 3882 11863 3938 11872
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3792 11552 3844 11558
rect 3792 11494 3844 11500
rect 3700 11212 3752 11218
rect 3700 11154 3752 11160
rect 3804 11098 3832 11494
rect 3896 11218 3924 11863
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3712 11070 3832 11098
rect 3712 8974 3740 11070
rect 3790 10976 3846 10985
rect 3790 10911 3846 10920
rect 3804 10538 3832 10911
rect 3792 10532 3844 10538
rect 3792 10474 3844 10480
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3896 10062 3924 10406
rect 3884 10056 3936 10062
rect 3884 9998 3936 10004
rect 3988 8974 4016 12406
rect 4172 12170 4200 12582
rect 4264 12170 4292 13382
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4252 12164 4304 12170
rect 4252 12106 4304 12112
rect 4066 11928 4122 11937
rect 4066 11863 4122 11872
rect 4252 11892 4304 11898
rect 4080 11830 4108 11863
rect 4252 11834 4304 11840
rect 4068 11824 4120 11830
rect 4068 11766 4120 11772
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4080 11150 4108 11630
rect 4160 11280 4212 11286
rect 4158 11248 4160 11257
rect 4212 11248 4214 11257
rect 4158 11183 4214 11192
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4172 10810 4200 11183
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4066 10160 4122 10169
rect 4172 10130 4200 10610
rect 4066 10095 4122 10104
rect 4160 10124 4212 10130
rect 4080 10062 4108 10095
rect 4160 10066 4212 10072
rect 4068 10056 4120 10062
rect 4068 9998 4120 10004
rect 4068 9376 4120 9382
rect 4068 9318 4120 9324
rect 3700 8968 3752 8974
rect 3700 8910 3752 8916
rect 3976 8968 4028 8974
rect 3976 8910 4028 8916
rect 3712 8022 3740 8910
rect 3988 8838 4016 8910
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3700 8016 3752 8022
rect 3700 7958 3752 7964
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3054 6151 3110 6160
rect 3148 6180 3200 6186
rect 2964 6112 3016 6118
rect 2964 6054 3016 6060
rect 2872 5092 2924 5098
rect 2872 5034 2924 5040
rect 2870 3904 2926 3913
rect 2870 3839 2926 3848
rect 2884 3126 2912 3839
rect 2976 3534 3004 6054
rect 3068 5778 3096 6151
rect 3528 6174 3648 6202
rect 3148 6122 3200 6128
rect 3516 6112 3568 6118
rect 3516 6054 3568 6060
rect 3174 6012 3482 6032
rect 3174 6010 3180 6012
rect 3236 6010 3260 6012
rect 3316 6010 3340 6012
rect 3396 6010 3420 6012
rect 3476 6010 3482 6012
rect 3236 5958 3238 6010
rect 3418 5958 3420 6010
rect 3174 5956 3180 5958
rect 3236 5956 3260 5958
rect 3316 5956 3340 5958
rect 3396 5956 3420 5958
rect 3476 5956 3482 5958
rect 3174 5936 3482 5956
rect 3056 5772 3108 5778
rect 3056 5714 3108 5720
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 2872 3120 2924 3126
rect 2872 3062 2924 3068
rect 2976 2514 3004 3130
rect 2964 2508 3016 2514
rect 2964 2450 3016 2456
rect 2872 2304 2924 2310
rect 2872 2246 2924 2252
rect 2884 2009 2912 2246
rect 2870 2000 2926 2009
rect 2870 1935 2926 1944
rect 3068 800 3096 5578
rect 3174 4924 3482 4944
rect 3174 4922 3180 4924
rect 3236 4922 3260 4924
rect 3316 4922 3340 4924
rect 3396 4922 3420 4924
rect 3476 4922 3482 4924
rect 3236 4870 3238 4922
rect 3418 4870 3420 4922
rect 3174 4868 3180 4870
rect 3236 4868 3260 4870
rect 3316 4868 3340 4870
rect 3396 4868 3420 4870
rect 3476 4868 3482 4870
rect 3174 4848 3482 4868
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3436 4214 3464 4422
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 3174 3836 3482 3856
rect 3174 3834 3180 3836
rect 3236 3834 3260 3836
rect 3316 3834 3340 3836
rect 3396 3834 3420 3836
rect 3476 3834 3482 3836
rect 3236 3782 3238 3834
rect 3418 3782 3420 3834
rect 3174 3780 3180 3782
rect 3236 3780 3260 3782
rect 3316 3780 3340 3782
rect 3396 3780 3420 3782
rect 3476 3780 3482 3782
rect 3174 3760 3482 3780
rect 3528 3194 3556 6054
rect 3620 3942 3648 6174
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3712 5001 3740 5646
rect 3698 4992 3754 5001
rect 3698 4927 3754 4936
rect 3700 4208 3752 4214
rect 3700 4150 3752 4156
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3712 3466 3740 4150
rect 3804 3641 3832 8774
rect 3988 8673 4016 8774
rect 3974 8664 4030 8673
rect 3974 8599 4030 8608
rect 4080 8362 4108 9318
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4172 8090 4200 9114
rect 4264 8566 4292 11834
rect 4356 11286 4384 14606
rect 5552 14346 5580 16400
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 5540 14340 5592 14346
rect 5540 14282 5592 14288
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 5398 14172 5706 14192
rect 5398 14170 5404 14172
rect 5460 14170 5484 14172
rect 5540 14170 5564 14172
rect 5620 14170 5644 14172
rect 5700 14170 5706 14172
rect 5460 14118 5462 14170
rect 5642 14118 5644 14170
rect 5398 14116 5404 14118
rect 5460 14116 5484 14118
rect 5540 14116 5564 14118
rect 5620 14116 5644 14118
rect 5700 14116 5706 14118
rect 5398 14096 5706 14116
rect 4988 14000 5040 14006
rect 5172 14000 5224 14006
rect 5040 13948 5172 13954
rect 4988 13942 5224 13948
rect 4896 13932 4948 13938
rect 5000 13926 5212 13942
rect 4896 13874 4948 13880
rect 4804 13864 4856 13870
rect 4804 13806 4856 13812
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4448 12986 4476 13670
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4526 13152 4582 13161
rect 4526 13087 4582 13096
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4344 11280 4396 11286
rect 4344 11222 4396 11228
rect 4342 10704 4398 10713
rect 4342 10639 4344 10648
rect 4396 10639 4398 10648
rect 4344 10610 4396 10616
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 4356 9178 4384 10134
rect 4344 9172 4396 9178
rect 4344 9114 4396 9120
rect 4252 8560 4304 8566
rect 4250 8528 4252 8537
rect 4304 8528 4306 8537
rect 4250 8463 4306 8472
rect 4252 8424 4304 8430
rect 4252 8366 4304 8372
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3896 7313 3924 7686
rect 4264 7410 4292 8366
rect 4448 7886 4476 12922
rect 4540 12646 4568 13087
rect 4632 12782 4660 13330
rect 4816 12986 4844 13806
rect 4908 13530 4936 13874
rect 6920 13864 6972 13870
rect 6920 13806 6972 13812
rect 5172 13796 5224 13802
rect 5172 13738 5224 13744
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4896 13184 4948 13190
rect 4896 13126 4948 13132
rect 4804 12980 4856 12986
rect 4804 12922 4856 12928
rect 4712 12912 4764 12918
rect 4712 12854 4764 12860
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4528 12640 4580 12646
rect 4528 12582 4580 12588
rect 4724 12434 4752 12854
rect 4632 12406 4752 12434
rect 4804 12436 4856 12442
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4540 10713 4568 12106
rect 4632 11014 4660 12406
rect 4804 12378 4856 12384
rect 4816 12322 4844 12378
rect 4724 12294 4844 12322
rect 4724 11762 4752 12294
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4620 11008 4672 11014
rect 4620 10950 4672 10956
rect 4620 10736 4672 10742
rect 4526 10704 4582 10713
rect 4620 10678 4672 10684
rect 4526 10639 4582 10648
rect 4632 10248 4660 10678
rect 4540 10220 4660 10248
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 3882 7304 3938 7313
rect 3882 7239 3938 7248
rect 3882 6896 3938 6905
rect 3882 6831 3938 6840
rect 3896 6662 3924 6831
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 3988 6118 4016 6734
rect 4160 6724 4212 6730
rect 4160 6666 4212 6672
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3882 5944 3938 5953
rect 3882 5879 3938 5888
rect 3896 5302 3924 5879
rect 3988 5642 4016 6054
rect 3976 5636 4028 5642
rect 3976 5578 4028 5584
rect 4068 5636 4120 5642
rect 4068 5578 4120 5584
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3988 5030 4016 5578
rect 3976 5024 4028 5030
rect 3976 4966 4028 4972
rect 3882 4856 3938 4865
rect 3882 4791 3884 4800
rect 3936 4791 3938 4800
rect 3884 4762 3936 4768
rect 3882 4720 3938 4729
rect 3882 4655 3938 4664
rect 3896 4214 3924 4655
rect 3988 4622 4016 4966
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3884 4208 3936 4214
rect 3884 4150 3936 4156
rect 3988 4078 4016 4558
rect 3976 4072 4028 4078
rect 3976 4014 4028 4020
rect 3988 3913 4016 4014
rect 3974 3904 4030 3913
rect 3974 3839 4030 3848
rect 3974 3768 4030 3777
rect 3974 3703 4030 3712
rect 3790 3632 3846 3641
rect 3988 3602 4016 3703
rect 3976 3596 4028 3602
rect 3790 3567 3846 3576
rect 3896 3556 3976 3584
rect 3700 3460 3752 3466
rect 3700 3402 3752 3408
rect 3516 3188 3568 3194
rect 3516 3130 3568 3136
rect 3792 2984 3844 2990
rect 3792 2926 3844 2932
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3174 2748 3482 2768
rect 3174 2746 3180 2748
rect 3236 2746 3260 2748
rect 3316 2746 3340 2748
rect 3396 2746 3420 2748
rect 3476 2746 3482 2748
rect 3236 2694 3238 2746
rect 3418 2694 3420 2746
rect 3174 2692 3180 2694
rect 3236 2692 3260 2694
rect 3316 2692 3340 2694
rect 3396 2692 3420 2694
rect 3476 2692 3482 2694
rect 3174 2672 3482 2692
rect 3528 2310 3556 2790
rect 3804 2650 3832 2926
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 3896 2514 3924 3556
rect 3976 3538 4028 3544
rect 4080 2774 4108 5578
rect 4172 3738 4200 6666
rect 4540 6361 4568 10220
rect 4620 10124 4672 10130
rect 4620 10066 4672 10072
rect 4632 8294 4660 10066
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4632 6458 4660 7686
rect 4724 7342 4752 11698
rect 4804 10804 4856 10810
rect 4804 10746 4856 10752
rect 4816 10538 4844 10746
rect 4908 10742 4936 13126
rect 5080 12776 5132 12782
rect 5080 12718 5132 12724
rect 5092 12442 5120 12718
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 5184 12374 5212 13738
rect 5816 13728 5868 13734
rect 5816 13670 5868 13676
rect 6092 13728 6144 13734
rect 6092 13670 6144 13676
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 5276 13258 5304 13398
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5264 13252 5316 13258
rect 5264 13194 5316 13200
rect 5398 13084 5706 13104
rect 5398 13082 5404 13084
rect 5460 13082 5484 13084
rect 5540 13082 5564 13084
rect 5620 13082 5644 13084
rect 5700 13082 5706 13084
rect 5460 13030 5462 13082
rect 5642 13030 5644 13082
rect 5398 13028 5404 13030
rect 5460 13028 5484 13030
rect 5540 13028 5564 13030
rect 5620 13028 5644 13030
rect 5700 13028 5706 13030
rect 5398 13008 5706 13028
rect 5736 12714 5764 13330
rect 5828 13190 5856 13670
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5828 12986 5856 13126
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 6104 12850 6132 13670
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 6092 12844 6144 12850
rect 6092 12786 6144 12792
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5172 12368 5224 12374
rect 5172 12310 5224 12316
rect 5184 11762 5212 12310
rect 5736 12306 5764 12650
rect 5828 12646 5856 12786
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5264 12096 5316 12102
rect 5264 12038 5316 12044
rect 5724 12096 5776 12102
rect 5724 12038 5776 12044
rect 5172 11756 5224 11762
rect 5172 11698 5224 11704
rect 4988 11076 5040 11082
rect 4988 11018 5040 11024
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 5000 10538 5028 11018
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 4804 10532 4856 10538
rect 4804 10474 4856 10480
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 5000 10130 5028 10474
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4908 9926 4936 9998
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4908 9586 4936 9862
rect 4896 9580 4948 9586
rect 4896 9522 4948 9528
rect 5000 9042 5028 10066
rect 5092 9654 5120 10950
rect 5276 10062 5304 12038
rect 5398 11996 5706 12016
rect 5398 11994 5404 11996
rect 5460 11994 5484 11996
rect 5540 11994 5564 11996
rect 5620 11994 5644 11996
rect 5700 11994 5706 11996
rect 5460 11942 5462 11994
rect 5642 11942 5644 11994
rect 5398 11940 5404 11942
rect 5460 11940 5484 11942
rect 5540 11940 5564 11942
rect 5620 11940 5644 11942
rect 5700 11940 5706 11942
rect 5398 11920 5706 11940
rect 5736 11898 5764 12038
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 11082 5488 11494
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5398 10908 5706 10928
rect 5398 10906 5404 10908
rect 5460 10906 5484 10908
rect 5540 10906 5564 10908
rect 5620 10906 5644 10908
rect 5700 10906 5706 10908
rect 5460 10854 5462 10906
rect 5642 10854 5644 10906
rect 5398 10852 5404 10854
rect 5460 10852 5484 10854
rect 5540 10852 5564 10854
rect 5620 10852 5644 10854
rect 5700 10852 5706 10854
rect 5398 10832 5706 10852
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5264 10056 5316 10062
rect 5264 9998 5316 10004
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5092 8906 5120 9590
rect 5172 9580 5224 9586
rect 5172 9522 5224 9528
rect 5184 9382 5212 9522
rect 5172 9376 5224 9382
rect 5170 9344 5172 9353
rect 5224 9344 5226 9353
rect 5170 9279 5226 9288
rect 5080 8900 5132 8906
rect 5080 8842 5132 8848
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4816 7954 4844 8570
rect 4988 8492 5040 8498
rect 4988 8434 5040 8440
rect 4896 8084 4948 8090
rect 4896 8026 4948 8032
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4908 7834 4936 8026
rect 5000 8022 5028 8434
rect 5276 8378 5304 9998
rect 5398 9820 5706 9840
rect 5398 9818 5404 9820
rect 5460 9818 5484 9820
rect 5540 9818 5564 9820
rect 5620 9818 5644 9820
rect 5700 9818 5706 9820
rect 5460 9766 5462 9818
rect 5642 9766 5644 9818
rect 5398 9764 5404 9766
rect 5460 9764 5484 9766
rect 5540 9764 5564 9766
rect 5620 9764 5644 9766
rect 5700 9764 5706 9766
rect 5398 9744 5706 9764
rect 5736 8974 5764 10406
rect 5724 8968 5776 8974
rect 5630 8936 5686 8945
rect 5724 8910 5776 8916
rect 5630 8871 5686 8880
rect 5644 8820 5672 8871
rect 5644 8792 5764 8820
rect 5398 8732 5706 8752
rect 5398 8730 5404 8732
rect 5460 8730 5484 8732
rect 5540 8730 5564 8732
rect 5620 8730 5644 8732
rect 5700 8730 5706 8732
rect 5460 8678 5462 8730
rect 5642 8678 5644 8730
rect 5398 8676 5404 8678
rect 5460 8676 5484 8678
rect 5540 8676 5564 8678
rect 5620 8676 5644 8678
rect 5700 8676 5706 8678
rect 5398 8656 5706 8676
rect 5092 8350 5304 8378
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 4816 7806 4936 7834
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4620 6452 4672 6458
rect 4620 6394 4672 6400
rect 4526 6352 4582 6361
rect 4252 6316 4304 6322
rect 4724 6322 4752 7278
rect 4526 6287 4528 6296
rect 4252 6258 4304 6264
rect 4580 6287 4582 6296
rect 4712 6316 4764 6322
rect 4528 6258 4580 6264
rect 4712 6258 4764 6264
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4264 3602 4292 6258
rect 4540 6227 4568 6258
rect 4528 6112 4580 6118
rect 4342 6080 4398 6089
rect 4528 6054 4580 6060
rect 4342 6015 4398 6024
rect 4356 5370 4384 6015
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4448 5273 4476 5646
rect 4434 5264 4490 5273
rect 4434 5199 4490 5208
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4356 4282 4384 4490
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4252 3596 4304 3602
rect 4252 3538 4304 3544
rect 4158 3496 4214 3505
rect 4356 3482 4384 4218
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4448 4049 4476 4082
rect 4434 4040 4490 4049
rect 4434 3975 4490 3984
rect 4436 3664 4488 3670
rect 4434 3632 4436 3641
rect 4488 3632 4490 3641
rect 4434 3567 4490 3576
rect 4158 3431 4214 3440
rect 4264 3454 4384 3482
rect 4540 3482 4568 6054
rect 4712 5568 4764 5574
rect 4618 5536 4674 5545
rect 4712 5510 4764 5516
rect 4618 5471 4674 5480
rect 4632 3738 4660 5471
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4724 3670 4752 5510
rect 4816 5370 4844 7806
rect 5000 6866 5028 7958
rect 5092 7478 5120 8350
rect 5264 8288 5316 8294
rect 5264 8230 5316 8236
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5184 7478 5212 7890
rect 5276 7546 5304 8230
rect 5398 7644 5706 7664
rect 5398 7642 5404 7644
rect 5460 7642 5484 7644
rect 5540 7642 5564 7644
rect 5620 7642 5644 7644
rect 5700 7642 5706 7644
rect 5460 7590 5462 7642
rect 5642 7590 5644 7642
rect 5398 7588 5404 7590
rect 5460 7588 5484 7590
rect 5540 7588 5564 7590
rect 5620 7588 5644 7590
rect 5700 7588 5706 7590
rect 5398 7568 5706 7588
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5080 7472 5132 7478
rect 5080 7414 5132 7420
rect 5172 7472 5224 7478
rect 5172 7414 5224 7420
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5632 7472 5684 7478
rect 5632 7414 5684 7420
rect 4988 6860 5040 6866
rect 4988 6802 5040 6808
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4908 5846 4936 6598
rect 5000 6254 5028 6802
rect 4988 6248 5040 6254
rect 4988 6190 5040 6196
rect 5092 5953 5120 7414
rect 5264 7336 5316 7342
rect 5264 7278 5316 7284
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5184 6390 5212 7142
rect 5172 6384 5224 6390
rect 5172 6326 5224 6332
rect 5078 5944 5134 5953
rect 5078 5879 5134 5888
rect 4896 5840 4948 5846
rect 4896 5782 4948 5788
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4908 5250 4936 5782
rect 5092 5710 5120 5879
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 5080 5704 5132 5710
rect 5080 5646 5132 5652
rect 5000 5545 5028 5646
rect 4986 5536 5042 5545
rect 4986 5471 5042 5480
rect 4908 5222 5028 5250
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4816 4622 4844 4966
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4908 4282 4936 5102
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4802 3904 4858 3913
rect 4802 3839 4858 3848
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 4436 3460 4488 3466
rect 4172 3398 4200 3431
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 3988 2746 4108 2774
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 3516 2304 3568 2310
rect 3516 2246 3568 2252
rect 3882 2272 3938 2281
rect 3882 2207 3938 2216
rect 3896 1698 3924 2207
rect 3884 1692 3936 1698
rect 3884 1634 3936 1640
rect 3332 1488 3384 1494
rect 3330 1456 3332 1465
rect 3384 1456 3386 1465
rect 3330 1391 3386 1400
rect 3700 1284 3752 1290
rect 3700 1226 3752 1232
rect 2778 232 2834 241
rect 2778 167 2834 176
rect 3054 0 3110 800
rect 3712 649 3740 1226
rect 3988 800 4016 2746
rect 4264 2446 4292 3454
rect 4540 3454 4752 3482
rect 4436 3402 4488 3408
rect 4448 2854 4476 3402
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4632 3058 4660 3130
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4620 2916 4672 2922
rect 4620 2858 4672 2864
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 4342 2544 4398 2553
rect 4342 2479 4344 2488
rect 4396 2479 4398 2488
rect 4344 2450 4396 2456
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4632 2281 4660 2858
rect 4724 2417 4752 3454
rect 4816 3058 4844 3839
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4908 2582 4936 4082
rect 5000 3777 5028 5222
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4986 3768 5042 3777
rect 4986 3703 5042 3712
rect 5092 3194 5120 4422
rect 5184 3369 5212 5034
rect 5276 5030 5304 7278
rect 5552 6730 5580 7414
rect 5644 7177 5672 7414
rect 5630 7168 5686 7177
rect 5630 7103 5686 7112
rect 5630 6896 5686 6905
rect 5630 6831 5686 6840
rect 5644 6798 5672 6831
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5398 6556 5706 6576
rect 5398 6554 5404 6556
rect 5460 6554 5484 6556
rect 5540 6554 5564 6556
rect 5620 6554 5644 6556
rect 5700 6554 5706 6556
rect 5460 6502 5462 6554
rect 5642 6502 5644 6554
rect 5398 6500 5404 6502
rect 5460 6500 5484 6502
rect 5540 6500 5564 6502
rect 5620 6500 5644 6502
rect 5700 6500 5706 6502
rect 5398 6480 5706 6500
rect 5398 5468 5706 5488
rect 5398 5466 5404 5468
rect 5460 5466 5484 5468
rect 5540 5466 5564 5468
rect 5620 5466 5644 5468
rect 5700 5466 5706 5468
rect 5460 5414 5462 5466
rect 5642 5414 5644 5466
rect 5398 5412 5404 5414
rect 5460 5412 5484 5414
rect 5540 5412 5564 5414
rect 5620 5412 5644 5414
rect 5700 5412 5706 5414
rect 5398 5392 5706 5412
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5368 4468 5396 5170
rect 5276 4440 5396 4468
rect 5276 4010 5304 4440
rect 5398 4380 5706 4400
rect 5398 4378 5404 4380
rect 5460 4378 5484 4380
rect 5540 4378 5564 4380
rect 5620 4378 5644 4380
rect 5700 4378 5706 4380
rect 5460 4326 5462 4378
rect 5642 4326 5644 4378
rect 5398 4324 5404 4326
rect 5460 4324 5484 4326
rect 5540 4324 5564 4326
rect 5620 4324 5644 4326
rect 5700 4324 5706 4326
rect 5398 4304 5706 4324
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5264 4004 5316 4010
rect 5264 3946 5316 3952
rect 5262 3768 5318 3777
rect 5460 3738 5488 4082
rect 5262 3703 5318 3712
rect 5448 3732 5500 3738
rect 5276 3602 5304 3703
rect 5448 3674 5500 3680
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5736 3534 5764 8792
rect 5828 6458 5856 12582
rect 5920 12442 5948 12718
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 6276 11280 6328 11286
rect 6276 11222 6328 11228
rect 6092 11076 6144 11082
rect 6092 11018 6144 11024
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5920 8634 5948 10610
rect 5998 10024 6054 10033
rect 5998 9959 6000 9968
rect 6052 9959 6054 9968
rect 6000 9930 6052 9936
rect 6012 9722 6040 9930
rect 6000 9716 6052 9722
rect 6000 9658 6052 9664
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5908 7744 5960 7750
rect 5908 7686 5960 7692
rect 5816 6452 5868 6458
rect 5816 6394 5868 6400
rect 5920 5250 5948 7686
rect 6012 7002 6040 9454
rect 6104 8945 6132 11018
rect 6288 9674 6316 11222
rect 6380 11218 6408 13126
rect 6564 12714 6592 13330
rect 6932 13326 6960 13806
rect 6920 13320 6972 13326
rect 6920 13262 6972 13268
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 6552 12708 6604 12714
rect 6552 12650 6604 12656
rect 6736 12164 6788 12170
rect 6736 12106 6788 12112
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6564 11898 6592 12038
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 6748 11762 6776 12106
rect 6828 12096 6880 12102
rect 6932 12050 6960 13126
rect 7024 12850 7052 13126
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 7024 12306 7052 12786
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7012 12300 7064 12306
rect 7012 12242 7064 12248
rect 6880 12044 6960 12050
rect 6828 12038 6960 12044
rect 6840 12022 6960 12038
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6828 11688 6880 11694
rect 6932 11665 6960 12022
rect 7024 11694 7052 12242
rect 7116 12238 7144 12582
rect 7208 12434 7236 14214
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 7208 12406 7328 12434
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7208 11694 7236 12310
rect 7012 11688 7064 11694
rect 6828 11630 6880 11636
rect 6918 11656 6974 11665
rect 6736 11620 6788 11626
rect 6736 11562 6788 11568
rect 6644 11280 6696 11286
rect 6644 11222 6696 11228
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6380 10452 6408 10746
rect 6472 10742 6500 11018
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6460 10736 6512 10742
rect 6460 10678 6512 10684
rect 6472 10577 6500 10678
rect 6458 10568 6514 10577
rect 6458 10503 6514 10512
rect 6380 10424 6500 10452
rect 6288 9646 6408 9674
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 6196 8974 6224 9522
rect 6184 8968 6236 8974
rect 6090 8936 6146 8945
rect 6184 8910 6236 8916
rect 6090 8871 6146 8880
rect 6196 8498 6224 8910
rect 6184 8492 6236 8498
rect 6236 8452 6316 8480
rect 6184 8434 6236 8440
rect 6184 8356 6236 8362
rect 6184 8298 6236 8304
rect 6196 8090 6224 8298
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 6288 7886 6316 8452
rect 6380 8430 6408 9646
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6092 7812 6144 7818
rect 6092 7754 6144 7760
rect 6104 7274 6132 7754
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6196 7313 6224 7346
rect 6182 7304 6238 7313
rect 6092 7268 6144 7274
rect 6182 7239 6238 7248
rect 6276 7268 6328 7274
rect 6092 7210 6144 7216
rect 6276 7210 6328 7216
rect 6184 7200 6236 7206
rect 6184 7142 6236 7148
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 6196 6866 6224 7142
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6092 6656 6144 6662
rect 6092 6598 6144 6604
rect 6184 6656 6236 6662
rect 6184 6598 6236 6604
rect 6104 6458 6132 6598
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6196 6186 6224 6598
rect 6288 6254 6316 7210
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6184 6180 6236 6186
rect 6184 6122 6236 6128
rect 6092 5908 6144 5914
rect 6092 5850 6144 5856
rect 5828 5222 5948 5250
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5170 3360 5226 3369
rect 5170 3295 5226 3304
rect 5398 3292 5706 3312
rect 5398 3290 5404 3292
rect 5460 3290 5484 3292
rect 5540 3290 5564 3292
rect 5620 3290 5644 3292
rect 5700 3290 5706 3292
rect 5460 3238 5462 3290
rect 5642 3238 5644 3290
rect 5398 3236 5404 3238
rect 5460 3236 5484 3238
rect 5540 3236 5564 3238
rect 5620 3236 5644 3238
rect 5700 3236 5706 3238
rect 5398 3216 5706 3236
rect 5080 3188 5132 3194
rect 5080 3130 5132 3136
rect 5092 3058 5120 3130
rect 5538 3088 5594 3097
rect 5080 3052 5132 3058
rect 5538 3023 5540 3032
rect 5080 2994 5132 3000
rect 5592 3023 5594 3032
rect 5540 2994 5592 3000
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 4710 2408 4766 2417
rect 4710 2343 4766 2352
rect 5000 2310 5028 2586
rect 4712 2304 4764 2310
rect 4618 2272 4674 2281
rect 4712 2246 4764 2252
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 4988 2304 5040 2310
rect 4988 2246 5040 2252
rect 4618 2207 4674 2216
rect 4068 1896 4120 1902
rect 4066 1864 4068 1873
rect 4120 1864 4122 1873
rect 4066 1799 4122 1808
rect 4724 1170 4752 2246
rect 4816 2106 4844 2246
rect 4804 2100 4856 2106
rect 4804 2042 4856 2048
rect 5092 1766 5120 2994
rect 5540 2848 5592 2854
rect 5540 2790 5592 2796
rect 5552 2689 5580 2790
rect 5538 2680 5594 2689
rect 5538 2615 5594 2624
rect 5722 2544 5778 2553
rect 5722 2479 5778 2488
rect 5736 2446 5764 2479
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5398 2204 5706 2224
rect 5398 2202 5404 2204
rect 5460 2202 5484 2204
rect 5540 2202 5564 2204
rect 5620 2202 5644 2204
rect 5700 2202 5706 2204
rect 5460 2150 5462 2202
rect 5642 2150 5644 2202
rect 5398 2148 5404 2150
rect 5460 2148 5484 2150
rect 5540 2148 5564 2150
rect 5620 2148 5644 2150
rect 5700 2148 5706 2150
rect 5398 2128 5706 2148
rect 5736 1834 5764 2382
rect 5724 1828 5776 1834
rect 5724 1770 5776 1776
rect 5080 1760 5132 1766
rect 5080 1702 5132 1708
rect 5828 1290 5856 5222
rect 6000 5160 6052 5166
rect 6000 5102 6052 5108
rect 6012 4486 6040 5102
rect 6000 4480 6052 4486
rect 6000 4422 6052 4428
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5920 3194 5948 4014
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 5906 2544 5962 2553
rect 5906 2479 5962 2488
rect 5920 2310 5948 2479
rect 5908 2304 5960 2310
rect 5908 2246 5960 2252
rect 6012 1970 6040 4422
rect 6000 1964 6052 1970
rect 6000 1906 6052 1912
rect 5816 1284 5868 1290
rect 5816 1226 5868 1232
rect 4724 1142 4936 1170
rect 4068 1080 4120 1086
rect 4066 1048 4068 1057
rect 4120 1048 4122 1057
rect 4066 983 4122 992
rect 4908 800 4936 1142
rect 5828 870 5948 898
rect 5828 800 5856 870
rect 3698 640 3754 649
rect 3698 575 3754 584
rect 3974 0 4030 800
rect 4894 0 4950 800
rect 5814 0 5870 800
rect 5920 762 5948 870
rect 6104 762 6132 5850
rect 6196 3516 6224 6122
rect 6380 4214 6408 8230
rect 6472 8090 6500 10424
rect 6460 8084 6512 8090
rect 6460 8026 6512 8032
rect 6460 7200 6512 7206
rect 6460 7142 6512 7148
rect 6368 4208 6420 4214
rect 6368 4150 6420 4156
rect 6196 3488 6408 3516
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 6274 3360 6330 3369
rect 6196 3126 6224 3334
rect 6274 3295 6330 3304
rect 6184 3120 6236 3126
rect 6184 3062 6236 3068
rect 6184 2848 6236 2854
rect 6184 2790 6236 2796
rect 6196 2038 6224 2790
rect 6288 2650 6316 3295
rect 6380 2854 6408 3488
rect 6472 3058 6500 7142
rect 6564 5681 6592 10950
rect 6656 10810 6684 11222
rect 6748 11218 6776 11562
rect 6840 11354 6868 11630
rect 7012 11630 7064 11636
rect 7196 11688 7248 11694
rect 7196 11630 7248 11636
rect 6918 11591 6974 11600
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6736 11212 6788 11218
rect 6736 11154 6788 11160
rect 6828 11144 6880 11150
rect 6932 11121 6960 11591
rect 7196 11552 7248 11558
rect 7196 11494 7248 11500
rect 6828 11086 6880 11092
rect 6918 11112 6974 11121
rect 6644 10804 6696 10810
rect 6644 10746 6696 10752
rect 6840 10674 6868 11086
rect 6918 11047 6974 11056
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6920 11008 6972 11014
rect 6920 10950 6972 10956
rect 6932 10810 6960 10950
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6656 10266 6684 10610
rect 6840 10266 6868 10610
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 6642 10024 6698 10033
rect 6642 9959 6698 9968
rect 6656 7206 6684 9959
rect 6748 8566 6776 10066
rect 6840 9654 6868 10202
rect 6828 9648 6880 9654
rect 6828 9590 6880 9596
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6932 9110 6960 9522
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6932 8906 6960 9046
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6736 8560 6788 8566
rect 6736 8502 6788 8508
rect 6748 7410 6776 8502
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6644 7200 6696 7206
rect 6696 7160 6776 7188
rect 6644 7142 6696 7148
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6656 6225 6684 6258
rect 6642 6216 6698 6225
rect 6642 6151 6698 6160
rect 6550 5672 6606 5681
rect 6550 5607 6606 5616
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6564 4622 6592 5510
rect 6748 4622 6776 7160
rect 6840 6780 6868 8774
rect 6920 8628 6972 8634
rect 7024 8616 7052 11018
rect 7104 10600 7156 10606
rect 7104 10542 7156 10548
rect 7116 10266 7144 10542
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7104 9376 7156 9382
rect 7104 9318 7156 9324
rect 7116 8634 7144 9318
rect 6972 8588 7052 8616
rect 7104 8628 7156 8634
rect 6920 8570 6972 8576
rect 7104 8570 7156 8576
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6918 8392 6974 8401
rect 6918 8327 6920 8336
rect 6972 8327 6974 8336
rect 6920 8298 6972 8304
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6932 7698 6960 8026
rect 7024 7857 7052 8434
rect 7010 7848 7066 7857
rect 7010 7783 7066 7792
rect 7104 7744 7156 7750
rect 6932 7670 7052 7698
rect 7104 7686 7156 7692
rect 6918 7576 6974 7585
rect 6918 7511 6920 7520
rect 6972 7511 6974 7520
rect 6920 7482 6972 7488
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6932 7206 6960 7278
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6920 6792 6972 6798
rect 6840 6760 6920 6780
rect 6972 6760 6974 6769
rect 6840 6752 6918 6760
rect 6918 6695 6974 6704
rect 6920 6656 6972 6662
rect 6918 6624 6920 6633
rect 6972 6624 6974 6633
rect 6918 6559 6974 6568
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6932 5914 6960 6326
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7024 5794 7052 7670
rect 6932 5766 7052 5794
rect 6552 4616 6604 4622
rect 6736 4616 6788 4622
rect 6552 4558 6604 4564
rect 6656 4576 6736 4604
rect 6552 4072 6604 4078
rect 6550 4040 6552 4049
rect 6604 4040 6606 4049
rect 6550 3975 6606 3984
rect 6656 3670 6684 4576
rect 6736 4558 6788 4564
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6644 3664 6696 3670
rect 6644 3606 6696 3612
rect 6460 3052 6512 3058
rect 6460 2994 6512 3000
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6276 2644 6328 2650
rect 6276 2586 6328 2592
rect 6184 2032 6236 2038
rect 6184 1974 6236 1980
rect 6748 800 6776 3946
rect 6840 1902 6868 4422
rect 6932 3233 6960 5766
rect 7012 5160 7064 5166
rect 7012 5102 7064 5108
rect 6918 3224 6974 3233
rect 6918 3159 6974 3168
rect 6920 2848 6972 2854
rect 6920 2790 6972 2796
rect 6932 2446 6960 2790
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 6920 2304 6972 2310
rect 6918 2272 6920 2281
rect 6972 2272 6974 2281
rect 6918 2207 6974 2216
rect 6828 1896 6880 1902
rect 6828 1838 6880 1844
rect 5920 734 6132 762
rect 6734 0 6790 800
rect 7024 762 7052 5102
rect 7116 3058 7144 7686
rect 7208 5234 7236 11494
rect 7300 9654 7328 12406
rect 7392 12306 7420 12854
rect 7380 12300 7432 12306
rect 7380 12242 7432 12248
rect 7392 10742 7420 12242
rect 7484 11354 7512 15370
rect 7622 14716 7930 14736
rect 7622 14714 7628 14716
rect 7684 14714 7708 14716
rect 7764 14714 7788 14716
rect 7844 14714 7868 14716
rect 7924 14714 7930 14716
rect 7684 14662 7686 14714
rect 7866 14662 7868 14714
rect 7622 14660 7628 14662
rect 7684 14660 7708 14662
rect 7764 14660 7788 14662
rect 7844 14660 7868 14662
rect 7924 14660 7930 14662
rect 7622 14640 7930 14660
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7576 14006 7604 14214
rect 7564 14000 7616 14006
rect 7564 13942 7616 13948
rect 7622 13628 7930 13648
rect 7622 13626 7628 13628
rect 7684 13626 7708 13628
rect 7764 13626 7788 13628
rect 7844 13626 7868 13628
rect 7924 13626 7930 13628
rect 7684 13574 7686 13626
rect 7866 13574 7868 13626
rect 7622 13572 7628 13574
rect 7684 13572 7708 13574
rect 7764 13572 7788 13574
rect 7844 13572 7868 13574
rect 7924 13572 7930 13574
rect 7622 13552 7930 13572
rect 7840 13320 7892 13326
rect 7840 13262 7892 13268
rect 7852 12850 7880 13262
rect 8036 13258 8064 16510
rect 9954 16510 10272 16538
rect 9954 16400 10010 16510
rect 9220 15224 9272 15230
rect 9220 15166 9272 15172
rect 8484 13524 8536 13530
rect 8484 13466 8536 13472
rect 8496 13394 8524 13466
rect 8484 13388 8536 13394
rect 8484 13330 8536 13336
rect 8024 13252 8076 13258
rect 8024 13194 8076 13200
rect 8116 12912 8168 12918
rect 8116 12854 8168 12860
rect 7840 12844 7892 12850
rect 7840 12786 7892 12792
rect 7622 12540 7930 12560
rect 7622 12538 7628 12540
rect 7684 12538 7708 12540
rect 7764 12538 7788 12540
rect 7844 12538 7868 12540
rect 7924 12538 7930 12540
rect 7684 12486 7686 12538
rect 7866 12486 7868 12538
rect 7622 12484 7628 12486
rect 7684 12484 7708 12486
rect 7764 12484 7788 12486
rect 7844 12484 7868 12486
rect 7924 12484 7930 12486
rect 7622 12464 7930 12484
rect 8128 12434 8156 12854
rect 8392 12776 8444 12782
rect 8392 12718 8444 12724
rect 8036 12406 8156 12434
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7668 11694 7696 11834
rect 7656 11688 7708 11694
rect 7656 11630 7708 11636
rect 7622 11452 7930 11472
rect 7622 11450 7628 11452
rect 7684 11450 7708 11452
rect 7764 11450 7788 11452
rect 7844 11450 7868 11452
rect 7924 11450 7930 11452
rect 7684 11398 7686 11450
rect 7866 11398 7868 11450
rect 7622 11396 7628 11398
rect 7684 11396 7708 11398
rect 7764 11396 7788 11398
rect 7844 11396 7868 11398
rect 7924 11396 7930 11398
rect 7622 11376 7930 11396
rect 7472 11348 7524 11354
rect 7472 11290 7524 11296
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 7944 11082 7972 11222
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7380 10736 7432 10742
rect 7380 10678 7432 10684
rect 7472 10668 7524 10674
rect 7472 10610 7524 10616
rect 7484 10470 7512 10610
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7484 9722 7512 10406
rect 7622 10364 7930 10384
rect 7622 10362 7628 10364
rect 7684 10362 7708 10364
rect 7764 10362 7788 10364
rect 7844 10362 7868 10364
rect 7924 10362 7930 10364
rect 7684 10310 7686 10362
rect 7866 10310 7868 10362
rect 7622 10308 7628 10310
rect 7684 10308 7708 10310
rect 7764 10308 7788 10310
rect 7844 10308 7868 10310
rect 7924 10308 7930 10310
rect 7622 10288 7930 10308
rect 7564 10192 7616 10198
rect 7562 10160 7564 10169
rect 7748 10192 7800 10198
rect 7616 10160 7618 10169
rect 7748 10134 7800 10140
rect 7562 10095 7618 10104
rect 7760 9926 7788 10134
rect 8036 10130 8064 12406
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8220 11218 8248 11698
rect 8404 11626 8432 12718
rect 8392 11620 8444 11626
rect 8392 11562 8444 11568
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8128 10130 8156 11154
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8116 10124 8168 10130
rect 8116 10066 8168 10072
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7288 9648 7340 9654
rect 7288 9590 7340 9596
rect 7392 9382 7420 9658
rect 7380 9376 7432 9382
rect 7286 9344 7342 9353
rect 7342 9324 7380 9330
rect 7342 9318 7432 9324
rect 7342 9302 7420 9318
rect 7286 9279 7342 9288
rect 7392 9253 7420 9302
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7300 6934 7328 9114
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7392 7324 7420 8842
rect 7484 8430 7512 9658
rect 7622 9276 7930 9296
rect 7622 9274 7628 9276
rect 7684 9274 7708 9276
rect 7764 9274 7788 9276
rect 7844 9274 7868 9276
rect 7924 9274 7930 9276
rect 7684 9222 7686 9274
rect 7866 9222 7868 9274
rect 7622 9220 7628 9222
rect 7684 9220 7708 9222
rect 7764 9220 7788 9222
rect 7844 9220 7868 9222
rect 7924 9220 7930 9222
rect 7622 9200 7930 9220
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7622 8188 7930 8208
rect 7622 8186 7628 8188
rect 7684 8186 7708 8188
rect 7764 8186 7788 8188
rect 7844 8186 7868 8188
rect 7924 8186 7930 8188
rect 7684 8134 7686 8186
rect 7866 8134 7868 8186
rect 7622 8132 7628 8134
rect 7684 8132 7708 8134
rect 7764 8132 7788 8134
rect 7844 8132 7868 8134
rect 7924 8132 7930 8134
rect 7622 8112 7930 8132
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7760 7410 7788 7890
rect 7748 7404 7800 7410
rect 7748 7346 7800 7352
rect 7472 7336 7524 7342
rect 7392 7296 7472 7324
rect 7472 7278 7524 7284
rect 7378 7168 7434 7177
rect 7378 7103 7434 7112
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 7392 6798 7420 7103
rect 7622 7100 7930 7120
rect 7622 7098 7628 7100
rect 7684 7098 7708 7100
rect 7764 7098 7788 7100
rect 7844 7098 7868 7100
rect 7924 7098 7930 7100
rect 7684 7046 7686 7098
rect 7866 7046 7868 7098
rect 7622 7044 7628 7046
rect 7684 7044 7708 7046
rect 7764 7044 7788 7046
rect 7844 7044 7868 7046
rect 7924 7044 7930 7046
rect 7622 7024 7930 7044
rect 8036 6798 8064 10066
rect 8128 9586 8156 10066
rect 8220 9994 8248 11018
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8312 10810 8340 10950
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8312 10169 8340 10406
rect 8298 10160 8354 10169
rect 8298 10095 8354 10104
rect 8208 9988 8260 9994
rect 8208 9930 8260 9936
rect 8496 9674 8524 13330
rect 9036 13320 9088 13326
rect 9036 13262 9088 13268
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8956 12986 8984 13126
rect 8944 12980 8996 12986
rect 8944 12922 8996 12928
rect 9048 12714 9076 13262
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8760 12436 8812 12442
rect 8760 12378 8812 12384
rect 8772 11694 8800 12378
rect 8864 11898 8892 12582
rect 8944 12096 8996 12102
rect 8944 12038 8996 12044
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 8956 11830 8984 12038
rect 8944 11824 8996 11830
rect 8944 11766 8996 11772
rect 9232 11762 9260 15166
rect 9846 14172 10154 14192
rect 9846 14170 9852 14172
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 10148 14170 10154 14172
rect 9908 14118 9910 14170
rect 10090 14118 10092 14170
rect 9846 14116 9852 14118
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 10148 14116 10154 14118
rect 9846 14096 10154 14116
rect 9404 13728 9456 13734
rect 9404 13670 9456 13676
rect 9416 13394 9444 13670
rect 10244 13530 10272 16510
rect 11900 16510 12112 16538
rect 10508 14476 10560 14482
rect 10508 14418 10560 14424
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10232 13524 10284 13530
rect 10232 13466 10284 13472
rect 10520 13462 10548 14418
rect 10612 13734 10640 14418
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10600 13728 10652 13734
rect 10600 13670 10652 13676
rect 10508 13456 10560 13462
rect 10508 13398 10560 13404
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9312 13184 9364 13190
rect 9312 13126 9364 13132
rect 9324 12306 9352 13126
rect 9692 12918 9720 13330
rect 10416 13184 10468 13190
rect 10416 13126 10468 13132
rect 9846 13084 10154 13104
rect 9846 13082 9852 13084
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 10148 13082 10154 13084
rect 9908 13030 9910 13082
rect 10090 13030 10092 13082
rect 9846 13028 9852 13030
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 10148 13028 10154 13030
rect 9846 13008 10154 13028
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9600 12306 9628 12582
rect 9692 12374 9720 12854
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10244 12442 10272 12786
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9312 12300 9364 12306
rect 9312 12242 9364 12248
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9402 12200 9458 12209
rect 9402 12135 9458 12144
rect 9496 12164 9548 12170
rect 9416 11898 9444 12135
rect 9496 12106 9548 12112
rect 9404 11892 9456 11898
rect 9404 11834 9456 11840
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9220 11756 9272 11762
rect 9220 11698 9272 11704
rect 8760 11688 8812 11694
rect 8760 11630 8812 11636
rect 8850 11656 8906 11665
rect 8850 11591 8906 11600
rect 8864 11354 8892 11591
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8588 10810 8616 11086
rect 8864 11014 8892 11290
rect 9048 11014 9076 11698
rect 9416 11354 9444 11834
rect 9508 11762 9536 12106
rect 9496 11756 9548 11762
rect 9496 11698 9548 11704
rect 9692 11694 9720 12310
rect 10428 12238 10456 13126
rect 10520 12238 10548 13398
rect 10980 13326 11008 14010
rect 11900 13394 11928 16510
rect 12084 16402 12112 16510
rect 12162 16402 12218 17200
rect 12084 16400 12218 16402
rect 14370 16400 14426 17200
rect 16578 16538 16634 17200
rect 18050 16824 18106 16833
rect 18050 16759 18106 16768
rect 16578 16510 16896 16538
rect 15290 16416 15346 16425
rect 12084 16374 12204 16400
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 12070 14716 12378 14736
rect 12070 14714 12076 14716
rect 12132 14714 12156 14716
rect 12212 14714 12236 14716
rect 12292 14714 12316 14716
rect 12372 14714 12378 14716
rect 12132 14662 12134 14714
rect 12314 14662 12316 14714
rect 12070 14660 12076 14662
rect 12132 14660 12156 14662
rect 12212 14660 12236 14662
rect 12292 14660 12316 14662
rect 12372 14660 12378 14662
rect 12070 14640 12378 14660
rect 13084 14408 13136 14414
rect 13084 14350 13136 14356
rect 13096 14006 13124 14350
rect 13084 14000 13136 14006
rect 13084 13942 13136 13948
rect 12070 13628 12378 13648
rect 12070 13626 12076 13628
rect 12132 13626 12156 13628
rect 12212 13626 12236 13628
rect 12292 13626 12316 13628
rect 12372 13626 12378 13628
rect 12132 13574 12134 13626
rect 12314 13574 12316 13626
rect 12070 13572 12076 13574
rect 12132 13572 12156 13574
rect 12212 13572 12236 13574
rect 12292 13572 12316 13574
rect 12372 13572 12378 13574
rect 12070 13552 12378 13572
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 12164 13320 12216 13326
rect 12164 13262 12216 13268
rect 10968 12912 11020 12918
rect 10968 12854 11020 12860
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 10600 12096 10652 12102
rect 10600 12038 10652 12044
rect 10784 12096 10836 12102
rect 10784 12038 10836 12044
rect 9784 11898 9812 12038
rect 9846 11996 10154 12016
rect 9846 11994 9852 11996
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 10148 11994 10154 11996
rect 9908 11942 9910 11994
rect 10090 11942 10092 11994
rect 9846 11940 9852 11942
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 10148 11940 10154 11942
rect 9846 11920 10154 11940
rect 10506 11928 10562 11937
rect 9772 11892 9824 11898
rect 10506 11863 10562 11872
rect 9772 11834 9824 11840
rect 10520 11762 10548 11863
rect 10508 11756 10560 11762
rect 10152 11716 10364 11744
rect 9680 11688 9732 11694
rect 9680 11630 9732 11636
rect 10152 11626 10180 11716
rect 10336 11676 10364 11716
rect 10508 11698 10560 11704
rect 10416 11688 10468 11694
rect 10336 11648 10416 11676
rect 10416 11630 10468 11636
rect 10140 11620 10192 11626
rect 10140 11562 10192 11568
rect 10232 11620 10284 11626
rect 10232 11562 10284 11568
rect 9954 11384 10010 11393
rect 9404 11348 9456 11354
rect 10244 11354 10272 11562
rect 10506 11520 10562 11529
rect 10506 11455 10562 11464
rect 9954 11319 10010 11328
rect 10232 11348 10284 11354
rect 9404 11290 9456 11296
rect 9220 11280 9272 11286
rect 9220 11222 9272 11228
rect 9232 11082 9260 11222
rect 9968 11218 9996 11319
rect 10232 11290 10284 11296
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9220 11076 9272 11082
rect 9220 11018 9272 11024
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8850 10160 8906 10169
rect 8850 10095 8906 10104
rect 8864 9926 8892 10095
rect 9048 9926 9076 10950
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8852 9920 8904 9926
rect 8852 9862 8904 9868
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 8496 9646 8616 9674
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8392 9376 8444 9382
rect 8392 9318 8444 9324
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8116 8424 8168 8430
rect 8116 8366 8168 8372
rect 7380 6792 7432 6798
rect 7380 6734 7432 6740
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 6322 7420 6598
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7392 6118 7420 6258
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7380 6112 7432 6118
rect 7484 6089 7512 6190
rect 7944 6186 7972 6326
rect 7932 6180 7984 6186
rect 7932 6122 7984 6128
rect 7380 6054 7432 6060
rect 7470 6080 7526 6089
rect 7470 6015 7526 6024
rect 7622 6012 7930 6032
rect 7622 6010 7628 6012
rect 7684 6010 7708 6012
rect 7764 6010 7788 6012
rect 7844 6010 7868 6012
rect 7924 6010 7930 6012
rect 7684 5958 7686 6010
rect 7866 5958 7868 6010
rect 7622 5956 7628 5958
rect 7684 5956 7708 5958
rect 7764 5956 7788 5958
rect 7844 5956 7868 5958
rect 7924 5956 7930 5958
rect 7622 5936 7930 5956
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7196 5228 7248 5234
rect 7196 5170 7248 5176
rect 7194 4992 7250 5001
rect 7194 4927 7250 4936
rect 7208 4826 7236 4927
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7392 4690 7420 5850
rect 7472 5840 7524 5846
rect 8036 5794 8064 6734
rect 8128 6458 8156 8366
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 8114 6352 8170 6361
rect 8114 6287 8170 6296
rect 8128 6254 8156 6287
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 8220 5914 8248 6734
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 7524 5788 7604 5794
rect 7472 5782 7604 5788
rect 7484 5766 7604 5782
rect 8036 5766 8248 5794
rect 7472 5568 7524 5574
rect 7576 5545 7604 5766
rect 7472 5510 7524 5516
rect 7562 5536 7618 5545
rect 7484 5166 7512 5510
rect 7562 5471 7618 5480
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 8116 5092 8168 5098
rect 8116 5034 8168 5040
rect 7622 4924 7930 4944
rect 7622 4922 7628 4924
rect 7684 4922 7708 4924
rect 7764 4922 7788 4924
rect 7844 4922 7868 4924
rect 7924 4922 7930 4924
rect 7684 4870 7686 4922
rect 7866 4870 7868 4922
rect 7622 4868 7628 4870
rect 7684 4868 7708 4870
rect 7764 4868 7788 4870
rect 7844 4868 7868 4870
rect 7924 4868 7930 4870
rect 7622 4848 7930 4868
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7196 4480 7248 4486
rect 7196 4422 7248 4428
rect 7208 3942 7236 4422
rect 7392 4214 7420 4626
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7196 3936 7248 3942
rect 7248 3884 7328 3890
rect 7196 3878 7328 3884
rect 7208 3862 7328 3878
rect 7300 3602 7328 3862
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 7104 2848 7156 2854
rect 7104 2790 7156 2796
rect 7116 2514 7144 2790
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7208 1494 7236 3334
rect 7300 2854 7328 3538
rect 7380 3460 7432 3466
rect 7380 3402 7432 3408
rect 7392 3194 7420 3402
rect 7484 3369 7512 4422
rect 7622 3836 7930 3856
rect 7622 3834 7628 3836
rect 7684 3834 7708 3836
rect 7764 3834 7788 3836
rect 7844 3834 7868 3836
rect 7924 3834 7930 3836
rect 7684 3782 7686 3834
rect 7866 3782 7868 3834
rect 7622 3780 7628 3782
rect 7684 3780 7708 3782
rect 7764 3780 7788 3782
rect 7844 3780 7868 3782
rect 7924 3780 7930 3782
rect 7622 3760 7930 3780
rect 8036 3398 8064 4558
rect 8128 4486 8156 5034
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8220 4146 8248 5766
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8116 4072 8168 4078
rect 8116 4014 8168 4020
rect 8024 3392 8076 3398
rect 7470 3360 7526 3369
rect 8024 3334 8076 3340
rect 7470 3295 7526 3304
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 7378 3088 7434 3097
rect 7378 3023 7380 3032
rect 7432 3023 7434 3032
rect 7654 3088 7710 3097
rect 7654 3023 7656 3032
rect 7380 2994 7432 3000
rect 7708 3023 7710 3032
rect 7656 2994 7708 3000
rect 7564 2984 7616 2990
rect 7484 2932 7564 2938
rect 7484 2926 7616 2932
rect 7484 2910 7604 2926
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7484 2514 7512 2910
rect 7622 2748 7930 2768
rect 7622 2746 7628 2748
rect 7684 2746 7708 2748
rect 7764 2746 7788 2748
rect 7844 2746 7868 2748
rect 7924 2746 7930 2748
rect 7684 2694 7686 2746
rect 7866 2694 7868 2746
rect 7622 2692 7628 2694
rect 7684 2692 7708 2694
rect 7764 2692 7788 2694
rect 7844 2692 7868 2694
rect 7924 2692 7930 2694
rect 7622 2672 7930 2692
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7484 1698 7512 2246
rect 8128 1902 8156 4014
rect 8312 2514 8340 8502
rect 8404 7954 8432 9318
rect 8496 9178 8524 9454
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8588 9058 8616 9646
rect 8496 9030 8616 9058
rect 8496 8362 8524 9030
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8392 7200 8444 7206
rect 8392 7142 8444 7148
rect 8404 5710 8432 7142
rect 8496 6361 8524 8298
rect 8588 7954 8616 8570
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8588 7478 8616 7890
rect 8576 7472 8628 7478
rect 8680 7449 8708 9862
rect 8864 9382 8892 9862
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8852 9376 8904 9382
rect 8852 9318 8904 9324
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 8576 7414 8628 7420
rect 8666 7440 8722 7449
rect 8666 7375 8722 7384
rect 8772 6458 8800 8434
rect 8864 8294 8892 9318
rect 8956 9110 8984 9590
rect 8944 9104 8996 9110
rect 8944 9046 8996 9052
rect 8852 8288 8904 8294
rect 8852 8230 8904 8236
rect 9048 7313 9076 9862
rect 9128 9512 9180 9518
rect 9128 9454 9180 9460
rect 9140 9382 9168 9454
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9232 8022 9260 11018
rect 9846 10908 10154 10928
rect 9846 10906 9852 10908
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 10148 10906 10154 10908
rect 9908 10854 9910 10906
rect 10090 10854 10092 10906
rect 9846 10852 9852 10854
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 10148 10852 10154 10854
rect 9846 10832 10154 10852
rect 10048 10464 10100 10470
rect 10048 10406 10100 10412
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9312 10192 9364 10198
rect 9312 10134 9364 10140
rect 9324 9586 9352 10134
rect 9416 9994 9444 10202
rect 10060 10130 10088 10406
rect 10520 10169 10548 11455
rect 10612 11354 10640 12038
rect 10796 11898 10824 12038
rect 10784 11892 10836 11898
rect 10784 11834 10836 11840
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10796 11393 10824 11698
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10782 11384 10838 11393
rect 10600 11348 10652 11354
rect 10782 11319 10838 11328
rect 10600 11290 10652 11296
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 10704 10810 10732 11018
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10888 10674 10916 11630
rect 10876 10668 10928 10674
rect 10704 10628 10876 10656
rect 10506 10160 10562 10169
rect 10048 10124 10100 10130
rect 10506 10095 10562 10104
rect 10048 10066 10100 10072
rect 10230 10024 10286 10033
rect 9404 9988 9456 9994
rect 10230 9959 10232 9968
rect 9404 9930 9456 9936
rect 10284 9959 10286 9968
rect 10232 9930 10284 9936
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9600 9722 9628 9862
rect 9846 9820 10154 9840
rect 9846 9818 9852 9820
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 10148 9818 10154 9820
rect 9908 9766 9910 9818
rect 10090 9766 10092 9818
rect 9846 9764 9852 9766
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 10148 9764 10154 9766
rect 9846 9744 10154 9764
rect 10244 9722 10272 9930
rect 9588 9716 9640 9722
rect 9588 9658 9640 9664
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10520 9674 10548 10095
rect 10520 9646 10640 9674
rect 9312 9580 9364 9586
rect 9364 9540 9536 9568
rect 9312 9522 9364 9528
rect 9404 9104 9456 9110
rect 9404 9046 9456 9052
rect 9416 8838 9444 9046
rect 9404 8832 9456 8838
rect 9402 8800 9404 8809
rect 9456 8800 9458 8809
rect 9402 8735 9458 8744
rect 9220 8016 9272 8022
rect 9272 7964 9444 7970
rect 9220 7958 9444 7964
rect 9232 7942 9444 7958
rect 9416 7886 9444 7942
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9034 7304 9090 7313
rect 9034 7239 9090 7248
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8760 6452 8812 6458
rect 8760 6394 8812 6400
rect 8576 6384 8628 6390
rect 8482 6352 8538 6361
rect 8576 6326 8628 6332
rect 8482 6287 8538 6296
rect 8588 6168 8616 6326
rect 8496 6140 8616 6168
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8392 5296 8444 5302
rect 8392 5238 8444 5244
rect 8404 4282 8432 5238
rect 8496 5166 8524 6140
rect 8574 6080 8630 6089
rect 8574 6015 8630 6024
rect 8588 5574 8616 6015
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8484 5160 8536 5166
rect 8484 5102 8536 5108
rect 8588 4468 8616 5510
rect 8680 5370 8708 6394
rect 8772 5953 8800 6394
rect 8850 6352 8906 6361
rect 8850 6287 8906 6296
rect 8758 5944 8814 5953
rect 8864 5914 8892 6287
rect 8956 6254 8984 6870
rect 9508 6866 9536 9540
rect 9588 9376 9640 9382
rect 9588 9318 9640 9324
rect 10140 9376 10192 9382
rect 10192 9336 10272 9364
rect 10140 9318 10192 9324
rect 9600 9042 9628 9318
rect 9954 9072 10010 9081
rect 9588 9036 9640 9042
rect 10244 9042 10272 9336
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 9954 9007 10010 9016
rect 10232 9036 10284 9042
rect 9588 8978 9640 8984
rect 9968 8974 9996 9007
rect 10232 8978 10284 8984
rect 9956 8968 10008 8974
rect 9956 8910 10008 8916
rect 9588 8832 9640 8838
rect 9588 8774 9640 8780
rect 9600 7818 9628 8774
rect 9846 8732 10154 8752
rect 9846 8730 9852 8732
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 10148 8730 10154 8732
rect 9908 8678 9910 8730
rect 10090 8678 10092 8730
rect 9846 8676 9852 8678
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 10148 8676 10154 8678
rect 9846 8656 10154 8676
rect 10244 8498 10272 8978
rect 10520 8838 10548 9046
rect 10508 8832 10560 8838
rect 10506 8800 10508 8809
rect 10560 8800 10562 8809
rect 10506 8735 10562 8744
rect 9864 8492 9916 8498
rect 9864 8434 9916 8440
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9678 7984 9734 7993
rect 9678 7919 9680 7928
rect 9732 7919 9734 7928
rect 9680 7890 9732 7896
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9692 7750 9720 7890
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9784 7410 9812 8366
rect 9876 8022 9904 8434
rect 9864 8016 9916 8022
rect 9864 7958 9916 7964
rect 10508 7744 10560 7750
rect 10506 7712 10508 7721
rect 10560 7712 10562 7721
rect 9846 7644 10154 7664
rect 10506 7647 10562 7656
rect 9846 7642 9852 7644
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 10148 7642 10154 7644
rect 9908 7590 9910 7642
rect 10090 7590 10092 7642
rect 9846 7588 9852 7590
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 10148 7588 10154 7590
rect 9846 7568 10154 7588
rect 10520 7449 10548 7647
rect 10506 7440 10562 7449
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 10048 7404 10100 7410
rect 10506 7375 10562 7384
rect 10048 7346 10100 7352
rect 10060 7002 10088 7346
rect 10612 7324 10640 9646
rect 10520 7296 10640 7324
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8758 5879 8814 5888
rect 8852 5908 8904 5914
rect 8852 5850 8904 5856
rect 9048 5642 9076 6802
rect 9128 6724 9180 6730
rect 9128 6666 9180 6672
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 8760 5568 8812 5574
rect 8944 5568 8996 5574
rect 8760 5510 8812 5516
rect 8942 5536 8944 5545
rect 8996 5536 8998 5545
rect 8668 5364 8720 5370
rect 8668 5306 8720 5312
rect 8668 4480 8720 4486
rect 8588 4440 8668 4468
rect 8668 4422 8720 4428
rect 8392 4276 8444 4282
rect 8392 4218 8444 4224
rect 8576 4072 8628 4078
rect 8390 4040 8446 4049
rect 8390 3975 8392 3984
rect 8444 3975 8446 3984
rect 8574 4040 8576 4049
rect 8628 4040 8630 4049
rect 8680 4010 8708 4422
rect 8772 4282 8800 5510
rect 8942 5471 8998 5480
rect 9036 4616 9088 4622
rect 9036 4558 9088 4564
rect 8760 4276 8812 4282
rect 8760 4218 8812 4224
rect 8574 3975 8630 3984
rect 8668 4004 8720 4010
rect 8392 3946 8444 3952
rect 8668 3946 8720 3952
rect 9048 3738 9076 4558
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 8390 3496 8446 3505
rect 8390 3431 8446 3440
rect 8404 3398 8432 3431
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8484 2916 8536 2922
rect 8484 2858 8536 2864
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8116 1896 8168 1902
rect 8116 1838 8168 1844
rect 7472 1692 7524 1698
rect 7472 1634 7524 1640
rect 7196 1488 7248 1494
rect 7196 1430 7248 1436
rect 7484 870 7604 898
rect 7484 762 7512 870
rect 7576 800 7604 870
rect 8496 800 8524 2858
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8772 2446 8800 2790
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 9140 2106 9168 6666
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9232 5681 9260 6598
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9324 6089 9352 6190
rect 9310 6080 9366 6089
rect 9310 6015 9366 6024
rect 9218 5672 9274 5681
rect 9218 5607 9274 5616
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9312 4548 9364 4554
rect 9312 4490 9364 4496
rect 9218 4176 9274 4185
rect 9218 4111 9274 4120
rect 9232 4010 9260 4111
rect 9220 4004 9272 4010
rect 9220 3946 9272 3952
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9232 2514 9260 2790
rect 9324 2774 9352 4490
rect 9416 3602 9444 4966
rect 9508 4146 9536 6802
rect 9846 6556 10154 6576
rect 9846 6554 9852 6556
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 10148 6554 10154 6556
rect 9908 6502 9910 6554
rect 10090 6502 10092 6554
rect 9846 6500 9852 6502
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 10148 6500 10154 6502
rect 9846 6480 10154 6500
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 9600 5817 9628 6054
rect 9586 5808 9642 5817
rect 9586 5743 9642 5752
rect 9846 5468 10154 5488
rect 9846 5466 9852 5468
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 10148 5466 10154 5468
rect 9908 5414 9910 5466
rect 10090 5414 10092 5466
rect 9846 5412 9852 5414
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 10148 5412 10154 5414
rect 9846 5392 10154 5412
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9692 5250 9720 5306
rect 9600 5222 9720 5250
rect 10138 5264 10194 5273
rect 9772 5228 9824 5234
rect 9600 4622 9628 5222
rect 10138 5199 10194 5208
rect 9772 5170 9824 5176
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9496 4140 9548 4146
rect 9496 4082 9548 4088
rect 9508 4049 9536 4082
rect 9494 4040 9550 4049
rect 9494 3975 9550 3984
rect 9600 3738 9628 4558
rect 9692 4486 9720 5102
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9784 4026 9812 5170
rect 10152 4468 10180 5199
rect 10244 5166 10272 6054
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 10244 4622 10272 5102
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 10324 4480 10376 4486
rect 10152 4440 10272 4468
rect 9846 4380 10154 4400
rect 9846 4378 9852 4380
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 10148 4378 10154 4380
rect 9908 4326 9910 4378
rect 10090 4326 10092 4378
rect 9846 4324 9852 4326
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 10148 4324 10154 4326
rect 9846 4304 10154 4324
rect 9784 3998 9904 4026
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9404 3596 9456 3602
rect 9404 3538 9456 3544
rect 9692 3534 9720 3878
rect 9876 3738 9904 3998
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9680 3528 9732 3534
rect 9680 3470 9732 3476
rect 9846 3292 10154 3312
rect 9846 3290 9852 3292
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 10148 3290 10154 3292
rect 9908 3238 9910 3290
rect 10090 3238 10092 3290
rect 9846 3236 9852 3238
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 10148 3236 10154 3238
rect 9846 3216 10154 3236
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9324 2746 9444 2774
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9128 2100 9180 2106
rect 9128 2042 9180 2048
rect 9416 800 9444 2746
rect 9692 2446 9720 2994
rect 10244 2650 10272 4440
rect 10324 4422 10376 4428
rect 10336 4214 10364 4422
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10324 3936 10376 3942
rect 10324 3878 10376 3884
rect 10336 3602 10364 3878
rect 10324 3596 10376 3602
rect 10324 3538 10376 3544
rect 10428 3534 10456 6938
rect 10520 3777 10548 7296
rect 10704 5370 10732 10628
rect 10876 10610 10928 10616
rect 10980 10266 11008 12854
rect 12176 12782 12204 13262
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 12164 12776 12216 12782
rect 12216 12736 12480 12764
rect 12164 12718 12216 12724
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11072 10606 11100 12582
rect 11150 12336 11206 12345
rect 11150 12271 11206 12280
rect 11164 11234 11192 12271
rect 11336 12232 11388 12238
rect 11388 12192 11468 12220
rect 11336 12174 11388 12180
rect 11164 11218 11284 11234
rect 11164 11212 11296 11218
rect 11164 11206 11244 11212
rect 11164 10810 11192 11206
rect 11244 11154 11296 11160
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11060 10600 11112 10606
rect 11060 10542 11112 10548
rect 10968 10260 11020 10266
rect 10968 10202 11020 10208
rect 10784 10124 10836 10130
rect 10784 10066 10836 10072
rect 10796 9586 10824 10066
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10796 9042 10824 9522
rect 10888 9382 10916 9998
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10888 8634 10916 9318
rect 11336 8900 11388 8906
rect 11336 8842 11388 8848
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 10876 8628 10928 8634
rect 10928 8588 11100 8616
rect 10876 8570 10928 8576
rect 10966 8392 11022 8401
rect 10966 8327 11022 8336
rect 10980 7954 11008 8327
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10968 6996 11020 7002
rect 10968 6938 11020 6944
rect 10980 6497 11008 6938
rect 10966 6488 11022 6497
rect 10966 6423 11022 6432
rect 11072 5710 11100 8588
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11164 7857 11192 8298
rect 11256 7886 11284 8774
rect 11348 8566 11376 8842
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11244 7880 11296 7886
rect 11150 7848 11206 7857
rect 11244 7822 11296 7828
rect 11150 7783 11206 7792
rect 11348 6866 11376 8366
rect 11336 6860 11388 6866
rect 11336 6802 11388 6808
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11256 6361 11284 6734
rect 11242 6352 11298 6361
rect 11152 6316 11204 6322
rect 11348 6322 11376 6802
rect 11440 6746 11468 12192
rect 11520 12096 11572 12102
rect 11520 12038 11572 12044
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11532 11626 11560 12038
rect 11716 11694 11744 12038
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11520 11620 11572 11626
rect 11520 11562 11572 11568
rect 11716 11354 11744 11630
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11532 10674 11560 11086
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11532 10130 11560 10610
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11624 9024 11652 11086
rect 11808 10198 11836 12582
rect 12070 12540 12378 12560
rect 12070 12538 12076 12540
rect 12132 12538 12156 12540
rect 12212 12538 12236 12540
rect 12292 12538 12316 12540
rect 12372 12538 12378 12540
rect 12132 12486 12134 12538
rect 12314 12486 12316 12538
rect 12070 12484 12076 12486
rect 12132 12484 12156 12486
rect 12212 12484 12236 12486
rect 12292 12484 12316 12486
rect 12372 12484 12378 12486
rect 12070 12464 12378 12484
rect 12452 12238 12480 12736
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 11886 11928 11942 11937
rect 11886 11863 11888 11872
rect 11940 11863 11942 11872
rect 12438 11928 12494 11937
rect 12438 11863 12494 11872
rect 12532 11892 12584 11898
rect 11888 11834 11940 11840
rect 12070 11452 12378 11472
rect 12070 11450 12076 11452
rect 12132 11450 12156 11452
rect 12212 11450 12236 11452
rect 12292 11450 12316 11452
rect 12372 11450 12378 11452
rect 12132 11398 12134 11450
rect 12314 11398 12316 11450
rect 12070 11396 12076 11398
rect 12132 11396 12156 11398
rect 12212 11396 12236 11398
rect 12292 11396 12316 11398
rect 12372 11396 12378 11398
rect 11886 11384 11942 11393
rect 12070 11376 12378 11396
rect 11886 11319 11942 11328
rect 11900 11014 11928 11319
rect 12254 11112 12310 11121
rect 12254 11047 12256 11056
rect 12308 11047 12310 11056
rect 12256 11018 12308 11024
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 11624 8996 11836 9024
rect 11702 8936 11758 8945
rect 11702 8871 11704 8880
rect 11756 8871 11758 8880
rect 11704 8842 11756 8848
rect 11520 8832 11572 8838
rect 11520 8774 11572 8780
rect 11532 8537 11560 8774
rect 11716 8537 11744 8842
rect 11518 8528 11574 8537
rect 11518 8463 11574 8472
rect 11702 8528 11758 8537
rect 11702 8463 11758 8472
rect 11704 7948 11756 7954
rect 11704 7890 11756 7896
rect 11612 7812 11664 7818
rect 11612 7754 11664 7760
rect 11624 7342 11652 7754
rect 11716 7478 11744 7890
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 11808 7426 11836 8996
rect 11900 8945 11928 10950
rect 12070 10364 12378 10384
rect 12070 10362 12076 10364
rect 12132 10362 12156 10364
rect 12212 10362 12236 10364
rect 12292 10362 12316 10364
rect 12372 10362 12378 10364
rect 12132 10310 12134 10362
rect 12314 10310 12316 10362
rect 12070 10308 12076 10310
rect 12132 10308 12156 10310
rect 12212 10308 12236 10310
rect 12292 10308 12316 10310
rect 12372 10308 12378 10310
rect 12070 10288 12378 10308
rect 11980 10124 12032 10130
rect 11980 10066 12032 10072
rect 11992 9450 12020 10066
rect 12348 9920 12400 9926
rect 12348 9862 12400 9868
rect 12072 9512 12124 9518
rect 12070 9480 12072 9489
rect 12124 9480 12126 9489
rect 11980 9444 12032 9450
rect 12360 9450 12388 9862
rect 12070 9415 12126 9424
rect 12348 9444 12400 9450
rect 11980 9386 12032 9392
rect 12348 9386 12400 9392
rect 11992 8974 12020 9386
rect 12070 9276 12378 9296
rect 12070 9274 12076 9276
rect 12132 9274 12156 9276
rect 12212 9274 12236 9276
rect 12292 9274 12316 9276
rect 12372 9274 12378 9276
rect 12132 9222 12134 9274
rect 12314 9222 12316 9274
rect 12070 9220 12076 9222
rect 12132 9220 12156 9222
rect 12212 9220 12236 9222
rect 12292 9220 12316 9222
rect 12372 9220 12378 9222
rect 12070 9200 12378 9220
rect 11980 8968 12032 8974
rect 11886 8936 11942 8945
rect 11980 8910 12032 8916
rect 11886 8871 11942 8880
rect 12348 8832 12400 8838
rect 12452 8820 12480 11863
rect 12532 11834 12584 11840
rect 12544 11529 12572 11834
rect 12530 11520 12586 11529
rect 12530 11455 12586 11464
rect 12624 11280 12676 11286
rect 12624 11222 12676 11228
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12544 10470 12572 10542
rect 12532 10464 12584 10470
rect 12532 10406 12584 10412
rect 12544 9654 12572 10406
rect 12636 10062 12664 11222
rect 12900 11212 12952 11218
rect 12900 11154 12952 11160
rect 12808 11008 12860 11014
rect 12808 10950 12860 10956
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12728 10266 12756 10678
rect 12820 10266 12848 10950
rect 12912 10606 12940 11154
rect 13004 10674 13032 12174
rect 13096 11762 13124 12922
rect 13084 11756 13136 11762
rect 13084 11698 13136 11704
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 13096 11257 13124 11494
rect 13082 11248 13138 11257
rect 13082 11183 13138 11192
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12808 10260 12860 10266
rect 12808 10202 12860 10208
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12728 9908 12756 10202
rect 13004 10198 13032 10610
rect 12992 10192 13044 10198
rect 12992 10134 13044 10140
rect 13096 9926 13124 11183
rect 12636 9880 12756 9908
rect 12992 9920 13044 9926
rect 12532 9648 12584 9654
rect 12532 9590 12584 9596
rect 12400 8792 12480 8820
rect 12348 8774 12400 8780
rect 12070 8188 12378 8208
rect 12070 8186 12076 8188
rect 12132 8186 12156 8188
rect 12212 8186 12236 8188
rect 12292 8186 12316 8188
rect 12372 8186 12378 8188
rect 12132 8134 12134 8186
rect 12314 8134 12316 8186
rect 12070 8132 12076 8134
rect 12132 8132 12156 8134
rect 12212 8132 12236 8134
rect 12292 8132 12316 8134
rect 12372 8132 12378 8134
rect 12070 8112 12378 8132
rect 12452 8022 12480 8792
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12544 8090 12572 8434
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12440 8016 12492 8022
rect 12440 7958 12492 7964
rect 12636 7970 12664 9880
rect 12992 9862 13044 9868
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13004 9761 13032 9862
rect 12990 9752 13046 9761
rect 12990 9687 13046 9696
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 12728 9110 12756 9590
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12716 9104 12768 9110
rect 12820 9081 12848 9522
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13096 9178 13124 9454
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 12716 9046 12768 9052
rect 12806 9072 12862 9081
rect 12806 9007 12862 9016
rect 12820 8276 12848 9007
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12912 8634 12940 8842
rect 12990 8800 13046 8809
rect 12990 8735 13046 8744
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12912 8430 12940 8570
rect 13004 8498 13032 8735
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12820 8248 12940 8276
rect 12636 7942 12848 7970
rect 12532 7472 12584 7478
rect 11808 7398 11928 7426
rect 12532 7414 12584 7420
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11808 7002 11836 7278
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11900 6746 11928 7398
rect 12440 7336 12492 7342
rect 12440 7278 12492 7284
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11440 6718 11652 6746
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11242 6287 11298 6296
rect 11336 6316 11388 6322
rect 11152 6258 11204 6264
rect 11336 6258 11388 6264
rect 11060 5704 11112 5710
rect 11060 5646 11112 5652
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 10600 5296 10652 5302
rect 10600 5238 10652 5244
rect 10506 3768 10562 3777
rect 10506 3703 10562 3712
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10520 3194 10548 3703
rect 10612 3194 10640 5238
rect 10704 5098 10732 5306
rect 10980 5166 11008 5510
rect 10968 5160 11020 5166
rect 10968 5102 11020 5108
rect 10692 5092 10744 5098
rect 10692 5034 10744 5040
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10704 3738 10732 4762
rect 10980 4758 11008 5102
rect 11164 4826 11192 6258
rect 11348 5914 11376 6258
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10782 4176 10838 4185
rect 10782 4111 10784 4120
rect 10836 4111 10838 4120
rect 10784 4082 10836 4088
rect 10692 3732 10744 3738
rect 10692 3674 10744 3680
rect 10508 3188 10560 3194
rect 10508 3130 10560 3136
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 10232 2644 10284 2650
rect 10232 2586 10284 2592
rect 10230 2544 10286 2553
rect 9956 2508 10008 2514
rect 9784 2468 9956 2496
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9784 1766 9812 2468
rect 10230 2479 10286 2488
rect 9956 2450 10008 2456
rect 10244 2281 10272 2479
rect 10230 2272 10286 2281
rect 9846 2204 10154 2224
rect 10230 2207 10286 2216
rect 9846 2202 9852 2204
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 10148 2202 10154 2204
rect 9908 2150 9910 2202
rect 10090 2150 10092 2202
rect 9846 2148 9852 2150
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 10148 2148 10154 2150
rect 9846 2128 10154 2148
rect 9772 1760 9824 1766
rect 9772 1702 9824 1708
rect 10336 800 10364 3062
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10428 2038 10456 2994
rect 10796 2774 10824 4082
rect 10888 4010 10916 4558
rect 11152 4548 11204 4554
rect 11152 4490 11204 4496
rect 11060 4480 11112 4486
rect 11060 4422 11112 4428
rect 11072 4282 11100 4422
rect 11164 4282 11192 4490
rect 11060 4276 11112 4282
rect 11060 4218 11112 4224
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 10968 4072 11020 4078
rect 10968 4014 11020 4020
rect 10876 4004 10928 4010
rect 10876 3946 10928 3952
rect 10888 3602 10916 3946
rect 10980 3738 11008 4014
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 11058 3632 11114 3641
rect 10876 3596 10928 3602
rect 11058 3567 11060 3576
rect 10876 3538 10928 3544
rect 11112 3567 11114 3576
rect 11060 3538 11112 3544
rect 11058 3496 11114 3505
rect 11256 3482 11284 4966
rect 11058 3431 11060 3440
rect 11112 3431 11114 3440
rect 11164 3454 11284 3482
rect 11060 3402 11112 3408
rect 11164 3346 11192 3454
rect 11348 3398 11376 5578
rect 11440 3466 11468 6598
rect 11624 6458 11652 6718
rect 11808 6718 11928 6746
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11624 6322 11652 6394
rect 11612 6316 11664 6322
rect 11612 6258 11664 6264
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11532 4622 11560 5102
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11532 4078 11560 4558
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11532 3602 11560 4014
rect 11520 3596 11572 3602
rect 11520 3538 11572 3544
rect 11612 3528 11664 3534
rect 11808 3482 11836 6718
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11900 6458 11928 6598
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11888 5024 11940 5030
rect 11888 4966 11940 4972
rect 11900 4690 11928 4966
rect 11992 4808 12020 7142
rect 12070 7100 12378 7120
rect 12070 7098 12076 7100
rect 12132 7098 12156 7100
rect 12212 7098 12236 7100
rect 12292 7098 12316 7100
rect 12372 7098 12378 7100
rect 12132 7046 12134 7098
rect 12314 7046 12316 7098
rect 12070 7044 12076 7046
rect 12132 7044 12156 7046
rect 12212 7044 12236 7046
rect 12292 7044 12316 7046
rect 12372 7044 12378 7046
rect 12070 7024 12378 7044
rect 12452 6934 12480 7278
rect 12440 6928 12492 6934
rect 12440 6870 12492 6876
rect 12544 6798 12572 7414
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12728 7002 12756 7346
rect 12716 6996 12768 7002
rect 12716 6938 12768 6944
rect 12624 6928 12676 6934
rect 12624 6870 12676 6876
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12164 6656 12216 6662
rect 12164 6598 12216 6604
rect 12176 6458 12204 6598
rect 12164 6452 12216 6458
rect 12164 6394 12216 6400
rect 12544 6390 12572 6734
rect 12532 6384 12584 6390
rect 12532 6326 12584 6332
rect 12348 6316 12400 6322
rect 12348 6258 12400 6264
rect 12360 6225 12388 6258
rect 12346 6216 12402 6225
rect 12346 6151 12402 6160
rect 12070 6012 12378 6032
rect 12070 6010 12076 6012
rect 12132 6010 12156 6012
rect 12212 6010 12236 6012
rect 12292 6010 12316 6012
rect 12372 6010 12378 6012
rect 12132 5958 12134 6010
rect 12314 5958 12316 6010
rect 12070 5956 12076 5958
rect 12132 5956 12156 5958
rect 12212 5956 12236 5958
rect 12292 5956 12316 5958
rect 12372 5956 12378 5958
rect 12070 5936 12378 5956
rect 12636 5914 12664 6870
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12820 5250 12848 7942
rect 12912 7750 12940 8248
rect 13188 8090 13216 15302
rect 13268 15224 13320 15230
rect 13268 15166 13320 15172
rect 13280 11801 13308 15166
rect 14384 14362 14412 16400
rect 16578 16400 16634 16510
rect 15290 16351 15346 16360
rect 15198 16008 15254 16017
rect 15198 15943 15254 15952
rect 15212 15230 15240 15943
rect 15200 15224 15252 15230
rect 15200 15166 15252 15172
rect 15304 14482 15332 16351
rect 15934 15600 15990 15609
rect 15934 15535 15990 15544
rect 15292 14476 15344 14482
rect 15292 14418 15344 14424
rect 14200 14334 14412 14362
rect 14200 14006 14228 14334
rect 15672 14278 15700 14309
rect 15660 14272 15712 14278
rect 15658 14240 15660 14249
rect 15712 14240 15714 14249
rect 14294 14172 14602 14192
rect 15658 14175 15714 14184
rect 14294 14170 14300 14172
rect 14356 14170 14380 14172
rect 14436 14170 14460 14172
rect 14516 14170 14540 14172
rect 14596 14170 14602 14172
rect 14356 14118 14358 14170
rect 14538 14118 14540 14170
rect 14294 14116 14300 14118
rect 14356 14116 14380 14118
rect 14436 14116 14460 14118
rect 14516 14116 14540 14118
rect 14596 14116 14602 14118
rect 14294 14096 14602 14116
rect 15198 14104 15254 14113
rect 15198 14039 15200 14048
rect 15252 14039 15254 14048
rect 15200 14010 15252 14016
rect 14188 14000 14240 14006
rect 14188 13942 14240 13948
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13452 13864 13504 13870
rect 13452 13806 13504 13812
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13464 12345 13492 13806
rect 13556 12986 13584 13806
rect 13648 13530 13676 13874
rect 13726 13832 13782 13841
rect 13726 13767 13782 13776
rect 13636 13524 13688 13530
rect 13636 13466 13688 13472
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13450 12336 13506 12345
rect 13450 12271 13506 12280
rect 13464 12238 13492 12271
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13266 11792 13322 11801
rect 13266 11727 13322 11736
rect 13280 11558 13308 11727
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13280 11218 13308 11494
rect 13268 11212 13320 11218
rect 13268 11154 13320 11160
rect 13464 10010 13492 12174
rect 13556 11694 13584 12922
rect 13740 12209 13768 13767
rect 14740 13728 14792 13734
rect 14740 13670 14792 13676
rect 14752 13258 14780 13670
rect 15120 13394 15148 13942
rect 15568 13796 15620 13802
rect 15568 13738 15620 13744
rect 15108 13388 15160 13394
rect 15108 13330 15160 13336
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 14740 13252 14792 13258
rect 14740 13194 14792 13200
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13832 12782 13860 12854
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13726 12200 13782 12209
rect 13648 12158 13726 12186
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 13280 9982 13492 10010
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 12900 7744 12952 7750
rect 13188 7721 13216 8026
rect 12900 7686 12952 7692
rect 13174 7712 13230 7721
rect 12912 7002 12940 7686
rect 13174 7647 13230 7656
rect 13084 7268 13136 7274
rect 13084 7210 13136 7216
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 13096 6798 13124 7210
rect 13084 6792 13136 6798
rect 13084 6734 13136 6740
rect 13280 6662 13308 9982
rect 13360 9920 13412 9926
rect 13360 9862 13412 9868
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13372 7449 13400 9862
rect 13450 9480 13506 9489
rect 13450 9415 13452 9424
rect 13504 9415 13506 9424
rect 13452 9386 13504 9392
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13464 8090 13492 8502
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 13464 7834 13492 8026
rect 13556 7993 13584 9862
rect 13542 7984 13598 7993
rect 13542 7919 13598 7928
rect 13464 7806 13584 7834
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13358 7440 13414 7449
rect 13358 7375 13414 7384
rect 13464 6934 13492 7686
rect 13452 6928 13504 6934
rect 13452 6870 13504 6876
rect 13360 6860 13412 6866
rect 13360 6802 13412 6808
rect 13372 6730 13400 6802
rect 13556 6798 13584 7806
rect 13648 7546 13676 12158
rect 13726 12135 13782 12144
rect 14016 11762 14044 13126
rect 14294 13084 14602 13104
rect 14294 13082 14300 13084
rect 14356 13082 14380 13084
rect 14436 13082 14460 13084
rect 14516 13082 14540 13084
rect 14596 13082 14602 13084
rect 14356 13030 14358 13082
rect 14538 13030 14540 13082
rect 14294 13028 14300 13030
rect 14356 13028 14380 13030
rect 14436 13028 14460 13030
rect 14516 13028 14540 13030
rect 14596 13028 14602 13030
rect 14294 13008 14602 13028
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14568 12374 14596 12786
rect 14740 12436 14792 12442
rect 14844 12434 14872 12854
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 15028 12730 15056 12786
rect 14792 12406 14872 12434
rect 14936 12702 15056 12730
rect 15106 12744 15162 12753
rect 14740 12378 14792 12384
rect 14556 12368 14608 12374
rect 14556 12310 14608 12316
rect 14188 12164 14240 12170
rect 14188 12106 14240 12112
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14108 11898 14136 12038
rect 14200 11898 14228 12106
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14294 11996 14602 12016
rect 14294 11994 14300 11996
rect 14356 11994 14380 11996
rect 14436 11994 14460 11996
rect 14516 11994 14540 11996
rect 14596 11994 14602 11996
rect 14356 11942 14358 11994
rect 14538 11942 14540 11994
rect 14294 11940 14300 11942
rect 14356 11940 14380 11942
rect 14436 11940 14460 11942
rect 14516 11940 14540 11942
rect 14596 11940 14602 11942
rect 14294 11920 14602 11940
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14660 11830 14688 12038
rect 14648 11824 14700 11830
rect 14648 11766 14700 11772
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 13728 11212 13780 11218
rect 13728 11154 13780 11160
rect 13740 10470 13768 11154
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10130 13768 10406
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13740 9654 13768 10066
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13740 8634 13768 9454
rect 14016 9058 14044 11698
rect 14752 11694 14780 12378
rect 14936 12238 14964 12702
rect 15106 12679 15162 12688
rect 15120 12646 15148 12679
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 14924 12232 14976 12238
rect 15212 12186 15240 13262
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 14924 12174 14976 12180
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14464 11620 14516 11626
rect 14464 11562 14516 11568
rect 14096 11552 14148 11558
rect 14096 11494 14148 11500
rect 14108 11257 14136 11494
rect 14476 11354 14504 11562
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14094 11248 14150 11257
rect 14936 11218 14964 12174
rect 15120 12158 15240 12186
rect 15120 11778 15148 12158
rect 15200 12096 15252 12102
rect 15200 12038 15252 12044
rect 15212 11898 15240 12038
rect 15200 11892 15252 11898
rect 15200 11834 15252 11840
rect 15120 11750 15240 11778
rect 14094 11183 14150 11192
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 14096 11144 14148 11150
rect 14096 11086 14148 11092
rect 14108 10470 14136 11086
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14294 10908 14602 10928
rect 14294 10906 14300 10908
rect 14356 10906 14380 10908
rect 14436 10906 14460 10908
rect 14516 10906 14540 10908
rect 14596 10906 14602 10908
rect 14356 10854 14358 10906
rect 14538 10854 14540 10906
rect 14294 10852 14300 10854
rect 14356 10852 14380 10854
rect 14436 10852 14460 10854
rect 14516 10852 14540 10854
rect 14596 10852 14602 10854
rect 14294 10832 14602 10852
rect 14096 10464 14148 10470
rect 14096 10406 14148 10412
rect 14108 10198 14136 10406
rect 14096 10192 14148 10198
rect 14096 10134 14148 10140
rect 14844 9994 14872 10950
rect 14936 10742 14964 11154
rect 14924 10736 14976 10742
rect 14924 10678 14976 10684
rect 14936 10062 14964 10678
rect 15212 10470 15240 11750
rect 15304 11082 15332 13126
rect 15384 12640 15436 12646
rect 15384 12582 15436 12588
rect 15396 12306 15424 12582
rect 15384 12300 15436 12306
rect 15384 12242 15436 12248
rect 15580 11898 15608 13738
rect 15568 11892 15620 11898
rect 15568 11834 15620 11840
rect 15476 11824 15528 11830
rect 15476 11766 15528 11772
rect 15488 11626 15516 11766
rect 15580 11762 15608 11834
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15476 11620 15528 11626
rect 15476 11562 15528 11568
rect 15382 11248 15438 11257
rect 15382 11183 15438 11192
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15290 10976 15346 10985
rect 15290 10911 15346 10920
rect 15304 10674 15332 10911
rect 15396 10810 15424 11183
rect 15384 10804 15436 10810
rect 15384 10746 15436 10752
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15200 10464 15252 10470
rect 15200 10406 15252 10412
rect 15212 10130 15240 10406
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 14096 9580 14148 9586
rect 14096 9522 14148 9528
rect 14108 9178 14136 9522
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 14016 9030 14136 9058
rect 14200 9042 14228 9930
rect 14294 9820 14602 9840
rect 14294 9818 14300 9820
rect 14356 9818 14380 9820
rect 14436 9818 14460 9820
rect 14516 9818 14540 9820
rect 14596 9818 14602 9820
rect 14356 9766 14358 9818
rect 14538 9766 14540 9818
rect 14294 9764 14300 9766
rect 14356 9764 14380 9766
rect 14436 9764 14460 9766
rect 14516 9764 14540 9766
rect 14596 9764 14602 9766
rect 14294 9744 14602 9764
rect 14936 9722 14964 9998
rect 14648 9716 14700 9722
rect 14648 9658 14700 9664
rect 14924 9716 14976 9722
rect 14924 9658 14976 9664
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13832 8537 13860 8774
rect 13818 8528 13874 8537
rect 13874 8486 14044 8514
rect 13818 8463 13874 8472
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13924 7478 13952 7686
rect 13912 7472 13964 7478
rect 13912 7414 13964 7420
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13728 7336 13780 7342
rect 13728 7278 13780 7284
rect 13740 6866 13768 7278
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13832 6798 13860 7346
rect 13544 6792 13596 6798
rect 13820 6792 13872 6798
rect 13544 6734 13596 6740
rect 13818 6760 13820 6769
rect 13872 6760 13874 6769
rect 13360 6724 13412 6730
rect 13360 6666 13412 6672
rect 13636 6724 13688 6730
rect 13818 6695 13874 6704
rect 13636 6666 13688 6672
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13176 6316 13228 6322
rect 13176 6258 13228 6264
rect 13188 5370 13216 6258
rect 13280 5370 13308 6598
rect 13372 6254 13400 6666
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13648 6168 13676 6666
rect 13818 6488 13874 6497
rect 13818 6423 13874 6432
rect 13832 6390 13860 6423
rect 13820 6384 13872 6390
rect 13820 6326 13872 6332
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13728 6180 13780 6186
rect 13648 6140 13728 6168
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 13266 5264 13322 5273
rect 12820 5222 13216 5250
rect 13084 5092 13136 5098
rect 13084 5034 13136 5040
rect 12070 4924 12378 4944
rect 12070 4922 12076 4924
rect 12132 4922 12156 4924
rect 12212 4922 12236 4924
rect 12292 4922 12316 4924
rect 12372 4922 12378 4924
rect 12132 4870 12134 4922
rect 12314 4870 12316 4922
rect 12070 4868 12076 4870
rect 12132 4868 12156 4870
rect 12212 4868 12236 4870
rect 12292 4868 12316 4870
rect 12372 4868 12378 4870
rect 12070 4848 12378 4868
rect 11992 4780 12112 4808
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11980 4480 12032 4486
rect 11980 4422 12032 4428
rect 11992 4214 12020 4422
rect 11980 4208 12032 4214
rect 11980 4150 12032 4156
rect 12084 4026 12112 4780
rect 13096 4690 13124 5034
rect 13084 4684 13136 4690
rect 13084 4626 13136 4632
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 11992 3998 12112 4026
rect 11888 3664 11940 3670
rect 11888 3606 11940 3612
rect 11612 3470 11664 3476
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11520 3460 11572 3466
rect 11520 3402 11572 3408
rect 10980 3318 11192 3346
rect 11336 3392 11388 3398
rect 11532 3346 11560 3402
rect 11336 3334 11388 3340
rect 11440 3318 11560 3346
rect 10980 3058 11008 3318
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10612 2746 10824 2774
rect 10416 2032 10468 2038
rect 10416 1974 10468 1980
rect 10612 1834 10640 2746
rect 11072 2514 11100 2790
rect 11348 2650 11376 2926
rect 11336 2644 11388 2650
rect 11336 2586 11388 2592
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 11152 2508 11204 2514
rect 11152 2450 11204 2456
rect 10966 2408 11022 2417
rect 10966 2343 11022 2352
rect 10980 2310 11008 2343
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 11164 2106 11192 2450
rect 11440 2446 11468 3318
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11532 2514 11560 2994
rect 11520 2508 11572 2514
rect 11520 2450 11572 2456
rect 11428 2440 11480 2446
rect 11428 2382 11480 2388
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 11336 2100 11388 2106
rect 11336 2042 11388 2048
rect 11348 1902 11376 2042
rect 11336 1896 11388 1902
rect 11336 1838 11388 1844
rect 11440 1834 11468 2382
rect 11624 2310 11652 3470
rect 11716 3466 11836 3482
rect 11704 3460 11836 3466
rect 11756 3454 11836 3460
rect 11704 3402 11756 3408
rect 11900 3210 11928 3606
rect 11808 3182 11928 3210
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 10600 1828 10652 1834
rect 10600 1770 10652 1776
rect 11428 1828 11480 1834
rect 11428 1770 11480 1776
rect 11244 1216 11296 1222
rect 11244 1158 11296 1164
rect 11256 800 11284 1158
rect 11808 1086 11836 3182
rect 11888 3052 11940 3058
rect 11888 2994 11940 3000
rect 11900 2650 11928 2994
rect 11992 2650 12020 3998
rect 12360 3992 12388 4422
rect 12360 3964 12480 3992
rect 12070 3836 12378 3856
rect 12070 3834 12076 3836
rect 12132 3834 12156 3836
rect 12212 3834 12236 3836
rect 12292 3834 12316 3836
rect 12372 3834 12378 3836
rect 12132 3782 12134 3834
rect 12314 3782 12316 3834
rect 12070 3780 12076 3782
rect 12132 3780 12156 3782
rect 12212 3780 12236 3782
rect 12292 3780 12316 3782
rect 12372 3780 12378 3782
rect 12070 3760 12378 3780
rect 12452 3618 12480 3964
rect 12360 3590 12480 3618
rect 12072 3528 12124 3534
rect 12072 3470 12124 3476
rect 12084 3194 12112 3470
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12360 3058 12388 3590
rect 12348 3052 12400 3058
rect 12348 2994 12400 3000
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12070 2748 12378 2768
rect 12070 2746 12076 2748
rect 12132 2746 12156 2748
rect 12212 2746 12236 2748
rect 12292 2746 12316 2748
rect 12372 2746 12378 2748
rect 12132 2694 12134 2746
rect 12314 2694 12316 2746
rect 12070 2692 12076 2694
rect 12132 2692 12156 2694
rect 12212 2692 12236 2694
rect 12292 2692 12316 2694
rect 12372 2692 12378 2694
rect 12070 2672 12378 2692
rect 11888 2644 11940 2650
rect 11888 2586 11940 2592
rect 11980 2644 12032 2650
rect 11980 2586 12032 2592
rect 12348 2440 12400 2446
rect 12348 2382 12400 2388
rect 12360 1970 12388 2382
rect 12452 2310 12480 2790
rect 13188 2774 13216 5222
rect 13266 5199 13322 5208
rect 13360 5228 13412 5234
rect 13280 4146 13308 5199
rect 13360 5170 13412 5176
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 13372 3602 13400 5170
rect 13464 4282 13492 5170
rect 13556 5098 13584 5646
rect 13648 5574 13676 6140
rect 13728 6122 13780 6128
rect 13726 5808 13782 5817
rect 13726 5743 13782 5752
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13648 5166 13676 5510
rect 13740 5302 13768 5743
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13544 5092 13596 5098
rect 13544 5034 13596 5040
rect 13832 4706 13860 6190
rect 13912 5568 13964 5574
rect 13912 5510 13964 5516
rect 13556 4678 13860 4706
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13360 3596 13412 3602
rect 13360 3538 13412 3544
rect 13464 3534 13492 4082
rect 13556 4078 13584 4678
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13556 3738 13584 4014
rect 13832 3942 13860 4558
rect 13924 4486 13952 5510
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 13910 4176 13966 4185
rect 13910 4111 13966 4120
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13924 3738 13952 4111
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13912 3732 13964 3738
rect 13912 3674 13964 3680
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13912 3528 13964 3534
rect 13912 3470 13964 3476
rect 13464 3194 13492 3470
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13740 2854 13768 3470
rect 13924 3398 13952 3470
rect 14016 3398 14044 8486
rect 14108 7410 14136 9030
rect 14188 9036 14240 9042
rect 14188 8978 14240 8984
rect 14660 8838 14688 9658
rect 15396 9466 15424 10746
rect 15476 10464 15528 10470
rect 15476 10406 15528 10412
rect 15488 9926 15516 10406
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15212 9438 15424 9466
rect 14738 8936 14794 8945
rect 14738 8871 14740 8880
rect 14792 8871 14794 8880
rect 14740 8842 14792 8848
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14294 8732 14602 8752
rect 14294 8730 14300 8732
rect 14356 8730 14380 8732
rect 14436 8730 14460 8732
rect 14516 8730 14540 8732
rect 14596 8730 14602 8732
rect 14356 8678 14358 8730
rect 14538 8678 14540 8730
rect 14294 8676 14300 8678
rect 14356 8676 14380 8678
rect 14436 8676 14460 8678
rect 14516 8676 14540 8678
rect 14596 8676 14602 8678
rect 14294 8656 14602 8676
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 7954 14596 8230
rect 14660 7954 14688 8774
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14648 7948 14700 7954
rect 14648 7890 14700 7896
rect 14752 7834 14780 8842
rect 15108 8832 15160 8838
rect 15108 8774 15160 8780
rect 15014 8664 15070 8673
rect 15120 8634 15148 8774
rect 15014 8599 15070 8608
rect 15108 8628 15160 8634
rect 15028 8498 15056 8599
rect 15108 8570 15160 8576
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 14844 8294 14872 8434
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14832 8288 14884 8294
rect 14832 8230 14884 8236
rect 14660 7806 14780 7834
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14200 7546 14228 7686
rect 14294 7644 14602 7664
rect 14294 7642 14300 7644
rect 14356 7642 14380 7644
rect 14436 7642 14460 7644
rect 14516 7642 14540 7644
rect 14596 7642 14602 7644
rect 14356 7590 14358 7642
rect 14538 7590 14540 7642
rect 14294 7588 14300 7590
rect 14356 7588 14380 7590
rect 14436 7588 14460 7590
rect 14516 7588 14540 7590
rect 14596 7588 14602 7590
rect 14294 7568 14602 7588
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14096 7404 14148 7410
rect 14096 7346 14148 7352
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14108 5846 14136 6734
rect 14294 6556 14602 6576
rect 14294 6554 14300 6556
rect 14356 6554 14380 6556
rect 14436 6554 14460 6556
rect 14516 6554 14540 6556
rect 14596 6554 14602 6556
rect 14356 6502 14358 6554
rect 14538 6502 14540 6554
rect 14294 6500 14300 6502
rect 14356 6500 14380 6502
rect 14436 6500 14460 6502
rect 14516 6500 14540 6502
rect 14596 6500 14602 6502
rect 14294 6480 14602 6500
rect 14660 6322 14688 7806
rect 14832 7744 14884 7750
rect 14832 7686 14884 7692
rect 14740 7336 14792 7342
rect 14740 7278 14792 7284
rect 14752 6730 14780 7278
rect 14740 6724 14792 6730
rect 14740 6666 14792 6672
rect 14648 6316 14700 6322
rect 14648 6258 14700 6264
rect 14660 6202 14688 6258
rect 14200 6174 14688 6202
rect 14096 5840 14148 5846
rect 14096 5782 14148 5788
rect 14108 5166 14136 5782
rect 14096 5160 14148 5166
rect 14096 5102 14148 5108
rect 14108 4214 14136 5102
rect 14096 4208 14148 4214
rect 14096 4150 14148 4156
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 14004 3392 14056 3398
rect 14004 3334 14056 3340
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13188 2746 13676 2774
rect 12992 2576 13044 2582
rect 12990 2544 12992 2553
rect 13044 2544 13046 2553
rect 12990 2479 13046 2488
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 13648 2038 13676 2746
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13740 2106 13768 2246
rect 13728 2100 13780 2106
rect 13728 2042 13780 2048
rect 13636 2032 13688 2038
rect 13636 1974 13688 1980
rect 12348 1964 12400 1970
rect 12348 1906 12400 1912
rect 12164 1896 12216 1902
rect 12164 1838 12216 1844
rect 11796 1080 11848 1086
rect 11796 1022 11848 1028
rect 12176 800 12204 1838
rect 13084 1556 13136 1562
rect 13084 1498 13136 1504
rect 13096 800 13124 1498
rect 13924 800 13952 3130
rect 14004 3120 14056 3126
rect 14004 3062 14056 3068
rect 14016 2650 14044 3062
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14108 2514 14136 3470
rect 14200 3126 14228 6174
rect 14660 5930 14688 6174
rect 14660 5902 14780 5930
rect 14646 5808 14702 5817
rect 14752 5778 14780 5902
rect 14646 5743 14648 5752
rect 14700 5743 14702 5752
rect 14740 5772 14792 5778
rect 14648 5714 14700 5720
rect 14740 5714 14792 5720
rect 14372 5704 14424 5710
rect 14556 5704 14608 5710
rect 14424 5652 14556 5658
rect 14372 5646 14608 5652
rect 14384 5630 14596 5646
rect 14294 5468 14602 5488
rect 14294 5466 14300 5468
rect 14356 5466 14380 5468
rect 14436 5466 14460 5468
rect 14516 5466 14540 5468
rect 14596 5466 14602 5468
rect 14356 5414 14358 5466
rect 14538 5414 14540 5466
rect 14294 5412 14300 5414
rect 14356 5412 14380 5414
rect 14436 5412 14460 5414
rect 14516 5412 14540 5414
rect 14596 5412 14602 5414
rect 14294 5392 14602 5412
rect 14660 5302 14688 5714
rect 14740 5636 14792 5642
rect 14740 5578 14792 5584
rect 14648 5296 14700 5302
rect 14648 5238 14700 5244
rect 14372 5228 14424 5234
rect 14372 5170 14424 5176
rect 14384 5137 14412 5170
rect 14370 5128 14426 5137
rect 14370 5063 14426 5072
rect 14660 4690 14688 5238
rect 14648 4684 14700 4690
rect 14648 4626 14700 4632
rect 14648 4548 14700 4554
rect 14648 4490 14700 4496
rect 14294 4380 14602 4400
rect 14294 4378 14300 4380
rect 14356 4378 14380 4380
rect 14436 4378 14460 4380
rect 14516 4378 14540 4380
rect 14596 4378 14602 4380
rect 14356 4326 14358 4378
rect 14538 4326 14540 4378
rect 14294 4324 14300 4326
rect 14356 4324 14380 4326
rect 14436 4324 14460 4326
rect 14516 4324 14540 4326
rect 14596 4324 14602 4326
rect 14294 4304 14602 4324
rect 14280 3936 14332 3942
rect 14280 3878 14332 3884
rect 14292 3602 14320 3878
rect 14660 3738 14688 4490
rect 14648 3732 14700 3738
rect 14648 3674 14700 3680
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14294 3292 14602 3312
rect 14294 3290 14300 3292
rect 14356 3290 14380 3292
rect 14436 3290 14460 3292
rect 14516 3290 14540 3292
rect 14596 3290 14602 3292
rect 14356 3238 14358 3290
rect 14538 3238 14540 3290
rect 14294 3236 14300 3238
rect 14356 3236 14380 3238
rect 14436 3236 14460 3238
rect 14516 3236 14540 3238
rect 14596 3236 14602 3238
rect 14294 3216 14602 3236
rect 14188 3120 14240 3126
rect 14188 3062 14240 3068
rect 14752 2922 14780 5578
rect 14844 4570 14872 7686
rect 14936 7342 14964 8366
rect 14924 7336 14976 7342
rect 14924 7278 14976 7284
rect 14924 5568 14976 5574
rect 14924 5510 14976 5516
rect 14936 4758 14964 5510
rect 15028 5370 15056 8434
rect 15120 8362 15148 8434
rect 15108 8356 15160 8362
rect 15108 8298 15160 8304
rect 15212 6322 15240 9438
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15396 8362 15424 9318
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15384 8356 15436 8362
rect 15384 8298 15436 8304
rect 15292 8288 15344 8294
rect 15292 8230 15344 8236
rect 15304 7750 15332 8230
rect 15396 8022 15424 8298
rect 15384 8016 15436 8022
rect 15384 7958 15436 7964
rect 15292 7744 15344 7750
rect 15292 7686 15344 7692
rect 15488 6458 15516 8774
rect 15580 8634 15608 11698
rect 15672 10470 15700 14175
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15856 10810 15884 12718
rect 15948 12374 15976 15535
rect 16518 14716 16826 14736
rect 16518 14714 16524 14716
rect 16580 14714 16604 14716
rect 16660 14714 16684 14716
rect 16740 14714 16764 14716
rect 16820 14714 16826 14716
rect 16580 14662 16582 14714
rect 16762 14662 16764 14714
rect 16518 14660 16524 14662
rect 16580 14660 16604 14662
rect 16660 14660 16684 14662
rect 16740 14660 16764 14662
rect 16820 14660 16826 14662
rect 16518 14640 16826 14660
rect 16868 13870 16896 16510
rect 18064 15366 18092 16759
rect 18786 16400 18842 17200
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 18064 14498 18092 15302
rect 18064 14470 18184 14498
rect 18052 14340 18104 14346
rect 18052 14282 18104 14288
rect 18064 14074 18092 14282
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 16948 14000 17000 14006
rect 16948 13942 17000 13948
rect 17038 13968 17094 13977
rect 16856 13864 16908 13870
rect 16856 13806 16908 13812
rect 16518 13628 16826 13648
rect 16518 13626 16524 13628
rect 16580 13626 16604 13628
rect 16660 13626 16684 13628
rect 16740 13626 16764 13628
rect 16820 13626 16826 13628
rect 16580 13574 16582 13626
rect 16762 13574 16764 13626
rect 16518 13572 16524 13574
rect 16580 13572 16604 13574
rect 16660 13572 16684 13574
rect 16740 13572 16764 13574
rect 16820 13572 16826 13574
rect 16518 13552 16826 13572
rect 16868 13530 16896 13806
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16960 13462 16988 13942
rect 17038 13903 17094 13912
rect 17868 13932 17920 13938
rect 17052 13870 17080 13903
rect 17868 13874 17920 13880
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 16948 13456 17000 13462
rect 16948 13398 17000 13404
rect 17144 13258 17172 13738
rect 17132 13252 17184 13258
rect 17132 13194 17184 13200
rect 17880 13190 17908 13874
rect 18064 13326 18092 13874
rect 18052 13320 18104 13326
rect 18050 13288 18052 13297
rect 18104 13288 18106 13297
rect 18050 13223 18106 13232
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 17868 13184 17920 13190
rect 17868 13126 17920 13132
rect 16118 13016 16174 13025
rect 16118 12951 16174 12960
rect 15936 12368 15988 12374
rect 15934 12336 15936 12345
rect 15988 12336 15990 12345
rect 15934 12271 15990 12280
rect 16132 11830 16160 12951
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16518 12540 16826 12560
rect 16518 12538 16524 12540
rect 16580 12538 16604 12540
rect 16660 12538 16684 12540
rect 16740 12538 16764 12540
rect 16820 12538 16826 12540
rect 16580 12486 16582 12538
rect 16762 12486 16764 12538
rect 16518 12484 16524 12486
rect 16580 12484 16604 12486
rect 16660 12484 16684 12486
rect 16740 12484 16764 12486
rect 16820 12484 16826 12486
rect 16518 12464 16826 12484
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16120 11824 16172 11830
rect 16040 11784 16120 11812
rect 15844 10804 15896 10810
rect 15844 10746 15896 10752
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15844 10192 15896 10198
rect 15844 10134 15896 10140
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15660 9104 15712 9110
rect 15660 9046 15712 9052
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15476 6452 15528 6458
rect 15476 6394 15528 6400
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 15212 6168 15240 6258
rect 15384 6180 15436 6186
rect 15212 6140 15384 6168
rect 15384 6122 15436 6128
rect 15382 5808 15438 5817
rect 15200 5772 15252 5778
rect 15382 5743 15438 5752
rect 15200 5714 15252 5720
rect 15106 5672 15162 5681
rect 15106 5607 15162 5616
rect 15016 5364 15068 5370
rect 15016 5306 15068 5312
rect 15028 4758 15056 5306
rect 14924 4752 14976 4758
rect 14924 4694 14976 4700
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 14844 4542 14964 4570
rect 14832 4480 14884 4486
rect 14832 4422 14884 4428
rect 14844 4282 14872 4422
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14832 3052 14884 3058
rect 14936 3040 14964 4542
rect 14884 3012 14964 3040
rect 14832 2994 14884 3000
rect 15028 2938 15056 4694
rect 15120 4486 15148 5607
rect 15212 5137 15240 5714
rect 15396 5574 15424 5743
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15304 5370 15332 5510
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15198 5128 15254 5137
rect 15488 5114 15516 6394
rect 15198 5063 15254 5072
rect 15396 5086 15516 5114
rect 15212 4690 15240 5063
rect 15396 5030 15424 5086
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15200 4684 15252 4690
rect 15200 4626 15252 4632
rect 15108 4480 15160 4486
rect 15108 4422 15160 4428
rect 15212 4010 15240 4626
rect 15396 4486 15424 4762
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15476 4480 15528 4486
rect 15476 4422 15528 4428
rect 15290 4176 15346 4185
rect 15290 4111 15346 4120
rect 15384 4140 15436 4146
rect 15200 4004 15252 4010
rect 15200 3946 15252 3952
rect 15304 3058 15332 4111
rect 15384 4082 15436 4088
rect 15396 3738 15424 4082
rect 15384 3732 15436 3738
rect 15384 3674 15436 3680
rect 15488 3466 15516 4422
rect 15580 4162 15608 7686
rect 15672 4758 15700 9046
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 15672 4282 15700 4694
rect 15660 4276 15712 4282
rect 15660 4218 15712 4224
rect 15580 4134 15700 4162
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15476 3460 15528 3466
rect 15476 3402 15528 3408
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 15200 2984 15252 2990
rect 14740 2916 14792 2922
rect 14740 2858 14792 2864
rect 14832 2916 14884 2922
rect 15028 2910 15148 2938
rect 15200 2926 15252 2932
rect 14832 2858 14884 2864
rect 14752 2650 14780 2858
rect 14740 2644 14792 2650
rect 14740 2586 14792 2592
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14096 2372 14148 2378
rect 14096 2314 14148 2320
rect 14108 1902 14136 2314
rect 14294 2204 14602 2224
rect 14294 2202 14300 2204
rect 14356 2202 14380 2204
rect 14436 2202 14460 2204
rect 14516 2202 14540 2204
rect 14596 2202 14602 2204
rect 14356 2150 14358 2202
rect 14538 2150 14540 2202
rect 14294 2148 14300 2150
rect 14356 2148 14380 2150
rect 14436 2148 14460 2150
rect 14516 2148 14540 2150
rect 14596 2148 14602 2150
rect 14294 2128 14602 2148
rect 14660 1970 14688 2382
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14752 2106 14780 2246
rect 14740 2100 14792 2106
rect 14740 2042 14792 2048
rect 14648 1964 14700 1970
rect 14648 1906 14700 1912
rect 14096 1896 14148 1902
rect 14096 1838 14148 1844
rect 14844 800 14872 2858
rect 14924 2576 14976 2582
rect 14924 2518 14976 2524
rect 15016 2576 15068 2582
rect 15016 2518 15068 2524
rect 14936 2446 14964 2518
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15028 1222 15056 2518
rect 15120 2446 15148 2910
rect 15108 2440 15160 2446
rect 15108 2382 15160 2388
rect 15212 1562 15240 2926
rect 15474 2680 15530 2689
rect 15474 2615 15530 2624
rect 15488 2446 15516 2615
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 15580 2310 15608 4014
rect 15672 3738 15700 4134
rect 15660 3732 15712 3738
rect 15660 3674 15712 3680
rect 15672 3126 15700 3674
rect 15660 3120 15712 3126
rect 15660 3062 15712 3068
rect 15764 3058 15792 9862
rect 15856 9586 15884 10134
rect 15934 10024 15990 10033
rect 15934 9959 15990 9968
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 15856 9042 15884 9522
rect 15844 9036 15896 9042
rect 15844 8978 15896 8984
rect 15948 8022 15976 9959
rect 15936 8016 15988 8022
rect 15936 7958 15988 7964
rect 15948 7426 15976 7958
rect 15856 7398 15976 7426
rect 15856 6474 15884 7398
rect 15934 7304 15990 7313
rect 15934 7239 15990 7248
rect 15948 6798 15976 7239
rect 15936 6792 15988 6798
rect 15936 6734 15988 6740
rect 16040 6644 16068 11784
rect 16120 11766 16172 11772
rect 16212 11688 16264 11694
rect 16500 11665 16528 12038
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16212 11630 16264 11636
rect 16486 11656 16542 11665
rect 16120 11620 16172 11626
rect 16120 11562 16172 11568
rect 16132 10169 16160 11562
rect 16224 11529 16252 11630
rect 16486 11591 16542 11600
rect 16396 11552 16448 11558
rect 16210 11520 16266 11529
rect 16396 11494 16448 11500
rect 16210 11455 16266 11464
rect 16408 11286 16436 11494
rect 16518 11452 16826 11472
rect 16518 11450 16524 11452
rect 16580 11450 16604 11452
rect 16660 11450 16684 11452
rect 16740 11450 16764 11452
rect 16820 11450 16826 11452
rect 16580 11398 16582 11450
rect 16762 11398 16764 11450
rect 16518 11396 16524 11398
rect 16580 11396 16604 11398
rect 16660 11396 16684 11398
rect 16740 11396 16764 11398
rect 16820 11396 16826 11398
rect 16518 11376 16826 11396
rect 16396 11280 16448 11286
rect 16396 11222 16448 11228
rect 16304 10736 16356 10742
rect 16304 10678 16356 10684
rect 16316 10470 16344 10678
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16118 10160 16174 10169
rect 16118 10095 16174 10104
rect 16212 9376 16264 9382
rect 16212 9318 16264 9324
rect 16224 8906 16252 9318
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 16224 8809 16252 8842
rect 16316 8838 16344 10406
rect 16408 9024 16436 11222
rect 16868 11014 16896 11698
rect 16672 11008 16724 11014
rect 16856 11008 16908 11014
rect 16672 10950 16724 10956
rect 16854 10976 16856 10985
rect 16908 10976 16910 10985
rect 16684 10606 16712 10950
rect 16854 10911 16910 10920
rect 16868 10885 16896 10911
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 16518 10364 16826 10384
rect 16518 10362 16524 10364
rect 16580 10362 16604 10364
rect 16660 10362 16684 10364
rect 16740 10362 16764 10364
rect 16820 10362 16826 10364
rect 16580 10310 16582 10362
rect 16762 10310 16764 10362
rect 16518 10308 16524 10310
rect 16580 10308 16604 10310
rect 16660 10308 16684 10310
rect 16740 10308 16764 10310
rect 16820 10308 16826 10310
rect 16518 10288 16826 10308
rect 16868 10198 16896 10610
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16856 10192 16908 10198
rect 16856 10134 16908 10140
rect 16868 9674 16896 10134
rect 16960 10130 16988 10542
rect 16948 10124 17000 10130
rect 16948 10066 17000 10072
rect 16776 9646 16896 9674
rect 16776 9450 16804 9646
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16764 9444 16816 9450
rect 16764 9386 16816 9392
rect 16518 9276 16826 9296
rect 16518 9274 16524 9276
rect 16580 9274 16604 9276
rect 16660 9274 16684 9276
rect 16740 9274 16764 9276
rect 16820 9274 16826 9276
rect 16580 9222 16582 9274
rect 16762 9222 16764 9274
rect 16518 9220 16524 9222
rect 16580 9220 16604 9222
rect 16660 9220 16684 9222
rect 16740 9220 16764 9222
rect 16820 9220 16826 9222
rect 16518 9200 16826 9220
rect 16408 8996 16528 9024
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16304 8832 16356 8838
rect 16210 8800 16266 8809
rect 16304 8774 16356 8780
rect 16210 8735 16266 8744
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16132 7410 16160 8366
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16132 6866 16160 7346
rect 16224 6866 16252 8570
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 16316 7954 16344 8366
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 16120 6860 16172 6866
rect 16120 6802 16172 6808
rect 16212 6860 16264 6866
rect 16212 6802 16264 6808
rect 16120 6656 16172 6662
rect 16040 6616 16120 6644
rect 16120 6598 16172 6604
rect 15856 6446 16068 6474
rect 15844 6384 15896 6390
rect 15844 6326 15896 6332
rect 15934 6352 15990 6361
rect 15856 3738 15884 6326
rect 15934 6287 15936 6296
rect 15988 6287 15990 6296
rect 15936 6258 15988 6264
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15948 5302 15976 6054
rect 16040 5370 16068 6446
rect 16028 5364 16080 5370
rect 16028 5306 16080 5312
rect 15936 5296 15988 5302
rect 15936 5238 15988 5244
rect 15948 4622 15976 5238
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 16132 4146 16160 6598
rect 16224 6458 16252 6802
rect 16316 6730 16344 7754
rect 16408 7546 16436 8842
rect 16500 8673 16528 8996
rect 16868 8974 16896 9454
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16486 8664 16542 8673
rect 16486 8599 16488 8608
rect 16540 8599 16542 8608
rect 16488 8570 16540 8576
rect 16500 8539 16528 8570
rect 16684 8498 16712 8910
rect 16672 8492 16724 8498
rect 16672 8434 16724 8440
rect 16518 8188 16826 8208
rect 16518 8186 16524 8188
rect 16580 8186 16604 8188
rect 16660 8186 16684 8188
rect 16740 8186 16764 8188
rect 16820 8186 16826 8188
rect 16580 8134 16582 8186
rect 16762 8134 16764 8186
rect 16518 8132 16524 8134
rect 16580 8132 16604 8134
rect 16660 8132 16684 8134
rect 16740 8132 16764 8134
rect 16820 8132 16826 8134
rect 16518 8112 16826 8132
rect 16868 8090 16896 8910
rect 17052 8401 17080 12582
rect 17132 11824 17184 11830
rect 17132 11766 17184 11772
rect 17144 11626 17172 11766
rect 17132 11620 17184 11626
rect 17132 11562 17184 11568
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 17144 9178 17172 9862
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17038 8392 17094 8401
rect 17038 8327 17094 8336
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 16764 7948 16816 7954
rect 16764 7890 16816 7896
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 16776 7188 16804 7890
rect 16868 7478 16896 8026
rect 16946 7848 17002 7857
rect 16946 7783 17002 7792
rect 16856 7472 16908 7478
rect 16856 7414 16908 7420
rect 16776 7160 16896 7188
rect 16518 7100 16826 7120
rect 16518 7098 16524 7100
rect 16580 7098 16604 7100
rect 16660 7098 16684 7100
rect 16740 7098 16764 7100
rect 16820 7098 16826 7100
rect 16580 7046 16582 7098
rect 16762 7046 16764 7098
rect 16518 7044 16524 7046
rect 16580 7044 16604 7046
rect 16660 7044 16684 7046
rect 16740 7044 16764 7046
rect 16820 7044 16826 7046
rect 16518 7024 16826 7044
rect 16868 7002 16896 7160
rect 16856 6996 16908 7002
rect 16856 6938 16908 6944
rect 16304 6724 16356 6730
rect 16304 6666 16356 6672
rect 16212 6452 16264 6458
rect 16212 6394 16264 6400
rect 16316 5642 16344 6666
rect 16868 6390 16896 6938
rect 16856 6384 16908 6390
rect 16856 6326 16908 6332
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16856 6248 16908 6254
rect 16856 6190 16908 6196
rect 16304 5636 16356 5642
rect 16304 5578 16356 5584
rect 16316 5370 16344 5578
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16212 5296 16264 5302
rect 16212 5238 16264 5244
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 15936 4072 15988 4078
rect 15934 4040 15936 4049
rect 15988 4040 15990 4049
rect 15934 3975 15990 3984
rect 16028 4004 16080 4010
rect 16028 3946 16080 3952
rect 15844 3732 15896 3738
rect 15844 3674 15896 3680
rect 16040 3641 16068 3946
rect 16224 3670 16252 5238
rect 16302 4856 16358 4865
rect 16302 4791 16304 4800
rect 16356 4791 16358 4800
rect 16304 4762 16356 4768
rect 16408 4729 16436 6190
rect 16518 6012 16826 6032
rect 16518 6010 16524 6012
rect 16580 6010 16604 6012
rect 16660 6010 16684 6012
rect 16740 6010 16764 6012
rect 16820 6010 16826 6012
rect 16580 5958 16582 6010
rect 16762 5958 16764 6010
rect 16518 5956 16524 5958
rect 16580 5956 16604 5958
rect 16660 5956 16684 5958
rect 16740 5956 16764 5958
rect 16820 5956 16826 5958
rect 16518 5936 16826 5956
rect 16868 5846 16896 6190
rect 16856 5840 16908 5846
rect 16856 5782 16908 5788
rect 16672 5568 16724 5574
rect 16486 5536 16542 5545
rect 16672 5510 16724 5516
rect 16486 5471 16542 5480
rect 16500 5370 16528 5471
rect 16684 5370 16712 5510
rect 16854 5400 16910 5409
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16672 5364 16724 5370
rect 16854 5335 16856 5344
rect 16672 5306 16724 5312
rect 16908 5335 16910 5344
rect 16856 5306 16908 5312
rect 16518 4924 16826 4944
rect 16518 4922 16524 4924
rect 16580 4922 16604 4924
rect 16660 4922 16684 4924
rect 16740 4922 16764 4924
rect 16820 4922 16826 4924
rect 16580 4870 16582 4922
rect 16762 4870 16764 4922
rect 16518 4868 16524 4870
rect 16580 4868 16604 4870
rect 16660 4868 16684 4870
rect 16740 4868 16764 4870
rect 16820 4868 16826 4870
rect 16518 4848 16826 4868
rect 16960 4826 16988 7783
rect 17052 6322 17080 8327
rect 17236 7954 17264 13126
rect 18156 12986 18184 14470
rect 18512 14068 18564 14074
rect 18512 14010 18564 14016
rect 18418 13424 18474 13433
rect 18418 13359 18474 13368
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 17500 12844 17552 12850
rect 17500 12786 17552 12792
rect 18328 12844 18380 12850
rect 18328 12786 18380 12792
rect 17408 12232 17460 12238
rect 17408 12174 17460 12180
rect 17316 12164 17368 12170
rect 17316 12106 17368 12112
rect 17328 11694 17356 12106
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17328 11354 17356 11630
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17328 10674 17356 11290
rect 17420 11150 17448 12174
rect 17512 11898 17540 12786
rect 18144 12776 18196 12782
rect 18144 12718 18196 12724
rect 17776 12708 17828 12714
rect 17776 12650 17828 12656
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17604 10674 17632 12582
rect 17788 12238 17816 12650
rect 18156 12306 18184 12718
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 17776 12232 17828 12238
rect 17776 12174 17828 12180
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17788 11354 17816 11698
rect 17776 11348 17828 11354
rect 17776 11290 17828 11296
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17592 10668 17644 10674
rect 17592 10610 17644 10616
rect 17314 10568 17370 10577
rect 17314 10503 17370 10512
rect 17328 7993 17356 10503
rect 17500 10464 17552 10470
rect 17696 10441 17724 10950
rect 17500 10406 17552 10412
rect 17682 10432 17738 10441
rect 17512 10062 17540 10406
rect 17682 10367 17738 10376
rect 17500 10056 17552 10062
rect 17500 9998 17552 10004
rect 17788 9625 17816 11290
rect 17880 10810 17908 12038
rect 18156 11150 18184 12242
rect 18144 11144 18196 11150
rect 18144 11086 18196 11092
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17958 10704 18014 10713
rect 17958 10639 18014 10648
rect 17972 10062 18000 10639
rect 18156 10130 18184 11086
rect 18340 10810 18368 12786
rect 18432 12170 18460 13359
rect 18420 12164 18472 12170
rect 18420 12106 18472 12112
rect 18328 10804 18380 10810
rect 18328 10746 18380 10752
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 17960 10056 18012 10062
rect 17960 9998 18012 10004
rect 17972 9654 18000 9998
rect 18156 9722 18184 10066
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 17960 9648 18012 9654
rect 17774 9616 17830 9625
rect 17500 9580 17552 9586
rect 17960 9590 18012 9596
rect 17774 9551 17830 9560
rect 17500 9522 17552 9528
rect 17314 7984 17370 7993
rect 17224 7948 17276 7954
rect 17314 7919 17370 7928
rect 17408 7948 17460 7954
rect 17224 7890 17276 7896
rect 17408 7890 17460 7896
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17144 7410 17172 7822
rect 17314 7712 17370 7721
rect 17314 7647 17370 7656
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 17132 6792 17184 6798
rect 17132 6734 17184 6740
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17144 6118 17172 6734
rect 17328 6304 17356 7647
rect 17236 6276 17356 6304
rect 17132 6112 17184 6118
rect 17132 6054 17184 6060
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 16948 4820 17000 4826
rect 16948 4762 17000 4768
rect 16394 4720 16450 4729
rect 16394 4655 16450 4664
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16316 3738 16344 4082
rect 16304 3732 16356 3738
rect 16408 3720 16436 4558
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16868 4162 16896 4422
rect 16960 4282 16988 4762
rect 17052 4486 17080 5510
rect 17144 4554 17172 6054
rect 17132 4548 17184 4554
rect 17132 4490 17184 4496
rect 17040 4480 17092 4486
rect 17040 4422 17092 4428
rect 17052 4321 17080 4422
rect 17038 4312 17094 4321
rect 16948 4276 17000 4282
rect 17038 4247 17094 4256
rect 16948 4218 17000 4224
rect 17040 4208 17092 4214
rect 16868 4134 16988 4162
rect 17040 4150 17092 4156
rect 16960 4078 16988 4134
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 16948 4072 17000 4078
rect 16948 4014 17000 4020
rect 16518 3836 16826 3856
rect 16518 3834 16524 3836
rect 16580 3834 16604 3836
rect 16660 3834 16684 3836
rect 16740 3834 16764 3836
rect 16820 3834 16826 3836
rect 16580 3782 16582 3834
rect 16762 3782 16764 3834
rect 16518 3780 16524 3782
rect 16580 3780 16604 3782
rect 16660 3780 16684 3782
rect 16740 3780 16764 3782
rect 16820 3780 16826 3782
rect 16518 3760 16826 3780
rect 16408 3692 16620 3720
rect 16304 3674 16356 3680
rect 16212 3664 16264 3670
rect 16026 3632 16082 3641
rect 16212 3606 16264 3612
rect 16026 3567 16028 3576
rect 16080 3567 16082 3576
rect 16028 3538 16080 3544
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 16040 2990 16068 3538
rect 16224 3398 16252 3606
rect 16212 3392 16264 3398
rect 16212 3334 16264 3340
rect 16316 3126 16344 3674
rect 16592 3466 16620 3692
rect 16580 3460 16632 3466
rect 16580 3402 16632 3408
rect 16120 3120 16172 3126
rect 16120 3062 16172 3068
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 15568 2304 15620 2310
rect 15568 2246 15620 2252
rect 15200 1556 15252 1562
rect 15200 1498 15252 1504
rect 15016 1216 15068 1222
rect 15016 1158 15068 1164
rect 15764 800 15792 2790
rect 16132 2310 16160 3062
rect 16592 2922 16620 3402
rect 16868 3097 16896 4014
rect 16960 3602 16988 4014
rect 17052 3738 17080 4150
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 16948 3596 17000 3602
rect 16948 3538 17000 3544
rect 16946 3496 17002 3505
rect 16946 3431 16948 3440
rect 17000 3431 17002 3440
rect 16948 3402 17000 3408
rect 17038 3224 17094 3233
rect 17038 3159 17094 3168
rect 16854 3088 16910 3097
rect 17052 3058 17080 3159
rect 16854 3023 16910 3032
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16762 2952 16818 2961
rect 16304 2916 16356 2922
rect 16304 2858 16356 2864
rect 16580 2916 16632 2922
rect 16762 2887 16764 2896
rect 16580 2858 16632 2864
rect 16816 2887 16818 2896
rect 16764 2858 16816 2864
rect 16316 2650 16344 2858
rect 16946 2816 17002 2825
rect 16518 2748 16826 2768
rect 16946 2751 17002 2760
rect 16518 2746 16524 2748
rect 16580 2746 16604 2748
rect 16660 2746 16684 2748
rect 16740 2746 16764 2748
rect 16820 2746 16826 2748
rect 16580 2694 16582 2746
rect 16762 2694 16764 2746
rect 16518 2692 16524 2694
rect 16580 2692 16604 2694
rect 16660 2692 16684 2694
rect 16740 2692 16764 2694
rect 16820 2692 16826 2694
rect 16518 2672 16826 2692
rect 16304 2644 16356 2650
rect 16304 2586 16356 2592
rect 16672 2576 16724 2582
rect 16672 2518 16724 2524
rect 16684 2310 16712 2518
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 16132 2106 16160 2246
rect 16120 2100 16172 2106
rect 16120 2042 16172 2048
rect 16684 1834 16712 2246
rect 16672 1828 16724 1834
rect 16672 1770 16724 1776
rect 16684 870 16804 898
rect 16684 800 16712 870
rect 7024 734 7512 762
rect 7562 0 7618 800
rect 8482 0 8538 800
rect 9402 0 9458 800
rect 10322 0 10378 800
rect 11242 0 11298 800
rect 12162 0 12218 800
rect 13082 0 13138 800
rect 13910 0 13966 800
rect 14830 0 14886 800
rect 15750 0 15806 800
rect 16670 0 16726 800
rect 16776 762 16804 870
rect 16960 762 16988 2751
rect 17236 2650 17264 6276
rect 17314 6216 17370 6225
rect 17314 6151 17370 6160
rect 17328 5914 17356 6151
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17328 5710 17356 5850
rect 17316 5704 17368 5710
rect 17316 5646 17368 5652
rect 17316 5296 17368 5302
rect 17316 5238 17368 5244
rect 17328 4282 17356 5238
rect 17316 4276 17368 4282
rect 17316 4218 17368 4224
rect 17316 3732 17368 3738
rect 17316 3674 17368 3680
rect 17328 3058 17356 3674
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17224 2644 17276 2650
rect 17224 2586 17276 2592
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 17052 1970 17080 2246
rect 17236 2038 17264 2246
rect 17224 2032 17276 2038
rect 17224 1974 17276 1980
rect 17040 1964 17092 1970
rect 17040 1906 17092 1912
rect 17328 1873 17356 2790
rect 17314 1864 17370 1873
rect 17420 1850 17448 7890
rect 17512 7546 17540 9522
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17604 7954 17632 8774
rect 17788 8498 17816 9551
rect 17866 9208 17922 9217
rect 17866 9143 17922 9152
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17684 8016 17736 8022
rect 17684 7958 17736 7964
rect 17592 7948 17644 7954
rect 17592 7890 17644 7896
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17604 7410 17632 7890
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17500 7200 17552 7206
rect 17500 7142 17552 7148
rect 17512 7002 17540 7142
rect 17500 6996 17552 7002
rect 17500 6938 17552 6944
rect 17696 6882 17724 7958
rect 17774 7848 17830 7857
rect 17880 7818 17908 9143
rect 17972 8498 18000 9590
rect 18156 9042 18184 9658
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 17960 8492 18012 8498
rect 17960 8434 18012 8440
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17972 7886 18000 8298
rect 18064 8090 18092 8774
rect 18328 8356 18380 8362
rect 18328 8298 18380 8304
rect 18142 8256 18198 8265
rect 18142 8191 18198 8200
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17774 7783 17830 7792
rect 17868 7812 17920 7818
rect 17512 6854 17724 6882
rect 17512 3942 17540 6854
rect 17592 6792 17644 6798
rect 17592 6734 17644 6740
rect 17604 6322 17632 6734
rect 17788 6730 17816 7783
rect 17868 7754 17920 7760
rect 17880 7206 17908 7754
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17866 7032 17922 7041
rect 17866 6967 17922 6976
rect 17776 6724 17828 6730
rect 17776 6666 17828 6672
rect 17684 6656 17736 6662
rect 17682 6624 17684 6633
rect 17736 6624 17738 6633
rect 17682 6559 17738 6568
rect 17880 6458 17908 6967
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17684 6452 17736 6458
rect 17684 6394 17736 6400
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17592 6316 17644 6322
rect 17592 6258 17644 6264
rect 17696 5370 17724 6394
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17880 5574 17908 6258
rect 17972 5914 18000 6802
rect 18050 6760 18106 6769
rect 18050 6695 18106 6704
rect 18064 6304 18092 6695
rect 18156 6662 18184 8191
rect 18236 6928 18288 6934
rect 18236 6870 18288 6876
rect 18144 6656 18196 6662
rect 18144 6598 18196 6604
rect 18144 6316 18196 6322
rect 18064 6276 18144 6304
rect 18144 6258 18196 6264
rect 18050 6216 18106 6225
rect 18050 6151 18052 6160
rect 18104 6151 18106 6160
rect 18052 6122 18104 6128
rect 17960 5908 18012 5914
rect 17960 5850 18012 5856
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 18064 5273 18092 5510
rect 18050 5264 18106 5273
rect 18156 5234 18184 6258
rect 18248 5710 18276 6870
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18248 5370 18276 5646
rect 18236 5364 18288 5370
rect 18236 5306 18288 5312
rect 18050 5199 18106 5208
rect 18144 5228 18196 5234
rect 18144 5170 18196 5176
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17880 4049 17908 4422
rect 17866 4040 17922 4049
rect 17866 3975 17922 3984
rect 17500 3936 17552 3942
rect 17500 3878 17552 3884
rect 17512 3534 17540 3878
rect 17500 3528 17552 3534
rect 17500 3470 17552 3476
rect 17512 1970 17540 3470
rect 17972 3097 18000 4490
rect 18064 4457 18092 4966
rect 18340 4865 18368 8298
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18432 7449 18460 7482
rect 18418 7440 18474 7449
rect 18418 7375 18474 7384
rect 18420 7336 18472 7342
rect 18418 7304 18420 7313
rect 18472 7304 18474 7313
rect 18418 7239 18474 7248
rect 18432 6254 18460 7239
rect 18420 6248 18472 6254
rect 18420 6190 18472 6196
rect 18418 5672 18474 5681
rect 18418 5607 18474 5616
rect 18432 5574 18460 5607
rect 18420 5568 18472 5574
rect 18420 5510 18472 5516
rect 18326 4856 18382 4865
rect 18326 4791 18382 4800
rect 18326 4720 18382 4729
rect 18326 4655 18382 4664
rect 18340 4486 18368 4655
rect 18328 4480 18380 4486
rect 18050 4448 18106 4457
rect 18328 4422 18380 4428
rect 18050 4383 18106 4392
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18144 3664 18196 3670
rect 18144 3606 18196 3612
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18064 3233 18092 3334
rect 18050 3224 18106 3233
rect 18050 3159 18106 3168
rect 17958 3088 18014 3097
rect 17958 3023 18014 3032
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 17500 1964 17552 1970
rect 17500 1906 17552 1912
rect 17420 1822 17632 1850
rect 17314 1799 17370 1808
rect 17604 800 17632 1822
rect 17696 1465 17724 2790
rect 17972 2446 18000 3023
rect 18052 2848 18104 2854
rect 18052 2790 18104 2796
rect 18064 2689 18092 2790
rect 18050 2680 18106 2689
rect 18050 2615 18106 2624
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 17868 2304 17920 2310
rect 17868 2246 17920 2252
rect 17682 1456 17738 1465
rect 17682 1391 17738 1400
rect 17880 1057 17908 2246
rect 17866 1048 17922 1057
rect 17866 983 17922 992
rect 16776 734 16988 762
rect 17590 0 17646 800
rect 18156 649 18184 3606
rect 18248 3534 18276 3878
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18248 2582 18276 3470
rect 18340 3058 18368 4422
rect 18420 3664 18472 3670
rect 18418 3632 18420 3641
rect 18472 3632 18474 3641
rect 18418 3567 18474 3576
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 18236 2576 18288 2582
rect 18236 2518 18288 2524
rect 18236 2304 18288 2310
rect 18234 2272 18236 2281
rect 18288 2272 18290 2281
rect 18234 2207 18290 2216
rect 18524 800 18552 14010
rect 18800 14006 18828 16400
rect 18788 14000 18840 14006
rect 18788 13942 18840 13948
rect 18696 13252 18748 13258
rect 18696 13194 18748 13200
rect 18602 10024 18658 10033
rect 18602 9959 18604 9968
rect 18656 9959 18658 9968
rect 18604 9930 18656 9936
rect 18708 2922 18736 13194
rect 19432 3460 19484 3466
rect 19432 3402 19484 3408
rect 18696 2916 18748 2922
rect 18696 2858 18748 2864
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18142 640 18198 649
rect 18142 575 18198 584
rect 18510 0 18566 800
rect 18892 241 18920 2790
rect 19444 800 19472 3402
rect 18878 232 18934 241
rect 18878 167 18934 176
rect 19430 0 19486 800
<< via2 >>
rect 3698 16768 3754 16824
rect 3514 16360 3570 16416
rect 1582 15136 1638 15192
rect 2778 14728 2834 14784
rect 3180 14714 3236 14716
rect 3260 14714 3316 14716
rect 3340 14714 3396 14716
rect 3420 14714 3476 14716
rect 3180 14662 3226 14714
rect 3226 14662 3236 14714
rect 3260 14662 3290 14714
rect 3290 14662 3302 14714
rect 3302 14662 3316 14714
rect 3340 14662 3354 14714
rect 3354 14662 3366 14714
rect 3366 14662 3396 14714
rect 3420 14662 3430 14714
rect 3430 14662 3476 14714
rect 3180 14660 3236 14662
rect 3260 14660 3316 14662
rect 3340 14660 3396 14662
rect 3420 14660 3476 14662
rect 3180 13626 3236 13628
rect 3260 13626 3316 13628
rect 3340 13626 3396 13628
rect 3420 13626 3476 13628
rect 3180 13574 3226 13626
rect 3226 13574 3236 13626
rect 3260 13574 3290 13626
rect 3290 13574 3302 13626
rect 3302 13574 3316 13626
rect 3340 13574 3354 13626
rect 3354 13574 3366 13626
rect 3366 13574 3396 13626
rect 3420 13574 3430 13626
rect 3430 13574 3476 13626
rect 3180 13572 3236 13574
rect 3260 13572 3316 13574
rect 3340 13572 3396 13574
rect 3420 13572 3476 13574
rect 4066 15952 4122 16008
rect 3974 15544 4030 15600
rect 3790 13912 3846 13968
rect 3606 13232 3662 13288
rect 4066 14320 4122 14376
rect 4066 13368 4122 13424
rect 2134 12588 2136 12608
rect 2136 12588 2188 12608
rect 2188 12588 2190 12608
rect 1582 12416 1638 12472
rect 1306 9324 1308 9344
rect 1308 9324 1360 9344
rect 1360 9324 1362 9344
rect 1306 9288 1362 9324
rect 938 5072 994 5128
rect 938 2896 994 2952
rect 1490 8472 1546 8528
rect 1766 10784 1822 10840
rect 1674 7656 1730 7712
rect 1674 7404 1730 7440
rect 1674 7384 1676 7404
rect 1676 7384 1728 7404
rect 1728 7384 1730 7404
rect 1490 6432 1546 6488
rect 1398 6024 1454 6080
rect 2134 12552 2190 12588
rect 2042 9696 2098 9752
rect 2318 11328 2374 11384
rect 1858 7656 1914 7712
rect 1674 3984 1730 4040
rect 3180 12538 3236 12540
rect 3260 12538 3316 12540
rect 3340 12538 3396 12540
rect 3420 12538 3476 12540
rect 3180 12486 3226 12538
rect 3226 12486 3236 12538
rect 3260 12486 3290 12538
rect 3290 12486 3302 12538
rect 3302 12486 3316 12538
rect 3340 12486 3354 12538
rect 3354 12486 3366 12538
rect 3366 12486 3396 12538
rect 3420 12486 3430 12538
rect 3430 12486 3476 12538
rect 3180 12484 3236 12486
rect 3260 12484 3316 12486
rect 3340 12484 3396 12486
rect 3420 12484 3476 12486
rect 2410 6432 2466 6488
rect 2318 6160 2374 6216
rect 2134 3984 2190 4040
rect 2226 3304 2282 3360
rect 2318 2624 2374 2680
rect 3514 11772 3516 11792
rect 3516 11772 3568 11792
rect 3568 11772 3570 11792
rect 3514 11736 3570 11772
rect 3180 11450 3236 11452
rect 3260 11450 3316 11452
rect 3340 11450 3396 11452
rect 3420 11450 3476 11452
rect 3180 11398 3226 11450
rect 3226 11398 3236 11450
rect 3260 11398 3290 11450
rect 3290 11398 3302 11450
rect 3302 11398 3316 11450
rect 3340 11398 3354 11450
rect 3354 11398 3366 11450
rect 3366 11398 3396 11450
rect 3420 11398 3430 11450
rect 3430 11398 3476 11450
rect 3180 11396 3236 11398
rect 3260 11396 3316 11398
rect 3340 11396 3396 11398
rect 3420 11396 3476 11398
rect 3180 10362 3236 10364
rect 3260 10362 3316 10364
rect 3340 10362 3396 10364
rect 3420 10362 3476 10364
rect 3180 10310 3226 10362
rect 3226 10310 3236 10362
rect 3260 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3316 10362
rect 3340 10310 3354 10362
rect 3354 10310 3366 10362
rect 3366 10310 3396 10362
rect 3420 10310 3430 10362
rect 3430 10310 3476 10362
rect 3180 10308 3236 10310
rect 3260 10308 3316 10310
rect 3340 10308 3396 10310
rect 3420 10308 3476 10310
rect 3054 9696 3110 9752
rect 3180 9274 3236 9276
rect 3260 9274 3316 9276
rect 3340 9274 3396 9276
rect 3420 9274 3476 9276
rect 3180 9222 3226 9274
rect 3226 9222 3236 9274
rect 3260 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3316 9274
rect 3340 9222 3354 9274
rect 3354 9222 3366 9274
rect 3366 9222 3396 9274
rect 3420 9222 3430 9274
rect 3430 9222 3476 9274
rect 3180 9220 3236 9222
rect 3260 9220 3316 9222
rect 3340 9220 3396 9222
rect 3420 9220 3476 9222
rect 3514 8880 3570 8936
rect 2870 8064 2926 8120
rect 2686 6704 2742 6760
rect 3180 8186 3236 8188
rect 3260 8186 3316 8188
rect 3340 8186 3396 8188
rect 3420 8186 3476 8188
rect 3180 8134 3226 8186
rect 3226 8134 3236 8186
rect 3260 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3316 8186
rect 3340 8134 3354 8186
rect 3354 8134 3366 8186
rect 3366 8134 3396 8186
rect 3420 8134 3430 8186
rect 3430 8134 3476 8186
rect 3180 8132 3236 8134
rect 3260 8132 3316 8134
rect 3340 8132 3396 8134
rect 3420 8132 3476 8134
rect 3330 7692 3332 7712
rect 3332 7692 3384 7712
rect 3384 7692 3386 7712
rect 3330 7656 3386 7692
rect 3180 7098 3236 7100
rect 3260 7098 3316 7100
rect 3340 7098 3396 7100
rect 3420 7098 3476 7100
rect 3180 7046 3226 7098
rect 3226 7046 3236 7098
rect 3260 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3316 7098
rect 3340 7046 3354 7098
rect 3354 7046 3366 7098
rect 3366 7046 3396 7098
rect 3420 7046 3430 7098
rect 3430 7046 3476 7098
rect 3180 7044 3236 7046
rect 3260 7044 3316 7046
rect 3340 7044 3396 7046
rect 3420 7044 3476 7046
rect 3054 6160 3110 6216
rect 3882 11872 3938 11928
rect 3790 10920 3846 10976
rect 4066 11872 4122 11928
rect 4158 11228 4160 11248
rect 4160 11228 4212 11248
rect 4212 11228 4214 11248
rect 4158 11192 4214 11228
rect 4066 10104 4122 10160
rect 2870 3848 2926 3904
rect 3180 6010 3236 6012
rect 3260 6010 3316 6012
rect 3340 6010 3396 6012
rect 3420 6010 3476 6012
rect 3180 5958 3226 6010
rect 3226 5958 3236 6010
rect 3260 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3316 6010
rect 3340 5958 3354 6010
rect 3354 5958 3366 6010
rect 3366 5958 3396 6010
rect 3420 5958 3430 6010
rect 3430 5958 3476 6010
rect 3180 5956 3236 5958
rect 3260 5956 3316 5958
rect 3340 5956 3396 5958
rect 3420 5956 3476 5958
rect 2870 1944 2926 2000
rect 3180 4922 3236 4924
rect 3260 4922 3316 4924
rect 3340 4922 3396 4924
rect 3420 4922 3476 4924
rect 3180 4870 3226 4922
rect 3226 4870 3236 4922
rect 3260 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3316 4922
rect 3340 4870 3354 4922
rect 3354 4870 3366 4922
rect 3366 4870 3396 4922
rect 3420 4870 3430 4922
rect 3430 4870 3476 4922
rect 3180 4868 3236 4870
rect 3260 4868 3316 4870
rect 3340 4868 3396 4870
rect 3420 4868 3476 4870
rect 3180 3834 3236 3836
rect 3260 3834 3316 3836
rect 3340 3834 3396 3836
rect 3420 3834 3476 3836
rect 3180 3782 3226 3834
rect 3226 3782 3236 3834
rect 3260 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3316 3834
rect 3340 3782 3354 3834
rect 3354 3782 3366 3834
rect 3366 3782 3396 3834
rect 3420 3782 3430 3834
rect 3430 3782 3476 3834
rect 3180 3780 3236 3782
rect 3260 3780 3316 3782
rect 3340 3780 3396 3782
rect 3420 3780 3476 3782
rect 3698 4936 3754 4992
rect 3974 8608 4030 8664
rect 5404 14170 5460 14172
rect 5484 14170 5540 14172
rect 5564 14170 5620 14172
rect 5644 14170 5700 14172
rect 5404 14118 5450 14170
rect 5450 14118 5460 14170
rect 5484 14118 5514 14170
rect 5514 14118 5526 14170
rect 5526 14118 5540 14170
rect 5564 14118 5578 14170
rect 5578 14118 5590 14170
rect 5590 14118 5620 14170
rect 5644 14118 5654 14170
rect 5654 14118 5700 14170
rect 5404 14116 5460 14118
rect 5484 14116 5540 14118
rect 5564 14116 5620 14118
rect 5644 14116 5700 14118
rect 4526 13096 4582 13152
rect 4342 10668 4398 10704
rect 4342 10648 4344 10668
rect 4344 10648 4396 10668
rect 4396 10648 4398 10668
rect 4250 8508 4252 8528
rect 4252 8508 4304 8528
rect 4304 8508 4306 8528
rect 4250 8472 4306 8508
rect 4526 10648 4582 10704
rect 3882 7248 3938 7304
rect 3882 6840 3938 6896
rect 3882 5888 3938 5944
rect 3882 4820 3938 4856
rect 3882 4800 3884 4820
rect 3884 4800 3936 4820
rect 3936 4800 3938 4820
rect 3882 4664 3938 4720
rect 3974 3848 4030 3904
rect 3974 3712 4030 3768
rect 3790 3576 3846 3632
rect 3180 2746 3236 2748
rect 3260 2746 3316 2748
rect 3340 2746 3396 2748
rect 3420 2746 3476 2748
rect 3180 2694 3226 2746
rect 3226 2694 3236 2746
rect 3260 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3316 2746
rect 3340 2694 3354 2746
rect 3354 2694 3366 2746
rect 3366 2694 3396 2746
rect 3420 2694 3430 2746
rect 3430 2694 3476 2746
rect 3180 2692 3236 2694
rect 3260 2692 3316 2694
rect 3340 2692 3396 2694
rect 3420 2692 3476 2694
rect 5404 13082 5460 13084
rect 5484 13082 5540 13084
rect 5564 13082 5620 13084
rect 5644 13082 5700 13084
rect 5404 13030 5450 13082
rect 5450 13030 5460 13082
rect 5484 13030 5514 13082
rect 5514 13030 5526 13082
rect 5526 13030 5540 13082
rect 5564 13030 5578 13082
rect 5578 13030 5590 13082
rect 5590 13030 5620 13082
rect 5644 13030 5654 13082
rect 5654 13030 5700 13082
rect 5404 13028 5460 13030
rect 5484 13028 5540 13030
rect 5564 13028 5620 13030
rect 5644 13028 5700 13030
rect 5404 11994 5460 11996
rect 5484 11994 5540 11996
rect 5564 11994 5620 11996
rect 5644 11994 5700 11996
rect 5404 11942 5450 11994
rect 5450 11942 5460 11994
rect 5484 11942 5514 11994
rect 5514 11942 5526 11994
rect 5526 11942 5540 11994
rect 5564 11942 5578 11994
rect 5578 11942 5590 11994
rect 5590 11942 5620 11994
rect 5644 11942 5654 11994
rect 5654 11942 5700 11994
rect 5404 11940 5460 11942
rect 5484 11940 5540 11942
rect 5564 11940 5620 11942
rect 5644 11940 5700 11942
rect 5404 10906 5460 10908
rect 5484 10906 5540 10908
rect 5564 10906 5620 10908
rect 5644 10906 5700 10908
rect 5404 10854 5450 10906
rect 5450 10854 5460 10906
rect 5484 10854 5514 10906
rect 5514 10854 5526 10906
rect 5526 10854 5540 10906
rect 5564 10854 5578 10906
rect 5578 10854 5590 10906
rect 5590 10854 5620 10906
rect 5644 10854 5654 10906
rect 5654 10854 5700 10906
rect 5404 10852 5460 10854
rect 5484 10852 5540 10854
rect 5564 10852 5620 10854
rect 5644 10852 5700 10854
rect 5170 9324 5172 9344
rect 5172 9324 5224 9344
rect 5224 9324 5226 9344
rect 5170 9288 5226 9324
rect 5404 9818 5460 9820
rect 5484 9818 5540 9820
rect 5564 9818 5620 9820
rect 5644 9818 5700 9820
rect 5404 9766 5450 9818
rect 5450 9766 5460 9818
rect 5484 9766 5514 9818
rect 5514 9766 5526 9818
rect 5526 9766 5540 9818
rect 5564 9766 5578 9818
rect 5578 9766 5590 9818
rect 5590 9766 5620 9818
rect 5644 9766 5654 9818
rect 5654 9766 5700 9818
rect 5404 9764 5460 9766
rect 5484 9764 5540 9766
rect 5564 9764 5620 9766
rect 5644 9764 5700 9766
rect 5630 8880 5686 8936
rect 5404 8730 5460 8732
rect 5484 8730 5540 8732
rect 5564 8730 5620 8732
rect 5644 8730 5700 8732
rect 5404 8678 5450 8730
rect 5450 8678 5460 8730
rect 5484 8678 5514 8730
rect 5514 8678 5526 8730
rect 5526 8678 5540 8730
rect 5564 8678 5578 8730
rect 5578 8678 5590 8730
rect 5590 8678 5620 8730
rect 5644 8678 5654 8730
rect 5654 8678 5700 8730
rect 5404 8676 5460 8678
rect 5484 8676 5540 8678
rect 5564 8676 5620 8678
rect 5644 8676 5700 8678
rect 4526 6316 4582 6352
rect 4526 6296 4528 6316
rect 4528 6296 4580 6316
rect 4580 6296 4582 6316
rect 4342 6024 4398 6080
rect 4434 5208 4490 5264
rect 4158 3440 4214 3496
rect 4434 3984 4490 4040
rect 4434 3612 4436 3632
rect 4436 3612 4488 3632
rect 4488 3612 4490 3632
rect 4434 3576 4490 3612
rect 4618 5480 4674 5536
rect 5404 7642 5460 7644
rect 5484 7642 5540 7644
rect 5564 7642 5620 7644
rect 5644 7642 5700 7644
rect 5404 7590 5450 7642
rect 5450 7590 5460 7642
rect 5484 7590 5514 7642
rect 5514 7590 5526 7642
rect 5526 7590 5540 7642
rect 5564 7590 5578 7642
rect 5578 7590 5590 7642
rect 5590 7590 5620 7642
rect 5644 7590 5654 7642
rect 5654 7590 5700 7642
rect 5404 7588 5460 7590
rect 5484 7588 5540 7590
rect 5564 7588 5620 7590
rect 5644 7588 5700 7590
rect 5078 5888 5134 5944
rect 4986 5480 5042 5536
rect 4802 3848 4858 3904
rect 3882 2216 3938 2272
rect 3330 1436 3332 1456
rect 3332 1436 3384 1456
rect 3384 1436 3386 1456
rect 3330 1400 3386 1436
rect 2778 176 2834 232
rect 4342 2508 4398 2544
rect 4342 2488 4344 2508
rect 4344 2488 4396 2508
rect 4396 2488 4398 2508
rect 4986 3712 5042 3768
rect 5630 7112 5686 7168
rect 5630 6840 5686 6896
rect 5404 6554 5460 6556
rect 5484 6554 5540 6556
rect 5564 6554 5620 6556
rect 5644 6554 5700 6556
rect 5404 6502 5450 6554
rect 5450 6502 5460 6554
rect 5484 6502 5514 6554
rect 5514 6502 5526 6554
rect 5526 6502 5540 6554
rect 5564 6502 5578 6554
rect 5578 6502 5590 6554
rect 5590 6502 5620 6554
rect 5644 6502 5654 6554
rect 5654 6502 5700 6554
rect 5404 6500 5460 6502
rect 5484 6500 5540 6502
rect 5564 6500 5620 6502
rect 5644 6500 5700 6502
rect 5404 5466 5460 5468
rect 5484 5466 5540 5468
rect 5564 5466 5620 5468
rect 5644 5466 5700 5468
rect 5404 5414 5450 5466
rect 5450 5414 5460 5466
rect 5484 5414 5514 5466
rect 5514 5414 5526 5466
rect 5526 5414 5540 5466
rect 5564 5414 5578 5466
rect 5578 5414 5590 5466
rect 5590 5414 5620 5466
rect 5644 5414 5654 5466
rect 5654 5414 5700 5466
rect 5404 5412 5460 5414
rect 5484 5412 5540 5414
rect 5564 5412 5620 5414
rect 5644 5412 5700 5414
rect 5404 4378 5460 4380
rect 5484 4378 5540 4380
rect 5564 4378 5620 4380
rect 5644 4378 5700 4380
rect 5404 4326 5450 4378
rect 5450 4326 5460 4378
rect 5484 4326 5514 4378
rect 5514 4326 5526 4378
rect 5526 4326 5540 4378
rect 5564 4326 5578 4378
rect 5578 4326 5590 4378
rect 5590 4326 5620 4378
rect 5644 4326 5654 4378
rect 5654 4326 5700 4378
rect 5404 4324 5460 4326
rect 5484 4324 5540 4326
rect 5564 4324 5620 4326
rect 5644 4324 5700 4326
rect 5262 3712 5318 3768
rect 5998 9988 6054 10024
rect 5998 9968 6000 9988
rect 6000 9968 6052 9988
rect 6052 9968 6054 9988
rect 6458 10512 6514 10568
rect 6090 8880 6146 8936
rect 6182 7248 6238 7304
rect 5170 3304 5226 3360
rect 5404 3290 5460 3292
rect 5484 3290 5540 3292
rect 5564 3290 5620 3292
rect 5644 3290 5700 3292
rect 5404 3238 5450 3290
rect 5450 3238 5460 3290
rect 5484 3238 5514 3290
rect 5514 3238 5526 3290
rect 5526 3238 5540 3290
rect 5564 3238 5578 3290
rect 5578 3238 5590 3290
rect 5590 3238 5620 3290
rect 5644 3238 5654 3290
rect 5654 3238 5700 3290
rect 5404 3236 5460 3238
rect 5484 3236 5540 3238
rect 5564 3236 5620 3238
rect 5644 3236 5700 3238
rect 5538 3052 5594 3088
rect 5538 3032 5540 3052
rect 5540 3032 5592 3052
rect 5592 3032 5594 3052
rect 4710 2352 4766 2408
rect 4618 2216 4674 2272
rect 4066 1844 4068 1864
rect 4068 1844 4120 1864
rect 4120 1844 4122 1864
rect 4066 1808 4122 1844
rect 5538 2624 5594 2680
rect 5722 2488 5778 2544
rect 5404 2202 5460 2204
rect 5484 2202 5540 2204
rect 5564 2202 5620 2204
rect 5644 2202 5700 2204
rect 5404 2150 5450 2202
rect 5450 2150 5460 2202
rect 5484 2150 5514 2202
rect 5514 2150 5526 2202
rect 5526 2150 5540 2202
rect 5564 2150 5578 2202
rect 5578 2150 5590 2202
rect 5590 2150 5620 2202
rect 5644 2150 5654 2202
rect 5654 2150 5700 2202
rect 5404 2148 5460 2150
rect 5484 2148 5540 2150
rect 5564 2148 5620 2150
rect 5644 2148 5700 2150
rect 5906 2488 5962 2544
rect 4066 1028 4068 1048
rect 4068 1028 4120 1048
rect 4120 1028 4122 1048
rect 4066 992 4122 1028
rect 3698 584 3754 640
rect 6274 3304 6330 3360
rect 6918 11600 6974 11656
rect 6918 11056 6974 11112
rect 6642 9968 6698 10024
rect 6642 6160 6698 6216
rect 6550 5616 6606 5672
rect 6918 8356 6974 8392
rect 6918 8336 6920 8356
rect 6920 8336 6972 8356
rect 6972 8336 6974 8356
rect 7010 7792 7066 7848
rect 6918 7540 6974 7576
rect 6918 7520 6920 7540
rect 6920 7520 6972 7540
rect 6972 7520 6974 7540
rect 6918 6740 6920 6760
rect 6920 6740 6972 6760
rect 6972 6740 6974 6760
rect 6918 6704 6974 6740
rect 6918 6604 6920 6624
rect 6920 6604 6972 6624
rect 6972 6604 6974 6624
rect 6918 6568 6974 6604
rect 6550 4020 6552 4040
rect 6552 4020 6604 4040
rect 6604 4020 6606 4040
rect 6550 3984 6606 4020
rect 6918 3168 6974 3224
rect 6918 2252 6920 2272
rect 6920 2252 6972 2272
rect 6972 2252 6974 2272
rect 6918 2216 6974 2252
rect 7628 14714 7684 14716
rect 7708 14714 7764 14716
rect 7788 14714 7844 14716
rect 7868 14714 7924 14716
rect 7628 14662 7674 14714
rect 7674 14662 7684 14714
rect 7708 14662 7738 14714
rect 7738 14662 7750 14714
rect 7750 14662 7764 14714
rect 7788 14662 7802 14714
rect 7802 14662 7814 14714
rect 7814 14662 7844 14714
rect 7868 14662 7878 14714
rect 7878 14662 7924 14714
rect 7628 14660 7684 14662
rect 7708 14660 7764 14662
rect 7788 14660 7844 14662
rect 7868 14660 7924 14662
rect 7628 13626 7684 13628
rect 7708 13626 7764 13628
rect 7788 13626 7844 13628
rect 7868 13626 7924 13628
rect 7628 13574 7674 13626
rect 7674 13574 7684 13626
rect 7708 13574 7738 13626
rect 7738 13574 7750 13626
rect 7750 13574 7764 13626
rect 7788 13574 7802 13626
rect 7802 13574 7814 13626
rect 7814 13574 7844 13626
rect 7868 13574 7878 13626
rect 7878 13574 7924 13626
rect 7628 13572 7684 13574
rect 7708 13572 7764 13574
rect 7788 13572 7844 13574
rect 7868 13572 7924 13574
rect 7628 12538 7684 12540
rect 7708 12538 7764 12540
rect 7788 12538 7844 12540
rect 7868 12538 7924 12540
rect 7628 12486 7674 12538
rect 7674 12486 7684 12538
rect 7708 12486 7738 12538
rect 7738 12486 7750 12538
rect 7750 12486 7764 12538
rect 7788 12486 7802 12538
rect 7802 12486 7814 12538
rect 7814 12486 7844 12538
rect 7868 12486 7878 12538
rect 7878 12486 7924 12538
rect 7628 12484 7684 12486
rect 7708 12484 7764 12486
rect 7788 12484 7844 12486
rect 7868 12484 7924 12486
rect 7628 11450 7684 11452
rect 7708 11450 7764 11452
rect 7788 11450 7844 11452
rect 7868 11450 7924 11452
rect 7628 11398 7674 11450
rect 7674 11398 7684 11450
rect 7708 11398 7738 11450
rect 7738 11398 7750 11450
rect 7750 11398 7764 11450
rect 7788 11398 7802 11450
rect 7802 11398 7814 11450
rect 7814 11398 7844 11450
rect 7868 11398 7878 11450
rect 7878 11398 7924 11450
rect 7628 11396 7684 11398
rect 7708 11396 7764 11398
rect 7788 11396 7844 11398
rect 7868 11396 7924 11398
rect 7628 10362 7684 10364
rect 7708 10362 7764 10364
rect 7788 10362 7844 10364
rect 7868 10362 7924 10364
rect 7628 10310 7674 10362
rect 7674 10310 7684 10362
rect 7708 10310 7738 10362
rect 7738 10310 7750 10362
rect 7750 10310 7764 10362
rect 7788 10310 7802 10362
rect 7802 10310 7814 10362
rect 7814 10310 7844 10362
rect 7868 10310 7878 10362
rect 7878 10310 7924 10362
rect 7628 10308 7684 10310
rect 7708 10308 7764 10310
rect 7788 10308 7844 10310
rect 7868 10308 7924 10310
rect 7562 10140 7564 10160
rect 7564 10140 7616 10160
rect 7616 10140 7618 10160
rect 7562 10104 7618 10140
rect 7286 9288 7342 9344
rect 7628 9274 7684 9276
rect 7708 9274 7764 9276
rect 7788 9274 7844 9276
rect 7868 9274 7924 9276
rect 7628 9222 7674 9274
rect 7674 9222 7684 9274
rect 7708 9222 7738 9274
rect 7738 9222 7750 9274
rect 7750 9222 7764 9274
rect 7788 9222 7802 9274
rect 7802 9222 7814 9274
rect 7814 9222 7844 9274
rect 7868 9222 7878 9274
rect 7878 9222 7924 9274
rect 7628 9220 7684 9222
rect 7708 9220 7764 9222
rect 7788 9220 7844 9222
rect 7868 9220 7924 9222
rect 7628 8186 7684 8188
rect 7708 8186 7764 8188
rect 7788 8186 7844 8188
rect 7868 8186 7924 8188
rect 7628 8134 7674 8186
rect 7674 8134 7684 8186
rect 7708 8134 7738 8186
rect 7738 8134 7750 8186
rect 7750 8134 7764 8186
rect 7788 8134 7802 8186
rect 7802 8134 7814 8186
rect 7814 8134 7844 8186
rect 7868 8134 7878 8186
rect 7878 8134 7924 8186
rect 7628 8132 7684 8134
rect 7708 8132 7764 8134
rect 7788 8132 7844 8134
rect 7868 8132 7924 8134
rect 7378 7112 7434 7168
rect 7628 7098 7684 7100
rect 7708 7098 7764 7100
rect 7788 7098 7844 7100
rect 7868 7098 7924 7100
rect 7628 7046 7674 7098
rect 7674 7046 7684 7098
rect 7708 7046 7738 7098
rect 7738 7046 7750 7098
rect 7750 7046 7764 7098
rect 7788 7046 7802 7098
rect 7802 7046 7814 7098
rect 7814 7046 7844 7098
rect 7868 7046 7878 7098
rect 7878 7046 7924 7098
rect 7628 7044 7684 7046
rect 7708 7044 7764 7046
rect 7788 7044 7844 7046
rect 7868 7044 7924 7046
rect 8298 10104 8354 10160
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9898 14170
rect 9898 14118 9908 14170
rect 9932 14118 9962 14170
rect 9962 14118 9974 14170
rect 9974 14118 9988 14170
rect 10012 14118 10026 14170
rect 10026 14118 10038 14170
rect 10038 14118 10068 14170
rect 10092 14118 10102 14170
rect 10102 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9898 13082
rect 9898 13030 9908 13082
rect 9932 13030 9962 13082
rect 9962 13030 9974 13082
rect 9974 13030 9988 13082
rect 10012 13030 10026 13082
rect 10026 13030 10038 13082
rect 10038 13030 10068 13082
rect 10092 13030 10102 13082
rect 10102 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9402 12144 9458 12200
rect 8850 11600 8906 11656
rect 18050 16768 18106 16824
rect 12076 14714 12132 14716
rect 12156 14714 12212 14716
rect 12236 14714 12292 14716
rect 12316 14714 12372 14716
rect 12076 14662 12122 14714
rect 12122 14662 12132 14714
rect 12156 14662 12186 14714
rect 12186 14662 12198 14714
rect 12198 14662 12212 14714
rect 12236 14662 12250 14714
rect 12250 14662 12262 14714
rect 12262 14662 12292 14714
rect 12316 14662 12326 14714
rect 12326 14662 12372 14714
rect 12076 14660 12132 14662
rect 12156 14660 12212 14662
rect 12236 14660 12292 14662
rect 12316 14660 12372 14662
rect 12076 13626 12132 13628
rect 12156 13626 12212 13628
rect 12236 13626 12292 13628
rect 12316 13626 12372 13628
rect 12076 13574 12122 13626
rect 12122 13574 12132 13626
rect 12156 13574 12186 13626
rect 12186 13574 12198 13626
rect 12198 13574 12212 13626
rect 12236 13574 12250 13626
rect 12250 13574 12262 13626
rect 12262 13574 12292 13626
rect 12316 13574 12326 13626
rect 12326 13574 12372 13626
rect 12076 13572 12132 13574
rect 12156 13572 12212 13574
rect 12236 13572 12292 13574
rect 12316 13572 12372 13574
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9898 11994
rect 9898 11942 9908 11994
rect 9932 11942 9962 11994
rect 9962 11942 9974 11994
rect 9974 11942 9988 11994
rect 10012 11942 10026 11994
rect 10026 11942 10038 11994
rect 10038 11942 10068 11994
rect 10092 11942 10102 11994
rect 10102 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 10506 11872 10562 11928
rect 9954 11328 10010 11384
rect 10506 11464 10562 11520
rect 8850 10104 8906 10160
rect 7470 6024 7526 6080
rect 7628 6010 7684 6012
rect 7708 6010 7764 6012
rect 7788 6010 7844 6012
rect 7868 6010 7924 6012
rect 7628 5958 7674 6010
rect 7674 5958 7684 6010
rect 7708 5958 7738 6010
rect 7738 5958 7750 6010
rect 7750 5958 7764 6010
rect 7788 5958 7802 6010
rect 7802 5958 7814 6010
rect 7814 5958 7844 6010
rect 7868 5958 7878 6010
rect 7878 5958 7924 6010
rect 7628 5956 7684 5958
rect 7708 5956 7764 5958
rect 7788 5956 7844 5958
rect 7868 5956 7924 5958
rect 7194 4936 7250 4992
rect 8114 6296 8170 6352
rect 7562 5480 7618 5536
rect 7628 4922 7684 4924
rect 7708 4922 7764 4924
rect 7788 4922 7844 4924
rect 7868 4922 7924 4924
rect 7628 4870 7674 4922
rect 7674 4870 7684 4922
rect 7708 4870 7738 4922
rect 7738 4870 7750 4922
rect 7750 4870 7764 4922
rect 7788 4870 7802 4922
rect 7802 4870 7814 4922
rect 7814 4870 7844 4922
rect 7868 4870 7878 4922
rect 7878 4870 7924 4922
rect 7628 4868 7684 4870
rect 7708 4868 7764 4870
rect 7788 4868 7844 4870
rect 7868 4868 7924 4870
rect 7628 3834 7684 3836
rect 7708 3834 7764 3836
rect 7788 3834 7844 3836
rect 7868 3834 7924 3836
rect 7628 3782 7674 3834
rect 7674 3782 7684 3834
rect 7708 3782 7738 3834
rect 7738 3782 7750 3834
rect 7750 3782 7764 3834
rect 7788 3782 7802 3834
rect 7802 3782 7814 3834
rect 7814 3782 7844 3834
rect 7868 3782 7878 3834
rect 7878 3782 7924 3834
rect 7628 3780 7684 3782
rect 7708 3780 7764 3782
rect 7788 3780 7844 3782
rect 7868 3780 7924 3782
rect 7470 3304 7526 3360
rect 7378 3052 7434 3088
rect 7378 3032 7380 3052
rect 7380 3032 7432 3052
rect 7432 3032 7434 3052
rect 7654 3052 7710 3088
rect 7654 3032 7656 3052
rect 7656 3032 7708 3052
rect 7708 3032 7710 3052
rect 7628 2746 7684 2748
rect 7708 2746 7764 2748
rect 7788 2746 7844 2748
rect 7868 2746 7924 2748
rect 7628 2694 7674 2746
rect 7674 2694 7684 2746
rect 7708 2694 7738 2746
rect 7738 2694 7750 2746
rect 7750 2694 7764 2746
rect 7788 2694 7802 2746
rect 7802 2694 7814 2746
rect 7814 2694 7844 2746
rect 7868 2694 7878 2746
rect 7878 2694 7924 2746
rect 7628 2692 7684 2694
rect 7708 2692 7764 2694
rect 7788 2692 7844 2694
rect 7868 2692 7924 2694
rect 8666 7384 8722 7440
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9898 10906
rect 9898 10854 9908 10906
rect 9932 10854 9962 10906
rect 9962 10854 9974 10906
rect 9974 10854 9988 10906
rect 10012 10854 10026 10906
rect 10026 10854 10038 10906
rect 10038 10854 10068 10906
rect 10092 10854 10102 10906
rect 10102 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 10782 11328 10838 11384
rect 10506 10104 10562 10160
rect 10230 9988 10286 10024
rect 10230 9968 10232 9988
rect 10232 9968 10284 9988
rect 10284 9968 10286 9988
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9898 9818
rect 9898 9766 9908 9818
rect 9932 9766 9962 9818
rect 9962 9766 9974 9818
rect 9974 9766 9988 9818
rect 10012 9766 10026 9818
rect 10026 9766 10038 9818
rect 10038 9766 10068 9818
rect 10092 9766 10102 9818
rect 10102 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9402 8780 9404 8800
rect 9404 8780 9456 8800
rect 9456 8780 9458 8800
rect 9402 8744 9458 8780
rect 9034 7248 9090 7304
rect 8482 6296 8538 6352
rect 8574 6024 8630 6080
rect 8850 6296 8906 6352
rect 8758 5888 8814 5944
rect 9954 9016 10010 9072
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9898 8730
rect 9898 8678 9908 8730
rect 9932 8678 9962 8730
rect 9962 8678 9974 8730
rect 9974 8678 9988 8730
rect 10012 8678 10026 8730
rect 10026 8678 10038 8730
rect 10038 8678 10068 8730
rect 10092 8678 10102 8730
rect 10102 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 10506 8780 10508 8800
rect 10508 8780 10560 8800
rect 10560 8780 10562 8800
rect 10506 8744 10562 8780
rect 9678 7948 9734 7984
rect 9678 7928 9680 7948
rect 9680 7928 9732 7948
rect 9732 7928 9734 7948
rect 10506 7692 10508 7712
rect 10508 7692 10560 7712
rect 10560 7692 10562 7712
rect 10506 7656 10562 7692
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9898 7642
rect 9898 7590 9908 7642
rect 9932 7590 9962 7642
rect 9962 7590 9974 7642
rect 9974 7590 9988 7642
rect 10012 7590 10026 7642
rect 10026 7590 10038 7642
rect 10038 7590 10068 7642
rect 10092 7590 10102 7642
rect 10102 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 10506 7384 10562 7440
rect 8942 5516 8944 5536
rect 8944 5516 8996 5536
rect 8996 5516 8998 5536
rect 8390 4004 8446 4040
rect 8390 3984 8392 4004
rect 8392 3984 8444 4004
rect 8444 3984 8446 4004
rect 8574 4020 8576 4040
rect 8576 4020 8628 4040
rect 8628 4020 8630 4040
rect 8574 3984 8630 4020
rect 8942 5480 8998 5516
rect 8390 3440 8446 3496
rect 9310 6024 9366 6080
rect 9218 5616 9274 5672
rect 9218 4120 9274 4176
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9898 6554
rect 9898 6502 9908 6554
rect 9932 6502 9962 6554
rect 9962 6502 9974 6554
rect 9974 6502 9988 6554
rect 10012 6502 10026 6554
rect 10026 6502 10038 6554
rect 10038 6502 10068 6554
rect 10092 6502 10102 6554
rect 10102 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 9586 5752 9642 5808
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9898 5466
rect 9898 5414 9908 5466
rect 9932 5414 9962 5466
rect 9962 5414 9974 5466
rect 9974 5414 9988 5466
rect 10012 5414 10026 5466
rect 10026 5414 10038 5466
rect 10038 5414 10068 5466
rect 10092 5414 10102 5466
rect 10102 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 10138 5208 10194 5264
rect 9494 3984 9550 4040
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9898 4378
rect 9898 4326 9908 4378
rect 9932 4326 9962 4378
rect 9962 4326 9974 4378
rect 9974 4326 9988 4378
rect 10012 4326 10026 4378
rect 10026 4326 10038 4378
rect 10038 4326 10068 4378
rect 10092 4326 10102 4378
rect 10102 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9898 3290
rect 9898 3238 9908 3290
rect 9932 3238 9962 3290
rect 9962 3238 9974 3290
rect 9974 3238 9988 3290
rect 10012 3238 10026 3290
rect 10026 3238 10038 3290
rect 10038 3238 10068 3290
rect 10092 3238 10102 3290
rect 10102 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 11150 12280 11206 12336
rect 10966 8336 11022 8392
rect 10966 6432 11022 6488
rect 11150 7792 11206 7848
rect 11242 6296 11298 6352
rect 12076 12538 12132 12540
rect 12156 12538 12212 12540
rect 12236 12538 12292 12540
rect 12316 12538 12372 12540
rect 12076 12486 12122 12538
rect 12122 12486 12132 12538
rect 12156 12486 12186 12538
rect 12186 12486 12198 12538
rect 12198 12486 12212 12538
rect 12236 12486 12250 12538
rect 12250 12486 12262 12538
rect 12262 12486 12292 12538
rect 12316 12486 12326 12538
rect 12326 12486 12372 12538
rect 12076 12484 12132 12486
rect 12156 12484 12212 12486
rect 12236 12484 12292 12486
rect 12316 12484 12372 12486
rect 11886 11892 11942 11928
rect 11886 11872 11888 11892
rect 11888 11872 11940 11892
rect 11940 11872 11942 11892
rect 12438 11872 12494 11928
rect 12076 11450 12132 11452
rect 12156 11450 12212 11452
rect 12236 11450 12292 11452
rect 12316 11450 12372 11452
rect 12076 11398 12122 11450
rect 12122 11398 12132 11450
rect 12156 11398 12186 11450
rect 12186 11398 12198 11450
rect 12198 11398 12212 11450
rect 12236 11398 12250 11450
rect 12250 11398 12262 11450
rect 12262 11398 12292 11450
rect 12316 11398 12326 11450
rect 12326 11398 12372 11450
rect 12076 11396 12132 11398
rect 12156 11396 12212 11398
rect 12236 11396 12292 11398
rect 12316 11396 12372 11398
rect 11886 11328 11942 11384
rect 12254 11076 12310 11112
rect 12254 11056 12256 11076
rect 12256 11056 12308 11076
rect 12308 11056 12310 11076
rect 11702 8900 11758 8936
rect 11702 8880 11704 8900
rect 11704 8880 11756 8900
rect 11756 8880 11758 8900
rect 11518 8472 11574 8528
rect 11702 8472 11758 8528
rect 12076 10362 12132 10364
rect 12156 10362 12212 10364
rect 12236 10362 12292 10364
rect 12316 10362 12372 10364
rect 12076 10310 12122 10362
rect 12122 10310 12132 10362
rect 12156 10310 12186 10362
rect 12186 10310 12198 10362
rect 12198 10310 12212 10362
rect 12236 10310 12250 10362
rect 12250 10310 12262 10362
rect 12262 10310 12292 10362
rect 12316 10310 12326 10362
rect 12326 10310 12372 10362
rect 12076 10308 12132 10310
rect 12156 10308 12212 10310
rect 12236 10308 12292 10310
rect 12316 10308 12372 10310
rect 12070 9460 12072 9480
rect 12072 9460 12124 9480
rect 12124 9460 12126 9480
rect 12070 9424 12126 9460
rect 12076 9274 12132 9276
rect 12156 9274 12212 9276
rect 12236 9274 12292 9276
rect 12316 9274 12372 9276
rect 12076 9222 12122 9274
rect 12122 9222 12132 9274
rect 12156 9222 12186 9274
rect 12186 9222 12198 9274
rect 12198 9222 12212 9274
rect 12236 9222 12250 9274
rect 12250 9222 12262 9274
rect 12262 9222 12292 9274
rect 12316 9222 12326 9274
rect 12326 9222 12372 9274
rect 12076 9220 12132 9222
rect 12156 9220 12212 9222
rect 12236 9220 12292 9222
rect 12316 9220 12372 9222
rect 11886 8880 11942 8936
rect 12530 11464 12586 11520
rect 13082 11192 13138 11248
rect 12076 8186 12132 8188
rect 12156 8186 12212 8188
rect 12236 8186 12292 8188
rect 12316 8186 12372 8188
rect 12076 8134 12122 8186
rect 12122 8134 12132 8186
rect 12156 8134 12186 8186
rect 12186 8134 12198 8186
rect 12198 8134 12212 8186
rect 12236 8134 12250 8186
rect 12250 8134 12262 8186
rect 12262 8134 12292 8186
rect 12316 8134 12326 8186
rect 12326 8134 12372 8186
rect 12076 8132 12132 8134
rect 12156 8132 12212 8134
rect 12236 8132 12292 8134
rect 12316 8132 12372 8134
rect 12990 9696 13046 9752
rect 12806 9016 12862 9072
rect 12990 8744 13046 8800
rect 10506 3712 10562 3768
rect 10782 4140 10838 4176
rect 10782 4120 10784 4140
rect 10784 4120 10836 4140
rect 10836 4120 10838 4140
rect 10230 2488 10286 2544
rect 10230 2216 10286 2272
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9898 2202
rect 9898 2150 9908 2202
rect 9932 2150 9962 2202
rect 9962 2150 9974 2202
rect 9974 2150 9988 2202
rect 10012 2150 10026 2202
rect 10026 2150 10038 2202
rect 10038 2150 10068 2202
rect 10092 2150 10102 2202
rect 10102 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 11058 3596 11114 3632
rect 11058 3576 11060 3596
rect 11060 3576 11112 3596
rect 11112 3576 11114 3596
rect 11058 3460 11114 3496
rect 11058 3440 11060 3460
rect 11060 3440 11112 3460
rect 11112 3440 11114 3460
rect 12076 7098 12132 7100
rect 12156 7098 12212 7100
rect 12236 7098 12292 7100
rect 12316 7098 12372 7100
rect 12076 7046 12122 7098
rect 12122 7046 12132 7098
rect 12156 7046 12186 7098
rect 12186 7046 12198 7098
rect 12198 7046 12212 7098
rect 12236 7046 12250 7098
rect 12250 7046 12262 7098
rect 12262 7046 12292 7098
rect 12316 7046 12326 7098
rect 12326 7046 12372 7098
rect 12076 7044 12132 7046
rect 12156 7044 12212 7046
rect 12236 7044 12292 7046
rect 12316 7044 12372 7046
rect 12346 6160 12402 6216
rect 12076 6010 12132 6012
rect 12156 6010 12212 6012
rect 12236 6010 12292 6012
rect 12316 6010 12372 6012
rect 12076 5958 12122 6010
rect 12122 5958 12132 6010
rect 12156 5958 12186 6010
rect 12186 5958 12198 6010
rect 12198 5958 12212 6010
rect 12236 5958 12250 6010
rect 12250 5958 12262 6010
rect 12262 5958 12292 6010
rect 12316 5958 12326 6010
rect 12326 5958 12372 6010
rect 12076 5956 12132 5958
rect 12156 5956 12212 5958
rect 12236 5956 12292 5958
rect 12316 5956 12372 5958
rect 15290 16360 15346 16416
rect 15198 15952 15254 16008
rect 15934 15544 15990 15600
rect 15658 14220 15660 14240
rect 15660 14220 15712 14240
rect 15712 14220 15714 14240
rect 15658 14184 15714 14220
rect 14300 14170 14356 14172
rect 14380 14170 14436 14172
rect 14460 14170 14516 14172
rect 14540 14170 14596 14172
rect 14300 14118 14346 14170
rect 14346 14118 14356 14170
rect 14380 14118 14410 14170
rect 14410 14118 14422 14170
rect 14422 14118 14436 14170
rect 14460 14118 14474 14170
rect 14474 14118 14486 14170
rect 14486 14118 14516 14170
rect 14540 14118 14550 14170
rect 14550 14118 14596 14170
rect 14300 14116 14356 14118
rect 14380 14116 14436 14118
rect 14460 14116 14516 14118
rect 14540 14116 14596 14118
rect 15198 14068 15254 14104
rect 15198 14048 15200 14068
rect 15200 14048 15252 14068
rect 15252 14048 15254 14068
rect 13726 13776 13782 13832
rect 13450 12280 13506 12336
rect 13266 11736 13322 11792
rect 13174 7656 13230 7712
rect 13450 9444 13506 9480
rect 13450 9424 13452 9444
rect 13452 9424 13504 9444
rect 13504 9424 13506 9444
rect 13542 7928 13598 7984
rect 13358 7384 13414 7440
rect 13726 12144 13782 12200
rect 14300 13082 14356 13084
rect 14380 13082 14436 13084
rect 14460 13082 14516 13084
rect 14540 13082 14596 13084
rect 14300 13030 14346 13082
rect 14346 13030 14356 13082
rect 14380 13030 14410 13082
rect 14410 13030 14422 13082
rect 14422 13030 14436 13082
rect 14460 13030 14474 13082
rect 14474 13030 14486 13082
rect 14486 13030 14516 13082
rect 14540 13030 14550 13082
rect 14550 13030 14596 13082
rect 14300 13028 14356 13030
rect 14380 13028 14436 13030
rect 14460 13028 14516 13030
rect 14540 13028 14596 13030
rect 14300 11994 14356 11996
rect 14380 11994 14436 11996
rect 14460 11994 14516 11996
rect 14540 11994 14596 11996
rect 14300 11942 14346 11994
rect 14346 11942 14356 11994
rect 14380 11942 14410 11994
rect 14410 11942 14422 11994
rect 14422 11942 14436 11994
rect 14460 11942 14474 11994
rect 14474 11942 14486 11994
rect 14486 11942 14516 11994
rect 14540 11942 14550 11994
rect 14550 11942 14596 11994
rect 14300 11940 14356 11942
rect 14380 11940 14436 11942
rect 14460 11940 14516 11942
rect 14540 11940 14596 11942
rect 15106 12688 15162 12744
rect 14094 11192 14150 11248
rect 14300 10906 14356 10908
rect 14380 10906 14436 10908
rect 14460 10906 14516 10908
rect 14540 10906 14596 10908
rect 14300 10854 14346 10906
rect 14346 10854 14356 10906
rect 14380 10854 14410 10906
rect 14410 10854 14422 10906
rect 14422 10854 14436 10906
rect 14460 10854 14474 10906
rect 14474 10854 14486 10906
rect 14486 10854 14516 10906
rect 14540 10854 14550 10906
rect 14550 10854 14596 10906
rect 14300 10852 14356 10854
rect 14380 10852 14436 10854
rect 14460 10852 14516 10854
rect 14540 10852 14596 10854
rect 15382 11192 15438 11248
rect 15290 10920 15346 10976
rect 14300 9818 14356 9820
rect 14380 9818 14436 9820
rect 14460 9818 14516 9820
rect 14540 9818 14596 9820
rect 14300 9766 14346 9818
rect 14346 9766 14356 9818
rect 14380 9766 14410 9818
rect 14410 9766 14422 9818
rect 14422 9766 14436 9818
rect 14460 9766 14474 9818
rect 14474 9766 14486 9818
rect 14486 9766 14516 9818
rect 14540 9766 14550 9818
rect 14550 9766 14596 9818
rect 14300 9764 14356 9766
rect 14380 9764 14436 9766
rect 14460 9764 14516 9766
rect 14540 9764 14596 9766
rect 13818 8472 13874 8528
rect 13818 6740 13820 6760
rect 13820 6740 13872 6760
rect 13872 6740 13874 6760
rect 13818 6704 13874 6740
rect 13818 6432 13874 6488
rect 12076 4922 12132 4924
rect 12156 4922 12212 4924
rect 12236 4922 12292 4924
rect 12316 4922 12372 4924
rect 12076 4870 12122 4922
rect 12122 4870 12132 4922
rect 12156 4870 12186 4922
rect 12186 4870 12198 4922
rect 12198 4870 12212 4922
rect 12236 4870 12250 4922
rect 12250 4870 12262 4922
rect 12262 4870 12292 4922
rect 12316 4870 12326 4922
rect 12326 4870 12372 4922
rect 12076 4868 12132 4870
rect 12156 4868 12212 4870
rect 12236 4868 12292 4870
rect 12316 4868 12372 4870
rect 10966 2352 11022 2408
rect 12076 3834 12132 3836
rect 12156 3834 12212 3836
rect 12236 3834 12292 3836
rect 12316 3834 12372 3836
rect 12076 3782 12122 3834
rect 12122 3782 12132 3834
rect 12156 3782 12186 3834
rect 12186 3782 12198 3834
rect 12198 3782 12212 3834
rect 12236 3782 12250 3834
rect 12250 3782 12262 3834
rect 12262 3782 12292 3834
rect 12316 3782 12326 3834
rect 12326 3782 12372 3834
rect 12076 3780 12132 3782
rect 12156 3780 12212 3782
rect 12236 3780 12292 3782
rect 12316 3780 12372 3782
rect 12076 2746 12132 2748
rect 12156 2746 12212 2748
rect 12236 2746 12292 2748
rect 12316 2746 12372 2748
rect 12076 2694 12122 2746
rect 12122 2694 12132 2746
rect 12156 2694 12186 2746
rect 12186 2694 12198 2746
rect 12198 2694 12212 2746
rect 12236 2694 12250 2746
rect 12250 2694 12262 2746
rect 12262 2694 12292 2746
rect 12316 2694 12326 2746
rect 12326 2694 12372 2746
rect 12076 2692 12132 2694
rect 12156 2692 12212 2694
rect 12236 2692 12292 2694
rect 12316 2692 12372 2694
rect 13266 5208 13322 5264
rect 13726 5752 13782 5808
rect 13910 4120 13966 4176
rect 14738 8900 14794 8936
rect 14738 8880 14740 8900
rect 14740 8880 14792 8900
rect 14792 8880 14794 8900
rect 14300 8730 14356 8732
rect 14380 8730 14436 8732
rect 14460 8730 14516 8732
rect 14540 8730 14596 8732
rect 14300 8678 14346 8730
rect 14346 8678 14356 8730
rect 14380 8678 14410 8730
rect 14410 8678 14422 8730
rect 14422 8678 14436 8730
rect 14460 8678 14474 8730
rect 14474 8678 14486 8730
rect 14486 8678 14516 8730
rect 14540 8678 14550 8730
rect 14550 8678 14596 8730
rect 14300 8676 14356 8678
rect 14380 8676 14436 8678
rect 14460 8676 14516 8678
rect 14540 8676 14596 8678
rect 15014 8608 15070 8664
rect 14300 7642 14356 7644
rect 14380 7642 14436 7644
rect 14460 7642 14516 7644
rect 14540 7642 14596 7644
rect 14300 7590 14346 7642
rect 14346 7590 14356 7642
rect 14380 7590 14410 7642
rect 14410 7590 14422 7642
rect 14422 7590 14436 7642
rect 14460 7590 14474 7642
rect 14474 7590 14486 7642
rect 14486 7590 14516 7642
rect 14540 7590 14550 7642
rect 14550 7590 14596 7642
rect 14300 7588 14356 7590
rect 14380 7588 14436 7590
rect 14460 7588 14516 7590
rect 14540 7588 14596 7590
rect 14300 6554 14356 6556
rect 14380 6554 14436 6556
rect 14460 6554 14516 6556
rect 14540 6554 14596 6556
rect 14300 6502 14346 6554
rect 14346 6502 14356 6554
rect 14380 6502 14410 6554
rect 14410 6502 14422 6554
rect 14422 6502 14436 6554
rect 14460 6502 14474 6554
rect 14474 6502 14486 6554
rect 14486 6502 14516 6554
rect 14540 6502 14550 6554
rect 14550 6502 14596 6554
rect 14300 6500 14356 6502
rect 14380 6500 14436 6502
rect 14460 6500 14516 6502
rect 14540 6500 14596 6502
rect 12990 2524 12992 2544
rect 12992 2524 13044 2544
rect 13044 2524 13046 2544
rect 12990 2488 13046 2524
rect 14646 5772 14702 5808
rect 14646 5752 14648 5772
rect 14648 5752 14700 5772
rect 14700 5752 14702 5772
rect 14300 5466 14356 5468
rect 14380 5466 14436 5468
rect 14460 5466 14516 5468
rect 14540 5466 14596 5468
rect 14300 5414 14346 5466
rect 14346 5414 14356 5466
rect 14380 5414 14410 5466
rect 14410 5414 14422 5466
rect 14422 5414 14436 5466
rect 14460 5414 14474 5466
rect 14474 5414 14486 5466
rect 14486 5414 14516 5466
rect 14540 5414 14550 5466
rect 14550 5414 14596 5466
rect 14300 5412 14356 5414
rect 14380 5412 14436 5414
rect 14460 5412 14516 5414
rect 14540 5412 14596 5414
rect 14370 5072 14426 5128
rect 14300 4378 14356 4380
rect 14380 4378 14436 4380
rect 14460 4378 14516 4380
rect 14540 4378 14596 4380
rect 14300 4326 14346 4378
rect 14346 4326 14356 4378
rect 14380 4326 14410 4378
rect 14410 4326 14422 4378
rect 14422 4326 14436 4378
rect 14460 4326 14474 4378
rect 14474 4326 14486 4378
rect 14486 4326 14516 4378
rect 14540 4326 14550 4378
rect 14550 4326 14596 4378
rect 14300 4324 14356 4326
rect 14380 4324 14436 4326
rect 14460 4324 14516 4326
rect 14540 4324 14596 4326
rect 14300 3290 14356 3292
rect 14380 3290 14436 3292
rect 14460 3290 14516 3292
rect 14540 3290 14596 3292
rect 14300 3238 14346 3290
rect 14346 3238 14356 3290
rect 14380 3238 14410 3290
rect 14410 3238 14422 3290
rect 14422 3238 14436 3290
rect 14460 3238 14474 3290
rect 14474 3238 14486 3290
rect 14486 3238 14516 3290
rect 14540 3238 14550 3290
rect 14550 3238 14596 3290
rect 14300 3236 14356 3238
rect 14380 3236 14436 3238
rect 14460 3236 14516 3238
rect 14540 3236 14596 3238
rect 16524 14714 16580 14716
rect 16604 14714 16660 14716
rect 16684 14714 16740 14716
rect 16764 14714 16820 14716
rect 16524 14662 16570 14714
rect 16570 14662 16580 14714
rect 16604 14662 16634 14714
rect 16634 14662 16646 14714
rect 16646 14662 16660 14714
rect 16684 14662 16698 14714
rect 16698 14662 16710 14714
rect 16710 14662 16740 14714
rect 16764 14662 16774 14714
rect 16774 14662 16820 14714
rect 16524 14660 16580 14662
rect 16604 14660 16660 14662
rect 16684 14660 16740 14662
rect 16764 14660 16820 14662
rect 16524 13626 16580 13628
rect 16604 13626 16660 13628
rect 16684 13626 16740 13628
rect 16764 13626 16820 13628
rect 16524 13574 16570 13626
rect 16570 13574 16580 13626
rect 16604 13574 16634 13626
rect 16634 13574 16646 13626
rect 16646 13574 16660 13626
rect 16684 13574 16698 13626
rect 16698 13574 16710 13626
rect 16710 13574 16740 13626
rect 16764 13574 16774 13626
rect 16774 13574 16820 13626
rect 16524 13572 16580 13574
rect 16604 13572 16660 13574
rect 16684 13572 16740 13574
rect 16764 13572 16820 13574
rect 17038 13912 17094 13968
rect 18050 13268 18052 13288
rect 18052 13268 18104 13288
rect 18104 13268 18106 13288
rect 18050 13232 18106 13268
rect 16118 12960 16174 13016
rect 15934 12316 15936 12336
rect 15936 12316 15988 12336
rect 15988 12316 15990 12336
rect 15934 12280 15990 12316
rect 16524 12538 16580 12540
rect 16604 12538 16660 12540
rect 16684 12538 16740 12540
rect 16764 12538 16820 12540
rect 16524 12486 16570 12538
rect 16570 12486 16580 12538
rect 16604 12486 16634 12538
rect 16634 12486 16646 12538
rect 16646 12486 16660 12538
rect 16684 12486 16698 12538
rect 16698 12486 16710 12538
rect 16710 12486 16740 12538
rect 16764 12486 16774 12538
rect 16774 12486 16820 12538
rect 16524 12484 16580 12486
rect 16604 12484 16660 12486
rect 16684 12484 16740 12486
rect 16764 12484 16820 12486
rect 15382 5752 15438 5808
rect 15106 5616 15162 5672
rect 15198 5072 15254 5128
rect 15290 4120 15346 4176
rect 14300 2202 14356 2204
rect 14380 2202 14436 2204
rect 14460 2202 14516 2204
rect 14540 2202 14596 2204
rect 14300 2150 14346 2202
rect 14346 2150 14356 2202
rect 14380 2150 14410 2202
rect 14410 2150 14422 2202
rect 14422 2150 14436 2202
rect 14460 2150 14474 2202
rect 14474 2150 14486 2202
rect 14486 2150 14516 2202
rect 14540 2150 14550 2202
rect 14550 2150 14596 2202
rect 14300 2148 14356 2150
rect 14380 2148 14436 2150
rect 14460 2148 14516 2150
rect 14540 2148 14596 2150
rect 15474 2624 15530 2680
rect 15934 9968 15990 10024
rect 15934 7248 15990 7304
rect 16486 11600 16542 11656
rect 16210 11464 16266 11520
rect 16524 11450 16580 11452
rect 16604 11450 16660 11452
rect 16684 11450 16740 11452
rect 16764 11450 16820 11452
rect 16524 11398 16570 11450
rect 16570 11398 16580 11450
rect 16604 11398 16634 11450
rect 16634 11398 16646 11450
rect 16646 11398 16660 11450
rect 16684 11398 16698 11450
rect 16698 11398 16710 11450
rect 16710 11398 16740 11450
rect 16764 11398 16774 11450
rect 16774 11398 16820 11450
rect 16524 11396 16580 11398
rect 16604 11396 16660 11398
rect 16684 11396 16740 11398
rect 16764 11396 16820 11398
rect 16118 10104 16174 10160
rect 16854 10956 16856 10976
rect 16856 10956 16908 10976
rect 16908 10956 16910 10976
rect 16854 10920 16910 10956
rect 16524 10362 16580 10364
rect 16604 10362 16660 10364
rect 16684 10362 16740 10364
rect 16764 10362 16820 10364
rect 16524 10310 16570 10362
rect 16570 10310 16580 10362
rect 16604 10310 16634 10362
rect 16634 10310 16646 10362
rect 16646 10310 16660 10362
rect 16684 10310 16698 10362
rect 16698 10310 16710 10362
rect 16710 10310 16740 10362
rect 16764 10310 16774 10362
rect 16774 10310 16820 10362
rect 16524 10308 16580 10310
rect 16604 10308 16660 10310
rect 16684 10308 16740 10310
rect 16764 10308 16820 10310
rect 16524 9274 16580 9276
rect 16604 9274 16660 9276
rect 16684 9274 16740 9276
rect 16764 9274 16820 9276
rect 16524 9222 16570 9274
rect 16570 9222 16580 9274
rect 16604 9222 16634 9274
rect 16634 9222 16646 9274
rect 16646 9222 16660 9274
rect 16684 9222 16698 9274
rect 16698 9222 16710 9274
rect 16710 9222 16740 9274
rect 16764 9222 16774 9274
rect 16774 9222 16820 9274
rect 16524 9220 16580 9222
rect 16604 9220 16660 9222
rect 16684 9220 16740 9222
rect 16764 9220 16820 9222
rect 16210 8744 16266 8800
rect 15934 6316 15990 6352
rect 15934 6296 15936 6316
rect 15936 6296 15988 6316
rect 15988 6296 15990 6316
rect 16486 8628 16542 8664
rect 16486 8608 16488 8628
rect 16488 8608 16540 8628
rect 16540 8608 16542 8628
rect 16524 8186 16580 8188
rect 16604 8186 16660 8188
rect 16684 8186 16740 8188
rect 16764 8186 16820 8188
rect 16524 8134 16570 8186
rect 16570 8134 16580 8186
rect 16604 8134 16634 8186
rect 16634 8134 16646 8186
rect 16646 8134 16660 8186
rect 16684 8134 16698 8186
rect 16698 8134 16710 8186
rect 16710 8134 16740 8186
rect 16764 8134 16774 8186
rect 16774 8134 16820 8186
rect 16524 8132 16580 8134
rect 16604 8132 16660 8134
rect 16684 8132 16740 8134
rect 16764 8132 16820 8134
rect 17038 8336 17094 8392
rect 16946 7792 17002 7848
rect 16524 7098 16580 7100
rect 16604 7098 16660 7100
rect 16684 7098 16740 7100
rect 16764 7098 16820 7100
rect 16524 7046 16570 7098
rect 16570 7046 16580 7098
rect 16604 7046 16634 7098
rect 16634 7046 16646 7098
rect 16646 7046 16660 7098
rect 16684 7046 16698 7098
rect 16698 7046 16710 7098
rect 16710 7046 16740 7098
rect 16764 7046 16774 7098
rect 16774 7046 16820 7098
rect 16524 7044 16580 7046
rect 16604 7044 16660 7046
rect 16684 7044 16740 7046
rect 16764 7044 16820 7046
rect 15934 4020 15936 4040
rect 15936 4020 15988 4040
rect 15988 4020 15990 4040
rect 15934 3984 15990 4020
rect 16302 4820 16358 4856
rect 16302 4800 16304 4820
rect 16304 4800 16356 4820
rect 16356 4800 16358 4820
rect 16524 6010 16580 6012
rect 16604 6010 16660 6012
rect 16684 6010 16740 6012
rect 16764 6010 16820 6012
rect 16524 5958 16570 6010
rect 16570 5958 16580 6010
rect 16604 5958 16634 6010
rect 16634 5958 16646 6010
rect 16646 5958 16660 6010
rect 16684 5958 16698 6010
rect 16698 5958 16710 6010
rect 16710 5958 16740 6010
rect 16764 5958 16774 6010
rect 16774 5958 16820 6010
rect 16524 5956 16580 5958
rect 16604 5956 16660 5958
rect 16684 5956 16740 5958
rect 16764 5956 16820 5958
rect 16486 5480 16542 5536
rect 16854 5364 16910 5400
rect 16854 5344 16856 5364
rect 16856 5344 16908 5364
rect 16908 5344 16910 5364
rect 16524 4922 16580 4924
rect 16604 4922 16660 4924
rect 16684 4922 16740 4924
rect 16764 4922 16820 4924
rect 16524 4870 16570 4922
rect 16570 4870 16580 4922
rect 16604 4870 16634 4922
rect 16634 4870 16646 4922
rect 16646 4870 16660 4922
rect 16684 4870 16698 4922
rect 16698 4870 16710 4922
rect 16710 4870 16740 4922
rect 16764 4870 16774 4922
rect 16774 4870 16820 4922
rect 16524 4868 16580 4870
rect 16604 4868 16660 4870
rect 16684 4868 16740 4870
rect 16764 4868 16820 4870
rect 18418 13368 18474 13424
rect 17314 10512 17370 10568
rect 17682 10376 17738 10432
rect 17958 10648 18014 10704
rect 17774 9560 17830 9616
rect 17314 7928 17370 7984
rect 17314 7656 17370 7712
rect 16394 4664 16450 4720
rect 17038 4256 17094 4312
rect 16524 3834 16580 3836
rect 16604 3834 16660 3836
rect 16684 3834 16740 3836
rect 16764 3834 16820 3836
rect 16524 3782 16570 3834
rect 16570 3782 16580 3834
rect 16604 3782 16634 3834
rect 16634 3782 16646 3834
rect 16646 3782 16660 3834
rect 16684 3782 16698 3834
rect 16698 3782 16710 3834
rect 16710 3782 16740 3834
rect 16764 3782 16774 3834
rect 16774 3782 16820 3834
rect 16524 3780 16580 3782
rect 16604 3780 16660 3782
rect 16684 3780 16740 3782
rect 16764 3780 16820 3782
rect 16026 3596 16082 3632
rect 16026 3576 16028 3596
rect 16028 3576 16080 3596
rect 16080 3576 16082 3596
rect 16946 3460 17002 3496
rect 16946 3440 16948 3460
rect 16948 3440 17000 3460
rect 17000 3440 17002 3460
rect 17038 3168 17094 3224
rect 16854 3032 16910 3088
rect 16762 2916 16818 2952
rect 16762 2896 16764 2916
rect 16764 2896 16816 2916
rect 16816 2896 16818 2916
rect 16946 2760 17002 2816
rect 16524 2746 16580 2748
rect 16604 2746 16660 2748
rect 16684 2746 16740 2748
rect 16764 2746 16820 2748
rect 16524 2694 16570 2746
rect 16570 2694 16580 2746
rect 16604 2694 16634 2746
rect 16634 2694 16646 2746
rect 16646 2694 16660 2746
rect 16684 2694 16698 2746
rect 16698 2694 16710 2746
rect 16710 2694 16740 2746
rect 16764 2694 16774 2746
rect 16774 2694 16820 2746
rect 16524 2692 16580 2694
rect 16604 2692 16660 2694
rect 16684 2692 16740 2694
rect 16764 2692 16820 2694
rect 17314 6160 17370 6216
rect 17314 1808 17370 1864
rect 17866 9152 17922 9208
rect 17774 7792 17830 7848
rect 18142 8200 18198 8256
rect 17866 6976 17922 7032
rect 17682 6604 17684 6624
rect 17684 6604 17736 6624
rect 17736 6604 17738 6624
rect 17682 6568 17738 6604
rect 18050 6704 18106 6760
rect 18050 6180 18106 6216
rect 18050 6160 18052 6180
rect 18052 6160 18104 6180
rect 18104 6160 18106 6180
rect 18050 5208 18106 5264
rect 17866 3984 17922 4040
rect 18418 7384 18474 7440
rect 18418 7284 18420 7304
rect 18420 7284 18472 7304
rect 18472 7284 18474 7304
rect 18418 7248 18474 7284
rect 18418 5616 18474 5672
rect 18326 4800 18382 4856
rect 18326 4664 18382 4720
rect 18050 4392 18106 4448
rect 18050 3168 18106 3224
rect 17958 3032 18014 3088
rect 18050 2624 18106 2680
rect 17682 1400 17738 1456
rect 17866 992 17922 1048
rect 18418 3612 18420 3632
rect 18420 3612 18472 3632
rect 18472 3612 18474 3632
rect 18418 3576 18474 3612
rect 18234 2252 18236 2272
rect 18236 2252 18288 2272
rect 18288 2252 18290 2272
rect 18234 2216 18290 2252
rect 18602 9988 18658 10024
rect 18602 9968 18604 9988
rect 18604 9968 18656 9988
rect 18656 9968 18658 9988
rect 18142 584 18198 640
rect 18878 176 18934 232
<< metal3 >>
rect 0 16826 800 16856
rect 3693 16826 3759 16829
rect 0 16824 3759 16826
rect 0 16768 3698 16824
rect 3754 16768 3759 16824
rect 0 16766 3759 16768
rect 0 16736 800 16766
rect 3693 16763 3759 16766
rect 18045 16826 18111 16829
rect 19200 16826 20000 16856
rect 18045 16824 20000 16826
rect 18045 16768 18050 16824
rect 18106 16768 20000 16824
rect 18045 16766 20000 16768
rect 18045 16763 18111 16766
rect 19200 16736 20000 16766
rect 0 16418 800 16448
rect 3509 16418 3575 16421
rect 0 16416 3575 16418
rect 0 16360 3514 16416
rect 3570 16360 3575 16416
rect 0 16358 3575 16360
rect 0 16328 800 16358
rect 3509 16355 3575 16358
rect 15285 16418 15351 16421
rect 19200 16418 20000 16448
rect 15285 16416 20000 16418
rect 15285 16360 15290 16416
rect 15346 16360 20000 16416
rect 15285 16358 20000 16360
rect 15285 16355 15351 16358
rect 19200 16328 20000 16358
rect 0 16010 800 16040
rect 4061 16010 4127 16013
rect 0 16008 4127 16010
rect 0 15952 4066 16008
rect 4122 15952 4127 16008
rect 0 15950 4127 15952
rect 0 15920 800 15950
rect 4061 15947 4127 15950
rect 15193 16010 15259 16013
rect 19200 16010 20000 16040
rect 15193 16008 20000 16010
rect 15193 15952 15198 16008
rect 15254 15952 20000 16008
rect 15193 15950 20000 15952
rect 15193 15947 15259 15950
rect 19200 15920 20000 15950
rect 0 15602 800 15632
rect 3969 15602 4035 15605
rect 0 15600 4035 15602
rect 0 15544 3974 15600
rect 4030 15544 4035 15600
rect 0 15542 4035 15544
rect 0 15512 800 15542
rect 3969 15539 4035 15542
rect 15929 15602 15995 15605
rect 19200 15602 20000 15632
rect 15929 15600 20000 15602
rect 15929 15544 15934 15600
rect 15990 15544 20000 15600
rect 15929 15542 20000 15544
rect 15929 15539 15995 15542
rect 19200 15512 20000 15542
rect 0 15194 800 15224
rect 1577 15194 1643 15197
rect 0 15192 1643 15194
rect 0 15136 1582 15192
rect 1638 15136 1643 15192
rect 0 15134 1643 15136
rect 0 15104 800 15134
rect 1577 15131 1643 15134
rect 15510 15132 15516 15196
rect 15580 15194 15586 15196
rect 19200 15194 20000 15224
rect 15580 15134 20000 15194
rect 15580 15132 15586 15134
rect 19200 15104 20000 15134
rect 0 14786 800 14816
rect 2773 14786 2839 14789
rect 0 14784 2839 14786
rect 0 14728 2778 14784
rect 2834 14728 2839 14784
rect 0 14726 2839 14728
rect 0 14696 800 14726
rect 2773 14723 2839 14726
rect 17166 14724 17172 14788
rect 17236 14786 17242 14788
rect 19200 14786 20000 14816
rect 17236 14726 20000 14786
rect 17236 14724 17242 14726
rect 3168 14720 3488 14721
rect 3168 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3488 14720
rect 3168 14655 3488 14656
rect 7616 14720 7936 14721
rect 7616 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7936 14720
rect 7616 14655 7936 14656
rect 12064 14720 12384 14721
rect 12064 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12384 14720
rect 12064 14655 12384 14656
rect 16512 14720 16832 14721
rect 16512 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16832 14720
rect 19200 14696 20000 14726
rect 16512 14655 16832 14656
rect 0 14378 800 14408
rect 4061 14378 4127 14381
rect 0 14376 4127 14378
rect 0 14320 4066 14376
rect 4122 14320 4127 14376
rect 0 14318 4127 14320
rect 0 14288 800 14318
rect 4061 14315 4127 14318
rect 15653 14242 15719 14245
rect 19200 14242 20000 14272
rect 15653 14240 20000 14242
rect 15653 14184 15658 14240
rect 15714 14184 20000 14240
rect 15653 14182 20000 14184
rect 15653 14179 15719 14182
rect 5392 14176 5712 14177
rect 5392 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5712 14176
rect 5392 14111 5712 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 14288 14176 14608 14177
rect 14288 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14608 14176
rect 19200 14152 20000 14182
rect 14288 14111 14608 14112
rect 15193 14106 15259 14109
rect 17166 14106 17172 14108
rect 15193 14104 17172 14106
rect 15193 14048 15198 14104
rect 15254 14048 17172 14104
rect 15193 14046 17172 14048
rect 15193 14043 15259 14046
rect 17166 14044 17172 14046
rect 17236 14044 17242 14108
rect 0 13970 800 14000
rect 3785 13970 3851 13973
rect 17033 13972 17099 13973
rect 16982 13970 16988 13972
rect 0 13968 3851 13970
rect 0 13912 3790 13968
rect 3846 13912 3851 13968
rect 0 13910 3851 13912
rect 16942 13910 16988 13970
rect 17052 13968 17099 13972
rect 17094 13912 17099 13968
rect 0 13880 800 13910
rect 3785 13907 3851 13910
rect 16982 13908 16988 13910
rect 17052 13908 17099 13912
rect 17033 13907 17099 13908
rect 13721 13834 13787 13837
rect 19200 13834 20000 13864
rect 13721 13832 20000 13834
rect 13721 13776 13726 13832
rect 13782 13776 20000 13832
rect 13721 13774 20000 13776
rect 13721 13771 13787 13774
rect 19200 13744 20000 13774
rect 3168 13632 3488 13633
rect 0 13562 800 13592
rect 3168 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3488 13632
rect 3168 13567 3488 13568
rect 7616 13632 7936 13633
rect 7616 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7936 13632
rect 7616 13567 7936 13568
rect 12064 13632 12384 13633
rect 12064 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12384 13632
rect 12064 13567 12384 13568
rect 16512 13632 16832 13633
rect 16512 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16832 13632
rect 16512 13567 16832 13568
rect 0 13502 2790 13562
rect 0 13472 800 13502
rect 2730 13426 2790 13502
rect 4061 13426 4127 13429
rect 2730 13424 4127 13426
rect 2730 13368 4066 13424
rect 4122 13368 4127 13424
rect 2730 13366 4127 13368
rect 4061 13363 4127 13366
rect 18413 13426 18479 13429
rect 19200 13426 20000 13456
rect 18413 13424 20000 13426
rect 18413 13368 18418 13424
rect 18474 13368 20000 13424
rect 18413 13366 20000 13368
rect 18413 13363 18479 13366
rect 19200 13336 20000 13366
rect 3601 13290 3667 13293
rect 18045 13290 18111 13293
rect 3601 13288 18111 13290
rect 3601 13232 3606 13288
rect 3662 13232 18050 13288
rect 18106 13232 18111 13288
rect 3601 13230 18111 13232
rect 3601 13227 3667 13230
rect 18045 13227 18111 13230
rect 0 13154 800 13184
rect 4521 13154 4587 13157
rect 0 13152 4587 13154
rect 0 13096 4526 13152
rect 4582 13096 4587 13152
rect 0 13094 4587 13096
rect 0 13064 800 13094
rect 4521 13091 4587 13094
rect 5392 13088 5712 13089
rect 5392 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5712 13088
rect 5392 13023 5712 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 14288 13088 14608 13089
rect 14288 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14608 13088
rect 14288 13023 14608 13024
rect 16113 13018 16179 13021
rect 19200 13018 20000 13048
rect 16113 13016 20000 13018
rect 16113 12960 16118 13016
rect 16174 12960 20000 13016
rect 16113 12958 20000 12960
rect 16113 12955 16179 12958
rect 19200 12928 20000 12958
rect 0 12746 800 12776
rect 8518 12746 8524 12748
rect 0 12686 8524 12746
rect 0 12656 800 12686
rect 8518 12684 8524 12686
rect 8588 12684 8594 12748
rect 15101 12746 15167 12749
rect 15101 12744 17970 12746
rect 15101 12688 15106 12744
rect 15162 12688 17970 12744
rect 15101 12686 17970 12688
rect 15101 12683 15167 12686
rect 1894 12548 1900 12612
rect 1964 12610 1970 12612
rect 2129 12610 2195 12613
rect 1964 12608 2195 12610
rect 1964 12552 2134 12608
rect 2190 12552 2195 12608
rect 1964 12550 2195 12552
rect 17910 12610 17970 12686
rect 19200 12610 20000 12640
rect 17910 12550 20000 12610
rect 1964 12548 1970 12550
rect 2129 12547 2195 12550
rect 3168 12544 3488 12545
rect 3168 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3488 12544
rect 3168 12479 3488 12480
rect 7616 12544 7936 12545
rect 7616 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7936 12544
rect 7616 12479 7936 12480
rect 12064 12544 12384 12545
rect 12064 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12384 12544
rect 12064 12479 12384 12480
rect 16512 12544 16832 12545
rect 16512 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16832 12544
rect 19200 12520 20000 12550
rect 16512 12479 16832 12480
rect 1577 12474 1643 12477
rect 2446 12474 2452 12476
rect 1577 12472 2452 12474
rect 1577 12416 1582 12472
rect 1638 12416 2452 12472
rect 1577 12414 2452 12416
rect 1577 12411 1643 12414
rect 2446 12412 2452 12414
rect 2516 12412 2522 12476
rect 0 12338 800 12368
rect 11145 12338 11211 12341
rect 0 12336 11211 12338
rect 0 12280 11150 12336
rect 11206 12280 11211 12336
rect 0 12278 11211 12280
rect 0 12248 800 12278
rect 11145 12275 11211 12278
rect 13445 12338 13511 12341
rect 15929 12338 15995 12341
rect 13445 12336 15995 12338
rect 13445 12280 13450 12336
rect 13506 12280 15934 12336
rect 15990 12280 15995 12336
rect 13445 12278 15995 12280
rect 13445 12275 13511 12278
rect 15929 12275 15995 12278
rect 9397 12202 9463 12205
rect 13721 12202 13787 12205
rect 9397 12200 13787 12202
rect 9397 12144 9402 12200
rect 9458 12144 13726 12200
rect 13782 12144 13787 12200
rect 9397 12142 13787 12144
rect 9397 12139 9463 12142
rect 13721 12139 13787 12142
rect 16062 12140 16068 12204
rect 16132 12202 16138 12204
rect 19200 12202 20000 12232
rect 16132 12142 20000 12202
rect 16132 12140 16138 12142
rect 19200 12112 20000 12142
rect 5392 12000 5712 12001
rect 0 11930 800 11960
rect 5392 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5712 12000
rect 5392 11935 5712 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 14288 12000 14608 12001
rect 14288 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14608 12000
rect 14288 11935 14608 11936
rect 3877 11930 3943 11933
rect 0 11928 3943 11930
rect 0 11872 3882 11928
rect 3938 11872 3943 11928
rect 0 11870 3943 11872
rect 0 11840 800 11870
rect 3877 11867 3943 11870
rect 4061 11932 4127 11933
rect 4061 11928 4108 11932
rect 4172 11930 4178 11932
rect 10501 11930 10567 11933
rect 11881 11930 11947 11933
rect 4061 11872 4066 11928
rect 4061 11868 4108 11872
rect 4172 11870 4218 11930
rect 10501 11928 11947 11930
rect 10501 11872 10506 11928
rect 10562 11872 11886 11928
rect 11942 11872 11947 11928
rect 10501 11870 11947 11872
rect 4172 11868 4178 11870
rect 4061 11867 4127 11868
rect 10501 11867 10567 11870
rect 11881 11867 11947 11870
rect 12433 11930 12499 11933
rect 12433 11928 13554 11930
rect 12433 11872 12438 11928
rect 12494 11872 13554 11928
rect 12433 11870 13554 11872
rect 12433 11867 12499 11870
rect 3509 11794 3575 11797
rect 13261 11794 13327 11797
rect 3509 11792 13327 11794
rect 3509 11736 3514 11792
rect 3570 11736 13266 11792
rect 13322 11736 13327 11792
rect 3509 11734 13327 11736
rect 13494 11794 13554 11870
rect 16246 11794 16252 11796
rect 13494 11734 16252 11794
rect 3509 11731 3575 11734
rect 13261 11731 13327 11734
rect 16246 11732 16252 11734
rect 16316 11794 16322 11796
rect 19200 11794 20000 11824
rect 16316 11734 20000 11794
rect 16316 11732 16322 11734
rect 19200 11704 20000 11734
rect 6913 11658 6979 11661
rect 8845 11658 8911 11661
rect 16481 11658 16547 11661
rect 6913 11656 8218 11658
rect 6913 11600 6918 11656
rect 6974 11600 8218 11656
rect 6913 11598 8218 11600
rect 6913 11595 6979 11598
rect 8158 11522 8218 11598
rect 8845 11656 16547 11658
rect 8845 11600 8850 11656
rect 8906 11600 16486 11656
rect 16542 11600 16547 11656
rect 8845 11598 16547 11600
rect 8845 11595 8911 11598
rect 16481 11595 16547 11598
rect 10501 11522 10567 11525
rect 8158 11520 10567 11522
rect 8158 11464 10506 11520
rect 10562 11464 10567 11520
rect 8158 11462 10567 11464
rect 10501 11459 10567 11462
rect 12525 11522 12591 11525
rect 16205 11522 16271 11525
rect 12525 11520 16271 11522
rect 12525 11464 12530 11520
rect 12586 11464 16210 11520
rect 16266 11464 16271 11520
rect 12525 11462 16271 11464
rect 12525 11459 12591 11462
rect 16205 11459 16271 11462
rect 3168 11456 3488 11457
rect 0 11386 800 11416
rect 3168 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3488 11456
rect 3168 11391 3488 11392
rect 7616 11456 7936 11457
rect 7616 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7936 11456
rect 7616 11391 7936 11392
rect 12064 11456 12384 11457
rect 12064 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12384 11456
rect 12064 11391 12384 11392
rect 16512 11456 16832 11457
rect 16512 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16832 11456
rect 16512 11391 16832 11392
rect 2313 11386 2379 11389
rect 0 11384 2379 11386
rect 0 11328 2318 11384
rect 2374 11328 2379 11384
rect 0 11326 2379 11328
rect 0 11296 800 11326
rect 2313 11323 2379 11326
rect 9949 11386 10015 11389
rect 10777 11386 10843 11389
rect 11881 11386 11947 11389
rect 9949 11384 11947 11386
rect 9949 11328 9954 11384
rect 10010 11328 10782 11384
rect 10838 11328 11886 11384
rect 11942 11328 11947 11384
rect 9949 11326 11947 11328
rect 9949 11323 10015 11326
rect 10777 11323 10843 11326
rect 11881 11323 11947 11326
rect 4153 11250 4219 11253
rect 13077 11250 13143 11253
rect 4153 11248 13143 11250
rect 4153 11192 4158 11248
rect 4214 11192 13082 11248
rect 13138 11192 13143 11248
rect 4153 11190 13143 11192
rect 4153 11187 4219 11190
rect 13077 11187 13143 11190
rect 14089 11250 14155 11253
rect 15142 11250 15148 11252
rect 14089 11248 15148 11250
rect 14089 11192 14094 11248
rect 14150 11192 15148 11248
rect 14089 11190 15148 11192
rect 14089 11187 14155 11190
rect 15142 11188 15148 11190
rect 15212 11188 15218 11252
rect 15377 11250 15443 11253
rect 19200 11250 20000 11280
rect 15377 11248 20000 11250
rect 15377 11192 15382 11248
rect 15438 11192 20000 11248
rect 15377 11190 20000 11192
rect 15377 11187 15443 11190
rect 19200 11160 20000 11190
rect 6913 11114 6979 11117
rect 4110 11112 6979 11114
rect 4110 11056 6918 11112
rect 6974 11056 6979 11112
rect 4110 11054 6979 11056
rect 0 10978 800 11008
rect 3785 10978 3851 10981
rect 0 10976 3851 10978
rect 0 10920 3790 10976
rect 3846 10920 3851 10976
rect 0 10918 3851 10920
rect 0 10888 800 10918
rect 3785 10915 3851 10918
rect 1761 10844 1827 10845
rect 1710 10842 1716 10844
rect 1670 10782 1716 10842
rect 1780 10840 1827 10844
rect 1822 10784 1827 10840
rect 1710 10780 1716 10782
rect 1780 10780 1827 10784
rect 1761 10779 1827 10780
rect 0 10570 800 10600
rect 4110 10570 4170 11054
rect 6913 11051 6979 11054
rect 12249 11114 12315 11117
rect 16062 11114 16068 11116
rect 12249 11112 16068 11114
rect 12249 11056 12254 11112
rect 12310 11056 16068 11112
rect 12249 11054 16068 11056
rect 12249 11051 12315 11054
rect 16062 11052 16068 11054
rect 16132 11052 16138 11116
rect 15285 10978 15351 10981
rect 16849 10978 16915 10981
rect 15285 10976 16915 10978
rect 15285 10920 15290 10976
rect 15346 10920 16854 10976
rect 16910 10920 16915 10976
rect 15285 10918 16915 10920
rect 15285 10915 15351 10918
rect 16849 10915 16915 10918
rect 5392 10912 5712 10913
rect 5392 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5712 10912
rect 5392 10847 5712 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 14288 10912 14608 10913
rect 14288 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14608 10912
rect 14288 10847 14608 10848
rect 19200 10842 20000 10872
rect 18094 10782 20000 10842
rect 4337 10706 4403 10709
rect 4521 10706 4587 10709
rect 17953 10706 18019 10709
rect 4337 10704 18019 10706
rect 4337 10648 4342 10704
rect 4398 10648 4526 10704
rect 4582 10648 17958 10704
rect 18014 10648 18019 10704
rect 4337 10646 18019 10648
rect 4337 10643 4403 10646
rect 4521 10643 4587 10646
rect 17953 10643 18019 10646
rect 0 10510 4170 10570
rect 6453 10570 6519 10573
rect 17309 10570 17375 10573
rect 18094 10570 18154 10782
rect 19200 10752 20000 10782
rect 6453 10568 18154 10570
rect 6453 10512 6458 10568
rect 6514 10512 17314 10568
rect 17370 10512 18154 10568
rect 6453 10510 18154 10512
rect 0 10480 800 10510
rect 6453 10507 6519 10510
rect 17309 10507 17375 10510
rect 17677 10434 17743 10437
rect 19200 10434 20000 10464
rect 17677 10432 20000 10434
rect 17677 10376 17682 10432
rect 17738 10376 20000 10432
rect 17677 10374 20000 10376
rect 17677 10371 17743 10374
rect 3168 10368 3488 10369
rect 3168 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3488 10368
rect 3168 10303 3488 10304
rect 7616 10368 7936 10369
rect 7616 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7936 10368
rect 7616 10303 7936 10304
rect 12064 10368 12384 10369
rect 12064 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12384 10368
rect 12064 10303 12384 10304
rect 16512 10368 16832 10369
rect 16512 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16832 10368
rect 19200 10344 20000 10374
rect 16512 10303 16832 10304
rect 0 10162 800 10192
rect 4061 10162 4127 10165
rect 0 10160 4127 10162
rect 0 10104 4066 10160
rect 4122 10104 4127 10160
rect 0 10102 4127 10104
rect 0 10072 800 10102
rect 4061 10099 4127 10102
rect 7557 10162 7623 10165
rect 8293 10162 8359 10165
rect 7557 10160 8359 10162
rect 7557 10104 7562 10160
rect 7618 10104 8298 10160
rect 8354 10104 8359 10160
rect 7557 10102 8359 10104
rect 7557 10099 7623 10102
rect 8293 10099 8359 10102
rect 8518 10100 8524 10164
rect 8588 10162 8594 10164
rect 8845 10162 8911 10165
rect 8588 10160 8911 10162
rect 8588 10104 8850 10160
rect 8906 10104 8911 10160
rect 8588 10102 8911 10104
rect 8588 10100 8594 10102
rect 8845 10099 8911 10102
rect 10501 10162 10567 10165
rect 16113 10162 16179 10165
rect 10501 10160 16179 10162
rect 10501 10104 10506 10160
rect 10562 10104 16118 10160
rect 16174 10104 16179 10160
rect 10501 10102 16179 10104
rect 10501 10099 10567 10102
rect 16113 10099 16179 10102
rect 5993 10026 6059 10029
rect 6637 10026 6703 10029
rect 10225 10026 10291 10029
rect 5993 10024 10291 10026
rect 5993 9968 5998 10024
rect 6054 9968 6642 10024
rect 6698 9968 10230 10024
rect 10286 9968 10291 10024
rect 5993 9966 10291 9968
rect 5993 9963 6059 9966
rect 6637 9963 6703 9966
rect 10225 9963 10291 9966
rect 15929 10026 15995 10029
rect 18597 10026 18663 10029
rect 19200 10026 20000 10056
rect 15929 10024 20000 10026
rect 15929 9968 15934 10024
rect 15990 9968 18602 10024
rect 18658 9968 20000 10024
rect 15929 9966 20000 9968
rect 15929 9963 15995 9966
rect 18597 9963 18663 9966
rect 19200 9936 20000 9966
rect 5392 9824 5712 9825
rect 0 9754 800 9784
rect 5392 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5712 9824
rect 5392 9759 5712 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 14288 9824 14608 9825
rect 14288 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14608 9824
rect 14288 9759 14608 9760
rect 2037 9754 2103 9757
rect 3049 9754 3115 9757
rect 0 9752 3115 9754
rect 0 9696 2042 9752
rect 2098 9696 3054 9752
rect 3110 9696 3115 9752
rect 0 9694 3115 9696
rect 0 9664 800 9694
rect 2037 9691 2103 9694
rect 3049 9691 3115 9694
rect 12985 9754 13051 9757
rect 13118 9754 13124 9756
rect 12985 9752 13124 9754
rect 12985 9696 12990 9752
rect 13046 9696 13124 9752
rect 12985 9694 13124 9696
rect 12985 9691 13051 9694
rect 13118 9692 13124 9694
rect 13188 9692 13194 9756
rect 17769 9618 17835 9621
rect 19200 9618 20000 9648
rect 17769 9616 20000 9618
rect 17769 9560 17774 9616
rect 17830 9560 20000 9616
rect 17769 9558 20000 9560
rect 17769 9555 17835 9558
rect 19200 9528 20000 9558
rect 12065 9482 12131 9485
rect 13445 9482 13511 9485
rect 12065 9480 13511 9482
rect 12065 9424 12070 9480
rect 12126 9424 13450 9480
rect 13506 9424 13511 9480
rect 12065 9422 13511 9424
rect 12065 9419 12131 9422
rect 13445 9419 13511 9422
rect 0 9346 800 9376
rect 1301 9346 1367 9349
rect 5165 9348 5231 9349
rect 7281 9348 7347 9349
rect 5165 9346 5212 9348
rect 0 9344 1367 9346
rect 0 9288 1306 9344
rect 1362 9288 1367 9344
rect 0 9286 1367 9288
rect 5120 9344 5212 9346
rect 5120 9288 5170 9344
rect 5120 9286 5212 9288
rect 0 9256 800 9286
rect 1301 9283 1367 9286
rect 5165 9284 5212 9286
rect 5276 9284 5282 9348
rect 7230 9284 7236 9348
rect 7300 9346 7347 9348
rect 7300 9344 7392 9346
rect 7342 9288 7392 9344
rect 7300 9286 7392 9288
rect 7300 9284 7347 9286
rect 5165 9283 5231 9284
rect 7281 9283 7347 9284
rect 3168 9280 3488 9281
rect 3168 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3488 9280
rect 3168 9215 3488 9216
rect 7616 9280 7936 9281
rect 7616 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7936 9280
rect 7616 9215 7936 9216
rect 12064 9280 12384 9281
rect 12064 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12384 9280
rect 12064 9215 12384 9216
rect 16512 9280 16832 9281
rect 16512 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16832 9280
rect 16512 9215 16832 9216
rect 17861 9210 17927 9213
rect 19200 9210 20000 9240
rect 17861 9208 20000 9210
rect 17861 9152 17866 9208
rect 17922 9152 20000 9208
rect 17861 9150 20000 9152
rect 17861 9147 17927 9150
rect 19200 9120 20000 9150
rect 9949 9074 10015 9077
rect 12801 9074 12867 9077
rect 9949 9072 12867 9074
rect 9949 9016 9954 9072
rect 10010 9016 12806 9072
rect 12862 9016 12867 9072
rect 9949 9014 12867 9016
rect 9949 9011 10015 9014
rect 12801 9011 12867 9014
rect 0 8938 800 8968
rect 3509 8938 3575 8941
rect 0 8936 3575 8938
rect 0 8880 3514 8936
rect 3570 8880 3575 8936
rect 0 8878 3575 8880
rect 0 8848 800 8878
rect 3509 8875 3575 8878
rect 5625 8938 5691 8941
rect 6085 8938 6151 8941
rect 11697 8938 11763 8941
rect 5625 8936 11763 8938
rect 5625 8880 5630 8936
rect 5686 8880 6090 8936
rect 6146 8880 11702 8936
rect 11758 8880 11763 8936
rect 5625 8878 11763 8880
rect 5625 8875 5691 8878
rect 6085 8875 6151 8878
rect 11697 8875 11763 8878
rect 11881 8938 11947 8941
rect 14733 8938 14799 8941
rect 11881 8936 14799 8938
rect 11881 8880 11886 8936
rect 11942 8880 14738 8936
rect 14794 8880 14799 8936
rect 11881 8878 14799 8880
rect 11881 8875 11947 8878
rect 14733 8875 14799 8878
rect 7230 8740 7236 8804
rect 7300 8802 7306 8804
rect 9397 8802 9463 8805
rect 7300 8800 9463 8802
rect 7300 8744 9402 8800
rect 9458 8744 9463 8800
rect 7300 8742 9463 8744
rect 7300 8740 7306 8742
rect 9397 8739 9463 8742
rect 10501 8802 10567 8805
rect 12985 8802 13051 8805
rect 10501 8800 13051 8802
rect 10501 8744 10506 8800
rect 10562 8744 12990 8800
rect 13046 8744 13051 8800
rect 10501 8742 13051 8744
rect 10501 8739 10567 8742
rect 12985 8739 13051 8742
rect 16205 8802 16271 8805
rect 19200 8802 20000 8832
rect 16205 8800 20000 8802
rect 16205 8744 16210 8800
rect 16266 8744 20000 8800
rect 16205 8742 20000 8744
rect 16205 8739 16271 8742
rect 5392 8736 5712 8737
rect 5392 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5712 8736
rect 5392 8671 5712 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 14288 8736 14608 8737
rect 14288 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14608 8736
rect 19200 8712 20000 8742
rect 14288 8671 14608 8672
rect 2814 8604 2820 8668
rect 2884 8666 2890 8668
rect 3969 8666 4035 8669
rect 15009 8666 15075 8669
rect 16481 8666 16547 8669
rect 2884 8664 5274 8666
rect 2884 8608 3974 8664
rect 4030 8608 5274 8664
rect 2884 8606 5274 8608
rect 2884 8604 2890 8606
rect 3969 8603 4035 8606
rect 0 8530 800 8560
rect 1485 8530 1551 8533
rect 0 8528 1551 8530
rect 0 8472 1490 8528
rect 1546 8472 1551 8528
rect 0 8470 1551 8472
rect 0 8440 800 8470
rect 1485 8467 1551 8470
rect 4245 8530 4311 8533
rect 4470 8530 4476 8532
rect 4245 8528 4476 8530
rect 4245 8472 4250 8528
rect 4306 8472 4476 8528
rect 4245 8470 4476 8472
rect 4245 8467 4311 8470
rect 4470 8468 4476 8470
rect 4540 8468 4546 8532
rect 5214 8530 5274 8606
rect 15009 8664 16547 8666
rect 15009 8608 15014 8664
rect 15070 8608 16486 8664
rect 16542 8608 16547 8664
rect 15009 8606 16547 8608
rect 15009 8603 15075 8606
rect 16481 8603 16547 8606
rect 11513 8530 11579 8533
rect 5214 8528 11579 8530
rect 5214 8472 11518 8528
rect 11574 8472 11579 8528
rect 5214 8470 11579 8472
rect 11513 8467 11579 8470
rect 11697 8530 11763 8533
rect 13813 8530 13879 8533
rect 11697 8528 13879 8530
rect 11697 8472 11702 8528
rect 11758 8472 13818 8528
rect 13874 8472 13879 8528
rect 11697 8470 13879 8472
rect 11697 8467 11763 8470
rect 13813 8467 13879 8470
rect 2446 8332 2452 8396
rect 2516 8394 2522 8396
rect 6913 8394 6979 8397
rect 2516 8392 6979 8394
rect 2516 8336 6918 8392
rect 6974 8336 6979 8392
rect 2516 8334 6979 8336
rect 2516 8332 2522 8334
rect 6913 8331 6979 8334
rect 10961 8394 11027 8397
rect 17033 8394 17099 8397
rect 10961 8392 17099 8394
rect 10961 8336 10966 8392
rect 11022 8336 17038 8392
rect 17094 8336 17099 8392
rect 10961 8334 17099 8336
rect 10961 8331 11027 8334
rect 17033 8331 17099 8334
rect 18137 8258 18203 8261
rect 19200 8258 20000 8288
rect 18137 8256 20000 8258
rect 18137 8200 18142 8256
rect 18198 8200 20000 8256
rect 18137 8198 20000 8200
rect 18137 8195 18203 8198
rect 3168 8192 3488 8193
rect 0 8122 800 8152
rect 3168 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3488 8192
rect 3168 8127 3488 8128
rect 7616 8192 7936 8193
rect 7616 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7936 8192
rect 7616 8127 7936 8128
rect 12064 8192 12384 8193
rect 12064 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12384 8192
rect 12064 8127 12384 8128
rect 16512 8192 16832 8193
rect 16512 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16832 8192
rect 19200 8168 20000 8198
rect 16512 8127 16832 8128
rect 2865 8122 2931 8125
rect 0 8120 2931 8122
rect 0 8064 2870 8120
rect 2926 8064 2931 8120
rect 0 8062 2931 8064
rect 0 8032 800 8062
rect 2865 8059 2931 8062
rect 9673 7986 9739 7989
rect 13537 7986 13603 7989
rect 9673 7984 13603 7986
rect 9673 7928 9678 7984
rect 9734 7928 13542 7984
rect 13598 7928 13603 7984
rect 9673 7926 13603 7928
rect 9673 7923 9739 7926
rect 13537 7923 13603 7926
rect 17309 7984 17375 7989
rect 17309 7928 17314 7984
rect 17370 7928 17375 7984
rect 17309 7923 17375 7928
rect 7005 7850 7071 7853
rect 11145 7850 11211 7853
rect 16941 7850 17007 7853
rect 7005 7848 7114 7850
rect 7005 7792 7010 7848
rect 7066 7792 7114 7848
rect 7005 7787 7114 7792
rect 11145 7848 17007 7850
rect 11145 7792 11150 7848
rect 11206 7792 16946 7848
rect 17002 7792 17007 7848
rect 11145 7790 17007 7792
rect 11145 7787 11211 7790
rect 16941 7787 17007 7790
rect 0 7714 800 7744
rect 1669 7714 1735 7717
rect 0 7712 1735 7714
rect 0 7656 1674 7712
rect 1730 7656 1735 7712
rect 0 7654 1735 7656
rect 0 7624 800 7654
rect 1669 7651 1735 7654
rect 1853 7714 1919 7717
rect 2630 7714 2636 7716
rect 1853 7712 2636 7714
rect 1853 7656 1858 7712
rect 1914 7656 2636 7712
rect 1853 7654 2636 7656
rect 1853 7651 1919 7654
rect 2630 7652 2636 7654
rect 2700 7714 2706 7716
rect 3325 7714 3391 7717
rect 2700 7712 3391 7714
rect 2700 7656 3330 7712
rect 3386 7656 3391 7712
rect 2700 7654 3391 7656
rect 2700 7652 2706 7654
rect 3325 7651 3391 7654
rect 5392 7648 5712 7649
rect 5392 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5712 7648
rect 5392 7583 5712 7584
rect 6913 7578 6979 7581
rect 7054 7578 7114 7787
rect 17312 7717 17372 7923
rect 17769 7850 17835 7853
rect 19200 7850 20000 7880
rect 17769 7848 20000 7850
rect 17769 7792 17774 7848
rect 17830 7792 20000 7848
rect 17769 7790 20000 7792
rect 17769 7787 17835 7790
rect 19200 7760 20000 7790
rect 10501 7714 10567 7717
rect 13169 7714 13235 7717
rect 10501 7712 13235 7714
rect 10501 7656 10506 7712
rect 10562 7656 13174 7712
rect 13230 7656 13235 7712
rect 10501 7654 13235 7656
rect 10501 7651 10567 7654
rect 13169 7651 13235 7654
rect 17309 7712 17375 7717
rect 17309 7656 17314 7712
rect 17370 7656 17375 7712
rect 17309 7651 17375 7656
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 14288 7648 14608 7649
rect 14288 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14608 7648
rect 14288 7583 14608 7584
rect 6913 7576 7114 7578
rect 6913 7520 6918 7576
rect 6974 7520 7114 7576
rect 6913 7518 7114 7520
rect 6913 7515 6979 7518
rect 1669 7444 1735 7445
rect 1669 7442 1716 7444
rect 1624 7440 1716 7442
rect 1780 7442 1786 7444
rect 8661 7442 8727 7445
rect 10501 7442 10567 7445
rect 1780 7440 10567 7442
rect 1624 7384 1674 7440
rect 1780 7384 8666 7440
rect 8722 7384 10506 7440
rect 10562 7384 10567 7440
rect 1624 7382 1716 7384
rect 1669 7380 1716 7382
rect 1780 7382 10567 7384
rect 1780 7380 1786 7382
rect 1669 7379 1735 7380
rect 8661 7379 8727 7382
rect 10501 7379 10567 7382
rect 13353 7442 13419 7445
rect 18413 7442 18479 7445
rect 19200 7442 20000 7472
rect 13353 7440 16130 7442
rect 13353 7384 13358 7440
rect 13414 7384 16130 7440
rect 13353 7382 16130 7384
rect 13353 7379 13419 7382
rect 0 7306 800 7336
rect 3877 7306 3943 7309
rect 0 7304 3943 7306
rect 0 7248 3882 7304
rect 3938 7248 3943 7304
rect 0 7246 3943 7248
rect 0 7216 800 7246
rect 3877 7243 3943 7246
rect 6177 7306 6243 7309
rect 9029 7306 9095 7309
rect 15929 7306 15995 7309
rect 6177 7304 15995 7306
rect 6177 7248 6182 7304
rect 6238 7248 9034 7304
rect 9090 7248 15934 7304
rect 15990 7248 15995 7304
rect 6177 7246 15995 7248
rect 16070 7306 16130 7382
rect 18413 7440 20000 7442
rect 18413 7384 18418 7440
rect 18474 7384 20000 7440
rect 18413 7382 20000 7384
rect 18413 7379 18479 7382
rect 19200 7352 20000 7382
rect 18413 7306 18479 7309
rect 16070 7304 18479 7306
rect 16070 7248 18418 7304
rect 18474 7248 18479 7304
rect 16070 7246 18479 7248
rect 6177 7243 6243 7246
rect 9029 7243 9095 7246
rect 15929 7243 15995 7246
rect 18413 7243 18479 7246
rect 5625 7170 5691 7173
rect 7373 7170 7439 7173
rect 5625 7168 7439 7170
rect 5625 7112 5630 7168
rect 5686 7112 7378 7168
rect 7434 7112 7439 7168
rect 5625 7110 7439 7112
rect 5625 7107 5691 7110
rect 7373 7107 7439 7110
rect 3168 7104 3488 7105
rect 3168 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3488 7104
rect 3168 7039 3488 7040
rect 7616 7104 7936 7105
rect 7616 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7936 7104
rect 7616 7039 7936 7040
rect 12064 7104 12384 7105
rect 12064 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12384 7104
rect 12064 7039 12384 7040
rect 16512 7104 16832 7105
rect 16512 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16832 7104
rect 16512 7039 16832 7040
rect 17861 7034 17927 7037
rect 19200 7034 20000 7064
rect 17861 7032 20000 7034
rect 17861 6976 17866 7032
rect 17922 6976 20000 7032
rect 17861 6974 20000 6976
rect 17861 6971 17927 6974
rect 19200 6944 20000 6974
rect 0 6898 800 6928
rect 3877 6898 3943 6901
rect 0 6896 3943 6898
rect 0 6840 3882 6896
rect 3938 6840 3943 6896
rect 0 6838 3943 6840
rect 0 6808 800 6838
rect 3877 6835 3943 6838
rect 4102 6836 4108 6900
rect 4172 6898 4178 6900
rect 5625 6898 5691 6901
rect 8518 6898 8524 6900
rect 4172 6896 8524 6898
rect 4172 6840 5630 6896
rect 5686 6840 8524 6896
rect 4172 6838 8524 6840
rect 4172 6836 4178 6838
rect 5625 6835 5691 6838
rect 8518 6836 8524 6838
rect 8588 6898 8594 6900
rect 15510 6898 15516 6900
rect 8588 6838 15516 6898
rect 8588 6836 8594 6838
rect 15510 6836 15516 6838
rect 15580 6836 15586 6900
rect 2681 6762 2747 6765
rect 6913 6764 6979 6765
rect 6862 6762 6868 6764
rect 2681 6760 6868 6762
rect 6932 6762 6979 6764
rect 13813 6762 13879 6765
rect 18045 6762 18111 6765
rect 6932 6760 7024 6762
rect 2681 6704 2686 6760
rect 2742 6704 6868 6760
rect 6974 6704 7024 6760
rect 2681 6702 6868 6704
rect 2681 6699 2747 6702
rect 6862 6700 6868 6702
rect 6932 6702 7024 6704
rect 13813 6760 18111 6762
rect 13813 6704 13818 6760
rect 13874 6704 18050 6760
rect 18106 6704 18111 6760
rect 13813 6702 18111 6704
rect 6932 6700 6979 6702
rect 6913 6699 6979 6700
rect 13813 6699 13879 6702
rect 18045 6699 18111 6702
rect 6913 6626 6979 6629
rect 7230 6626 7236 6628
rect 6913 6624 7236 6626
rect 6913 6568 6918 6624
rect 6974 6568 7236 6624
rect 6913 6566 7236 6568
rect 6913 6563 6979 6566
rect 7230 6564 7236 6566
rect 7300 6564 7306 6628
rect 17677 6626 17743 6629
rect 19200 6626 20000 6656
rect 17677 6624 20000 6626
rect 17677 6568 17682 6624
rect 17738 6568 20000 6624
rect 17677 6566 20000 6568
rect 17677 6563 17743 6566
rect 5392 6560 5712 6561
rect 0 6490 800 6520
rect 5392 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5712 6560
rect 5392 6495 5712 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 14288 6560 14608 6561
rect 14288 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14608 6560
rect 19200 6536 20000 6566
rect 14288 6495 14608 6496
rect 1485 6490 1551 6493
rect 0 6488 1551 6490
rect 0 6432 1490 6488
rect 1546 6432 1551 6488
rect 0 6430 1551 6432
rect 0 6400 800 6430
rect 1485 6427 1551 6430
rect 2405 6492 2471 6493
rect 2405 6488 2452 6492
rect 2516 6490 2522 6492
rect 10961 6490 11027 6493
rect 13813 6490 13879 6493
rect 2405 6432 2410 6488
rect 2405 6428 2452 6432
rect 2516 6430 2562 6490
rect 10961 6488 13879 6490
rect 10961 6432 10966 6488
rect 11022 6432 13818 6488
rect 13874 6432 13879 6488
rect 10961 6430 13879 6432
rect 2516 6428 2522 6430
rect 2405 6427 2471 6428
rect 10961 6427 11027 6430
rect 13813 6427 13879 6430
rect 4521 6354 4587 6357
rect 7230 6354 7236 6356
rect 4521 6352 7236 6354
rect 4521 6296 4526 6352
rect 4582 6296 7236 6352
rect 4521 6294 7236 6296
rect 4521 6291 4587 6294
rect 7230 6292 7236 6294
rect 7300 6292 7306 6356
rect 8109 6354 8175 6357
rect 8477 6354 8543 6357
rect 8845 6354 8911 6357
rect 8109 6352 8911 6354
rect 8109 6296 8114 6352
rect 8170 6296 8482 6352
rect 8538 6296 8850 6352
rect 8906 6296 8911 6352
rect 8109 6294 8911 6296
rect 8109 6291 8175 6294
rect 8477 6291 8543 6294
rect 8845 6291 8911 6294
rect 11237 6354 11303 6357
rect 15929 6354 15995 6357
rect 11237 6352 15995 6354
rect 11237 6296 11242 6352
rect 11298 6296 15934 6352
rect 15990 6296 15995 6352
rect 11237 6294 15995 6296
rect 11237 6291 11303 6294
rect 15929 6291 15995 6294
rect 2313 6218 2379 6221
rect 3049 6218 3115 6221
rect 2313 6216 3115 6218
rect 2313 6160 2318 6216
rect 2374 6160 3054 6216
rect 3110 6160 3115 6216
rect 2313 6158 3115 6160
rect 2313 6155 2379 6158
rect 3049 6155 3115 6158
rect 6637 6218 6703 6221
rect 10910 6218 10916 6220
rect 6637 6216 10916 6218
rect 6637 6160 6642 6216
rect 6698 6160 10916 6216
rect 6637 6158 10916 6160
rect 6637 6155 6703 6158
rect 10910 6156 10916 6158
rect 10980 6156 10986 6220
rect 12341 6218 12407 6221
rect 17309 6218 17375 6221
rect 12341 6216 17375 6218
rect 12341 6160 12346 6216
rect 12402 6160 17314 6216
rect 17370 6160 17375 6216
rect 12341 6158 17375 6160
rect 12341 6155 12407 6158
rect 17309 6155 17375 6158
rect 18045 6218 18111 6221
rect 19200 6218 20000 6248
rect 18045 6216 20000 6218
rect 18045 6160 18050 6216
rect 18106 6160 20000 6216
rect 18045 6158 20000 6160
rect 18045 6155 18111 6158
rect 19200 6128 20000 6158
rect 0 6082 800 6112
rect 1393 6082 1459 6085
rect 0 6080 1459 6082
rect 0 6024 1398 6080
rect 1454 6024 1459 6080
rect 0 6022 1459 6024
rect 0 5992 800 6022
rect 1393 6019 1459 6022
rect 4337 6082 4403 6085
rect 7465 6082 7531 6085
rect 4337 6080 7531 6082
rect 4337 6024 4342 6080
rect 4398 6024 7470 6080
rect 7526 6024 7531 6080
rect 4337 6022 7531 6024
rect 4337 6019 4403 6022
rect 7465 6019 7531 6022
rect 8569 6082 8635 6085
rect 9305 6082 9371 6085
rect 8569 6080 9371 6082
rect 8569 6024 8574 6080
rect 8630 6024 9310 6080
rect 9366 6024 9371 6080
rect 8569 6022 9371 6024
rect 8569 6019 8635 6022
rect 9305 6019 9371 6022
rect 3168 6016 3488 6017
rect 3168 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3488 6016
rect 3168 5951 3488 5952
rect 7616 6016 7936 6017
rect 7616 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7936 6016
rect 7616 5951 7936 5952
rect 12064 6016 12384 6017
rect 12064 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12384 6016
rect 12064 5951 12384 5952
rect 16512 6016 16832 6017
rect 16512 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16832 6016
rect 16512 5951 16832 5952
rect 3877 5946 3943 5949
rect 5073 5946 5139 5949
rect 3877 5944 5139 5946
rect 3877 5888 3882 5944
rect 3938 5888 5078 5944
rect 5134 5888 5139 5944
rect 3877 5886 5139 5888
rect 3877 5883 3943 5886
rect 5073 5883 5139 5886
rect 8753 5946 8819 5949
rect 8753 5944 9874 5946
rect 8753 5888 8758 5944
rect 8814 5888 9874 5944
rect 8753 5886 9874 5888
rect 8753 5883 8819 5886
rect 9581 5810 9647 5813
rect 4110 5808 9647 5810
rect 4110 5752 9586 5808
rect 9642 5752 9647 5808
rect 4110 5750 9647 5752
rect 0 5538 800 5568
rect 4110 5538 4170 5750
rect 9581 5747 9647 5750
rect 4654 5612 4660 5676
rect 4724 5674 4730 5676
rect 6545 5674 6611 5677
rect 4724 5672 6611 5674
rect 4724 5616 6550 5672
rect 6606 5616 6611 5672
rect 4724 5614 6611 5616
rect 4724 5612 4730 5614
rect 6545 5611 6611 5614
rect 8334 5612 8340 5676
rect 8404 5674 8410 5676
rect 9213 5674 9279 5677
rect 8404 5672 9279 5674
rect 8404 5616 9218 5672
rect 9274 5616 9279 5672
rect 8404 5614 9279 5616
rect 9814 5674 9874 5886
rect 13721 5810 13787 5813
rect 14641 5810 14707 5813
rect 13721 5808 14707 5810
rect 13721 5752 13726 5808
rect 13782 5752 14646 5808
rect 14702 5752 14707 5808
rect 13721 5750 14707 5752
rect 13721 5747 13787 5750
rect 14641 5747 14707 5750
rect 15377 5810 15443 5813
rect 15510 5810 15516 5812
rect 15377 5808 15516 5810
rect 15377 5752 15382 5808
rect 15438 5752 15516 5808
rect 15377 5750 15516 5752
rect 15377 5747 15443 5750
rect 15510 5748 15516 5750
rect 15580 5748 15586 5812
rect 15101 5674 15167 5677
rect 9814 5672 15167 5674
rect 9814 5616 15106 5672
rect 15162 5616 15167 5672
rect 9814 5614 15167 5616
rect 8404 5612 8410 5614
rect 9213 5611 9279 5614
rect 15101 5611 15167 5614
rect 18413 5674 18479 5677
rect 19200 5674 20000 5704
rect 18413 5672 20000 5674
rect 18413 5616 18418 5672
rect 18474 5616 20000 5672
rect 18413 5614 20000 5616
rect 18413 5611 18479 5614
rect 19200 5584 20000 5614
rect 0 5478 4170 5538
rect 4613 5538 4679 5541
rect 4981 5538 5047 5541
rect 4613 5536 5047 5538
rect 4613 5480 4618 5536
rect 4674 5480 4986 5536
rect 5042 5480 5047 5536
rect 4613 5478 5047 5480
rect 0 5448 800 5478
rect 4613 5475 4679 5478
rect 4981 5475 5047 5478
rect 7557 5538 7623 5541
rect 8937 5538 9003 5541
rect 7557 5536 9003 5538
rect 7557 5480 7562 5536
rect 7618 5480 8942 5536
rect 8998 5480 9003 5536
rect 7557 5478 9003 5480
rect 7557 5475 7623 5478
rect 8937 5475 9003 5478
rect 16062 5476 16068 5540
rect 16132 5538 16138 5540
rect 16481 5538 16547 5541
rect 16132 5536 16547 5538
rect 16132 5480 16486 5536
rect 16542 5480 16547 5536
rect 16132 5478 16547 5480
rect 16132 5476 16138 5478
rect 16481 5475 16547 5478
rect 5392 5472 5712 5473
rect 5392 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5712 5472
rect 5392 5407 5712 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 14288 5472 14608 5473
rect 14288 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14608 5472
rect 14288 5407 14608 5408
rect 16849 5402 16915 5405
rect 17166 5402 17172 5404
rect 14782 5400 17172 5402
rect 14782 5344 16854 5400
rect 16910 5344 17172 5400
rect 14782 5342 17172 5344
rect 4429 5266 4495 5269
rect 10133 5266 10199 5269
rect 4429 5264 10199 5266
rect 4429 5208 4434 5264
rect 4490 5208 10138 5264
rect 10194 5208 10199 5264
rect 4429 5206 10199 5208
rect 4429 5203 4495 5206
rect 10133 5203 10199 5206
rect 13261 5266 13327 5269
rect 14782 5266 14842 5342
rect 16849 5339 16915 5342
rect 17166 5340 17172 5342
rect 17236 5340 17242 5404
rect 13261 5264 14842 5266
rect 13261 5208 13266 5264
rect 13322 5208 14842 5264
rect 13261 5206 14842 5208
rect 18045 5266 18111 5269
rect 19200 5266 20000 5296
rect 18045 5264 20000 5266
rect 18045 5208 18050 5264
rect 18106 5208 20000 5264
rect 18045 5206 20000 5208
rect 13261 5203 13327 5206
rect 18045 5203 18111 5206
rect 19200 5176 20000 5206
rect 0 5130 800 5160
rect 933 5130 999 5133
rect 0 5128 999 5130
rect 0 5072 938 5128
rect 994 5072 999 5128
rect 0 5070 999 5072
rect 0 5040 800 5070
rect 933 5067 999 5070
rect 14365 5130 14431 5133
rect 15193 5130 15259 5133
rect 14365 5128 15259 5130
rect 14365 5072 14370 5128
rect 14426 5072 15198 5128
rect 15254 5072 15259 5128
rect 14365 5070 15259 5072
rect 14365 5067 14431 5070
rect 15193 5067 15259 5070
rect 3693 4994 3759 4997
rect 7189 4994 7255 4997
rect 3693 4992 7255 4994
rect 3693 4936 3698 4992
rect 3754 4936 7194 4992
rect 7250 4936 7255 4992
rect 3693 4934 7255 4936
rect 3693 4931 3759 4934
rect 7189 4931 7255 4934
rect 3168 4928 3488 4929
rect 3168 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3488 4928
rect 3168 4863 3488 4864
rect 7616 4928 7936 4929
rect 7616 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7936 4928
rect 7616 4863 7936 4864
rect 12064 4928 12384 4929
rect 12064 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12384 4928
rect 12064 4863 12384 4864
rect 16512 4928 16832 4929
rect 16512 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16832 4928
rect 16512 4863 16832 4864
rect 3877 4858 3943 4861
rect 16297 4860 16363 4861
rect 4102 4858 4108 4860
rect 3877 4856 4108 4858
rect 3877 4800 3882 4856
rect 3938 4800 4108 4856
rect 3877 4798 4108 4800
rect 3877 4795 3943 4798
rect 4102 4796 4108 4798
rect 4172 4796 4178 4860
rect 16246 4796 16252 4860
rect 16316 4858 16363 4860
rect 18321 4858 18387 4861
rect 19200 4858 20000 4888
rect 16316 4856 16408 4858
rect 16358 4800 16408 4856
rect 16316 4798 16408 4800
rect 18321 4856 20000 4858
rect 18321 4800 18326 4856
rect 18382 4800 20000 4856
rect 18321 4798 20000 4800
rect 16316 4796 16363 4798
rect 16297 4795 16363 4796
rect 18321 4795 18387 4798
rect 19200 4768 20000 4798
rect 0 4722 800 4752
rect 3877 4722 3943 4725
rect 0 4720 3943 4722
rect 0 4664 3882 4720
rect 3938 4664 3943 4720
rect 0 4662 3943 4664
rect 0 4632 800 4662
rect 3877 4659 3943 4662
rect 16389 4722 16455 4725
rect 18321 4722 18387 4725
rect 16389 4720 18387 4722
rect 16389 4664 16394 4720
rect 16450 4664 18326 4720
rect 18382 4664 18387 4720
rect 16389 4662 18387 4664
rect 16389 4659 16455 4662
rect 18321 4659 18387 4662
rect 18045 4450 18111 4453
rect 19200 4450 20000 4480
rect 18045 4448 20000 4450
rect 18045 4392 18050 4448
rect 18106 4392 20000 4448
rect 18045 4390 20000 4392
rect 18045 4387 18111 4390
rect 5392 4384 5712 4385
rect 0 4314 800 4344
rect 5392 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5712 4384
rect 5392 4319 5712 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 14288 4384 14608 4385
rect 14288 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14608 4384
rect 19200 4360 20000 4390
rect 14288 4319 14608 4320
rect 17033 4314 17099 4317
rect 0 4254 2790 4314
rect 0 4224 800 4254
rect 2730 4178 2790 4254
rect 14966 4312 17099 4314
rect 14966 4256 17038 4312
rect 17094 4256 17099 4312
rect 14966 4254 17099 4256
rect 9213 4178 9279 4181
rect 2730 4176 9279 4178
rect 2730 4120 9218 4176
rect 9274 4120 9279 4176
rect 2730 4118 9279 4120
rect 9213 4115 9279 4118
rect 10777 4178 10843 4181
rect 13905 4178 13971 4181
rect 14966 4178 15026 4254
rect 17033 4251 17099 4254
rect 10777 4176 15026 4178
rect 10777 4120 10782 4176
rect 10838 4120 13910 4176
rect 13966 4120 15026 4176
rect 10777 4118 15026 4120
rect 10777 4115 10843 4118
rect 13905 4115 13971 4118
rect 15142 4116 15148 4180
rect 15212 4178 15218 4180
rect 15285 4178 15351 4181
rect 15212 4176 15351 4178
rect 15212 4120 15290 4176
rect 15346 4120 15351 4176
rect 15212 4118 15351 4120
rect 15212 4116 15218 4118
rect 15285 4115 15351 4118
rect 1669 4044 1735 4045
rect 1669 4040 1716 4044
rect 1780 4042 1786 4044
rect 2129 4042 2195 4045
rect 2630 4042 2636 4044
rect 1669 3984 1674 4040
rect 1669 3980 1716 3984
rect 1780 3982 1826 4042
rect 2129 4040 2636 4042
rect 2129 3984 2134 4040
rect 2190 3984 2636 4040
rect 2129 3982 2636 3984
rect 1780 3980 1786 3982
rect 1669 3979 1735 3980
rect 2129 3979 2195 3982
rect 2630 3980 2636 3982
rect 2700 3980 2706 4044
rect 4429 4042 4495 4045
rect 4654 4042 4660 4044
rect 4429 4040 4660 4042
rect 4429 3984 4434 4040
rect 4490 3984 4660 4040
rect 4429 3982 4660 3984
rect 4429 3979 4495 3982
rect 4654 3980 4660 3982
rect 4724 3980 4730 4044
rect 6545 4042 6611 4045
rect 8385 4042 8451 4045
rect 8569 4044 8635 4045
rect 6545 4040 8451 4042
rect 6545 3984 6550 4040
rect 6606 3984 8390 4040
rect 8446 3984 8451 4040
rect 6545 3982 8451 3984
rect 6545 3979 6611 3982
rect 8385 3979 8451 3982
rect 8518 3980 8524 4044
rect 8588 4042 8635 4044
rect 9489 4042 9555 4045
rect 15929 4042 15995 4045
rect 8588 4040 8680 4042
rect 8630 3984 8680 4040
rect 8588 3982 8680 3984
rect 9489 4040 15995 4042
rect 9489 3984 9494 4040
rect 9550 3984 15934 4040
rect 15990 3984 15995 4040
rect 9489 3982 15995 3984
rect 8588 3980 8635 3982
rect 8569 3979 8635 3980
rect 9489 3979 9555 3982
rect 15929 3979 15995 3982
rect 17861 4042 17927 4045
rect 19200 4042 20000 4072
rect 17861 4040 20000 4042
rect 17861 3984 17866 4040
rect 17922 3984 20000 4040
rect 17861 3982 20000 3984
rect 17861 3979 17927 3982
rect 19200 3952 20000 3982
rect 0 3906 800 3936
rect 2865 3906 2931 3909
rect 0 3904 2931 3906
rect 0 3848 2870 3904
rect 2926 3848 2931 3904
rect 0 3846 2931 3848
rect 0 3816 800 3846
rect 2865 3843 2931 3846
rect 3969 3906 4035 3909
rect 4797 3906 4863 3909
rect 3969 3904 4863 3906
rect 3969 3848 3974 3904
rect 4030 3848 4802 3904
rect 4858 3848 4863 3904
rect 3969 3846 4863 3848
rect 3969 3843 4035 3846
rect 4797 3843 4863 3846
rect 3168 3840 3488 3841
rect 3168 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3488 3840
rect 3168 3775 3488 3776
rect 7616 3840 7936 3841
rect 7616 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7936 3840
rect 7616 3775 7936 3776
rect 12064 3840 12384 3841
rect 12064 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12384 3840
rect 12064 3775 12384 3776
rect 16512 3840 16832 3841
rect 16512 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16832 3840
rect 16512 3775 16832 3776
rect 3969 3770 4035 3773
rect 4981 3770 5047 3773
rect 5257 3770 5323 3773
rect 3969 3768 5323 3770
rect 3969 3712 3974 3768
rect 4030 3712 4986 3768
rect 5042 3712 5262 3768
rect 5318 3712 5323 3768
rect 3969 3710 5323 3712
rect 3969 3707 4035 3710
rect 4981 3707 5047 3710
rect 5257 3707 5323 3710
rect 10501 3770 10567 3773
rect 10501 3768 11346 3770
rect 10501 3712 10506 3768
rect 10562 3712 11346 3768
rect 10501 3710 11346 3712
rect 10501 3707 10567 3710
rect 3785 3634 3851 3637
rect 1902 3632 3851 3634
rect 1902 3576 3790 3632
rect 3846 3576 3851 3632
rect 1902 3574 3851 3576
rect 0 3498 800 3528
rect 1902 3498 1962 3574
rect 3785 3571 3851 3574
rect 4429 3634 4495 3637
rect 11053 3634 11119 3637
rect 4429 3632 11119 3634
rect 4429 3576 4434 3632
rect 4490 3576 11058 3632
rect 11114 3576 11119 3632
rect 4429 3574 11119 3576
rect 11286 3634 11346 3710
rect 16021 3634 16087 3637
rect 11286 3632 16087 3634
rect 11286 3576 16026 3632
rect 16082 3576 16087 3632
rect 11286 3574 16087 3576
rect 4429 3571 4495 3574
rect 11053 3571 11119 3574
rect 16021 3571 16087 3574
rect 18413 3634 18479 3637
rect 19200 3634 20000 3664
rect 18413 3632 20000 3634
rect 18413 3576 18418 3632
rect 18474 3576 20000 3632
rect 18413 3574 20000 3576
rect 18413 3571 18479 3574
rect 19200 3544 20000 3574
rect 0 3438 1962 3498
rect 4153 3498 4219 3501
rect 5206 3498 5212 3500
rect 4153 3496 5212 3498
rect 4153 3440 4158 3496
rect 4214 3440 5212 3496
rect 4153 3438 5212 3440
rect 0 3408 800 3438
rect 4153 3435 4219 3438
rect 5206 3436 5212 3438
rect 5276 3498 5282 3500
rect 8385 3498 8451 3501
rect 5276 3496 8451 3498
rect 5276 3440 8390 3496
rect 8446 3440 8451 3496
rect 5276 3438 8451 3440
rect 5276 3436 5282 3438
rect 8385 3435 8451 3438
rect 11053 3498 11119 3501
rect 16941 3498 17007 3501
rect 11053 3496 17007 3498
rect 11053 3440 11058 3496
rect 11114 3440 16946 3496
rect 17002 3440 17007 3496
rect 11053 3438 17007 3440
rect 11053 3435 11119 3438
rect 16941 3435 17007 3438
rect 2221 3362 2287 3365
rect 5165 3362 5231 3365
rect 2221 3360 5231 3362
rect 2221 3304 2226 3360
rect 2282 3304 5170 3360
rect 5226 3304 5231 3360
rect 2221 3302 5231 3304
rect 2221 3299 2287 3302
rect 5165 3299 5231 3302
rect 6269 3362 6335 3365
rect 7465 3362 7531 3365
rect 6269 3360 7531 3362
rect 6269 3304 6274 3360
rect 6330 3304 7470 3360
rect 7526 3304 7531 3360
rect 6269 3302 7531 3304
rect 6269 3299 6335 3302
rect 7465 3299 7531 3302
rect 5392 3296 5712 3297
rect 5392 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5712 3296
rect 5392 3231 5712 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 14288 3296 14608 3297
rect 14288 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14608 3296
rect 14288 3231 14608 3232
rect 6913 3226 6979 3229
rect 17033 3228 17099 3229
rect 6913 3224 7666 3226
rect 6913 3168 6918 3224
rect 6974 3168 7666 3224
rect 6913 3166 7666 3168
rect 6913 3163 6979 3166
rect 0 3090 800 3120
rect 7606 3093 7666 3166
rect 16982 3164 16988 3228
rect 17052 3226 17099 3228
rect 18045 3226 18111 3229
rect 19200 3226 20000 3256
rect 17052 3224 17144 3226
rect 17094 3168 17144 3224
rect 17052 3166 17144 3168
rect 18045 3224 20000 3226
rect 18045 3168 18050 3224
rect 18106 3168 20000 3224
rect 18045 3166 20000 3168
rect 17052 3164 17099 3166
rect 17033 3163 17099 3164
rect 18045 3163 18111 3166
rect 19200 3136 20000 3166
rect 5533 3090 5599 3093
rect 0 3088 5599 3090
rect 0 3032 5538 3088
rect 5594 3032 5599 3088
rect 0 3030 5599 3032
rect 0 3000 800 3030
rect 5533 3027 5599 3030
rect 7230 3028 7236 3092
rect 7300 3090 7306 3092
rect 7373 3090 7439 3093
rect 7300 3088 7439 3090
rect 7300 3032 7378 3088
rect 7434 3032 7439 3088
rect 7300 3030 7439 3032
rect 7606 3090 7715 3093
rect 16849 3090 16915 3093
rect 17953 3090 18019 3093
rect 7606 3088 18019 3090
rect 7606 3032 7654 3088
rect 7710 3032 16854 3088
rect 16910 3032 17958 3088
rect 18014 3032 18019 3088
rect 7606 3030 18019 3032
rect 7300 3028 7306 3030
rect 7373 3027 7439 3030
rect 7649 3027 7715 3030
rect 16849 3027 16915 3030
rect 17953 3027 18019 3030
rect 933 2954 999 2957
rect 16757 2954 16823 2957
rect 933 2952 16823 2954
rect 933 2896 938 2952
rect 994 2896 16762 2952
rect 16818 2896 16823 2952
rect 933 2894 16823 2896
rect 933 2891 999 2894
rect 16757 2891 16823 2894
rect 16941 2820 17007 2821
rect 16941 2816 16988 2820
rect 17052 2818 17058 2820
rect 16941 2760 16946 2816
rect 16941 2756 16988 2760
rect 17052 2758 17098 2818
rect 17052 2756 17058 2758
rect 16941 2755 17007 2756
rect 3168 2752 3488 2753
rect 0 2682 800 2712
rect 3168 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3488 2752
rect 3168 2687 3488 2688
rect 7616 2752 7936 2753
rect 7616 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7936 2752
rect 7616 2687 7936 2688
rect 12064 2752 12384 2753
rect 12064 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12384 2752
rect 12064 2687 12384 2688
rect 16512 2752 16832 2753
rect 16512 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16832 2752
rect 16512 2687 16832 2688
rect 2313 2682 2379 2685
rect 2814 2682 2820 2684
rect 0 2622 2146 2682
rect 0 2592 800 2622
rect 2086 2410 2146 2622
rect 2313 2680 2820 2682
rect 2313 2624 2318 2680
rect 2374 2624 2820 2680
rect 2313 2622 2820 2624
rect 2313 2619 2379 2622
rect 2814 2620 2820 2622
rect 2884 2620 2890 2684
rect 5533 2682 5599 2685
rect 5533 2680 6010 2682
rect 5533 2624 5538 2680
rect 5594 2624 6010 2680
rect 5533 2622 6010 2624
rect 5533 2619 5599 2622
rect 5950 2549 6010 2622
rect 13118 2620 13124 2684
rect 13188 2682 13194 2684
rect 15469 2682 15535 2685
rect 13188 2680 15535 2682
rect 13188 2624 15474 2680
rect 15530 2624 15535 2680
rect 13188 2622 15535 2624
rect 13188 2620 13194 2622
rect 15469 2619 15535 2622
rect 18045 2682 18111 2685
rect 19200 2682 20000 2712
rect 18045 2680 20000 2682
rect 18045 2624 18050 2680
rect 18106 2624 20000 2680
rect 18045 2622 20000 2624
rect 18045 2619 18111 2622
rect 19200 2592 20000 2622
rect 3918 2484 3924 2548
rect 3988 2546 3994 2548
rect 4337 2546 4403 2549
rect 3988 2544 4403 2546
rect 3988 2488 4342 2544
rect 4398 2488 4403 2544
rect 3988 2486 4403 2488
rect 3988 2484 3994 2486
rect 4337 2483 4403 2486
rect 4654 2484 4660 2548
rect 4724 2546 4730 2548
rect 5717 2546 5783 2549
rect 4724 2544 5783 2546
rect 4724 2488 5722 2544
rect 5778 2488 5783 2544
rect 4724 2486 5783 2488
rect 4724 2484 4730 2486
rect 5717 2483 5783 2486
rect 5901 2546 6010 2549
rect 10225 2546 10291 2549
rect 5901 2544 10291 2546
rect 5901 2488 5906 2544
rect 5962 2488 10230 2544
rect 10286 2488 10291 2544
rect 5901 2486 10291 2488
rect 5901 2483 5967 2486
rect 10225 2483 10291 2486
rect 10910 2484 10916 2548
rect 10980 2546 10986 2548
rect 12985 2546 13051 2549
rect 10980 2544 13051 2546
rect 10980 2488 12990 2544
rect 13046 2488 13051 2544
rect 10980 2486 13051 2488
rect 10980 2484 10986 2486
rect 12985 2483 13051 2486
rect 4705 2410 4771 2413
rect 10961 2410 11027 2413
rect 16246 2410 16252 2412
rect 2086 2408 4771 2410
rect 2086 2352 4710 2408
rect 4766 2352 4771 2408
rect 2086 2350 4771 2352
rect 4705 2347 4771 2350
rect 5214 2408 11027 2410
rect 5214 2352 10966 2408
rect 11022 2352 11027 2408
rect 5214 2350 11027 2352
rect 0 2274 800 2304
rect 3877 2274 3943 2277
rect 0 2272 3943 2274
rect 0 2216 3882 2272
rect 3938 2216 3943 2272
rect 0 2214 3943 2216
rect 0 2184 800 2214
rect 3877 2211 3943 2214
rect 4613 2274 4679 2277
rect 5214 2274 5274 2350
rect 10961 2347 11027 2350
rect 12390 2350 16252 2410
rect 6913 2276 6979 2277
rect 6862 2274 6868 2276
rect 4613 2272 5274 2274
rect 4613 2216 4618 2272
rect 4674 2216 5274 2272
rect 4613 2214 5274 2216
rect 6822 2214 6868 2274
rect 6932 2272 6979 2276
rect 6974 2216 6979 2272
rect 4613 2211 4679 2214
rect 6862 2212 6868 2214
rect 6932 2212 6979 2216
rect 6913 2211 6979 2212
rect 10225 2274 10291 2277
rect 12390 2274 12450 2350
rect 16246 2348 16252 2350
rect 16316 2348 16322 2412
rect 10225 2272 12450 2274
rect 10225 2216 10230 2272
rect 10286 2216 12450 2272
rect 10225 2214 12450 2216
rect 18229 2274 18295 2277
rect 19200 2274 20000 2304
rect 18229 2272 20000 2274
rect 18229 2216 18234 2272
rect 18290 2216 20000 2272
rect 18229 2214 20000 2216
rect 10225 2211 10291 2214
rect 18229 2211 18295 2214
rect 5392 2208 5712 2209
rect 5392 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5712 2208
rect 5392 2143 5712 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 14288 2208 14608 2209
rect 14288 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14608 2208
rect 19200 2184 20000 2214
rect 14288 2143 14608 2144
rect 2865 2002 2931 2005
rect 8334 2002 8340 2004
rect 2865 2000 8340 2002
rect 2865 1944 2870 2000
rect 2926 1944 8340 2000
rect 2865 1942 8340 1944
rect 2865 1939 2931 1942
rect 8334 1940 8340 1942
rect 8404 1940 8410 2004
rect 0 1866 800 1896
rect 4061 1866 4127 1869
rect 0 1864 4127 1866
rect 0 1808 4066 1864
rect 4122 1808 4127 1864
rect 0 1806 4127 1808
rect 0 1776 800 1806
rect 4061 1803 4127 1806
rect 17309 1866 17375 1869
rect 19200 1866 20000 1896
rect 17309 1864 20000 1866
rect 17309 1808 17314 1864
rect 17370 1808 20000 1864
rect 17309 1806 20000 1808
rect 17309 1803 17375 1806
rect 19200 1776 20000 1806
rect 0 1458 800 1488
rect 3325 1458 3391 1461
rect 0 1456 3391 1458
rect 0 1400 3330 1456
rect 3386 1400 3391 1456
rect 0 1398 3391 1400
rect 0 1368 800 1398
rect 3325 1395 3391 1398
rect 17677 1458 17743 1461
rect 19200 1458 20000 1488
rect 17677 1456 20000 1458
rect 17677 1400 17682 1456
rect 17738 1400 20000 1456
rect 17677 1398 20000 1400
rect 17677 1395 17743 1398
rect 19200 1368 20000 1398
rect 0 1050 800 1080
rect 4061 1050 4127 1053
rect 0 1048 4127 1050
rect 0 992 4066 1048
rect 4122 992 4127 1048
rect 0 990 4127 992
rect 0 960 800 990
rect 4061 987 4127 990
rect 17861 1050 17927 1053
rect 19200 1050 20000 1080
rect 17861 1048 20000 1050
rect 17861 992 17866 1048
rect 17922 992 20000 1048
rect 17861 990 20000 992
rect 17861 987 17927 990
rect 19200 960 20000 990
rect 0 642 800 672
rect 3693 642 3759 645
rect 0 640 3759 642
rect 0 584 3698 640
rect 3754 584 3759 640
rect 0 582 3759 584
rect 0 552 800 582
rect 3693 579 3759 582
rect 18137 642 18203 645
rect 19200 642 20000 672
rect 18137 640 20000 642
rect 18137 584 18142 640
rect 18198 584 20000 640
rect 18137 582 20000 584
rect 18137 579 18203 582
rect 19200 552 20000 582
rect 0 234 800 264
rect 2773 234 2839 237
rect 0 232 2839 234
rect 0 176 2778 232
rect 2834 176 2839 232
rect 0 174 2839 176
rect 0 144 800 174
rect 2773 171 2839 174
rect 18873 234 18939 237
rect 19200 234 20000 264
rect 18873 232 20000 234
rect 18873 176 18878 232
rect 18934 176 20000 232
rect 18873 174 20000 176
rect 18873 171 18939 174
rect 19200 144 20000 174
<< via3 >>
rect 15516 15132 15580 15196
rect 17172 14724 17236 14788
rect 3176 14716 3240 14720
rect 3176 14660 3180 14716
rect 3180 14660 3236 14716
rect 3236 14660 3240 14716
rect 3176 14656 3240 14660
rect 3256 14716 3320 14720
rect 3256 14660 3260 14716
rect 3260 14660 3316 14716
rect 3316 14660 3320 14716
rect 3256 14656 3320 14660
rect 3336 14716 3400 14720
rect 3336 14660 3340 14716
rect 3340 14660 3396 14716
rect 3396 14660 3400 14716
rect 3336 14656 3400 14660
rect 3416 14716 3480 14720
rect 3416 14660 3420 14716
rect 3420 14660 3476 14716
rect 3476 14660 3480 14716
rect 3416 14656 3480 14660
rect 7624 14716 7688 14720
rect 7624 14660 7628 14716
rect 7628 14660 7684 14716
rect 7684 14660 7688 14716
rect 7624 14656 7688 14660
rect 7704 14716 7768 14720
rect 7704 14660 7708 14716
rect 7708 14660 7764 14716
rect 7764 14660 7768 14716
rect 7704 14656 7768 14660
rect 7784 14716 7848 14720
rect 7784 14660 7788 14716
rect 7788 14660 7844 14716
rect 7844 14660 7848 14716
rect 7784 14656 7848 14660
rect 7864 14716 7928 14720
rect 7864 14660 7868 14716
rect 7868 14660 7924 14716
rect 7924 14660 7928 14716
rect 7864 14656 7928 14660
rect 12072 14716 12136 14720
rect 12072 14660 12076 14716
rect 12076 14660 12132 14716
rect 12132 14660 12136 14716
rect 12072 14656 12136 14660
rect 12152 14716 12216 14720
rect 12152 14660 12156 14716
rect 12156 14660 12212 14716
rect 12212 14660 12216 14716
rect 12152 14656 12216 14660
rect 12232 14716 12296 14720
rect 12232 14660 12236 14716
rect 12236 14660 12292 14716
rect 12292 14660 12296 14716
rect 12232 14656 12296 14660
rect 12312 14716 12376 14720
rect 12312 14660 12316 14716
rect 12316 14660 12372 14716
rect 12372 14660 12376 14716
rect 12312 14656 12376 14660
rect 16520 14716 16584 14720
rect 16520 14660 16524 14716
rect 16524 14660 16580 14716
rect 16580 14660 16584 14716
rect 16520 14656 16584 14660
rect 16600 14716 16664 14720
rect 16600 14660 16604 14716
rect 16604 14660 16660 14716
rect 16660 14660 16664 14716
rect 16600 14656 16664 14660
rect 16680 14716 16744 14720
rect 16680 14660 16684 14716
rect 16684 14660 16740 14716
rect 16740 14660 16744 14716
rect 16680 14656 16744 14660
rect 16760 14716 16824 14720
rect 16760 14660 16764 14716
rect 16764 14660 16820 14716
rect 16820 14660 16824 14716
rect 16760 14656 16824 14660
rect 5400 14172 5464 14176
rect 5400 14116 5404 14172
rect 5404 14116 5460 14172
rect 5460 14116 5464 14172
rect 5400 14112 5464 14116
rect 5480 14172 5544 14176
rect 5480 14116 5484 14172
rect 5484 14116 5540 14172
rect 5540 14116 5544 14172
rect 5480 14112 5544 14116
rect 5560 14172 5624 14176
rect 5560 14116 5564 14172
rect 5564 14116 5620 14172
rect 5620 14116 5624 14172
rect 5560 14112 5624 14116
rect 5640 14172 5704 14176
rect 5640 14116 5644 14172
rect 5644 14116 5700 14172
rect 5700 14116 5704 14172
rect 5640 14112 5704 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 14296 14172 14360 14176
rect 14296 14116 14300 14172
rect 14300 14116 14356 14172
rect 14356 14116 14360 14172
rect 14296 14112 14360 14116
rect 14376 14172 14440 14176
rect 14376 14116 14380 14172
rect 14380 14116 14436 14172
rect 14436 14116 14440 14172
rect 14376 14112 14440 14116
rect 14456 14172 14520 14176
rect 14456 14116 14460 14172
rect 14460 14116 14516 14172
rect 14516 14116 14520 14172
rect 14456 14112 14520 14116
rect 14536 14172 14600 14176
rect 14536 14116 14540 14172
rect 14540 14116 14596 14172
rect 14596 14116 14600 14172
rect 14536 14112 14600 14116
rect 17172 14044 17236 14108
rect 16988 13968 17052 13972
rect 16988 13912 17038 13968
rect 17038 13912 17052 13968
rect 16988 13908 17052 13912
rect 3176 13628 3240 13632
rect 3176 13572 3180 13628
rect 3180 13572 3236 13628
rect 3236 13572 3240 13628
rect 3176 13568 3240 13572
rect 3256 13628 3320 13632
rect 3256 13572 3260 13628
rect 3260 13572 3316 13628
rect 3316 13572 3320 13628
rect 3256 13568 3320 13572
rect 3336 13628 3400 13632
rect 3336 13572 3340 13628
rect 3340 13572 3396 13628
rect 3396 13572 3400 13628
rect 3336 13568 3400 13572
rect 3416 13628 3480 13632
rect 3416 13572 3420 13628
rect 3420 13572 3476 13628
rect 3476 13572 3480 13628
rect 3416 13568 3480 13572
rect 7624 13628 7688 13632
rect 7624 13572 7628 13628
rect 7628 13572 7684 13628
rect 7684 13572 7688 13628
rect 7624 13568 7688 13572
rect 7704 13628 7768 13632
rect 7704 13572 7708 13628
rect 7708 13572 7764 13628
rect 7764 13572 7768 13628
rect 7704 13568 7768 13572
rect 7784 13628 7848 13632
rect 7784 13572 7788 13628
rect 7788 13572 7844 13628
rect 7844 13572 7848 13628
rect 7784 13568 7848 13572
rect 7864 13628 7928 13632
rect 7864 13572 7868 13628
rect 7868 13572 7924 13628
rect 7924 13572 7928 13628
rect 7864 13568 7928 13572
rect 12072 13628 12136 13632
rect 12072 13572 12076 13628
rect 12076 13572 12132 13628
rect 12132 13572 12136 13628
rect 12072 13568 12136 13572
rect 12152 13628 12216 13632
rect 12152 13572 12156 13628
rect 12156 13572 12212 13628
rect 12212 13572 12216 13628
rect 12152 13568 12216 13572
rect 12232 13628 12296 13632
rect 12232 13572 12236 13628
rect 12236 13572 12292 13628
rect 12292 13572 12296 13628
rect 12232 13568 12296 13572
rect 12312 13628 12376 13632
rect 12312 13572 12316 13628
rect 12316 13572 12372 13628
rect 12372 13572 12376 13628
rect 12312 13568 12376 13572
rect 16520 13628 16584 13632
rect 16520 13572 16524 13628
rect 16524 13572 16580 13628
rect 16580 13572 16584 13628
rect 16520 13568 16584 13572
rect 16600 13628 16664 13632
rect 16600 13572 16604 13628
rect 16604 13572 16660 13628
rect 16660 13572 16664 13628
rect 16600 13568 16664 13572
rect 16680 13628 16744 13632
rect 16680 13572 16684 13628
rect 16684 13572 16740 13628
rect 16740 13572 16744 13628
rect 16680 13568 16744 13572
rect 16760 13628 16824 13632
rect 16760 13572 16764 13628
rect 16764 13572 16820 13628
rect 16820 13572 16824 13628
rect 16760 13568 16824 13572
rect 5400 13084 5464 13088
rect 5400 13028 5404 13084
rect 5404 13028 5460 13084
rect 5460 13028 5464 13084
rect 5400 13024 5464 13028
rect 5480 13084 5544 13088
rect 5480 13028 5484 13084
rect 5484 13028 5540 13084
rect 5540 13028 5544 13084
rect 5480 13024 5544 13028
rect 5560 13084 5624 13088
rect 5560 13028 5564 13084
rect 5564 13028 5620 13084
rect 5620 13028 5624 13084
rect 5560 13024 5624 13028
rect 5640 13084 5704 13088
rect 5640 13028 5644 13084
rect 5644 13028 5700 13084
rect 5700 13028 5704 13084
rect 5640 13024 5704 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 14296 13084 14360 13088
rect 14296 13028 14300 13084
rect 14300 13028 14356 13084
rect 14356 13028 14360 13084
rect 14296 13024 14360 13028
rect 14376 13084 14440 13088
rect 14376 13028 14380 13084
rect 14380 13028 14436 13084
rect 14436 13028 14440 13084
rect 14376 13024 14440 13028
rect 14456 13084 14520 13088
rect 14456 13028 14460 13084
rect 14460 13028 14516 13084
rect 14516 13028 14520 13084
rect 14456 13024 14520 13028
rect 14536 13084 14600 13088
rect 14536 13028 14540 13084
rect 14540 13028 14596 13084
rect 14596 13028 14600 13084
rect 14536 13024 14600 13028
rect 8524 12684 8588 12748
rect 1900 12548 1964 12612
rect 3176 12540 3240 12544
rect 3176 12484 3180 12540
rect 3180 12484 3236 12540
rect 3236 12484 3240 12540
rect 3176 12480 3240 12484
rect 3256 12540 3320 12544
rect 3256 12484 3260 12540
rect 3260 12484 3316 12540
rect 3316 12484 3320 12540
rect 3256 12480 3320 12484
rect 3336 12540 3400 12544
rect 3336 12484 3340 12540
rect 3340 12484 3396 12540
rect 3396 12484 3400 12540
rect 3336 12480 3400 12484
rect 3416 12540 3480 12544
rect 3416 12484 3420 12540
rect 3420 12484 3476 12540
rect 3476 12484 3480 12540
rect 3416 12480 3480 12484
rect 7624 12540 7688 12544
rect 7624 12484 7628 12540
rect 7628 12484 7684 12540
rect 7684 12484 7688 12540
rect 7624 12480 7688 12484
rect 7704 12540 7768 12544
rect 7704 12484 7708 12540
rect 7708 12484 7764 12540
rect 7764 12484 7768 12540
rect 7704 12480 7768 12484
rect 7784 12540 7848 12544
rect 7784 12484 7788 12540
rect 7788 12484 7844 12540
rect 7844 12484 7848 12540
rect 7784 12480 7848 12484
rect 7864 12540 7928 12544
rect 7864 12484 7868 12540
rect 7868 12484 7924 12540
rect 7924 12484 7928 12540
rect 7864 12480 7928 12484
rect 12072 12540 12136 12544
rect 12072 12484 12076 12540
rect 12076 12484 12132 12540
rect 12132 12484 12136 12540
rect 12072 12480 12136 12484
rect 12152 12540 12216 12544
rect 12152 12484 12156 12540
rect 12156 12484 12212 12540
rect 12212 12484 12216 12540
rect 12152 12480 12216 12484
rect 12232 12540 12296 12544
rect 12232 12484 12236 12540
rect 12236 12484 12292 12540
rect 12292 12484 12296 12540
rect 12232 12480 12296 12484
rect 12312 12540 12376 12544
rect 12312 12484 12316 12540
rect 12316 12484 12372 12540
rect 12372 12484 12376 12540
rect 12312 12480 12376 12484
rect 16520 12540 16584 12544
rect 16520 12484 16524 12540
rect 16524 12484 16580 12540
rect 16580 12484 16584 12540
rect 16520 12480 16584 12484
rect 16600 12540 16664 12544
rect 16600 12484 16604 12540
rect 16604 12484 16660 12540
rect 16660 12484 16664 12540
rect 16600 12480 16664 12484
rect 16680 12540 16744 12544
rect 16680 12484 16684 12540
rect 16684 12484 16740 12540
rect 16740 12484 16744 12540
rect 16680 12480 16744 12484
rect 16760 12540 16824 12544
rect 16760 12484 16764 12540
rect 16764 12484 16820 12540
rect 16820 12484 16824 12540
rect 16760 12480 16824 12484
rect 2452 12412 2516 12476
rect 16068 12140 16132 12204
rect 5400 11996 5464 12000
rect 5400 11940 5404 11996
rect 5404 11940 5460 11996
rect 5460 11940 5464 11996
rect 5400 11936 5464 11940
rect 5480 11996 5544 12000
rect 5480 11940 5484 11996
rect 5484 11940 5540 11996
rect 5540 11940 5544 11996
rect 5480 11936 5544 11940
rect 5560 11996 5624 12000
rect 5560 11940 5564 11996
rect 5564 11940 5620 11996
rect 5620 11940 5624 11996
rect 5560 11936 5624 11940
rect 5640 11996 5704 12000
rect 5640 11940 5644 11996
rect 5644 11940 5700 11996
rect 5700 11940 5704 11996
rect 5640 11936 5704 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 14296 11996 14360 12000
rect 14296 11940 14300 11996
rect 14300 11940 14356 11996
rect 14356 11940 14360 11996
rect 14296 11936 14360 11940
rect 14376 11996 14440 12000
rect 14376 11940 14380 11996
rect 14380 11940 14436 11996
rect 14436 11940 14440 11996
rect 14376 11936 14440 11940
rect 14456 11996 14520 12000
rect 14456 11940 14460 11996
rect 14460 11940 14516 11996
rect 14516 11940 14520 11996
rect 14456 11936 14520 11940
rect 14536 11996 14600 12000
rect 14536 11940 14540 11996
rect 14540 11940 14596 11996
rect 14596 11940 14600 11996
rect 14536 11936 14600 11940
rect 4108 11928 4172 11932
rect 4108 11872 4122 11928
rect 4122 11872 4172 11928
rect 4108 11868 4172 11872
rect 16252 11732 16316 11796
rect 3176 11452 3240 11456
rect 3176 11396 3180 11452
rect 3180 11396 3236 11452
rect 3236 11396 3240 11452
rect 3176 11392 3240 11396
rect 3256 11452 3320 11456
rect 3256 11396 3260 11452
rect 3260 11396 3316 11452
rect 3316 11396 3320 11452
rect 3256 11392 3320 11396
rect 3336 11452 3400 11456
rect 3336 11396 3340 11452
rect 3340 11396 3396 11452
rect 3396 11396 3400 11452
rect 3336 11392 3400 11396
rect 3416 11452 3480 11456
rect 3416 11396 3420 11452
rect 3420 11396 3476 11452
rect 3476 11396 3480 11452
rect 3416 11392 3480 11396
rect 7624 11452 7688 11456
rect 7624 11396 7628 11452
rect 7628 11396 7684 11452
rect 7684 11396 7688 11452
rect 7624 11392 7688 11396
rect 7704 11452 7768 11456
rect 7704 11396 7708 11452
rect 7708 11396 7764 11452
rect 7764 11396 7768 11452
rect 7704 11392 7768 11396
rect 7784 11452 7848 11456
rect 7784 11396 7788 11452
rect 7788 11396 7844 11452
rect 7844 11396 7848 11452
rect 7784 11392 7848 11396
rect 7864 11452 7928 11456
rect 7864 11396 7868 11452
rect 7868 11396 7924 11452
rect 7924 11396 7928 11452
rect 7864 11392 7928 11396
rect 12072 11452 12136 11456
rect 12072 11396 12076 11452
rect 12076 11396 12132 11452
rect 12132 11396 12136 11452
rect 12072 11392 12136 11396
rect 12152 11452 12216 11456
rect 12152 11396 12156 11452
rect 12156 11396 12212 11452
rect 12212 11396 12216 11452
rect 12152 11392 12216 11396
rect 12232 11452 12296 11456
rect 12232 11396 12236 11452
rect 12236 11396 12292 11452
rect 12292 11396 12296 11452
rect 12232 11392 12296 11396
rect 12312 11452 12376 11456
rect 12312 11396 12316 11452
rect 12316 11396 12372 11452
rect 12372 11396 12376 11452
rect 12312 11392 12376 11396
rect 16520 11452 16584 11456
rect 16520 11396 16524 11452
rect 16524 11396 16580 11452
rect 16580 11396 16584 11452
rect 16520 11392 16584 11396
rect 16600 11452 16664 11456
rect 16600 11396 16604 11452
rect 16604 11396 16660 11452
rect 16660 11396 16664 11452
rect 16600 11392 16664 11396
rect 16680 11452 16744 11456
rect 16680 11396 16684 11452
rect 16684 11396 16740 11452
rect 16740 11396 16744 11452
rect 16680 11392 16744 11396
rect 16760 11452 16824 11456
rect 16760 11396 16764 11452
rect 16764 11396 16820 11452
rect 16820 11396 16824 11452
rect 16760 11392 16824 11396
rect 15148 11188 15212 11252
rect 1716 10840 1780 10844
rect 1716 10784 1766 10840
rect 1766 10784 1780 10840
rect 1716 10780 1780 10784
rect 16068 11052 16132 11116
rect 5400 10908 5464 10912
rect 5400 10852 5404 10908
rect 5404 10852 5460 10908
rect 5460 10852 5464 10908
rect 5400 10848 5464 10852
rect 5480 10908 5544 10912
rect 5480 10852 5484 10908
rect 5484 10852 5540 10908
rect 5540 10852 5544 10908
rect 5480 10848 5544 10852
rect 5560 10908 5624 10912
rect 5560 10852 5564 10908
rect 5564 10852 5620 10908
rect 5620 10852 5624 10908
rect 5560 10848 5624 10852
rect 5640 10908 5704 10912
rect 5640 10852 5644 10908
rect 5644 10852 5700 10908
rect 5700 10852 5704 10908
rect 5640 10848 5704 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 14296 10908 14360 10912
rect 14296 10852 14300 10908
rect 14300 10852 14356 10908
rect 14356 10852 14360 10908
rect 14296 10848 14360 10852
rect 14376 10908 14440 10912
rect 14376 10852 14380 10908
rect 14380 10852 14436 10908
rect 14436 10852 14440 10908
rect 14376 10848 14440 10852
rect 14456 10908 14520 10912
rect 14456 10852 14460 10908
rect 14460 10852 14516 10908
rect 14516 10852 14520 10908
rect 14456 10848 14520 10852
rect 14536 10908 14600 10912
rect 14536 10852 14540 10908
rect 14540 10852 14596 10908
rect 14596 10852 14600 10908
rect 14536 10848 14600 10852
rect 3176 10364 3240 10368
rect 3176 10308 3180 10364
rect 3180 10308 3236 10364
rect 3236 10308 3240 10364
rect 3176 10304 3240 10308
rect 3256 10364 3320 10368
rect 3256 10308 3260 10364
rect 3260 10308 3316 10364
rect 3316 10308 3320 10364
rect 3256 10304 3320 10308
rect 3336 10364 3400 10368
rect 3336 10308 3340 10364
rect 3340 10308 3396 10364
rect 3396 10308 3400 10364
rect 3336 10304 3400 10308
rect 3416 10364 3480 10368
rect 3416 10308 3420 10364
rect 3420 10308 3476 10364
rect 3476 10308 3480 10364
rect 3416 10304 3480 10308
rect 7624 10364 7688 10368
rect 7624 10308 7628 10364
rect 7628 10308 7684 10364
rect 7684 10308 7688 10364
rect 7624 10304 7688 10308
rect 7704 10364 7768 10368
rect 7704 10308 7708 10364
rect 7708 10308 7764 10364
rect 7764 10308 7768 10364
rect 7704 10304 7768 10308
rect 7784 10364 7848 10368
rect 7784 10308 7788 10364
rect 7788 10308 7844 10364
rect 7844 10308 7848 10364
rect 7784 10304 7848 10308
rect 7864 10364 7928 10368
rect 7864 10308 7868 10364
rect 7868 10308 7924 10364
rect 7924 10308 7928 10364
rect 7864 10304 7928 10308
rect 12072 10364 12136 10368
rect 12072 10308 12076 10364
rect 12076 10308 12132 10364
rect 12132 10308 12136 10364
rect 12072 10304 12136 10308
rect 12152 10364 12216 10368
rect 12152 10308 12156 10364
rect 12156 10308 12212 10364
rect 12212 10308 12216 10364
rect 12152 10304 12216 10308
rect 12232 10364 12296 10368
rect 12232 10308 12236 10364
rect 12236 10308 12292 10364
rect 12292 10308 12296 10364
rect 12232 10304 12296 10308
rect 12312 10364 12376 10368
rect 12312 10308 12316 10364
rect 12316 10308 12372 10364
rect 12372 10308 12376 10364
rect 12312 10304 12376 10308
rect 16520 10364 16584 10368
rect 16520 10308 16524 10364
rect 16524 10308 16580 10364
rect 16580 10308 16584 10364
rect 16520 10304 16584 10308
rect 16600 10364 16664 10368
rect 16600 10308 16604 10364
rect 16604 10308 16660 10364
rect 16660 10308 16664 10364
rect 16600 10304 16664 10308
rect 16680 10364 16744 10368
rect 16680 10308 16684 10364
rect 16684 10308 16740 10364
rect 16740 10308 16744 10364
rect 16680 10304 16744 10308
rect 16760 10364 16824 10368
rect 16760 10308 16764 10364
rect 16764 10308 16820 10364
rect 16820 10308 16824 10364
rect 16760 10304 16824 10308
rect 8524 10100 8588 10164
rect 5400 9820 5464 9824
rect 5400 9764 5404 9820
rect 5404 9764 5460 9820
rect 5460 9764 5464 9820
rect 5400 9760 5464 9764
rect 5480 9820 5544 9824
rect 5480 9764 5484 9820
rect 5484 9764 5540 9820
rect 5540 9764 5544 9820
rect 5480 9760 5544 9764
rect 5560 9820 5624 9824
rect 5560 9764 5564 9820
rect 5564 9764 5620 9820
rect 5620 9764 5624 9820
rect 5560 9760 5624 9764
rect 5640 9820 5704 9824
rect 5640 9764 5644 9820
rect 5644 9764 5700 9820
rect 5700 9764 5704 9820
rect 5640 9760 5704 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 14296 9820 14360 9824
rect 14296 9764 14300 9820
rect 14300 9764 14356 9820
rect 14356 9764 14360 9820
rect 14296 9760 14360 9764
rect 14376 9820 14440 9824
rect 14376 9764 14380 9820
rect 14380 9764 14436 9820
rect 14436 9764 14440 9820
rect 14376 9760 14440 9764
rect 14456 9820 14520 9824
rect 14456 9764 14460 9820
rect 14460 9764 14516 9820
rect 14516 9764 14520 9820
rect 14456 9760 14520 9764
rect 14536 9820 14600 9824
rect 14536 9764 14540 9820
rect 14540 9764 14596 9820
rect 14596 9764 14600 9820
rect 14536 9760 14600 9764
rect 13124 9692 13188 9756
rect 5212 9344 5276 9348
rect 5212 9288 5226 9344
rect 5226 9288 5276 9344
rect 5212 9284 5276 9288
rect 7236 9344 7300 9348
rect 7236 9288 7286 9344
rect 7286 9288 7300 9344
rect 7236 9284 7300 9288
rect 3176 9276 3240 9280
rect 3176 9220 3180 9276
rect 3180 9220 3236 9276
rect 3236 9220 3240 9276
rect 3176 9216 3240 9220
rect 3256 9276 3320 9280
rect 3256 9220 3260 9276
rect 3260 9220 3316 9276
rect 3316 9220 3320 9276
rect 3256 9216 3320 9220
rect 3336 9276 3400 9280
rect 3336 9220 3340 9276
rect 3340 9220 3396 9276
rect 3396 9220 3400 9276
rect 3336 9216 3400 9220
rect 3416 9276 3480 9280
rect 3416 9220 3420 9276
rect 3420 9220 3476 9276
rect 3476 9220 3480 9276
rect 3416 9216 3480 9220
rect 7624 9276 7688 9280
rect 7624 9220 7628 9276
rect 7628 9220 7684 9276
rect 7684 9220 7688 9276
rect 7624 9216 7688 9220
rect 7704 9276 7768 9280
rect 7704 9220 7708 9276
rect 7708 9220 7764 9276
rect 7764 9220 7768 9276
rect 7704 9216 7768 9220
rect 7784 9276 7848 9280
rect 7784 9220 7788 9276
rect 7788 9220 7844 9276
rect 7844 9220 7848 9276
rect 7784 9216 7848 9220
rect 7864 9276 7928 9280
rect 7864 9220 7868 9276
rect 7868 9220 7924 9276
rect 7924 9220 7928 9276
rect 7864 9216 7928 9220
rect 12072 9276 12136 9280
rect 12072 9220 12076 9276
rect 12076 9220 12132 9276
rect 12132 9220 12136 9276
rect 12072 9216 12136 9220
rect 12152 9276 12216 9280
rect 12152 9220 12156 9276
rect 12156 9220 12212 9276
rect 12212 9220 12216 9276
rect 12152 9216 12216 9220
rect 12232 9276 12296 9280
rect 12232 9220 12236 9276
rect 12236 9220 12292 9276
rect 12292 9220 12296 9276
rect 12232 9216 12296 9220
rect 12312 9276 12376 9280
rect 12312 9220 12316 9276
rect 12316 9220 12372 9276
rect 12372 9220 12376 9276
rect 12312 9216 12376 9220
rect 16520 9276 16584 9280
rect 16520 9220 16524 9276
rect 16524 9220 16580 9276
rect 16580 9220 16584 9276
rect 16520 9216 16584 9220
rect 16600 9276 16664 9280
rect 16600 9220 16604 9276
rect 16604 9220 16660 9276
rect 16660 9220 16664 9276
rect 16600 9216 16664 9220
rect 16680 9276 16744 9280
rect 16680 9220 16684 9276
rect 16684 9220 16740 9276
rect 16740 9220 16744 9276
rect 16680 9216 16744 9220
rect 16760 9276 16824 9280
rect 16760 9220 16764 9276
rect 16764 9220 16820 9276
rect 16820 9220 16824 9276
rect 16760 9216 16824 9220
rect 7236 8740 7300 8804
rect 5400 8732 5464 8736
rect 5400 8676 5404 8732
rect 5404 8676 5460 8732
rect 5460 8676 5464 8732
rect 5400 8672 5464 8676
rect 5480 8732 5544 8736
rect 5480 8676 5484 8732
rect 5484 8676 5540 8732
rect 5540 8676 5544 8732
rect 5480 8672 5544 8676
rect 5560 8732 5624 8736
rect 5560 8676 5564 8732
rect 5564 8676 5620 8732
rect 5620 8676 5624 8732
rect 5560 8672 5624 8676
rect 5640 8732 5704 8736
rect 5640 8676 5644 8732
rect 5644 8676 5700 8732
rect 5700 8676 5704 8732
rect 5640 8672 5704 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 14296 8732 14360 8736
rect 14296 8676 14300 8732
rect 14300 8676 14356 8732
rect 14356 8676 14360 8732
rect 14296 8672 14360 8676
rect 14376 8732 14440 8736
rect 14376 8676 14380 8732
rect 14380 8676 14436 8732
rect 14436 8676 14440 8732
rect 14376 8672 14440 8676
rect 14456 8732 14520 8736
rect 14456 8676 14460 8732
rect 14460 8676 14516 8732
rect 14516 8676 14520 8732
rect 14456 8672 14520 8676
rect 14536 8732 14600 8736
rect 14536 8676 14540 8732
rect 14540 8676 14596 8732
rect 14596 8676 14600 8732
rect 14536 8672 14600 8676
rect 2820 8604 2884 8668
rect 4476 8468 4540 8532
rect 2452 8332 2516 8396
rect 3176 8188 3240 8192
rect 3176 8132 3180 8188
rect 3180 8132 3236 8188
rect 3236 8132 3240 8188
rect 3176 8128 3240 8132
rect 3256 8188 3320 8192
rect 3256 8132 3260 8188
rect 3260 8132 3316 8188
rect 3316 8132 3320 8188
rect 3256 8128 3320 8132
rect 3336 8188 3400 8192
rect 3336 8132 3340 8188
rect 3340 8132 3396 8188
rect 3396 8132 3400 8188
rect 3336 8128 3400 8132
rect 3416 8188 3480 8192
rect 3416 8132 3420 8188
rect 3420 8132 3476 8188
rect 3476 8132 3480 8188
rect 3416 8128 3480 8132
rect 7624 8188 7688 8192
rect 7624 8132 7628 8188
rect 7628 8132 7684 8188
rect 7684 8132 7688 8188
rect 7624 8128 7688 8132
rect 7704 8188 7768 8192
rect 7704 8132 7708 8188
rect 7708 8132 7764 8188
rect 7764 8132 7768 8188
rect 7704 8128 7768 8132
rect 7784 8188 7848 8192
rect 7784 8132 7788 8188
rect 7788 8132 7844 8188
rect 7844 8132 7848 8188
rect 7784 8128 7848 8132
rect 7864 8188 7928 8192
rect 7864 8132 7868 8188
rect 7868 8132 7924 8188
rect 7924 8132 7928 8188
rect 7864 8128 7928 8132
rect 12072 8188 12136 8192
rect 12072 8132 12076 8188
rect 12076 8132 12132 8188
rect 12132 8132 12136 8188
rect 12072 8128 12136 8132
rect 12152 8188 12216 8192
rect 12152 8132 12156 8188
rect 12156 8132 12212 8188
rect 12212 8132 12216 8188
rect 12152 8128 12216 8132
rect 12232 8188 12296 8192
rect 12232 8132 12236 8188
rect 12236 8132 12292 8188
rect 12292 8132 12296 8188
rect 12232 8128 12296 8132
rect 12312 8188 12376 8192
rect 12312 8132 12316 8188
rect 12316 8132 12372 8188
rect 12372 8132 12376 8188
rect 12312 8128 12376 8132
rect 16520 8188 16584 8192
rect 16520 8132 16524 8188
rect 16524 8132 16580 8188
rect 16580 8132 16584 8188
rect 16520 8128 16584 8132
rect 16600 8188 16664 8192
rect 16600 8132 16604 8188
rect 16604 8132 16660 8188
rect 16660 8132 16664 8188
rect 16600 8128 16664 8132
rect 16680 8188 16744 8192
rect 16680 8132 16684 8188
rect 16684 8132 16740 8188
rect 16740 8132 16744 8188
rect 16680 8128 16744 8132
rect 16760 8188 16824 8192
rect 16760 8132 16764 8188
rect 16764 8132 16820 8188
rect 16820 8132 16824 8188
rect 16760 8128 16824 8132
rect 2636 7652 2700 7716
rect 5400 7644 5464 7648
rect 5400 7588 5404 7644
rect 5404 7588 5460 7644
rect 5460 7588 5464 7644
rect 5400 7584 5464 7588
rect 5480 7644 5544 7648
rect 5480 7588 5484 7644
rect 5484 7588 5540 7644
rect 5540 7588 5544 7644
rect 5480 7584 5544 7588
rect 5560 7644 5624 7648
rect 5560 7588 5564 7644
rect 5564 7588 5620 7644
rect 5620 7588 5624 7644
rect 5560 7584 5624 7588
rect 5640 7644 5704 7648
rect 5640 7588 5644 7644
rect 5644 7588 5700 7644
rect 5700 7588 5704 7644
rect 5640 7584 5704 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 14296 7644 14360 7648
rect 14296 7588 14300 7644
rect 14300 7588 14356 7644
rect 14356 7588 14360 7644
rect 14296 7584 14360 7588
rect 14376 7644 14440 7648
rect 14376 7588 14380 7644
rect 14380 7588 14436 7644
rect 14436 7588 14440 7644
rect 14376 7584 14440 7588
rect 14456 7644 14520 7648
rect 14456 7588 14460 7644
rect 14460 7588 14516 7644
rect 14516 7588 14520 7644
rect 14456 7584 14520 7588
rect 14536 7644 14600 7648
rect 14536 7588 14540 7644
rect 14540 7588 14596 7644
rect 14596 7588 14600 7644
rect 14536 7584 14600 7588
rect 1716 7440 1780 7444
rect 1716 7384 1730 7440
rect 1730 7384 1780 7440
rect 1716 7380 1780 7384
rect 3176 7100 3240 7104
rect 3176 7044 3180 7100
rect 3180 7044 3236 7100
rect 3236 7044 3240 7100
rect 3176 7040 3240 7044
rect 3256 7100 3320 7104
rect 3256 7044 3260 7100
rect 3260 7044 3316 7100
rect 3316 7044 3320 7100
rect 3256 7040 3320 7044
rect 3336 7100 3400 7104
rect 3336 7044 3340 7100
rect 3340 7044 3396 7100
rect 3396 7044 3400 7100
rect 3336 7040 3400 7044
rect 3416 7100 3480 7104
rect 3416 7044 3420 7100
rect 3420 7044 3476 7100
rect 3476 7044 3480 7100
rect 3416 7040 3480 7044
rect 7624 7100 7688 7104
rect 7624 7044 7628 7100
rect 7628 7044 7684 7100
rect 7684 7044 7688 7100
rect 7624 7040 7688 7044
rect 7704 7100 7768 7104
rect 7704 7044 7708 7100
rect 7708 7044 7764 7100
rect 7764 7044 7768 7100
rect 7704 7040 7768 7044
rect 7784 7100 7848 7104
rect 7784 7044 7788 7100
rect 7788 7044 7844 7100
rect 7844 7044 7848 7100
rect 7784 7040 7848 7044
rect 7864 7100 7928 7104
rect 7864 7044 7868 7100
rect 7868 7044 7924 7100
rect 7924 7044 7928 7100
rect 7864 7040 7928 7044
rect 12072 7100 12136 7104
rect 12072 7044 12076 7100
rect 12076 7044 12132 7100
rect 12132 7044 12136 7100
rect 12072 7040 12136 7044
rect 12152 7100 12216 7104
rect 12152 7044 12156 7100
rect 12156 7044 12212 7100
rect 12212 7044 12216 7100
rect 12152 7040 12216 7044
rect 12232 7100 12296 7104
rect 12232 7044 12236 7100
rect 12236 7044 12292 7100
rect 12292 7044 12296 7100
rect 12232 7040 12296 7044
rect 12312 7100 12376 7104
rect 12312 7044 12316 7100
rect 12316 7044 12372 7100
rect 12372 7044 12376 7100
rect 12312 7040 12376 7044
rect 16520 7100 16584 7104
rect 16520 7044 16524 7100
rect 16524 7044 16580 7100
rect 16580 7044 16584 7100
rect 16520 7040 16584 7044
rect 16600 7100 16664 7104
rect 16600 7044 16604 7100
rect 16604 7044 16660 7100
rect 16660 7044 16664 7100
rect 16600 7040 16664 7044
rect 16680 7100 16744 7104
rect 16680 7044 16684 7100
rect 16684 7044 16740 7100
rect 16740 7044 16744 7100
rect 16680 7040 16744 7044
rect 16760 7100 16824 7104
rect 16760 7044 16764 7100
rect 16764 7044 16820 7100
rect 16820 7044 16824 7100
rect 16760 7040 16824 7044
rect 4108 6836 4172 6900
rect 8524 6836 8588 6900
rect 15516 6836 15580 6900
rect 6868 6760 6932 6764
rect 6868 6704 6918 6760
rect 6918 6704 6932 6760
rect 6868 6700 6932 6704
rect 7236 6564 7300 6628
rect 5400 6556 5464 6560
rect 5400 6500 5404 6556
rect 5404 6500 5460 6556
rect 5460 6500 5464 6556
rect 5400 6496 5464 6500
rect 5480 6556 5544 6560
rect 5480 6500 5484 6556
rect 5484 6500 5540 6556
rect 5540 6500 5544 6556
rect 5480 6496 5544 6500
rect 5560 6556 5624 6560
rect 5560 6500 5564 6556
rect 5564 6500 5620 6556
rect 5620 6500 5624 6556
rect 5560 6496 5624 6500
rect 5640 6556 5704 6560
rect 5640 6500 5644 6556
rect 5644 6500 5700 6556
rect 5700 6500 5704 6556
rect 5640 6496 5704 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 14296 6556 14360 6560
rect 14296 6500 14300 6556
rect 14300 6500 14356 6556
rect 14356 6500 14360 6556
rect 14296 6496 14360 6500
rect 14376 6556 14440 6560
rect 14376 6500 14380 6556
rect 14380 6500 14436 6556
rect 14436 6500 14440 6556
rect 14376 6496 14440 6500
rect 14456 6556 14520 6560
rect 14456 6500 14460 6556
rect 14460 6500 14516 6556
rect 14516 6500 14520 6556
rect 14456 6496 14520 6500
rect 14536 6556 14600 6560
rect 14536 6500 14540 6556
rect 14540 6500 14596 6556
rect 14596 6500 14600 6556
rect 14536 6496 14600 6500
rect 2452 6488 2516 6492
rect 2452 6432 2466 6488
rect 2466 6432 2516 6488
rect 2452 6428 2516 6432
rect 7236 6292 7300 6356
rect 10916 6156 10980 6220
rect 3176 6012 3240 6016
rect 3176 5956 3180 6012
rect 3180 5956 3236 6012
rect 3236 5956 3240 6012
rect 3176 5952 3240 5956
rect 3256 6012 3320 6016
rect 3256 5956 3260 6012
rect 3260 5956 3316 6012
rect 3316 5956 3320 6012
rect 3256 5952 3320 5956
rect 3336 6012 3400 6016
rect 3336 5956 3340 6012
rect 3340 5956 3396 6012
rect 3396 5956 3400 6012
rect 3336 5952 3400 5956
rect 3416 6012 3480 6016
rect 3416 5956 3420 6012
rect 3420 5956 3476 6012
rect 3476 5956 3480 6012
rect 3416 5952 3480 5956
rect 7624 6012 7688 6016
rect 7624 5956 7628 6012
rect 7628 5956 7684 6012
rect 7684 5956 7688 6012
rect 7624 5952 7688 5956
rect 7704 6012 7768 6016
rect 7704 5956 7708 6012
rect 7708 5956 7764 6012
rect 7764 5956 7768 6012
rect 7704 5952 7768 5956
rect 7784 6012 7848 6016
rect 7784 5956 7788 6012
rect 7788 5956 7844 6012
rect 7844 5956 7848 6012
rect 7784 5952 7848 5956
rect 7864 6012 7928 6016
rect 7864 5956 7868 6012
rect 7868 5956 7924 6012
rect 7924 5956 7928 6012
rect 7864 5952 7928 5956
rect 12072 6012 12136 6016
rect 12072 5956 12076 6012
rect 12076 5956 12132 6012
rect 12132 5956 12136 6012
rect 12072 5952 12136 5956
rect 12152 6012 12216 6016
rect 12152 5956 12156 6012
rect 12156 5956 12212 6012
rect 12212 5956 12216 6012
rect 12152 5952 12216 5956
rect 12232 6012 12296 6016
rect 12232 5956 12236 6012
rect 12236 5956 12292 6012
rect 12292 5956 12296 6012
rect 12232 5952 12296 5956
rect 12312 6012 12376 6016
rect 12312 5956 12316 6012
rect 12316 5956 12372 6012
rect 12372 5956 12376 6012
rect 12312 5952 12376 5956
rect 16520 6012 16584 6016
rect 16520 5956 16524 6012
rect 16524 5956 16580 6012
rect 16580 5956 16584 6012
rect 16520 5952 16584 5956
rect 16600 6012 16664 6016
rect 16600 5956 16604 6012
rect 16604 5956 16660 6012
rect 16660 5956 16664 6012
rect 16600 5952 16664 5956
rect 16680 6012 16744 6016
rect 16680 5956 16684 6012
rect 16684 5956 16740 6012
rect 16740 5956 16744 6012
rect 16680 5952 16744 5956
rect 16760 6012 16824 6016
rect 16760 5956 16764 6012
rect 16764 5956 16820 6012
rect 16820 5956 16824 6012
rect 16760 5952 16824 5956
rect 4660 5612 4724 5676
rect 8340 5612 8404 5676
rect 15516 5748 15580 5812
rect 16068 5476 16132 5540
rect 5400 5468 5464 5472
rect 5400 5412 5404 5468
rect 5404 5412 5460 5468
rect 5460 5412 5464 5468
rect 5400 5408 5464 5412
rect 5480 5468 5544 5472
rect 5480 5412 5484 5468
rect 5484 5412 5540 5468
rect 5540 5412 5544 5468
rect 5480 5408 5544 5412
rect 5560 5468 5624 5472
rect 5560 5412 5564 5468
rect 5564 5412 5620 5468
rect 5620 5412 5624 5468
rect 5560 5408 5624 5412
rect 5640 5468 5704 5472
rect 5640 5412 5644 5468
rect 5644 5412 5700 5468
rect 5700 5412 5704 5468
rect 5640 5408 5704 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 14296 5468 14360 5472
rect 14296 5412 14300 5468
rect 14300 5412 14356 5468
rect 14356 5412 14360 5468
rect 14296 5408 14360 5412
rect 14376 5468 14440 5472
rect 14376 5412 14380 5468
rect 14380 5412 14436 5468
rect 14436 5412 14440 5468
rect 14376 5408 14440 5412
rect 14456 5468 14520 5472
rect 14456 5412 14460 5468
rect 14460 5412 14516 5468
rect 14516 5412 14520 5468
rect 14456 5408 14520 5412
rect 14536 5468 14600 5472
rect 14536 5412 14540 5468
rect 14540 5412 14596 5468
rect 14596 5412 14600 5468
rect 14536 5408 14600 5412
rect 17172 5340 17236 5404
rect 3176 4924 3240 4928
rect 3176 4868 3180 4924
rect 3180 4868 3236 4924
rect 3236 4868 3240 4924
rect 3176 4864 3240 4868
rect 3256 4924 3320 4928
rect 3256 4868 3260 4924
rect 3260 4868 3316 4924
rect 3316 4868 3320 4924
rect 3256 4864 3320 4868
rect 3336 4924 3400 4928
rect 3336 4868 3340 4924
rect 3340 4868 3396 4924
rect 3396 4868 3400 4924
rect 3336 4864 3400 4868
rect 3416 4924 3480 4928
rect 3416 4868 3420 4924
rect 3420 4868 3476 4924
rect 3476 4868 3480 4924
rect 3416 4864 3480 4868
rect 7624 4924 7688 4928
rect 7624 4868 7628 4924
rect 7628 4868 7684 4924
rect 7684 4868 7688 4924
rect 7624 4864 7688 4868
rect 7704 4924 7768 4928
rect 7704 4868 7708 4924
rect 7708 4868 7764 4924
rect 7764 4868 7768 4924
rect 7704 4864 7768 4868
rect 7784 4924 7848 4928
rect 7784 4868 7788 4924
rect 7788 4868 7844 4924
rect 7844 4868 7848 4924
rect 7784 4864 7848 4868
rect 7864 4924 7928 4928
rect 7864 4868 7868 4924
rect 7868 4868 7924 4924
rect 7924 4868 7928 4924
rect 7864 4864 7928 4868
rect 12072 4924 12136 4928
rect 12072 4868 12076 4924
rect 12076 4868 12132 4924
rect 12132 4868 12136 4924
rect 12072 4864 12136 4868
rect 12152 4924 12216 4928
rect 12152 4868 12156 4924
rect 12156 4868 12212 4924
rect 12212 4868 12216 4924
rect 12152 4864 12216 4868
rect 12232 4924 12296 4928
rect 12232 4868 12236 4924
rect 12236 4868 12292 4924
rect 12292 4868 12296 4924
rect 12232 4864 12296 4868
rect 12312 4924 12376 4928
rect 12312 4868 12316 4924
rect 12316 4868 12372 4924
rect 12372 4868 12376 4924
rect 12312 4864 12376 4868
rect 16520 4924 16584 4928
rect 16520 4868 16524 4924
rect 16524 4868 16580 4924
rect 16580 4868 16584 4924
rect 16520 4864 16584 4868
rect 16600 4924 16664 4928
rect 16600 4868 16604 4924
rect 16604 4868 16660 4924
rect 16660 4868 16664 4924
rect 16600 4864 16664 4868
rect 16680 4924 16744 4928
rect 16680 4868 16684 4924
rect 16684 4868 16740 4924
rect 16740 4868 16744 4924
rect 16680 4864 16744 4868
rect 16760 4924 16824 4928
rect 16760 4868 16764 4924
rect 16764 4868 16820 4924
rect 16820 4868 16824 4924
rect 16760 4864 16824 4868
rect 4108 4796 4172 4860
rect 16252 4856 16316 4860
rect 16252 4800 16302 4856
rect 16302 4800 16316 4856
rect 16252 4796 16316 4800
rect 5400 4380 5464 4384
rect 5400 4324 5404 4380
rect 5404 4324 5460 4380
rect 5460 4324 5464 4380
rect 5400 4320 5464 4324
rect 5480 4380 5544 4384
rect 5480 4324 5484 4380
rect 5484 4324 5540 4380
rect 5540 4324 5544 4380
rect 5480 4320 5544 4324
rect 5560 4380 5624 4384
rect 5560 4324 5564 4380
rect 5564 4324 5620 4380
rect 5620 4324 5624 4380
rect 5560 4320 5624 4324
rect 5640 4380 5704 4384
rect 5640 4324 5644 4380
rect 5644 4324 5700 4380
rect 5700 4324 5704 4380
rect 5640 4320 5704 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 14296 4380 14360 4384
rect 14296 4324 14300 4380
rect 14300 4324 14356 4380
rect 14356 4324 14360 4380
rect 14296 4320 14360 4324
rect 14376 4380 14440 4384
rect 14376 4324 14380 4380
rect 14380 4324 14436 4380
rect 14436 4324 14440 4380
rect 14376 4320 14440 4324
rect 14456 4380 14520 4384
rect 14456 4324 14460 4380
rect 14460 4324 14516 4380
rect 14516 4324 14520 4380
rect 14456 4320 14520 4324
rect 14536 4380 14600 4384
rect 14536 4324 14540 4380
rect 14540 4324 14596 4380
rect 14596 4324 14600 4380
rect 14536 4320 14600 4324
rect 15148 4116 15212 4180
rect 1716 4040 1780 4044
rect 1716 3984 1730 4040
rect 1730 3984 1780 4040
rect 1716 3980 1780 3984
rect 2636 3980 2700 4044
rect 4660 3980 4724 4044
rect 8524 4040 8588 4044
rect 8524 3984 8574 4040
rect 8574 3984 8588 4040
rect 8524 3980 8588 3984
rect 3176 3836 3240 3840
rect 3176 3780 3180 3836
rect 3180 3780 3236 3836
rect 3236 3780 3240 3836
rect 3176 3776 3240 3780
rect 3256 3836 3320 3840
rect 3256 3780 3260 3836
rect 3260 3780 3316 3836
rect 3316 3780 3320 3836
rect 3256 3776 3320 3780
rect 3336 3836 3400 3840
rect 3336 3780 3340 3836
rect 3340 3780 3396 3836
rect 3396 3780 3400 3836
rect 3336 3776 3400 3780
rect 3416 3836 3480 3840
rect 3416 3780 3420 3836
rect 3420 3780 3476 3836
rect 3476 3780 3480 3836
rect 3416 3776 3480 3780
rect 7624 3836 7688 3840
rect 7624 3780 7628 3836
rect 7628 3780 7684 3836
rect 7684 3780 7688 3836
rect 7624 3776 7688 3780
rect 7704 3836 7768 3840
rect 7704 3780 7708 3836
rect 7708 3780 7764 3836
rect 7764 3780 7768 3836
rect 7704 3776 7768 3780
rect 7784 3836 7848 3840
rect 7784 3780 7788 3836
rect 7788 3780 7844 3836
rect 7844 3780 7848 3836
rect 7784 3776 7848 3780
rect 7864 3836 7928 3840
rect 7864 3780 7868 3836
rect 7868 3780 7924 3836
rect 7924 3780 7928 3836
rect 7864 3776 7928 3780
rect 12072 3836 12136 3840
rect 12072 3780 12076 3836
rect 12076 3780 12132 3836
rect 12132 3780 12136 3836
rect 12072 3776 12136 3780
rect 12152 3836 12216 3840
rect 12152 3780 12156 3836
rect 12156 3780 12212 3836
rect 12212 3780 12216 3836
rect 12152 3776 12216 3780
rect 12232 3836 12296 3840
rect 12232 3780 12236 3836
rect 12236 3780 12292 3836
rect 12292 3780 12296 3836
rect 12232 3776 12296 3780
rect 12312 3836 12376 3840
rect 12312 3780 12316 3836
rect 12316 3780 12372 3836
rect 12372 3780 12376 3836
rect 12312 3776 12376 3780
rect 16520 3836 16584 3840
rect 16520 3780 16524 3836
rect 16524 3780 16580 3836
rect 16580 3780 16584 3836
rect 16520 3776 16584 3780
rect 16600 3836 16664 3840
rect 16600 3780 16604 3836
rect 16604 3780 16660 3836
rect 16660 3780 16664 3836
rect 16600 3776 16664 3780
rect 16680 3836 16744 3840
rect 16680 3780 16684 3836
rect 16684 3780 16740 3836
rect 16740 3780 16744 3836
rect 16680 3776 16744 3780
rect 16760 3836 16824 3840
rect 16760 3780 16764 3836
rect 16764 3780 16820 3836
rect 16820 3780 16824 3836
rect 16760 3776 16824 3780
rect 5212 3436 5276 3500
rect 5400 3292 5464 3296
rect 5400 3236 5404 3292
rect 5404 3236 5460 3292
rect 5460 3236 5464 3292
rect 5400 3232 5464 3236
rect 5480 3292 5544 3296
rect 5480 3236 5484 3292
rect 5484 3236 5540 3292
rect 5540 3236 5544 3292
rect 5480 3232 5544 3236
rect 5560 3292 5624 3296
rect 5560 3236 5564 3292
rect 5564 3236 5620 3292
rect 5620 3236 5624 3292
rect 5560 3232 5624 3236
rect 5640 3292 5704 3296
rect 5640 3236 5644 3292
rect 5644 3236 5700 3292
rect 5700 3236 5704 3292
rect 5640 3232 5704 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 14296 3292 14360 3296
rect 14296 3236 14300 3292
rect 14300 3236 14356 3292
rect 14356 3236 14360 3292
rect 14296 3232 14360 3236
rect 14376 3292 14440 3296
rect 14376 3236 14380 3292
rect 14380 3236 14436 3292
rect 14436 3236 14440 3292
rect 14376 3232 14440 3236
rect 14456 3292 14520 3296
rect 14456 3236 14460 3292
rect 14460 3236 14516 3292
rect 14516 3236 14520 3292
rect 14456 3232 14520 3236
rect 14536 3292 14600 3296
rect 14536 3236 14540 3292
rect 14540 3236 14596 3292
rect 14596 3236 14600 3292
rect 14536 3232 14600 3236
rect 16988 3224 17052 3228
rect 16988 3168 17038 3224
rect 17038 3168 17052 3224
rect 16988 3164 17052 3168
rect 7236 3028 7300 3092
rect 16988 2816 17052 2820
rect 16988 2760 17002 2816
rect 17002 2760 17052 2816
rect 16988 2756 17052 2760
rect 3176 2748 3240 2752
rect 3176 2692 3180 2748
rect 3180 2692 3236 2748
rect 3236 2692 3240 2748
rect 3176 2688 3240 2692
rect 3256 2748 3320 2752
rect 3256 2692 3260 2748
rect 3260 2692 3316 2748
rect 3316 2692 3320 2748
rect 3256 2688 3320 2692
rect 3336 2748 3400 2752
rect 3336 2692 3340 2748
rect 3340 2692 3396 2748
rect 3396 2692 3400 2748
rect 3336 2688 3400 2692
rect 3416 2748 3480 2752
rect 3416 2692 3420 2748
rect 3420 2692 3476 2748
rect 3476 2692 3480 2748
rect 3416 2688 3480 2692
rect 7624 2748 7688 2752
rect 7624 2692 7628 2748
rect 7628 2692 7684 2748
rect 7684 2692 7688 2748
rect 7624 2688 7688 2692
rect 7704 2748 7768 2752
rect 7704 2692 7708 2748
rect 7708 2692 7764 2748
rect 7764 2692 7768 2748
rect 7704 2688 7768 2692
rect 7784 2748 7848 2752
rect 7784 2692 7788 2748
rect 7788 2692 7844 2748
rect 7844 2692 7848 2748
rect 7784 2688 7848 2692
rect 7864 2748 7928 2752
rect 7864 2692 7868 2748
rect 7868 2692 7924 2748
rect 7924 2692 7928 2748
rect 7864 2688 7928 2692
rect 12072 2748 12136 2752
rect 12072 2692 12076 2748
rect 12076 2692 12132 2748
rect 12132 2692 12136 2748
rect 12072 2688 12136 2692
rect 12152 2748 12216 2752
rect 12152 2692 12156 2748
rect 12156 2692 12212 2748
rect 12212 2692 12216 2748
rect 12152 2688 12216 2692
rect 12232 2748 12296 2752
rect 12232 2692 12236 2748
rect 12236 2692 12292 2748
rect 12292 2692 12296 2748
rect 12232 2688 12296 2692
rect 12312 2748 12376 2752
rect 12312 2692 12316 2748
rect 12316 2692 12372 2748
rect 12372 2692 12376 2748
rect 12312 2688 12376 2692
rect 16520 2748 16584 2752
rect 16520 2692 16524 2748
rect 16524 2692 16580 2748
rect 16580 2692 16584 2748
rect 16520 2688 16584 2692
rect 16600 2748 16664 2752
rect 16600 2692 16604 2748
rect 16604 2692 16660 2748
rect 16660 2692 16664 2748
rect 16600 2688 16664 2692
rect 16680 2748 16744 2752
rect 16680 2692 16684 2748
rect 16684 2692 16740 2748
rect 16740 2692 16744 2748
rect 16680 2688 16744 2692
rect 16760 2748 16824 2752
rect 16760 2692 16764 2748
rect 16764 2692 16820 2748
rect 16820 2692 16824 2748
rect 16760 2688 16824 2692
rect 2820 2620 2884 2684
rect 13124 2620 13188 2684
rect 3924 2484 3988 2548
rect 4660 2484 4724 2548
rect 10916 2484 10980 2548
rect 6868 2272 6932 2276
rect 6868 2216 6918 2272
rect 6918 2216 6932 2272
rect 6868 2212 6932 2216
rect 16252 2348 16316 2412
rect 5400 2204 5464 2208
rect 5400 2148 5404 2204
rect 5404 2148 5460 2204
rect 5460 2148 5464 2204
rect 5400 2144 5464 2148
rect 5480 2204 5544 2208
rect 5480 2148 5484 2204
rect 5484 2148 5540 2204
rect 5540 2148 5544 2204
rect 5480 2144 5544 2148
rect 5560 2204 5624 2208
rect 5560 2148 5564 2204
rect 5564 2148 5620 2204
rect 5620 2148 5624 2204
rect 5560 2144 5624 2148
rect 5640 2204 5704 2208
rect 5640 2148 5644 2204
rect 5644 2148 5700 2204
rect 5700 2148 5704 2204
rect 5640 2144 5704 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 14296 2204 14360 2208
rect 14296 2148 14300 2204
rect 14300 2148 14356 2204
rect 14356 2148 14360 2204
rect 14296 2144 14360 2148
rect 14376 2204 14440 2208
rect 14376 2148 14380 2204
rect 14380 2148 14436 2204
rect 14436 2148 14440 2204
rect 14376 2144 14440 2148
rect 14456 2204 14520 2208
rect 14456 2148 14460 2204
rect 14460 2148 14516 2204
rect 14516 2148 14520 2204
rect 14456 2144 14520 2148
rect 14536 2204 14600 2208
rect 14536 2148 14540 2204
rect 14540 2148 14596 2204
rect 14596 2148 14600 2204
rect 14536 2144 14600 2148
rect 8340 1940 8404 2004
<< metal4 >>
rect 15515 15196 15581 15197
rect 15515 15132 15516 15196
rect 15580 15132 15581 15196
rect 15515 15131 15581 15132
rect 3168 14720 3488 14736
rect 3168 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3488 14720
rect 3168 13632 3488 14656
rect 3168 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3488 13632
rect 1899 12612 1965 12613
rect 1899 12548 1900 12612
rect 1964 12548 1965 12612
rect 1899 12547 1965 12548
rect 1715 10844 1781 10845
rect 1715 10780 1716 10844
rect 1780 10780 1781 10844
rect 1715 10779 1781 10780
rect 1718 7445 1778 10779
rect 1715 7444 1781 7445
rect 1715 7380 1716 7444
rect 1780 7380 1781 7444
rect 1715 7379 1781 7380
rect 1902 6930 1962 12547
rect 3168 12544 3488 13568
rect 3168 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3488 12544
rect 2451 12476 2517 12477
rect 2451 12412 2452 12476
rect 2516 12412 2517 12476
rect 2451 12411 2517 12412
rect 2454 8397 2514 12411
rect 3168 11456 3488 12480
rect 5392 14176 5712 14736
rect 5392 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5712 14176
rect 5392 13088 5712 14112
rect 5392 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5712 13088
rect 5392 12000 5712 13024
rect 5392 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5712 12000
rect 4107 11932 4173 11933
rect 4107 11868 4108 11932
rect 4172 11868 4173 11932
rect 4107 11867 4173 11868
rect 3168 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3488 11456
rect 3168 10368 3488 11392
rect 3168 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3488 10368
rect 3168 9280 3488 10304
rect 3168 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3488 9280
rect 2819 8668 2885 8669
rect 2819 8604 2820 8668
rect 2884 8604 2885 8668
rect 2819 8603 2885 8604
rect 2451 8396 2517 8397
rect 2451 8332 2452 8396
rect 2516 8332 2517 8396
rect 2451 8331 2517 8332
rect 1718 6870 1962 6930
rect 1718 4045 1778 6870
rect 2454 6493 2514 8331
rect 2635 7716 2701 7717
rect 2635 7652 2636 7716
rect 2700 7652 2701 7716
rect 2635 7651 2701 7652
rect 2451 6492 2517 6493
rect 2451 6428 2452 6492
rect 2516 6428 2517 6492
rect 2451 6427 2517 6428
rect 2638 4045 2698 7651
rect 1715 4044 1781 4045
rect 1715 3980 1716 4044
rect 1780 3980 1781 4044
rect 1715 3979 1781 3980
rect 2635 4044 2701 4045
rect 2635 3980 2636 4044
rect 2700 3980 2701 4044
rect 2635 3979 2701 3980
rect 2822 2685 2882 8603
rect 3168 8192 3488 9216
rect 3168 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3488 8192
rect 3168 7104 3488 8128
rect 3168 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3488 7104
rect 3168 6016 3488 7040
rect 4110 6901 4170 11867
rect 5392 10912 5712 11936
rect 5392 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5712 10912
rect 5392 9824 5712 10848
rect 5392 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5712 9824
rect 5211 9348 5277 9349
rect 5211 9284 5212 9348
rect 5276 9284 5277 9348
rect 5211 9283 5277 9284
rect 4475 8532 4541 8533
rect 4475 8468 4476 8532
rect 4540 8468 4541 8532
rect 4475 8467 4541 8468
rect 4107 6900 4173 6901
rect 4107 6836 4108 6900
rect 4172 6836 4173 6900
rect 4107 6835 4173 6836
rect 3168 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3488 6016
rect 3168 4928 3488 5952
rect 3168 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3488 4928
rect 3168 3840 3488 4864
rect 4110 4861 4170 6835
rect 4107 4860 4173 4861
rect 4107 4796 4108 4860
rect 4172 4796 4173 4860
rect 4107 4795 4173 4796
rect 3168 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3488 3840
rect 3168 2752 3488 3776
rect 4110 2790 4170 4795
rect 3168 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3488 2752
rect 2819 2684 2885 2685
rect 2819 2620 2820 2684
rect 2884 2620 2885 2684
rect 2819 2619 2885 2620
rect 3168 2128 3488 2688
rect 3926 2730 4170 2790
rect 4478 2790 4538 8467
rect 4659 5676 4725 5677
rect 4659 5612 4660 5676
rect 4724 5612 4725 5676
rect 4659 5611 4725 5612
rect 4662 4045 4722 5611
rect 4659 4044 4725 4045
rect 4659 3980 4660 4044
rect 4724 3980 4725 4044
rect 4659 3979 4725 3980
rect 5214 3501 5274 9283
rect 5392 8736 5712 9760
rect 7616 14720 7936 14736
rect 7616 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7936 14720
rect 7616 13632 7936 14656
rect 7616 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7936 13632
rect 7616 12544 7936 13568
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 8523 12748 8589 12749
rect 8523 12684 8524 12748
rect 8588 12684 8589 12748
rect 8523 12683 8589 12684
rect 7616 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7936 12544
rect 7616 11456 7936 12480
rect 7616 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7936 11456
rect 7616 10368 7936 11392
rect 7616 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7936 10368
rect 7235 9348 7301 9349
rect 7235 9284 7236 9348
rect 7300 9284 7301 9348
rect 7235 9283 7301 9284
rect 7238 8805 7298 9283
rect 7616 9280 7936 10304
rect 8526 10165 8586 12683
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 8523 10164 8589 10165
rect 8523 10100 8524 10164
rect 8588 10100 8589 10164
rect 8523 10099 8589 10100
rect 7616 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7936 9280
rect 7235 8804 7301 8805
rect 7235 8740 7236 8804
rect 7300 8740 7301 8804
rect 7235 8739 7301 8740
rect 5392 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5712 8736
rect 5392 7648 5712 8672
rect 5392 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5712 7648
rect 5392 6560 5712 7584
rect 6867 6764 6933 6765
rect 6867 6700 6868 6764
rect 6932 6700 6933 6764
rect 6867 6699 6933 6700
rect 5392 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5712 6560
rect 5392 5472 5712 6496
rect 5392 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5712 5472
rect 5392 4384 5712 5408
rect 5392 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5712 4384
rect 5211 3500 5277 3501
rect 5211 3436 5212 3500
rect 5276 3436 5277 3500
rect 5211 3435 5277 3436
rect 5392 3296 5712 4320
rect 5392 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5712 3296
rect 4478 2730 4722 2790
rect 3926 2549 3986 2730
rect 4662 2549 4722 2730
rect 3923 2548 3989 2549
rect 3923 2484 3924 2548
rect 3988 2484 3989 2548
rect 3923 2483 3989 2484
rect 4659 2548 4725 2549
rect 4659 2484 4660 2548
rect 4724 2484 4725 2548
rect 4659 2483 4725 2484
rect 5392 2208 5712 3232
rect 6870 2277 6930 6699
rect 7238 6629 7298 8739
rect 7616 8192 7936 9216
rect 7616 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7936 8192
rect 7616 7104 7936 8128
rect 7616 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7936 7104
rect 7235 6628 7301 6629
rect 7235 6564 7236 6628
rect 7300 6564 7301 6628
rect 7235 6563 7301 6564
rect 7235 6356 7301 6357
rect 7235 6292 7236 6356
rect 7300 6292 7301 6356
rect 7235 6291 7301 6292
rect 7238 3093 7298 6291
rect 7616 6016 7936 7040
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 8523 6900 8589 6901
rect 8523 6836 8524 6900
rect 8588 6836 8589 6900
rect 8523 6835 8589 6836
rect 7616 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7936 6016
rect 7616 4928 7936 5952
rect 8339 5676 8405 5677
rect 8339 5612 8340 5676
rect 8404 5612 8405 5676
rect 8339 5611 8405 5612
rect 7616 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7936 4928
rect 7616 3840 7936 4864
rect 7616 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7936 3840
rect 7235 3092 7301 3093
rect 7235 3028 7236 3092
rect 7300 3028 7301 3092
rect 7235 3027 7301 3028
rect 7616 2752 7936 3776
rect 7616 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7936 2752
rect 6867 2276 6933 2277
rect 6867 2212 6868 2276
rect 6932 2212 6933 2276
rect 6867 2211 6933 2212
rect 5392 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5712 2208
rect 5392 2128 5712 2144
rect 7616 2128 7936 2688
rect 8342 2005 8402 5611
rect 8526 4045 8586 6835
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 12064 14720 12384 14736
rect 12064 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12384 14720
rect 12064 13632 12384 14656
rect 12064 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12384 13632
rect 12064 12544 12384 13568
rect 12064 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12384 12544
rect 12064 11456 12384 12480
rect 12064 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12384 11456
rect 12064 10368 12384 11392
rect 12064 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12384 10368
rect 12064 9280 12384 10304
rect 14288 14176 14608 14736
rect 14288 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14608 14176
rect 14288 13088 14608 14112
rect 14288 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14608 13088
rect 14288 12000 14608 13024
rect 14288 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14608 12000
rect 14288 10912 14608 11936
rect 15147 11252 15213 11253
rect 15147 11188 15148 11252
rect 15212 11188 15213 11252
rect 15147 11187 15213 11188
rect 14288 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14608 10912
rect 14288 9824 14608 10848
rect 14288 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14608 9824
rect 13123 9756 13189 9757
rect 13123 9692 13124 9756
rect 13188 9692 13189 9756
rect 13123 9691 13189 9692
rect 12064 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12384 9280
rect 12064 8192 12384 9216
rect 12064 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12384 8192
rect 12064 7104 12384 8128
rect 12064 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12384 7104
rect 10915 6220 10981 6221
rect 10915 6156 10916 6220
rect 10980 6156 10981 6220
rect 10915 6155 10981 6156
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 8523 4044 8589 4045
rect 8523 3980 8524 4044
rect 8588 3980 8589 4044
rect 8523 3979 8589 3980
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 10918 2549 10978 6155
rect 12064 6016 12384 7040
rect 12064 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12384 6016
rect 12064 4928 12384 5952
rect 12064 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12384 4928
rect 12064 3840 12384 4864
rect 12064 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12384 3840
rect 12064 2752 12384 3776
rect 12064 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12384 2752
rect 10915 2548 10981 2549
rect 10915 2484 10916 2548
rect 10980 2484 10981 2548
rect 10915 2483 10981 2484
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12064 2128 12384 2688
rect 13126 2685 13186 9691
rect 14288 8736 14608 9760
rect 14288 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14608 8736
rect 14288 7648 14608 8672
rect 14288 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14608 7648
rect 14288 6560 14608 7584
rect 14288 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14608 6560
rect 14288 5472 14608 6496
rect 14288 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14608 5472
rect 14288 4384 14608 5408
rect 14288 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14608 4384
rect 14288 3296 14608 4320
rect 15150 4181 15210 11187
rect 15518 6901 15578 15131
rect 17171 14788 17237 14789
rect 16512 14720 16832 14736
rect 17171 14724 17172 14788
rect 17236 14724 17237 14788
rect 17171 14723 17237 14724
rect 16512 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16832 14720
rect 16512 13632 16832 14656
rect 17174 14109 17234 14723
rect 17171 14108 17237 14109
rect 17171 14044 17172 14108
rect 17236 14044 17237 14108
rect 17171 14043 17237 14044
rect 16987 13972 17053 13973
rect 16987 13908 16988 13972
rect 17052 13908 17053 13972
rect 16987 13907 17053 13908
rect 16512 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16832 13632
rect 16512 12544 16832 13568
rect 16512 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16832 12544
rect 16067 12204 16133 12205
rect 16067 12140 16068 12204
rect 16132 12140 16133 12204
rect 16067 12139 16133 12140
rect 16070 11117 16130 12139
rect 16251 11796 16317 11797
rect 16251 11732 16252 11796
rect 16316 11732 16317 11796
rect 16251 11731 16317 11732
rect 16067 11116 16133 11117
rect 16067 11052 16068 11116
rect 16132 11052 16133 11116
rect 16067 11051 16133 11052
rect 15515 6900 15581 6901
rect 15515 6836 15516 6900
rect 15580 6836 15581 6900
rect 15515 6835 15581 6836
rect 15518 5813 15578 6835
rect 15515 5812 15581 5813
rect 15515 5748 15516 5812
rect 15580 5748 15581 5812
rect 15515 5747 15581 5748
rect 16070 5541 16130 11051
rect 16067 5540 16133 5541
rect 16067 5476 16068 5540
rect 16132 5476 16133 5540
rect 16067 5475 16133 5476
rect 15147 4180 15213 4181
rect 15147 4116 15148 4180
rect 15212 4116 15213 4180
rect 15147 4115 15213 4116
rect 14288 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14608 3296
rect 13123 2684 13189 2685
rect 13123 2620 13124 2684
rect 13188 2620 13189 2684
rect 13123 2619 13189 2620
rect 14288 2208 14608 3232
rect 16070 2790 16130 5475
rect 16254 4861 16314 11731
rect 16512 11456 16832 12480
rect 16512 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16832 11456
rect 16512 10368 16832 11392
rect 16512 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16832 10368
rect 16512 9280 16832 10304
rect 16512 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16832 9280
rect 16512 8192 16832 9216
rect 16512 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16832 8192
rect 16512 7104 16832 8128
rect 16512 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16832 7104
rect 16512 6016 16832 7040
rect 16512 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16832 6016
rect 16512 4928 16832 5952
rect 16512 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16832 4928
rect 16251 4860 16317 4861
rect 16251 4796 16252 4860
rect 16316 4796 16317 4860
rect 16251 4795 16317 4796
rect 16512 3840 16832 4864
rect 16512 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16832 3840
rect 16070 2730 16314 2790
rect 16254 2413 16314 2730
rect 16512 2752 16832 3776
rect 16990 3229 17050 13907
rect 17174 5405 17234 14043
rect 17171 5404 17237 5405
rect 17171 5340 17172 5404
rect 17236 5340 17237 5404
rect 17171 5339 17237 5340
rect 16987 3228 17053 3229
rect 16987 3164 16988 3228
rect 17052 3164 17053 3228
rect 16987 3163 17053 3164
rect 16990 2821 17050 3163
rect 16987 2820 17053 2821
rect 16987 2756 16988 2820
rect 17052 2756 17053 2820
rect 16987 2755 17053 2756
rect 16512 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16832 2752
rect 16251 2412 16317 2413
rect 16251 2348 16252 2412
rect 16316 2348 16317 2412
rect 16251 2347 16317 2348
rect 14288 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14608 2208
rect 14288 2128 14608 2144
rect 16512 2128 16832 2688
rect 8339 2004 8405 2005
rect 8339 1940 8340 2004
rect 8404 1940 8405 2004
rect 8339 1939 8405 1940
use sky130_fd_sc_hd__diode_2  ANTENNA__34__A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18216 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1649977179
transform 1 0 6440 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1649977179
transform 1 0 15640 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform 1 0 16560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1649977179
transform 1 0 16008 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform 1 0 17204 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform -1 0 4140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform 1 0 4416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform 1 0 4140 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform -1 0 16100 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1649977179
transform -1 0 16284 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform -1 0 1656 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform -1 0 11684 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform 1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1649977179
transform 1 0 1932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform 1 0 3864 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform 1 0 4232 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1649977179
transform 1 0 1932 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1649977179
transform 1 0 1748 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1649977179
transform -1 0 18400 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1649977179
transform 1 0 17388 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1649977179
transform 1 0 17480 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1649977179
transform 1 0 17940 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1649977179
transform -1 0 17756 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1649977179
transform -1 0 18584 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1649977179
transform -1 0 18492 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform 1 0 17664 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1649977179
transform -1 0 17848 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform -1 0 18492 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1649977179
transform 1 0 17296 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform -1 0 18584 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform 1 0 17480 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1649977179
transform 1 0 17296 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1649977179
transform -1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform -1 0 17848 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1649977179
transform -1 0 17848 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1649977179
transform -1 0 17664 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_0_S_in_A
timestamp 1649977179
transform -1 0 17112 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 16192 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform -1 0 1564 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform -1 0 2944 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 13708 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform -1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 11592 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform -1 0 16744 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 16652 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE_B_N
timestamp 1649977179
transform 1 0 13064 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE_A
timestamp 1649977179
transform -1 0 16836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7360 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 7176 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 7360 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6164 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 8096 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4416 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 6164 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6808 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4876 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 5244 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 4232 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6348 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 3680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4048 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 2760 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 2576 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 1748 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 2392 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 2392 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7452 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 2760 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 1564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 17204 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 16836 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 17296 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 1564 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 2576 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16008 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 17020 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 17204 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16836 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17020 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 16192 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16744 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 17020 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 5152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 2208 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 17020 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 16836 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7820 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4600 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11960 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11132 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 12512 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12144 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10948 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 10488 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9384 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 9752 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9384 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9384 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 9016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 9016 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9200 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12788 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12144 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 9752 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 15824 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 13616 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 13156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18400 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 16284 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 16376 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 17112 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 16468 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 16652 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16192 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 15824 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 16008 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11776 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13708 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 12328 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 13984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13524 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 15364 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 15732 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12604 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12880 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15916 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 16284 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 16376 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 16744 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 16928 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 17112 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12512 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17296 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 18492 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 18584 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 18216 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 17296 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 18308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 18400 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 18032 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 18308 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 18492 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 18124 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 16008 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14996 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 15732 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_179
timestamp 1649977179
transform 1 0 17572 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_128
timestamp 1649977179
transform 1 0 12880 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_96
timestamp 1649977179
transform 1 0 9936 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_119
timestamp 1649977179
transform 1 0 12052 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_78
timestamp 1649977179
transform 1 0 8280 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_92
timestamp 1649977179
transform 1 0 9568 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_135
timestamp 1649977179
transform 1 0 13524 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1649977179
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_67
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_122
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_82
timestamp 1649977179
transform 1 0 8648 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_140
timestamp 1649977179
transform 1 0 13984 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_173 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17020 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_179
timestamp 1649977179
transform 1 0 17572 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_169
timestamp 1649977179
transform 1 0 16652 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_175
timestamp 1649977179
transform 1 0 17204 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_115
timestamp 1649977179
transform 1 0 11684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_175
timestamp 1649977179
transform 1 0 17204 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_112
timestamp 1649977179
transform 1 0 11408 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_18
timestamp 1649977179
transform 1 0 2760 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_157
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_19
timestamp 1649977179
transform 1 0 2852 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_189
timestamp 1649977179
transform 1 0 18492 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_143
timestamp 1649977179
transform 1 0 14260 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1649977179
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_33
timestamp 1649977179
transform 1 0 4140 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_87
timestamp 1649977179
transform 1 0 9108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_106
timestamp 1649977179
transform 1 0 10856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_163 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_34
timestamp 1649977179
transform 1 0 4232 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_54
timestamp 1649977179
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_89
timestamp 1649977179
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_108
timestamp 1649977179
transform 1 0 11040 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_75
timestamp 1649977179
transform 1 0 8004 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_126 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12696 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_130
timestamp 1649977179
transform 1 0 13064 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_189
timestamp 1649977179
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_11
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_45
timestamp 1649977179
transform 1 0 5244 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_123 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12420 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_127
timestamp 1649977179
transform 1 0 12788 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_161
timestamp 1649977179
transform 1 0 15916 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_13
timestamp 1649977179
transform 1 0 2300 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1649977179
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_119
timestamp 1649977179
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_136
timestamp 1649977179
transform 1 0 13616 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_153
timestamp 1649977179
transform 1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_164
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_175
timestamp 1649977179
transform 1 0 17204 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_178
timestamp 1649977179
transform 1 0 17480 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1649977179
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_20_104
timestamp 1649977179
transform 1 0 10672 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_110
timestamp 1649977179
transform 1 0 11224 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_117
timestamp 1649977179
transform 1 0 11868 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_123
timestamp 1649977179
transform 1 0 12420 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1649977179
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_154
timestamp 1649977179
transform 1 0 15272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_158
timestamp 1649977179
transform 1 0 15640 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_162
timestamp 1649977179
transform 1 0 16008 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_166
timestamp 1649977179
transform 1 0 16376 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_171 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16836 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_179
timestamp 1649977179
transform 1 0 17572 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_182
timestamp 1649977179
transform 1 0 17848 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_186
timestamp 1649977179
transform 1 0 18216 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_35
timestamp 1649977179
transform 1 0 4324 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_46
timestamp 1649977179
transform 1 0 5336 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_52
timestamp 1649977179
transform 1 0 5888 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_61
timestamp 1649977179
transform 1 0 6716 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_64
timestamp 1649977179
transform 1 0 6992 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_76
timestamp 1649977179
transform 1 0 8096 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_88
timestamp 1649977179
transform 1 0 9200 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_96
timestamp 1649977179
transform 1 0 9936 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1649977179
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_129
timestamp 1649977179
transform 1 0 12972 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_57
timestamp 1649977179
transform 1 0 6348 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_69
timestamp 1649977179
transform 1 0 7452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1649977179
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_113
timestamp 1649977179
transform 1 0 11500 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_125
timestamp 1649977179
transform 1 0 12604 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1649977179
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_169
timestamp 1649977179
transform 1 0 16652 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_181
timestamp 1649977179
transform 1 0 17756 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 16560 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _17_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _18_
timestamp 1649977179
transform -1 0 7912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _19_
timestamp 1649977179
transform 1 0 8372 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _20_
timestamp 1649977179
transform -1 0 9292 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _21_
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _22_
timestamp 1649977179
transform 1 0 11868 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _23_
timestamp 1649977179
transform -1 0 6072 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _24_
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _25_
timestamp 1649977179
transform 1 0 6808 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _26_
timestamp 1649977179
transform 1 0 15548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _27_
timestamp 1649977179
transform 1 0 13984 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _28_
timestamp 1649977179
transform 1 0 16376 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _29_
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _30_
timestamp 1649977179
transform 1 0 18308 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _31_
timestamp 1649977179
transform -1 0 13156 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _32_
timestamp 1649977179
transform -1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _33_
timestamp 1649977179
transform 1 0 5428 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _34_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18216 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _35_
timestamp 1649977179
transform 1 0 17848 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _36_
timestamp 1649977179
transform -1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _37_
timestamp 1649977179
transform -1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _38_
timestamp 1649977179
transform -1 0 12052 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _39_
timestamp 1649977179
transform -1 0 7912 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _40_
timestamp 1649977179
transform -1 0 7268 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _41_
timestamp 1649977179
transform -1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _42_
timestamp 1649977179
transform -1 0 4600 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _43_
timestamp 1649977179
transform -1 0 6716 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _44_
timestamp 1649977179
transform -1 0 4140 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _45_
timestamp 1649977179
transform -1 0 4784 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _46_
timestamp 1649977179
transform -1 0 9568 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _47_
timestamp 1649977179
transform -1 0 8280 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _48_
timestamp 1649977179
transform -1 0 2024 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _49_
timestamp 1649977179
transform -1 0 9844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _50_
timestamp 1649977179
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _51_
timestamp 1649977179
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _52_
timestamp 1649977179
transform -1 0 5704 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _53_
timestamp 1649977179
transform -1 0 4140 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _54_
timestamp 1649977179
transform -1 0 1932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _55_
timestamp 1649977179
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _56_
timestamp 1649977179
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _57_
timestamp 1649977179
transform 1 0 18216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _58_
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _59_
timestamp 1649977179
transform 1 0 17664 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _60_
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _61_
timestamp 1649977179
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _62_
timestamp 1649977179
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _63_
timestamp 1649977179
transform 1 0 17848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _64_
timestamp 1649977179
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _65_
timestamp 1649977179
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _66_
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _67_
timestamp 1649977179
transform 1 0 17848 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _68_
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _69_
timestamp 1649977179
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _70_
timestamp 1649977179
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _71_
timestamp 1649977179
transform 1 0 17848 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _72_
timestamp 1649977179
transform 1 0 17480 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _73_
timestamp 1649977179
transform 1 0 18216 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _74_
timestamp 1649977179
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _75_
timestamp 1649977179
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _76_
timestamp 1649977179
transform 1 0 17848 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9568 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk_0_S_in
timestamp 1649977179
transform -1 0 7544 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk_0_S_in
timestamp 1649977179
transform -1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk_0_S_in
timestamp 1649977179
transform 1 0 7820 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 2576 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 5244 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform -1 0 12236 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform -1 0 14812 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 10396 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14168 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1649977179
transform -1 0 6256 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1649977179
transform 1 0 8096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1649977179
transform 1 0 7728 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1649977179
transform 1 0 13248 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1649977179
transform 1 0 10120 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1649977179
transform -1 0 2208 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1649977179
transform 1 0 15732 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1649977179
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1649977179
transform 1 0 14076 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1649977179
transform 1 0 11868 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1649977179
transform 1 0 10396 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1649977179
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1649977179
transform 1 0 15272 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1649977179
transform 1 0 12328 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1649977179
transform -1 0 18216 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1649977179
transform 1 0 14904 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1649977179
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1649977179
transform -1 0 15272 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1649977179
transform 1 0 13064 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1649977179
transform 1 0 1472 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1649977179
transform 1 0 2944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1649977179
transform -1 0 17480 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1649977179
transform 1 0 15732 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1649977179
transform 1 0 9752 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15732 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13248 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_4  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 15364 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13984 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8464 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7912 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2760 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4048 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5796 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3680 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 2852 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 1932 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 3404 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 2852 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 1564 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 4232 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 3864 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3036 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 1472 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2208 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4048 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 3956 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4784 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7912 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8556 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6900 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8832 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 6440 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6256 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5152 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8096 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11040 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12420 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10396 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7360 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8648 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11132 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 9568 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 9936 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11316 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11040 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12144 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13616 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14076 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11408 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13800 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12972 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15824 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 15088 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16100 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16836 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18124 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15916 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14904 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17480 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15180 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12144 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6164 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5336 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5152 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 5152 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 5336 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_bottom_ipin_0.sky130_fd_sc_hd__buf_4_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11316 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4324 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4416 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3864 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2852 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2576 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2024 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2024 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 1932 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2944 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2576 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3772 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2208 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 1748 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1932 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 2760 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4600 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 2852 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform -1 0 4876 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5244 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10856 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3588 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11316 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5152 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2852 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10580 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2576 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4416 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6532 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7912 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6992 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8648 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8372 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6992 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform -1 0 6256 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7820 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5704 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6532 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6900 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7636 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6624 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6532 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4600 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10580 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9752 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10120 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8924 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9292 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8924 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6992 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10396 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9568 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform -1 0 9660 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8004 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9568 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 10212 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform -1 0 11040 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7912 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 11040 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6992 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10396 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9568 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11040 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 9568 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9016 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15088 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14904 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14904 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14904 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12420 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 12328 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14444 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1649977179
transform 1 0 13616 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12788 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1649977179
transform 1 0 11960 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13156 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12696 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11500 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13800 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12328 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13432 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13064 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1649977179
transform 1 0 13156 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12604 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12328 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1649977179
transform -1 0 13064 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14628 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15456 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1649977179
transform 1 0 15548 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1649977179
transform -1 0 13984 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1649977179
transform -1 0 14628 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14260 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18308 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17572 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17204 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1649977179
transform -1 0 18308 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17572 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16376 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17480 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15364 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1649977179
transform 1 0 15180 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1649977179
transform -1 0 13984 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1649977179
transform -1 0 14168 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__buf_4  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8832 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1649977179
transform -1 0 3588 0 1 6528
box -38 -48 590 592
<< labels >>
rlabel metal2 s 1122 16400 1178 17200 6 IO_ISOL_N
port 0 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 SC_IN_BOT
port 1 nsew signal input
rlabel metal2 s 3330 16400 3386 17200 6 SC_IN_TOP
port 2 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 SC_OUT_BOT
port 3 nsew signal tristate
rlabel metal2 s 5538 16400 5594 17200 6 SC_OUT_TOP
port 4 nsew signal tristate
rlabel metal4 s 5392 2128 5712 14736 6 VGND
port 5 nsew ground input
rlabel metal4 s 9840 2128 10160 14736 6 VGND
port 5 nsew ground input
rlabel metal4 s 14288 2128 14608 14736 6 VGND
port 5 nsew ground input
rlabel metal4 s 3168 2128 3488 14736 6 VPWR
port 6 nsew power input
rlabel metal4 s 7616 2128 7936 14736 6 VPWR
port 6 nsew power input
rlabel metal4 s 12064 2128 12384 14736 6 VPWR
port 6 nsew power input
rlabel metal4 s 16512 2128 16832 14736 6 VPWR
port 6 nsew power input
rlabel metal2 s 1214 0 1270 800 6 bottom_grid_pin_0_
port 7 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 bottom_grid_pin_10_
port 8 nsew signal tristate
rlabel metal2 s 11242 0 11298 800 6 bottom_grid_pin_11_
port 9 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 bottom_grid_pin_12_
port 10 nsew signal tristate
rlabel metal2 s 13082 0 13138 800 6 bottom_grid_pin_13_
port 11 nsew signal tristate
rlabel metal2 s 13910 0 13966 800 6 bottom_grid_pin_14_
port 12 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 bottom_grid_pin_15_
port 13 nsew signal tristate
rlabel metal2 s 2134 0 2190 800 6 bottom_grid_pin_1_
port 14 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 bottom_grid_pin_2_
port 15 nsew signal tristate
rlabel metal2 s 3974 0 4030 800 6 bottom_grid_pin_3_
port 16 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 bottom_grid_pin_4_
port 17 nsew signal tristate
rlabel metal2 s 5814 0 5870 800 6 bottom_grid_pin_5_
port 18 nsew signal tristate
rlabel metal2 s 6734 0 6790 800 6 bottom_grid_pin_6_
port 19 nsew signal tristate
rlabel metal2 s 7562 0 7618 800 6 bottom_grid_pin_7_
port 20 nsew signal tristate
rlabel metal2 s 8482 0 8538 800 6 bottom_grid_pin_8_
port 21 nsew signal tristate
rlabel metal2 s 9402 0 9458 800 6 bottom_grid_pin_9_
port 22 nsew signal tristate
rlabel metal2 s 15750 0 15806 800 6 bottom_width_0_height_0__pin_0_
port 23 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 bottom_width_0_height_0__pin_1_lower
port 24 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 bottom_width_0_height_0__pin_1_upper
port 25 nsew signal tristate
rlabel metal2 s 7746 16400 7802 17200 6 ccff_head
port 26 nsew signal input
rlabel metal2 s 9954 16400 10010 17200 6 ccff_tail
port 27 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 chanx_left_in[0]
port 28 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_in[10]
port 29 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 chanx_left_in[11]
port 30 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 chanx_left_in[12]
port 31 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 chanx_left_in[13]
port 32 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 chanx_left_in[14]
port 33 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 chanx_left_in[15]
port 34 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 chanx_left_in[16]
port 35 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 chanx_left_in[17]
port 36 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 chanx_left_in[18]
port 37 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 chanx_left_in[19]
port 38 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 chanx_left_in[1]
port 39 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[2]
port 40 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[3]
port 41 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 chanx_left_in[4]
port 42 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[5]
port 43 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[6]
port 44 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[7]
port 45 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[8]
port 46 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[9]
port 47 nsew signal input
rlabel metal3 s 0 552 800 672 6 chanx_left_out[0]
port 48 nsew signal tristate
rlabel metal3 s 0 4632 800 4752 6 chanx_left_out[10]
port 49 nsew signal tristate
rlabel metal3 s 0 5040 800 5160 6 chanx_left_out[11]
port 50 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 chanx_left_out[12]
port 51 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 chanx_left_out[13]
port 52 nsew signal tristate
rlabel metal3 s 0 6400 800 6520 6 chanx_left_out[14]
port 53 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 chanx_left_out[15]
port 54 nsew signal tristate
rlabel metal3 s 0 7216 800 7336 6 chanx_left_out[16]
port 55 nsew signal tristate
rlabel metal3 s 0 7624 800 7744 6 chanx_left_out[17]
port 56 nsew signal tristate
rlabel metal3 s 0 8032 800 8152 6 chanx_left_out[18]
port 57 nsew signal tristate
rlabel metal3 s 0 8440 800 8560 6 chanx_left_out[19]
port 58 nsew signal tristate
rlabel metal3 s 0 960 800 1080 6 chanx_left_out[1]
port 59 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 chanx_left_out[2]
port 60 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 chanx_left_out[3]
port 61 nsew signal tristate
rlabel metal3 s 0 2184 800 2304 6 chanx_left_out[4]
port 62 nsew signal tristate
rlabel metal3 s 0 2592 800 2712 6 chanx_left_out[5]
port 63 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 chanx_left_out[6]
port 64 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 chanx_left_out[7]
port 65 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 chanx_left_out[8]
port 66 nsew signal tristate
rlabel metal3 s 0 4224 800 4344 6 chanx_left_out[9]
port 67 nsew signal tristate
rlabel metal3 s 19200 8712 20000 8832 6 chanx_right_in[0]
port 68 nsew signal input
rlabel metal3 s 19200 12928 20000 13048 6 chanx_right_in[10]
port 69 nsew signal input
rlabel metal3 s 19200 13336 20000 13456 6 chanx_right_in[11]
port 70 nsew signal input
rlabel metal3 s 19200 13744 20000 13864 6 chanx_right_in[12]
port 71 nsew signal input
rlabel metal3 s 19200 14152 20000 14272 6 chanx_right_in[13]
port 72 nsew signal input
rlabel metal3 s 19200 14696 20000 14816 6 chanx_right_in[14]
port 73 nsew signal input
rlabel metal3 s 19200 15104 20000 15224 6 chanx_right_in[15]
port 74 nsew signal input
rlabel metal3 s 19200 15512 20000 15632 6 chanx_right_in[16]
port 75 nsew signal input
rlabel metal3 s 19200 15920 20000 16040 6 chanx_right_in[17]
port 76 nsew signal input
rlabel metal3 s 19200 16328 20000 16448 6 chanx_right_in[18]
port 77 nsew signal input
rlabel metal3 s 19200 16736 20000 16856 6 chanx_right_in[19]
port 78 nsew signal input
rlabel metal3 s 19200 9120 20000 9240 6 chanx_right_in[1]
port 79 nsew signal input
rlabel metal3 s 19200 9528 20000 9648 6 chanx_right_in[2]
port 80 nsew signal input
rlabel metal3 s 19200 9936 20000 10056 6 chanx_right_in[3]
port 81 nsew signal input
rlabel metal3 s 19200 10344 20000 10464 6 chanx_right_in[4]
port 82 nsew signal input
rlabel metal3 s 19200 10752 20000 10872 6 chanx_right_in[5]
port 83 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 chanx_right_in[6]
port 84 nsew signal input
rlabel metal3 s 19200 11704 20000 11824 6 chanx_right_in[7]
port 85 nsew signal input
rlabel metal3 s 19200 12112 20000 12232 6 chanx_right_in[8]
port 86 nsew signal input
rlabel metal3 s 19200 12520 20000 12640 6 chanx_right_in[9]
port 87 nsew signal input
rlabel metal3 s 19200 144 20000 264 6 chanx_right_out[0]
port 88 nsew signal tristate
rlabel metal3 s 19200 4360 20000 4480 6 chanx_right_out[10]
port 89 nsew signal tristate
rlabel metal3 s 19200 4768 20000 4888 6 chanx_right_out[11]
port 90 nsew signal tristate
rlabel metal3 s 19200 5176 20000 5296 6 chanx_right_out[12]
port 91 nsew signal tristate
rlabel metal3 s 19200 5584 20000 5704 6 chanx_right_out[13]
port 92 nsew signal tristate
rlabel metal3 s 19200 6128 20000 6248 6 chanx_right_out[14]
port 93 nsew signal tristate
rlabel metal3 s 19200 6536 20000 6656 6 chanx_right_out[15]
port 94 nsew signal tristate
rlabel metal3 s 19200 6944 20000 7064 6 chanx_right_out[16]
port 95 nsew signal tristate
rlabel metal3 s 19200 7352 20000 7472 6 chanx_right_out[17]
port 96 nsew signal tristate
rlabel metal3 s 19200 7760 20000 7880 6 chanx_right_out[18]
port 97 nsew signal tristate
rlabel metal3 s 19200 8168 20000 8288 6 chanx_right_out[19]
port 98 nsew signal tristate
rlabel metal3 s 19200 552 20000 672 6 chanx_right_out[1]
port 99 nsew signal tristate
rlabel metal3 s 19200 960 20000 1080 6 chanx_right_out[2]
port 100 nsew signal tristate
rlabel metal3 s 19200 1368 20000 1488 6 chanx_right_out[3]
port 101 nsew signal tristate
rlabel metal3 s 19200 1776 20000 1896 6 chanx_right_out[4]
port 102 nsew signal tristate
rlabel metal3 s 19200 2184 20000 2304 6 chanx_right_out[5]
port 103 nsew signal tristate
rlabel metal3 s 19200 2592 20000 2712 6 chanx_right_out[6]
port 104 nsew signal tristate
rlabel metal3 s 19200 3136 20000 3256 6 chanx_right_out[7]
port 105 nsew signal tristate
rlabel metal3 s 19200 3544 20000 3664 6 chanx_right_out[8]
port 106 nsew signal tristate
rlabel metal3 s 19200 3952 20000 4072 6 chanx_right_out[9]
port 107 nsew signal tristate
rlabel metal2 s 14370 16400 14426 17200 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 108 nsew signal tristate
rlabel metal2 s 16578 16400 16634 17200 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 109 nsew signal input
rlabel metal2 s 18786 16400 18842 17200 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 110 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 prog_clk_0_S_in
port 111 nsew signal input
rlabel metal3 s 0 144 800 264 6 prog_clk_0_W_out
port 112 nsew signal tristate
rlabel metal2 s 12162 16400 12218 17200 6 top_grid_pin_0_
port 113 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
