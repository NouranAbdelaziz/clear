* NGSPICE file created from sb_2__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt sb_2__1_ VGND VPWR bottom_left_grid_pin_42_ bottom_left_grid_pin_43_ bottom_left_grid_pin_44_
+ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_ bottom_left_grid_pin_47_ bottom_left_grid_pin_48_
+ bottom_left_grid_pin_49_ bottom_right_grid_pin_1_ ccff_head ccff_tail chanx_left_in[0]
+ chanx_left_in[10] chanx_left_in[11] chanx_left_in[12] chanx_left_in[13] chanx_left_in[14]
+ chanx_left_in[15] chanx_left_in[16] chanx_left_in[17] chanx_left_in[18] chanx_left_in[19]
+ chanx_left_in[1] chanx_left_in[2] chanx_left_in[3] chanx_left_in[4] chanx_left_in[5]
+ chanx_left_in[6] chanx_left_in[7] chanx_left_in[8] chanx_left_in[9] chanx_left_out[0]
+ chanx_left_out[10] chanx_left_out[11] chanx_left_out[12] chanx_left_out[13] chanx_left_out[14]
+ chanx_left_out[15] chanx_left_out[16] chanx_left_out[17] chanx_left_out[18] chanx_left_out[19]
+ chanx_left_out[1] chanx_left_out[2] chanx_left_out[3] chanx_left_out[4] chanx_left_out[5]
+ chanx_left_out[6] chanx_left_out[7] chanx_left_out[8] chanx_left_out[9] chany_bottom_in[0]
+ chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13]
+ chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17]
+ chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3]
+ chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8]
+ chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12]
+ chany_top_in[13] chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17]
+ chany_top_in[18] chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3]
+ chany_top_in[4] chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8]
+ chany_top_in[9] chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12]
+ chany_top_out[13] chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17]
+ chany_top_out[18] chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3]
+ chany_top_out[4] chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8]
+ chany_top_out[9] left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_
+ left_bottom_grid_pin_37_ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_
+ left_bottom_grid_pin_41_ prog_clk_0_N_in top_left_grid_pin_42_ top_left_grid_pin_43_
+ top_left_grid_pin_44_ top_left_grid_pin_45_ top_left_grid_pin_46_ top_left_grid_pin_47_
+ top_left_grid_pin_48_ top_left_grid_pin_49_ top_right_grid_pin_1_
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold42/X VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_3.mux_l1_in_1_ input3/X input1/X hold34/A VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__124__A _124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__119__A _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input55_A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_114_ _114_/A VGND VGND VPWR VPWR _114_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_17.mux_l1_in_0_ _104_/A _095_/A mux_bottom_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__dfxtp_1
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_20_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input18_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput97 _083_/X VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
XFILLER_16_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _087_/A sky130_fd_sc_hd__clkbuf_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_input85_A top_left_grid_pin_48_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_3.mux_l1_in_0_ _100_/A _091_/A hold34/A VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_33.mux_l2_in_1__179 VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_1_/A0
+ mux_bottom_track_33.mux_l2_in_1__179/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_0.mux_l1_in_0__A1 input79/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input48_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _070_/A sky130_fd_sc_hd__clkbuf_1
X_113_ _113_/A VGND VGND VPWR VPWR _113_/X sky130_fd_sc_hd__clkbuf_1
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_left_track_31.sky130_fd_sc_hd__buf_4_0_ mux_left_track_31.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__clkbuf_1
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_20_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold24/X VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__dfxtp_1
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_7.mux_l1_in_3_ mux_left_track_7.mux_l1_in_3_/A0 input78/X mux_left_track_7.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput98 _084_/X VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
XFILLER_16_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input30_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__clkbuf_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_15.mux_l3_in_0_ mux_left_track_15.mux_l2_in_1_/X mux_left_track_15.mux_l2_in_0_/X
+ hold42/A VGND VGND VPWR VPWR mux_left_track_15.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_3_ mux_top_track_0.mux_l2_in_3_/A0 input16/X mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_26_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input78_A left_bottom_grid_pin_41_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_19.sky130_fd_sc_hd__buf_4_0_ mux_left_track_19.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _075_/A sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_15.mux_l2_in_1_ mux_left_track_15.mux_l2_in_1_/A0 input74/X hold11/A
+ VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_7.mux_l3_in_0_ mux_left_track_7.mux_l2_in_1_/X mux_left_track_7.mux_l2_in_0_/X
+ hold28/A VGND VGND VPWR VPWR mux_left_track_7.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_0.mux_l4_in_0_ mux_top_track_0.mux_l3_in_1_/X mux_top_track_0.mux_l3_in_0_/X
+ hold22/A VGND VGND VPWR VPWR mux_top_track_0.mux_l4_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__dfxtp_1
X_112_ _112_/A VGND VGND VPWR VPWR _112_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_7.mux_l2_in_1_ mux_left_track_7.mux_l1_in_3_/X mux_left_track_7.mux_l1_in_2_/X
+ mux_left_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input60_A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ hold14/X VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_0.mux_l3_in_1_ mux_top_track_0.mux_l2_in_3_/X mux_top_track_0.mux_l2_in_2_/X
+ mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__dfxtp_1
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold35/X VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_7.mux_l1_in_2_ input76/X input74/X mux_left_track_7.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xoutput99 _085_/X VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
Xoutput88 output88/A VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_2
XFILLER_25_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input23_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_2_ input28/X input11/X mux_top_track_0.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ hold34/X VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_15.mux_l2_in_0_ input41/X mux_left_track_15.mux_l1_in_0_/X hold11/A
+ VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xprog_clk_0_FTB00 prog_clk_0_N_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_9.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
X_111_ _111_/A VGND VGND VPWR VPWR _111_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input53_A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_7.mux_l2_in_0_ mux_left_track_7.mux_l1_in_1_/X mux_left_track_7.mux_l1_in_0_/X
+ mux_left_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_0.mux_l3_in_0_ mux_top_track_0.mux_l2_in_1_/X mux_top_track_0.mux_l2_in_0_/X
+ mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_19_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_16.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput89 _066_/X VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
XFILLER_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_7.mux_l1_in_1_ _079_/A _113_/A mux_left_track_7.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_1_ _119_/A mux_top_track_0.mux_l1_in_2_/X mux_top_track_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input16_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xrepeater150 repeater150/A VGND VGND VPWR VPWR repeater150/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input8_A bottom_left_grid_pin_49_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold30/X VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input83_A top_left_grid_pin_46_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_0.mux_l1_in_2_ _109_/A input87/X mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_16.sky130_fd_sc_hd__buf_4_0_ mux_top_track_16.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _114_/A sky130_fd_sc_hd__clkbuf_1
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold25/X VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_15.mux_l1_in_0_ _119_/A _099_/A hold45/A VGND VGND VPWR VPWR mux_left_track_15.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_110_ _110_/A VGND VGND VPWR VPWR _110_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input46_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_4_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ hold4/X VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_9.mux_l2_in_3_ mux_bottom_track_9.mux_l2_in_3_/A0 input20/X mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_0.sky130_fd_sc_hd__buf_4_0_ mux_top_track_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _106_/A sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_7.mux_l1_in_0_ input44/X _093_/A mux_left_track_7.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_0.mux_l2_in_0_ mux_top_track_0.mux_l1_in_1_/X mux_top_track_0.mux_l1_in_0_/X
+ mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_1.mux_l1_in_1__A1 _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xrepeater151 repeater152/X VGND VGND VPWR VPWR repeater151/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_0.mux_l1_in_1_ input85/X input83/X mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.mux_l4_in_0_ mux_bottom_track_9.mux_l3_in_1_/X mux_bottom_track_9.mux_l3_in_0_/X
+ hold38/A VGND VGND VPWR VPWR mux_bottom_track_9.mux_l4_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_21.mux_l1_in_1_/S VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_39.mux_l2_in_0__164 VGND VGND VPWR VPWR mux_left_track_39.mux_l2_in_0_/A0
+ mux_left_track_39.mux_l2_in_0__164/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A0 _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input76_A left_bottom_grid_pin_39_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__091__A _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold15/X VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_9.mux_l3_in_1_ mux_bottom_track_9.mux_l2_in_3_/X mux_bottom_track_9.mux_l2_in_2_/X
+ mux_bottom_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_input39_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_bottom_track_9.mux_l2_in_2_ input13/X input25/X mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_39.mux_l2_in_0_ mux_left_track_39.mux_l2_in_0_/A0 mux_left_track_39.mux_l1_in_0_/X
+ output88/A VGND VGND VPWR VPWR mux_left_track_39.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xrepeater152 repeater152/A VGND VGND VPWR VPWR repeater152/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A0 _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_33.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _102_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input21_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_25.mux_l3_in_0_ mux_bottom_track_25.mux_l2_in_1_/X mux_bottom_track_25.mux_l2_in_0_/X
+ hold40/A VGND VGND VPWR VPWR mux_bottom_track_25.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_15.mux_l1_in_0__A0 _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__089__A _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input69_A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold26/X VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_0.mux_l1_in_0_ input81/X input79/X mux_top_track_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_17.mux_l1_in_0__A1 _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_25.mux_l2_in_1_ mux_bottom_track_25.mux_l2_in_1_/A0 mux_bottom_track_25.mux_l1_in_2_/X
+ mux_bottom_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.mux_l3_in_0_ mux_bottom_track_9.mux_l2_in_1_/X mux_bottom_track_9.mux_l2_in_0_/X
+ mux_bottom_track_9.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_9.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_17.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
X_099_ _099_/A VGND VGND VPWR VPWR _099_/X sky130_fd_sc_hd__clkbuf_1
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_mux_top_track_4.mux_l1_in_2__A1 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_3.mux_l1_in_2__A0 input76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input51_A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_25.mux_l1_in_2_ input15/X input27/X mux_bottom_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA__097__A _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l2_in_1_ input8/X input4/X mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_23.mux_l1_in_0__A0 _124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A0 _124_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_bottom_track_25.mux_l1_in_0__A1 _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input14_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_1__157 VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/A0
+ mux_left_track_25.mux_l1_in_1__157/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_15.mux_l1_in_0__A1 _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input6_A bottom_left_grid_pin_47_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_39.mux_l1_in_0_ input78/X input62/X hold20/A VGND VGND VPWR VPWR mux_left_track_39.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input81_A top_left_grid_pin_44_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A1 _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ mux_bottom_track_25.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold38/X VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_24_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_098_ _098_/A VGND VGND VPWR VPWR _098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_13.mux_l2_in_1__A1 input73/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_3.mux_l1_in_2__A1 input74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_24.mux_l1_in_1__A0 _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input44_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_bottom_track_25.mux_l1_in_1_ input6/X input2/X mux_bottom_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_9.mux_l2_in_0_ input9/X mux_bottom_track_9.mux_l1_in_0_/X mux_bottom_track_9.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_31.mux_l1_in_0__A0 input74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_33.mux_l1_in_0__A1 _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_16.mux_l1_in_1__A1 _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_16.mux_l1_in_3_ mux_top_track_16.mux_l1_in_3_/A0 input19/X mux_top_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_23.mux_l1_in_0__A1 _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _068_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_16.mux_l1_in_3__169 VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_3_/A0
+ mux_top_track_16.mux_l1_in_3__169/LO sky130_fd_sc_hd__conb_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_16.mux_l3_in_0_ mux_top_track_16.mux_l2_in_1_/X mux_top_track_16.mux_l2_in_0_/X
+ hold29/A VGND VGND VPWR VPWR mux_top_track_16.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_21.sky130_fd_sc_hd__buf_4_0_ mux_left_track_21.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _076_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input74_A left_bottom_grid_pin_37_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_5__A0 input26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_3.mux_l1_in_3_ mux_left_track_3.mux_l1_in_3_/A0 input78/X mux_left_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_5.mux_l2_in_3__180 VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_3_/A0
+ mux_bottom_track_5.mux_l2_in_3__180/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_11.mux_l3_in_0_ mux_left_track_11.mux_l2_in_1_/X mux_left_track_11.mux_l2_in_0_/X
+ hold5/A VGND VGND VPWR VPWR mux_left_track_11.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.mux_l2_in_1_ mux_top_track_16.mux_l1_in_3_/X mux_top_track_16.mux_l1_in_2_/X
+ mux_top_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_097_ _097_/A VGND VGND VPWR VPWR _097_/X sky130_fd_sc_hd__clkbuf_1
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_left_track_15.sky130_fd_sc_hd__buf_4_0_ mux_left_track_15.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _073_/A sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_24.mux_l1_in_1__A1 _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_bottom_track_25.mux_l1_in_0_ _105_/A _096_/A mux_bottom_track_25.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input37_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_139 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_11.mux_l2_in_1_ mux_left_track_11.mux_l2_in_1_/A0 _079_/A mux_left_track_11.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_16.mux_l1_in_2_ input12/X input24/X mux_top_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ hold43/A VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_9.mux_l1_in_0_ _103_/A _093_/A hold25/A VGND VGND VPWR VPWR mux_bottom_track_9.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _090_/A sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_13.mux_l2_in_1_/S VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_3.mux_l2_in_1_ mux_left_track_3.mux_l1_in_3_/X mux_left_track_3.mux_l1_in_2_/X
+ hold9/A VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input67_A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__100__A _100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_4.mux_l1_in_5__A1 _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l1_in_2_ input76/X input74/X mux_left_track_3.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_32.mux_l1_in_1__A1 _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_16.mux_l2_in_0_ mux_top_track_16.mux_l1_in_1_/X mux_top_track_16.mux_l1_in_0_/X
+ mux_top_track_16.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_16.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_096_ _096_/A VGND VGND VPWR VPWR _096_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__dfxtp_1
XFILLER_6_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ repeater149/X VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_27_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_bottom_track_5.mux_l1_in_6_ input19/X input12/X repeater152/A VGND VGND VPWR
+ VPWR mux_bottom_track_5.mux_l1_in_6_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_17.mux_l1_in_1__A1 input75/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_079_ _079_/A VGND VGND VPWR VPWR _079_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_37.sky130_fd_sc_hd__buf_4_0_ mux_left_track_37.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _084_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_16.mux_l1_in_1_ _124_/A _115_/A mux_top_track_16.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_16.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_11.mux_l2_in_0_ input33/X mux_left_track_11.mux_l1_in_0_/X mux_left_track_11.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__103__A _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_7.mux_l1_in_1__A1 _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_3__A1 input20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ hold33/X VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ hold44/X VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ hold9/A VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input12_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_3__A1 input77/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input4_A bottom_left_grid_pin_45_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_3.mux_l1_in_1_ _079_/A _111_/A mux_left_track_3.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA__111__A _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_1__A1 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_095_ _095_/A VGND VGND VPWR VPWR _095_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_7.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_6_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ hold17/X VGND VGND VPWR VPWR repeater150/A sky130_fd_sc_hd__dfxtp_1
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_27_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_5.mux_l1_in_5_ input24/X input8/X repeater152/X VGND VGND VPWR VPWR
+ mux_bottom_track_5.mux_l1_in_5_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_078_ _078_/A VGND VGND VPWR VPWR _078_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_7.mux_l1_in_3__166 VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_3_/A0
+ mux_left_track_7.mux_l1_in_3__166/LO sky130_fd_sc_hd__conb_1
Xmux_top_track_16.mux_l1_in_0_ input84/X input80/X mux_top_track_16.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_16.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input42_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ hold5/X VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_11.mux_l1_in_0_ _116_/A _096_/A hold18/A VGND VGND VPWR VPWR mux_left_track_11.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_192 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_23.mux_l2_in_0_ mux_left_track_23.mux_l1_in_1_/X mux_left_track_23.mux_l1_in_0_/X
+ hold36/A VGND VGND VPWR VPWR mux_left_track_23.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_37.mux_l2_in_0__163 VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/A0
+ mux_left_track_37.mux_l2_in_0__163/LO sky130_fd_sc_hd__conb_1
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__109__A _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_5.mux_l2_in_3_ mux_bottom_track_5.mux_l2_in_3_/A0 mux_bottom_track_5.mux_l1_in_6_/X
+ mux_bottom_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_3_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_23.mux_l1_in_1_ mux_left_track_23.mux_l1_in_1_/A0 input78/X mux_left_track_23.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l1_in_0_ input31/X _091_/A mux_left_track_3.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_19.mux_l1_in_1_/S VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_094_ _094_/A VGND VGND VPWR VPWR _094_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ hold48/X VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input72_A left_bottom_grid_pin_35_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_bottom_track_5.mux_l1_in_4_ input7/X input6/X repeater151/X VGND VGND VPWR VPWR
+ mux_bottom_track_5.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
X_077_ _077_/A VGND VGND VPWR VPWR _077_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_5.mux_l4_in_0_ mux_bottom_track_5.mux_l3_in_1_/X mux_bottom_track_5.mux_l3_in_0_/X
+ hold15/A VGND VGND VPWR VPWR mux_bottom_track_5.mux_l4_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA__117__A _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A0 _100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input35_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput80 top_left_grid_pin_43_ VGND VGND VPWR VPWR input80/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_29.mux_l1_in_0__A0 input73/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_5.mux_l3_in_1_ mux_bottom_track_5.mux_l2_in_3_/X mux_bottom_track_5.mux_l2_in_2_/X
+ mux_bottom_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_8.mux_l2_in_3__A1 input20/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_19.mux_l1_in_1__154 VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_1_/A0
+ mux_left_track_19.mux_l1_in_1__154/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_5.mux_l2_in_2_ mux_bottom_track_5.mux_l1_in_5_/X mux_bottom_track_5.mux_l1_in_4_/X
+ mux_bottom_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__125__A _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input65_A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_23.mux_l1_in_0_ _124_/A _104_/A mux_left_track_23.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_left_track_23.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold19/X VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_093_ _093_/A VGND VGND VPWR VPWR _093_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_35.mux_l2_in_0_ mux_left_track_35.mux_l2_in_0_/A0 mux_left_track_35.mux_l1_in_0_/X
+ hold37/A VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_5.mux_l1_in_3_ input5/X input4/X repeater151/X VGND VGND VPWR VPWR
+ mux_bottom_track_5.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xinput1 bottom_left_grid_pin_42_ VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_076_ _076_/A VGND VGND VPWR VPWR _076_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold1/X VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_37.mux_l1_in_0__A0 input77/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input28_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_bottom_track_3.mux_l1_in_0__A1 _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput70 chany_top_in[9] VGND VGND VPWR VPWR _096_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput81 top_left_grid_pin_44_ VGND VGND VPWR VPWR input81/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l2_in_1__A1 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _094_/A sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_23.mux_l1_in_1__156 VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_1_/A0
+ mux_left_track_23.mux_l1_in_1__156/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ mux_bottom_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_5.mux_l2_in_1_ mux_bottom_track_5.mux_l1_in_3_/X mux_bottom_track_5.mux_l1_in_2_/X
+ mux_bottom_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input10_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l3_in_1_/S VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_input2_A bottom_left_grid_pin_43_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input58_A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_092_ _092_/A VGND VGND VPWR VPWR _092_/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_5.mux_l1_in_2_ input3/X input2/X repeater151/X VGND VGND VPWR VPWR
+ mux_bottom_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 bottom_left_grid_pin_43_ VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_075_ _075_/A VGND VGND VPWR VPWR _075_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_0.mux_l2_in_3__168 VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_3_/A0
+ mux_top_track_0.mux_l2_in_3__168/LO sky130_fd_sc_hd__conb_1
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ hold31/X VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_35.mux_l1_in_0_ input76/X input68/X hold24/A VGND VGND VPWR VPWR mux_left_track_35.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_24_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xrepeater149 repeater150/X VGND VGND VPWR VPWR repeater149/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput60 chany_top_in[18] VGND VGND VPWR VPWR _105_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput82 top_left_grid_pin_45_ VGND VGND VPWR VPWR input82/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput71 left_bottom_grid_pin_34_ VGND VGND VPWR VPWR input71/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input40_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_33.mux_l3_in_0_ mux_bottom_track_33.mux_l2_in_1_/X mux_bottom_track_33.mux_l2_in_0_/X
+ hold44/A VGND VGND VPWR VPWR mux_bottom_track_33.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold41/X VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_top_track_0.mux_l1_in_2__A0 _109_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _066_/A sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_33.mux_l2_in_1_ mux_bottom_track_33.mux_l2_in_1_/A0 mux_bottom_track_33.mux_l1_in_2_/X
+ mux_bottom_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_25.mux_l2_in_1__177 VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_1_/A0
+ mux_bottom_track_25.mux_l2_in_1__177/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_0.mux_l2_in_1__A0 _119_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_091_ _091_/A VGND VGND VPWR VPWR _091_/X sky130_fd_sc_hd__clkbuf_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 bottom_left_grid_pin_44_ VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input70_A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_074_ _074_/A VGND VGND VPWR VPWR _074_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_11.mux_l1_in_0__A0 _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_5.mux_l1_in_1_ input1/X input9/X repeater152/X VGND VGND VPWR VPWR
+ mux_bottom_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_33.mux_l1_in_2_ input16/X input28/X mux_bottom_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput83 top_left_grid_pin_46_ VGND VGND VPWR VPWR input83/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_N_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput61 chany_top_in[19] VGND VGND VPWR VPWR input61/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_top_track_2.mux_l1_in_0__A1 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput50 chany_bottom_in[9] VGND VGND VPWR VPWR _116_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput72 left_bottom_grid_pin_35_ VGND VGND VPWR VPWR _079_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_20_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input33_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_109_ _109_/A VGND VGND VPWR VPWR _109_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold37/X VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_11.sky130_fd_sc_hd__buf_4_0_ mux_left_track_11.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _071_/A sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_17.mux_l1_in_3__176 VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_3_/A0
+ mux_bottom_track_17.mux_l1_in_3__176/LO sky130_fd_sc_hd__conb_1
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ repeater151/X VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_33.mux_l2_in_0_ mux_bottom_track_33.mux_l1_in_1_/X mux_bottom_track_33.mux_l1_in_0_/X
+ mux_bottom_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_090_ _090_/A VGND VGND VPWR VPWR _090_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_15.mux_l2_in_1__185 VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_1_/A0
+ mux_left_track_15.mux_l2_in_1__185/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _088_/A sky130_fd_sc_hd__clkbuf_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 bottom_left_grid_pin_45_ VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_5.mux_l1_in_0_ _101_/A _092_/A repeater152/X VGND VGND VPWR VPWR
+ mux_bottom_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_33.mux_l1_in_1_ input11/X input7/X mux_bottom_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_073_ _073_/A VGND VGND VPWR VPWR _073_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input63_A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_11.mux_l1_in_0__A1 _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_125_ _125_/A VGND VGND VPWR VPWR _125_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput51 chany_top_in[0] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_1
Xinput84 top_left_grid_pin_47_ VGND VGND VPWR VPWR input84/X sky130_fd_sc_hd__clkbuf_1
Xinput62 chany_top_in[1] VGND VGND VPWR VPWR input62/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_24.mux_l1_in_3_ mux_top_track_24.mux_l1_in_3_/A0 input18/X mux_top_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xinput40 chany_bottom_in[18] VGND VGND VPWR VPWR _125_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput73 left_bottom_grid_pin_36_ VGND VGND VPWR VPWR input73/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input26_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_108_ _108_/A VGND VGND VPWR VPWR _108_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _082_/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_24.mux_l3_in_0_ mux_top_track_24.mux_l2_in_1_/X mux_top_track_24.mux_l2_in_0_/X
+ hold3/A VGND VGND VPWR VPWR mux_top_track_24.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ hold23/X VGND VGND VPWR VPWR repeater152/A sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_2.mux_l2_in_3_ mux_top_track_2.mux_l2_in_3_/A0 input15/X mux_top_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xinput5 bottom_left_grid_pin_46_ VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XFILLER_27_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_24.mux_l2_in_1_ mux_top_track_24.mux_l1_in_3_/X mux_top_track_24.mux_l1_in_2_/X
+ mux_top_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_33.mux_l1_in_0_ input3/X _097_/A mux_bottom_track_33.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input56_A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_072_ _072_/A VGND VGND VPWR VPWR _072_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_8.mux_l2_in_3__174 VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_3_/A0
+ mux_top_track_8.mux_l2_in_3__174/LO sky130_fd_sc_hd__conb_1
XFILLER_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_5.mux_l1_in_3__165 VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_3_/A0
+ mux_left_track_5.mux_l1_in_3__165/LO sky130_fd_sc_hd__conb_1
X_124_ _124_/A VGND VGND VPWR VPWR _124_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_9.mux_l3_in_0_ mux_left_track_9.mux_l2_in_1_/X mux_left_track_9.mux_l2_in_0_/X
+ hold12/A VGND VGND VPWR VPWR mux_left_track_9.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
Xinput85 top_left_grid_pin_48_ VGND VGND VPWR VPWR input85/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput52 chany_top_in[10] VGND VGND VPWR VPWR _097_/A sky130_fd_sc_hd__clkbuf_2
Xinput63 chany_top_in[2] VGND VGND VPWR VPWR _089_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_2.mux_l4_in_0_ mux_top_track_2.mux_l3_in_1_/X mux_top_track_2.mux_l3_in_0_/X
+ hold17/A VGND VGND VPWR VPWR mux_top_track_2.mux_l4_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_24.mux_l1_in_2_ input30/X input23/X mux_top_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xinput30 chanx_left_in[9] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_1
Xinput41 chany_bottom_in[19] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_1
Xinput74 left_bottom_grid_pin_37_ VGND VGND VPWR VPWR input74/X sky130_fd_sc_hd__clkbuf_2
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A0 _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_107_ _107_/A VGND VGND VPWR VPWR _107_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input19_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_35.mux_l2_in_0__162 VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/A0
+ mux_left_track_35.mux_l2_in_0__162/LO sky130_fd_sc_hd__conb_1
XFILLER_26_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_9.mux_l2_in_1_ mux_left_track_9.mux_l2_in_1_/A0 input71/X mux_left_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l3_in_1_ mux_top_track_2.mux_l2_in_3_/X mux_top_track_2.mux_l2_in_2_/X
+ mux_top_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input86_A top_left_grid_pin_49_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_2.mux_l2_in_2_ input27/X _120_/A mux_top_track_2.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA__092__A _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_23.mux_l1_in_1_/S VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_13.mux_l2_in_0__A0 input37/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l2_in_0_ mux_top_track_24.mux_l1_in_1_/X mux_top_track_24.mux_l1_in_0_/X
+ mux_top_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_10_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 bottom_left_grid_pin_47_ VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_071_ _071_/A VGND VGND VPWR VPWR _071_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_167 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input49_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l1_in_1_/X mux_left_track_17.mux_l1_in_0_/X
+ hold19/A VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xoutput140 _107_/X VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
XFILLER_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_123_ _123_/A VGND VGND VPWR VPWR _123_/X sky130_fd_sc_hd__clkbuf_1
Xinput20 chanx_left_in[18] VGND VGND VPWR VPWR input20/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_24.mux_l1_in_1_ _125_/A _116_/A mux_top_track_24.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_24.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xinput31 chany_bottom_in[0] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput64 chany_top_in[3] VGND VGND VPWR VPWR input64/X sky130_fd_sc_hd__clkbuf_1
Xinput53 chany_top_in[11] VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__clkbuf_1
Xinput86 top_left_grid_pin_49_ VGND VGND VPWR VPWR input86/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput75 left_bottom_grid_pin_38_ VGND VGND VPWR VPWR input75/X sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA_mux_bottom_track_9.mux_l1_in_0__A1 _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput42 chany_bottom_in[1] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_1
X_106_ _106_/A VGND VGND VPWR VPWR _106_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_17.mux_l1_in_1_ mux_left_track_17.mux_l1_in_1_/A0 input75/X mux_left_track_17.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_1.mux_l2_in_3_ mux_bottom_track_1.mux_l2_in_3_/A0 input17/X mux_bottom_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_2.mux_l2_in_2__A1 _120_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l2_in_0_ _115_/A mux_left_track_9.mux_l1_in_0_/X mux_left_track_9.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l3_in_0_ mux_top_track_2.mux_l2_in_1_/X mux_top_track_2.mux_l2_in_0_/X
+ mux_top_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA__095__A _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input31_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l2_in_1__167 VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_1_/A0
+ mux_left_track_9.mux_l2_in_1__167/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_1__153 VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_1_/A0
+ mux_left_track_17.mux_l1_in_1__153/LO sky130_fd_sc_hd__conb_1
XFILLER_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input79_A top_left_grid_pin_42_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_1.mux_l4_in_0_ mux_bottom_track_1.mux_l3_in_1_/X mux_bottom_track_1.mux_l3_in_0_/X
+ hold30/A VGND VGND VPWR VPWR mux_bottom_track_1.mux_l4_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_1_ _111_/A input86/X mux_top_track_2.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_2.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_3.mux_l1_in_1__A1 _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 bottom_left_grid_pin_48_ VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ hold10/X VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
X_070_ _070_/A VGND VGND VPWR VPWR _070_/X sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l3_in_1_/S VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_24.sky130_fd_sc_hd__buf_4_0_ mux_top_track_24.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _118_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_179 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_1.mux_l3_in_1_ mux_bottom_track_1.mux_l2_in_3_/X mux_bottom_track_1.mux_l2_in_2_/X
+ mux_bottom_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput130 _116_/X VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
Xoutput141 _108_/X VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_1.mux_l1_in_3__A1 input77/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_122_ _122_/A VGND VGND VPWR VPWR _122_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input61_A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_24.mux_l1_in_0_ input85/X input81/X mux_top_track_24.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_16.mux_l1_in_0__A1 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput87 top_right_grid_pin_1_ VGND VGND VPWR VPWR input87/X sky130_fd_sc_hd__clkbuf_1
Xinput54 chany_top_in[12] VGND VGND VPWR VPWR _099_/A sky130_fd_sc_hd__clkbuf_2
Xinput65 chany_top_in[4] VGND VGND VPWR VPWR _091_/A sky130_fd_sc_hd__clkbuf_2
Xinput21 chanx_left_in[19] VGND VGND VPWR VPWR input21/X sky130_fd_sc_hd__clkbuf_1
Xinput32 chany_bottom_in[10] VGND VGND VPWR VPWR _117_/A sky130_fd_sc_hd__clkbuf_2
Xinput43 chany_bottom_in[2] VGND VGND VPWR VPWR _109_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput76 left_bottom_grid_pin_39_ VGND VGND VPWR VPWR input76/X sky130_fd_sc_hd__clkbuf_2
Xinput10 ccff_head VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ hold16/X VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_32.mux_l2_in_1__172 VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/A0
+ mux_top_track_32.mux_l2_in_1__172/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_1.mux_l2_in_2_ input29/X input22/X mux_bottom_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
X_105_ _105_/A VGND VGND VPWR VPWR _105_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_21.mux_l1_in_1__155 VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_1_/A0
+ mux_left_track_21.mux_l1_in_1__155/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_17.mux_l1_in_0_ _120_/A _100_/A mux_left_track_17.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_top_track_8.mux_l1_in_0__A0 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_29.mux_l2_in_0_ mux_left_track_29.mux_l2_in_0_/A0 mux_left_track_29.mux_l1_in_0_/X
+ hold31/A VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_21.mux_l1_in_1__A1 input77/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_31.mux_l2_in_0_ mux_left_track_31.mux_l2_in_0_/A0 mux_left_track_31.mux_l1_in_0_/X
+ hold39/A VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input24_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_9.mux_l1_in_0_ input48/X _095_/A hold46/A VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_top_track_4.mux_l1_in_4__A0 _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_2.sky130_fd_sc_hd__buf_4_0_ mux_top_track_2.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _107_/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_2.mux_l2_in_0_ input84/X mux_top_track_2.mux_l1_in_0_/X mux_top_track_2.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 bottom_left_grid_pin_49_ VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_0__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput131 _117_/X VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
Xoutput142 _109_/X VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 _120_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_24.mux_l1_in_3__171 VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_3_/A0
+ mux_top_track_24.mux_l1_in_3__171/LO sky130_fd_sc_hd__conb_1
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ mux_bottom_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput120 _087_/X VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
X_121_ _121_/A VGND VGND VPWR VPWR _121_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input54_A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput66 chany_top_in[5] VGND VGND VPWR VPWR _092_/A sky130_fd_sc_hd__clkbuf_2
Xinput55 chany_top_in[13] VGND VGND VPWR VPWR _100_/A sky130_fd_sc_hd__clkbuf_2
Xinput44 chany_bottom_in[3] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_1
Xinput33 chany_bottom_in[11] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
Xinput77 left_bottom_grid_pin_40_ VGND VGND VPWR VPWR input77/X sky130_fd_sc_hd__clkbuf_2
Xinput22 chanx_left_in[1] VGND VGND VPWR VPWR input22/X sky130_fd_sc_hd__clkbuf_1
Xinput11 chanx_left_in[0] VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ hold32/X VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_top_track_8.mux_l1_in_0__A1 input79/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_bottom_track_17.mux_l1_in_2__A1 input26/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_104_ _104_/A VGND VGND VPWR VPWR _104_/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_1.mux_l2_in_1_ input8/X mux_bottom_track_1.mux_l1_in_2_/X mux_bottom_track_1.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input17_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_2__A0 input75/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input9_A bottom_right_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_1.mux_l1_in_2_ input6/X input4/X mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_29.mux_l1_in_0_ input73/X input61/X hold16/A VGND VGND VPWR VPWR mux_left_track_29.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_31.mux_l1_in_0_ input74/X input57/X hold1/A VGND VGND VPWR VPWR mux_left_track_31.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 _125_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input84_A top_left_grid_pin_47_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ hold9/X VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__dfxtp_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 bottom_right_grid_pin_1_ VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__clkbuf_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_0.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_track_0.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
Xoutput132 _118_/X VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
Xoutput143 _110_/X VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
XANTENNA_mux_left_track_17.mux_l1_in_0__A1 _100_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_top_track_2.mux_l1_in_0_ input82/X input80/X hold7/A VGND VGND VPWR VPWR mux_top_track_2.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput110 _096_/X VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
Xoutput121 _088_/X VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
X_120_ _120_/A VGND VGND VPWR VPWR _120_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input47_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput67 chany_top_in[6] VGND VGND VPWR VPWR _093_/A sky130_fd_sc_hd__clkbuf_2
Xinput56 chany_top_in[14] VGND VGND VPWR VPWR _101_/A sky130_fd_sc_hd__clkbuf_2
Xinput23 chanx_left_in[2] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_1
Xinput34 chany_bottom_in[12] VGND VGND VPWR VPWR _119_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput45 chany_bottom_in[4] VGND VGND VPWR VPWR _111_/A sky130_fd_sc_hd__clkbuf_2
Xinput78 left_bottom_grid_pin_41_ VGND VGND VPWR VPWR input78/X sky130_fd_sc_hd__clkbuf_2
Xinput12 chanx_left_in[10] VGND VGND VPWR VPWR input12/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_103_ _103_/A VGND VGND VPWR VPWR _103_/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_7.mux_l1_in_0__A1 _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_9.mux_l2_in_2__A1 input25/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_mux_left_track_15.mux_l2_in_1__A1 input74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_1__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_3_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 input73/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_1.mux_l1_in_1_ input2/X input9/X mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 input75/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold11/X VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_13.mux_l2_in_1__184 VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_1_/A0
+ mux_left_track_13.mux_l2_in_1__184/LO sky130_fd_sc_hd__conb_1
XANTENNA__101__A _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input77_A left_bottom_grid_pin_40_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_25.mux_l1_in_0__A1 _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_3.mux_l1_in_3_/S VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dfxtp_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ input10/X VGND VGND VPWR VPWR mux_top_track_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_17_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput133 _119_/X VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
Xoutput144 _111_/X VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
Xoutput100 _067_/X VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
XFILLER_15_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput111 _097_/X VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
Xoutput122 _089_/X VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
XANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A mux_top_track_32.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput79 top_left_grid_pin_42_ VGND VGND VPWR VPWR input79/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput57 chany_top_in[15] VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_1
Xinput68 chany_top_in[7] VGND VGND VPWR VPWR input68/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput24 chanx_left_in[3] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_1
Xinput13 chanx_left_in[11] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_1
Xinput35 chany_bottom_in[13] VGND VGND VPWR VPWR _120_/A sky130_fd_sc_hd__clkbuf_2
Xinput46 chany_bottom_in[5] VGND VGND VPWR VPWR _112_/A sky130_fd_sc_hd__clkbuf_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_9.mux_l2_in_1_/S VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l4_in_0_/X VGND
+ VGND VPWR VPWR _086_/A sky130_fd_sc_hd__clkbuf_1
X_102_ _102_/A VGND VGND VPWR VPWR _102_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_31_206 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__104__A _104_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_1.mux_l1_in_0_ _099_/A _089_/A mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input22_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ hold45/X VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ hold8/X VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_7.sky130_fd_sc_hd__buf_4_0_ mux_left_track_7.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _069_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__112__A _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_161 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput134 _120_/X VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
Xoutput145 _112_/X VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
Xoutput101 _068_/X VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
Xclkbuf_0_mem_bottom_track_1.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_bottom_track_1.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
Xoutput112 _098_/X VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
Xoutput123 _090_/X VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
XFILLER_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_164 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput14 chanx_left_in[12] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_1
Xinput25 chanx_left_in[4] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
Xinput36 chany_bottom_in[14] VGND VGND VPWR VPWR _121_/A sky130_fd_sc_hd__clkbuf_2
Xinput58 chany_top_in[16] VGND VGND VPWR VPWR _103_/A sky130_fd_sc_hd__clkbuf_2
Xinput69 chany_top_in[8] VGND VGND VPWR VPWR _095_/A sky130_fd_sc_hd__clkbuf_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ hold46/X VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xinput47 chany_bottom_in[6] VGND VGND VPWR VPWR _113_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA_input52_A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_9.mux_l2_in_0__A0 _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_101_ _101_/A VGND VGND VPWR VPWR _101_/X sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_2__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
Xmux_left_track_23.sky130_fd_sc_hd__buf_4_0_ mux_left_track_23.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_5.mux_l1_in_3_ mux_left_track_5.mux_l1_in_3_/A0 input77/X mux_left_track_5.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_33.mux_l2_in_0__161 VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/A0
+ mux_left_track_33.mux_l2_in_0__161/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_13.mux_l3_in_0_ mux_left_track_13.mux_l2_in_1_/X mux_left_track_13.mux_l2_in_0_/X
+ hold13/A VGND VGND VPWR VPWR mux_left_track_13.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_8.mux_l2_in_2__A1 input25/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__120__A _120_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _074_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input15_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__115__A _115_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_19.mux_l1_in_1__A1 input76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_13.mux_l2_in_1_ mux_left_track_13.mux_l2_in_1_/A0 input73/X mux_left_track_13.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ hold13/X VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ hold48/A VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input7_A bottom_left_grid_pin_48_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_173 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input82_A top_left_grid_pin_45_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput135 _121_/X VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
Xoutput146 _113_/X VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
Xoutput102 _069_/X VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
Xoutput113 _099_/X VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
Xoutput124 _091_/X VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l1_in_3_/X mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xinput59 chany_top_in[17] VGND VGND VPWR VPWR _104_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__123__A _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput15 chanx_left_in[13] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_176 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput48 chany_bottom_in[7] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_7.mux_l1_in_3__A1 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput37 chany_bottom_in[15] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
Xinput26 chanx_left_in[5] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_1
X_100_ _100_/A VGND VGND VPWR VPWR _100_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ hold28/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_input45_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_2_ input75/X input73/X mux_left_track_5.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_top_track_32.mux_l3_in_0_ mux_top_track_32.mux_l2_in_1_/X mux_top_track_32.mux_l2_in_0_/X
+ hold2/A VGND VGND VPWR VPWR mux_top_track_32.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l2_in_3_ mux_top_track_8.mux_l2_in_3_/A0 input20/X mux_top_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_3.mux_l2_in_3__178 VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_3_/A0
+ mux_bottom_track_3.mux_l2_in_3__178/LO sky130_fd_sc_hd__conb_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l3_in_1_/S VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_13.mux_l2_in_0_ input37/X mux_left_track_13.mux_l1_in_0_/X mux_left_track_13.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_39.sky130_fd_sc_hd__buf_4_0_ mux_left_track_39.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _085_/A sky130_fd_sc_hd__clkbuf_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_32.mux_l2_in_1_ mux_top_track_32.mux_l2_in_1_/A0 mux_top_track_32.mux_l1_in_2_/X
+ mux_top_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input75_A left_bottom_grid_pin_38_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput136 _122_/X VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
Xoutput147 _114_/X VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
Xoutput103 _070_/X VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
Xclkbuf_3_3__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
Xoutput125 _092_/X VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
Xoutput114 _100_/X VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l4_in_0_ mux_top_track_8.mux_l3_in_1_/X mux_top_track_8.mux_l3_in_0_/X
+ hold4/A VGND VGND VPWR VPWR mux_top_track_8.mux_l4_in_0_/X sky130_fd_sc_hd__mux2_1
Xinput16 chanx_left_in[14] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_top_track_32.mux_l1_in_2_ input17/X input29/X mux_top_track_32.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xinput38 chany_bottom_in[16] VGND VGND VPWR VPWR _123_/A sky130_fd_sc_hd__clkbuf_2
Xinput49 chany_bottom_in[8] VGND VGND VPWR VPWR _115_/A sky130_fd_sc_hd__clkbuf_2
Xinput27 chanx_left_in[6] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input38_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_1_ input71/X _112_/A mux_left_track_5.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_top_track_8.mux_l3_in_1_ mux_top_track_8.mux_l2_in_3_/X mux_top_track_8.mux_l2_in_2_/X
+ mux_top_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold47/X VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__dfxtp_1
XFILLER_22_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_top_track_8.mux_l2_in_2_ input13/X input25/X mux_top_track_8.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_30_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input20_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A0 _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_32.mux_l2_in_0_ mux_top_track_32.mux_l1_in_1_/X mux_top_track_32.mux_l1_in_0_/X
+ mux_top_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput137 _123_/X VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
Xoutput148 _115_/X VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
XANTENNA_input68_A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput104 _071_/X VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
Xmux_left_track_13.mux_l1_in_0_ _117_/A _097_/A hold33/A VGND VGND VPWR VPWR mux_left_track_13.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l1_in_3__182 VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_3_/A0
+ mux_left_track_1.mux_l1_in_3__182/LO sky130_fd_sc_hd__conb_1
Xoutput126 _093_/X VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
Xoutput115 _101_/X VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ hold32/A VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xinput17 chanx_left_in[15] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_32.mux_l1_in_1_ input22/X _117_/A mux_top_track_32.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_top_track_32.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xinput39 chany_bottom_in[17] VGND VGND VPWR VPWR _124_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput28 chanx_left_in[7] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_5.mux_l1_in_0_ input42/X _092_/A mux_left_track_5.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_25.mux_l1_in_1_ mux_left_track_25.mux_l1_in_1_/A0 input71/X mux_left_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_170 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_089_ _089_/A VGND VGND VPWR VPWR _089_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold39/X VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__dfxtp_1
Xmux_top_track_8.mux_l3_in_0_ mux_top_track_8.mux_l2_in_1_/X mux_top_track_8.mux_l2_in_0_/X
+ mux_top_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_0.mux_l1_in_1__A1 input83/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input50_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_8.mux_l2_in_1_ _123_/A _113_/A mux_top_track_8.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_top_track_8.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_39.mux_l1_in_0__A0 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XANTENNA_input13_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_bottom_track_5.mux_l1_in_0__A1 _092_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold20/X VGND VGND VPWR VPWR output88/A sky130_fd_sc_hd__dfxtp_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input5_A bottom_left_grid_pin_46_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput138 _124_/X VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
Xoutput105 _072_/X VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
Xoutput127 _094_/X VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
Xoutput116 _102_/X VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input80_A top_left_grid_pin_43_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput18 chanx_left_in[16] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput29 chanx_left_in[8] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_32.mux_l1_in_0_ input86/X input82/X mux_top_track_32.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_0_ _125_/A _105_/A mux_left_track_25.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_182 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_088_ _088_/A VGND VGND VPWR VPWR _088_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_37.mux_l2_in_0_ mux_left_track_37.mux_l2_in_0_/A0 mux_left_track_37.mux_l1_in_0_/X
+ hold21/A VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input43_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_8.mux_l2_in_0_ input87/X mux_top_track_8.mux_l1_in_0_/X mux_top_track_8.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold2/X VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l3_in_0_/X
+ VGND VGND VPWR VPWR _098_/A sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold21/X VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_11.mux_l2_in_1__183 VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_1_/A0
+ mux_left_track_11.mux_l2_in_1__183/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_top_track_4.mux_l1_in_0__A0 input80/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.sky130_fd_sc_hd__buf_4_0_ mux_top_track_8.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _110_/A sky130_fd_sc_hd__clkbuf_1
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput139 _125_/X VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
Xoutput106 _073_/X VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
XFILLER_23_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput128 _095_/X VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
Xoutput117 _103_/X VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 chanx_left_in[17] VGND VGND VPWR VPWR input19/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input73_A left_bottom_grid_pin_36_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_087_ _087_/A VGND VGND VPWR VPWR _087_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_2.mux_l2_in_1__A0 _111_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_5__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_16_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input36_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0__A0 _117_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_37.mux_l1_in_0_ input77/X input64/X hold41/A VGND VGND VPWR VPWR mux_left_track_37.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_1.mux_l2_in_3__175 VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_3_/A0
+ mux_bottom_track_1.mux_l2_in_3__175/LO sky130_fd_sc_hd__conb_1
XFILLER_30_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_208 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_top_track_4.mux_l1_in_0__A1 input79/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_8.mux_l1_in_0_ input83/X input79/X hold6/A VGND VGND VPWR VPWR mux_top_track_8.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput129 _106_/X VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
Xoutput107 _074_/X VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
Xmux_left_track_3.mux_l1_in_3__159 VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_3_/A0
+ mux_left_track_3.mux_l1_in_3__159/LO sky130_fd_sc_hd__conb_1
Xoutput118 _104_/X VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_1.mux_l1_in_2__A0 input75/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l2_in_1_/S VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_input66_A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_086_ _086_/A VGND VGND VPWR VPWR _086_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_31.mux_l2_in_0__160 VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/A0
+ mux_left_track_31.mux_l2_in_0__160/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _067_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_21.mux_l1_in_0__A0 _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_069_ _069_/A VGND VGND VPWR VPWR _069_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input29_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_13.mux_l1_in_0__A1 _097_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l1_in_6_ input21/X input14/X repeater150/A VGND VGND VPWR VPWR
+ mux_top_track_4.mux_l1_in_6_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_3.mux_l1_in_0__A1 _091_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_top_track_4.mux_l2_in_3__173 VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_3_/A0
+ mux_top_track_4.mux_l2_in_3__173/LO sky130_fd_sc_hd__conb_1
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__093__A _093_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput108 _075_/X VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
Xoutput90 _076_/X VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
Xmux_left_track_1.mux_l1_in_3_ mux_left_track_1.mux_l1_in_3_/A0 input77/X mux_left_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xoutput119 _105_/X VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input11_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_13.sky130_fd_sc_hd__buf_4_0_ mux_left_track_13.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _072_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_1.mux_l1_in_2__A1 input73/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_32.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_top_track_32.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input3_A bottom_left_grid_pin_44_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input59_A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_6__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_13_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_25.mux_l1_in_1_/S VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_085_ _085_/A VGND VGND VPWR VPWR _085_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_21.mux_l1_in_0__A1 _103_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ hold8/A VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
X_068_ _068_/A VGND VGND VPWR VPWR _068_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l1_in_5_ input26/X _121_/A repeater150/X VGND VGND VPWR VPWR
+ mux_top_track_4.mux_l1_in_5_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input41_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__096__A _096_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_1_ mux_left_track_1.mux_l1_in_3_/X mux_left_track_1.mux_l1_in_2_/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_1.mux_l1_in_2_ input75/X input73/X mux_left_track_1.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xoutput109 _086_/X VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
XFILLER_1_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_194 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput91 _077_/X VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ hold3/X VGND VGND VPWR VPWR mux_top_track_32.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__099__A _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_084_ _084_/A VGND VGND VPWR VPWR _084_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ hold36/X VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_35.sky130_fd_sc_hd__buf_4_0_ mux_left_track_35.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _083_/A sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l3_in_1_/S VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input71_A left_bottom_grid_pin_34_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_39.mux_l2_in_0__S output88/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.mux_l2_in_3_ mux_top_track_4.mux_l2_in_3_/A0 mux_top_track_4.mux_l1_in_6_/X
+ mux_top_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_3_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_left_track_29.sky130_fd_sc_hd__buf_4_0_ mux_left_track_29.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _080_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_15.mux_l2_in_0__A0 input41/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_067_ _067_/A VGND VGND VPWR VPWR _067_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 input71/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.mux_l2_in_3__181 VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_3_/A0
+ mux_bottom_track_9.mux_l2_in_3__181/LO sky130_fd_sc_hd__conb_1
X_119_ _119_/A VGND VGND VPWR VPWR _119_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_4.mux_l1_in_4_ _112_/A input87/X repeater150/X VGND VGND VPWR VPWR
+ mux_top_track_4.mux_l1_in_4_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ mux_left_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input34_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l4_in_0_ mux_top_track_4.mux_l3_in_1_/X mux_top_track_4.mux_l3_in_0_/X
+ hold27/A VGND VGND VPWR VPWR mux_top_track_4.mux_l4_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_33.mux_l2_in_1_/S VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__dfxtp_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_7__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
Xmux_left_track_1.mux_l1_in_1_ input71/X _109_/A mux_left_track_1.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput92 _078_/X VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_4.mux_l3_in_1_ mux_top_track_4.mux_l2_in_3_/X mux_top_track_4.mux_l2_in_2_/X
+ mux_top_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input64_A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_083_ _083_/A VGND VGND VPWR VPWR _083_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_top_track_4.mux_l2_in_2_ mux_top_track_4.mux_l1_in_5_/X mux_top_track_4.mux_l1_in_4_/X
+ mux_top_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_2_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_2.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_2.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_21_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_066_ _066_/A VGND VGND VPWR VPWR _066_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_5.mux_l1_in_1__A1 _112_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_29.mux_l2_in_0__158 VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/A0
+ mux_left_track_29.mux_l2_in_0__158/LO sky130_fd_sc_hd__conb_1
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_118_ _118_/A VGND VGND VPWR VPWR _118_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_19.mux_l2_in_0_ mux_left_track_19.mux_l1_in_1_/X mux_left_track_19.mux_l1_in_0_/X
+ hold26/A VGND VGND VPWR VPWR mux_left_track_19.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l1_in_3_ input86/X input85/X repeater149/X VGND VGND VPWR VPWR
+ mux_top_track_4.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input27_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_21.mux_l2_in_0_ mux_left_track_21.mux_l1_in_1_/X mux_left_track_21.mux_l1_in_0_/X
+ hold10/A VGND VGND VPWR VPWR mux_left_track_21.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l3_in_1_/S VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_3.mux_l1_in_3__A1 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_11.mux_l2_in_1_/S VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_26_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_33.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_33.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_19.mux_l1_in_1_ mux_left_track_19.mux_l1_in_1_/A0 input76/X mux_left_track_19.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_3.mux_l2_in_3_ mux_bottom_track_3.mux_l2_in_3_/A0 input18/X mux_bottom_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_21.mux_l1_in_1_ mux_left_track_21.mux_l1_in_1_/A0 input77/X mux_left_track_21.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xoutput93 _079_/X VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
Xmux_left_track_1.mux_l1_in_0_ _089_/A input51/X mux_left_track_1.mux_l1_in_3_/S VGND
+ VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_23.mux_l1_in_1__A1 input78/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_top_track_4.mux_l3_in_0_ mux_top_track_4.mux_l2_in_1_/X mux_top_track_4.mux_l2_in_0_/X
+ mux_top_track_4.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input57_A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_082_ _082_/A VGND VGND VPWR VPWR _082_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_10_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_input1_A bottom_left_grid_pin_42_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_32.sky130_fd_sc_hd__buf_4_0_ mux_top_track_32.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _122_/A sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_4.mux_l2_in_1_ mux_top_track_4.mux_l1_in_3_/X mux_top_track_4.mux_l1_in_2_/X
+ mux_top_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ hold7/X VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_3.mux_l4_in_0_ mux_bottom_track_3.mux_l3_in_1_/X mux_bottom_track_3.mux_l3_in_0_/X
+ hold23/A VGND VGND VPWR VPWR mux_bottom_track_3.mux_l4_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_top_track_8.mux_l2_in_1__A0 _123_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_117_ _117_/A VGND VGND VPWR VPWR _117_/X sky130_fd_sc_hd__clkbuf_1
Xmux_top_track_4.mux_l1_in_2_ input84/X input83/X repeater150/X VGND VGND VPWR VPWR
+ mux_top_track_4.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l3_in_1_ mux_bottom_track_3.mux_l2_in_3_/X mux_bottom_track_3.mux_l2_in_2_/X
+ mux_bottom_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_output88_A output88/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_19.mux_l1_in_0__A0 _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_8.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_8.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_29_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ hold18/X VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_3_ mux_bottom_track_17.mux_l1_in_3_/A0 input21/X mux_bottom_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_3_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold40/X VGND VGND VPWR VPWR mux_bottom_track_33.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_19.mux_l1_in_0_ _121_/A _101_/A mux_left_track_19.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_left_track_19.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_top_track_2.mux_l2_in_3__170 VGND VGND VPWR VPWR mux_top_track_2.mux_l2_in_3_/A0
+ mux_top_track_2.mux_l2_in_3__170/LO sky130_fd_sc_hd__conb_1
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_2_ input30/X input23/X mux_bottom_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input87_A top_right_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput94 _080_/X VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
Xmux_left_track_21.mux_l1_in_0_ _123_/A _103_/A mux_left_track_21.mux_l1_in_1_/S VGND
+ VGND VPWR VPWR mux_left_track_21.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l2_in_1_/S VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l2_in_0_/A0 mux_left_track_33.mux_l1_in_0_/X
+ hold35/A VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_17.mux_l3_in_0_ mux_bottom_track_17.mux_l2_in_1_/X mux_bottom_track_17.mux_l2_in_0_/X
+ hold14/A VGND VGND VPWR VPWR mux_bottom_track_17.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_7.mux_l1_in_2__A0 input76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_081_ _081_/A VGND VGND VPWR VPWR _081_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_33_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l2_in_0_ mux_top_track_4.mux_l1_in_1_/X mux_top_track_4.mux_l1_in_0_/X
+ mux_top_track_4.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_top_track_4.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ hold22/X VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A0 _099_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_top_track_4.sky130_fd_sc_hd__buf_4_0_ mux_top_track_4.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR _108_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_top_track_8.mux_l2_in_1__A1 _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_17.mux_l2_in_1_ mux_bottom_track_17.mux_l1_in_3_/X mux_bottom_track_17.mux_l1_in_2_/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xmux_top_track_4.mux_l1_in_1_ input82/X input81/X repeater149/X VGND VGND VPWR VPWR
+ mux_top_track_4.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ mux_bottom_track_3.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_116_ _116_/A VGND VGND VPWR VPWR _116_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_mux_left_track_19.mux_l1_in_0__A1 _101_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__105__A _105_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ hold6/X VGND VGND VPWR VPWR mux_top_track_8.mux_l2_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_2_ input14/X input26/X mux_bottom_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ hold12/X VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_input32_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_3.mux_l2_in_1_ input7/X input5/X mux_bottom_track_3.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xoutput95 _081_/X VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
XFILLER_25_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ mux_top_track_24.mux_l1_in_3_/S VGND VGND VPWR VPWR mux_top_track_24.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_9.mux_l1_in_0__A1 _095_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__113__A _113_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_17.mux_l1_in_1_/S VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_mux_left_track_7.mux_l1_in_2__A1 input74/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_35.mux_l1_in_0__A0 input76/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_080_ _080_/A VGND VGND VPWR VPWR _080_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ hold43/X VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_33.mux_l1_in_0_ input75/X input53/X hold47/A VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_mux_bottom_track_1.mux_l1_in_0__A1 _089_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input62_A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l1_in_1_/X mux_bottom_track_17.mux_l1_in_0_/X
+ mux_bottom_track_17.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_2_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_top_track_4.mux_l1_in_0_ input80/X input79/X repeater149/X VGND VGND VPWR VPWR
+ mux_top_track_4.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA__121__A _121_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_115_ _115_/A VGND VGND VPWR VPWR _115_/X sky130_fd_sc_hd__clkbuf_1
Xmem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ hold27/X VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l1_in_1_ input5/X input1/X mux_bottom_track_17.mux_l1_in_3_/S
+ VGND VGND VPWR VPWR mux_bottom_track_17.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA__116__A _116_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input25_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_19_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ hold29/X VGND VGND VPWR VPWR mux_top_track_24.mux_l1_in_3_/S sky130_fd_sc_hd__dfxtp_1
Xoutput96 _082_/X VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

