magic
tech sky130A
magscale 1 2
timestamp 1650625948
<< viali >>
rect 3433 14569 3467 14603
rect 5733 14569 5767 14603
rect 7021 14569 7055 14603
rect 7389 14569 7423 14603
rect 8033 14569 8067 14603
rect 8677 14569 8711 14603
rect 9321 14569 9355 14603
rect 9965 14569 9999 14603
rect 10609 14569 10643 14603
rect 12265 14569 12299 14603
rect 12541 14569 12575 14603
rect 13185 14569 13219 14603
rect 6561 14501 6595 14535
rect 7849 14501 7883 14535
rect 8217 14501 8251 14535
rect 11713 14501 11747 14535
rect 1961 14433 1995 14467
rect 3157 14433 3191 14467
rect 4629 14433 4663 14467
rect 5273 14433 5307 14467
rect 14657 14433 14691 14467
rect 16773 14433 16807 14467
rect 17969 14433 18003 14467
rect 2237 14365 2271 14399
rect 2881 14365 2915 14399
rect 3617 14365 3651 14399
rect 4353 14365 4387 14399
rect 5549 14365 5583 14399
rect 5917 14365 5951 14399
rect 6009 14365 6043 14399
rect 6377 14365 6411 14399
rect 6837 14365 6871 14399
rect 7573 14365 7607 14399
rect 9137 14365 9171 14399
rect 9413 14365 9447 14399
rect 10057 14365 10091 14399
rect 10701 14365 10735 14399
rect 11529 14365 11563 14399
rect 11805 14365 11839 14399
rect 12173 14365 12207 14399
rect 12633 14365 12667 14399
rect 13277 14365 13311 14399
rect 14105 14365 14139 14399
rect 14381 14365 14415 14399
rect 15301 14365 15335 14399
rect 15577 14365 15611 14399
rect 16497 14365 16531 14399
rect 17049 14365 17083 14399
rect 17693 14365 17727 14399
rect 6193 14229 6227 14263
rect 7665 14229 7699 14263
rect 8953 14229 8987 14263
rect 9597 14229 9631 14263
rect 10241 14229 10275 14263
rect 10885 14229 10919 14263
rect 11989 14229 12023 14263
rect 12817 14229 12851 14263
rect 13461 14229 13495 14263
rect 14289 14229 14323 14263
rect 16267 14229 16301 14263
rect 2927 14025 2961 14059
rect 4353 14025 4387 14059
rect 4997 14025 5031 14059
rect 5365 14025 5399 14059
rect 6009 14025 6043 14059
rect 6561 14025 6595 14059
rect 7481 14025 7515 14059
rect 13645 14025 13679 14059
rect 14473 14025 14507 14059
rect 15209 14025 15243 14059
rect 15025 13957 15059 13991
rect 2237 13889 2271 13923
rect 3157 13889 3191 13923
rect 4537 13889 4571 13923
rect 4813 13889 4847 13923
rect 5181 13889 5215 13923
rect 5549 13889 5583 13923
rect 5917 13889 5951 13923
rect 6193 13889 6227 13923
rect 6377 13889 6411 13923
rect 6837 13889 6871 13923
rect 7021 13889 7055 13923
rect 7389 13889 7423 13923
rect 13829 13889 13863 13923
rect 14657 13889 14691 13923
rect 15485 13889 15519 13923
rect 16221 13889 16255 13923
rect 16497 13889 16531 13923
rect 1961 13821 1995 13855
rect 3801 13821 3835 13855
rect 4077 13821 4111 13855
rect 7113 13821 7147 13855
rect 16773 13821 16807 13855
rect 17049 13821 17083 13855
rect 17693 13821 17727 13855
rect 17969 13821 18003 13855
rect 5733 13753 5767 13787
rect 15301 13753 15335 13787
rect 4629 13685 4663 13719
rect 6653 13685 6687 13719
rect 3341 13481 3375 13515
rect 5457 13481 5491 13515
rect 5733 13481 5767 13515
rect 6837 13481 6871 13515
rect 15761 13481 15795 13515
rect 16405 13481 16439 13515
rect 16681 13481 16715 13515
rect 6009 13413 6043 13447
rect 6653 13413 6687 13447
rect 16313 13413 16347 13447
rect 3893 13345 3927 13379
rect 17601 13345 17635 13379
rect 1961 13277 1995 13311
rect 2237 13277 2271 13311
rect 2881 13277 2915 13311
rect 3157 13277 3191 13311
rect 3525 13277 3559 13311
rect 4629 13277 4663 13311
rect 5641 13277 5675 13311
rect 5917 13277 5951 13311
rect 6193 13277 6227 13311
rect 15945 13277 15979 13311
rect 17325 13277 17359 13311
rect 17693 13277 17727 13311
rect 17969 13277 18003 13311
rect 4169 13209 4203 13243
rect 6377 13209 6411 13243
rect 6561 13209 6595 13243
rect 16129 13209 16163 13243
rect 4077 13141 4111 13175
rect 4537 13141 4571 13175
rect 5273 13141 5307 13175
rect 5181 12937 5215 12971
rect 5917 12937 5951 12971
rect 16957 12937 16991 12971
rect 3608 12869 3642 12903
rect 6009 12869 6043 12903
rect 17233 12869 17267 12903
rect 17509 12869 17543 12903
rect 3157 12801 3191 12835
rect 3341 12801 3375 12835
rect 6377 12801 6411 12835
rect 1961 12733 1995 12767
rect 2237 12733 2271 12767
rect 2881 12733 2915 12767
rect 5273 12733 5307 12767
rect 5365 12733 5399 12767
rect 5733 12733 5767 12767
rect 16865 12733 16899 12767
rect 17693 12733 17727 12767
rect 17969 12733 18003 12767
rect 4721 12665 4755 12699
rect 17325 12665 17359 12699
rect 4813 12597 4847 12631
rect 4537 12393 4571 12427
rect 4905 12393 4939 12427
rect 17233 12393 17267 12427
rect 2237 12257 2271 12291
rect 2973 12257 3007 12291
rect 3893 12257 3927 12291
rect 17969 12257 18003 12291
rect 1961 12189 1995 12223
rect 3249 12189 3283 12223
rect 5089 12189 5123 12223
rect 5356 12189 5390 12223
rect 7757 12189 7791 12223
rect 16865 12189 16899 12223
rect 17601 12189 17635 12223
rect 17693 12189 17727 12223
rect 2789 12121 2823 12155
rect 3617 12121 3651 12155
rect 4169 12121 4203 12155
rect 8585 12121 8619 12155
rect 2329 12053 2363 12087
rect 2697 12053 2731 12087
rect 3341 12053 3375 12087
rect 4077 12053 4111 12087
rect 4629 12053 4663 12087
rect 6469 12053 6503 12087
rect 16957 12053 16991 12087
rect 17417 12053 17451 12087
rect 2421 11849 2455 11883
rect 3433 11849 3467 11883
rect 6622 11781 6656 11815
rect 17049 11781 17083 11815
rect 1961 11713 1995 11747
rect 2789 11713 2823 11747
rect 3525 11713 3559 11747
rect 5006 11713 5040 11747
rect 5273 11713 5307 11747
rect 6377 11713 6411 11747
rect 8401 11713 8435 11747
rect 17233 11713 17267 11747
rect 17509 11713 17543 11747
rect 17693 11713 17727 11747
rect 2237 11645 2271 11679
rect 2881 11645 2915 11679
rect 3065 11645 3099 11679
rect 17969 11645 18003 11679
rect 3709 11577 3743 11611
rect 16405 11577 16439 11611
rect 16865 11577 16899 11611
rect 3893 11509 3927 11543
rect 7757 11509 7791 11543
rect 9045 11509 9079 11543
rect 16129 11509 16163 11543
rect 17417 11509 17451 11543
rect 2513 11305 2547 11339
rect 3433 11305 3467 11339
rect 3801 11305 3835 11339
rect 4353 11305 4387 11339
rect 12265 11305 12299 11339
rect 17233 11305 17267 11339
rect 3617 11237 3651 11271
rect 4537 11237 4571 11271
rect 6561 11237 6595 11271
rect 15761 11237 15795 11271
rect 16037 11237 16071 11271
rect 2973 11169 3007 11203
rect 3065 11169 3099 11203
rect 4169 11169 4203 11203
rect 5181 11169 5215 11203
rect 6101 11169 6135 11203
rect 17969 11169 18003 11203
rect 1961 11101 1995 11135
rect 2237 11101 2271 11135
rect 3985 11101 4019 11135
rect 4905 11101 4939 11135
rect 5825 11101 5859 11135
rect 8125 11101 8159 11135
rect 10333 11101 10367 11135
rect 11897 11101 11931 11135
rect 13921 11101 13955 11135
rect 15485 11101 15519 11135
rect 15945 11101 15979 11135
rect 17601 11101 17635 11135
rect 17693 11101 17727 11135
rect 2881 11033 2915 11067
rect 5917 11033 5951 11067
rect 7858 11033 7892 11067
rect 10088 11033 10122 11067
rect 11652 11033 11686 11067
rect 13654 11033 13688 11067
rect 16497 11033 16531 11067
rect 16957 11033 16991 11067
rect 2421 10965 2455 10999
rect 4997 10965 5031 10999
rect 5457 10965 5491 10999
rect 6285 10965 6319 10999
rect 6745 10965 6779 10999
rect 8953 10965 8987 10999
rect 10517 10965 10551 10999
rect 12541 10965 12575 10999
rect 16221 10965 16255 10999
rect 16681 10965 16715 10999
rect 17141 10965 17175 10999
rect 17417 10965 17451 10999
rect 1961 10761 1995 10795
rect 2513 10761 2547 10795
rect 4629 10761 4663 10795
rect 5089 10761 5123 10795
rect 5457 10761 5491 10795
rect 5825 10761 5859 10795
rect 8401 10761 8435 10795
rect 11897 10761 11931 10795
rect 12357 10761 12391 10795
rect 12725 10761 12759 10795
rect 12817 10761 12851 10795
rect 13185 10761 13219 10795
rect 13553 10761 13587 10795
rect 14289 10761 14323 10795
rect 3626 10693 3660 10727
rect 4997 10693 5031 10727
rect 7288 10693 7322 10727
rect 14657 10693 14691 10727
rect 16681 10693 16715 10727
rect 17141 10693 17175 10727
rect 1593 10625 1627 10659
rect 2053 10625 2087 10659
rect 5917 10625 5951 10659
rect 7021 10625 7055 10659
rect 9045 10625 9079 10659
rect 10425 10625 10459 10659
rect 13645 10625 13679 10659
rect 14013 10625 14047 10659
rect 15577 10625 15611 10659
rect 15669 10625 15703 10659
rect 17233 10625 17267 10659
rect 1869 10557 1903 10591
rect 3893 10557 3927 10591
rect 5273 10557 5307 10591
rect 6101 10557 6135 10591
rect 10517 10557 10551 10591
rect 10701 10557 10735 10591
rect 11161 10557 11195 10591
rect 11989 10557 12023 10591
rect 12081 10557 12115 10591
rect 12909 10557 12943 10591
rect 13737 10557 13771 10591
rect 15761 10557 15795 10591
rect 16957 10557 16991 10591
rect 17693 10557 17727 10591
rect 17969 10557 18003 10591
rect 4077 10489 4111 10523
rect 9689 10489 9723 10523
rect 14841 10489 14875 10523
rect 15209 10489 15243 10523
rect 16037 10489 16071 10523
rect 16497 10489 16531 10523
rect 1409 10421 1443 10455
rect 2421 10421 2455 10455
rect 10057 10421 10091 10455
rect 11529 10421 11563 10455
rect 15025 10421 15059 10455
rect 16313 10421 16347 10455
rect 17601 10421 17635 10455
rect 2789 10217 2823 10251
rect 4629 10217 4663 10251
rect 4813 10217 4847 10251
rect 10517 10217 10551 10251
rect 11345 10217 11379 10251
rect 12173 10217 12207 10251
rect 17049 10217 17083 10251
rect 4445 10149 4479 10183
rect 6469 10149 6503 10183
rect 9597 10149 9631 10183
rect 2053 10081 2087 10115
rect 3433 10081 3467 10115
rect 5273 10081 5307 10115
rect 5457 10081 5491 10115
rect 6193 10081 6227 10115
rect 6929 10081 6963 10115
rect 7021 10081 7055 10115
rect 10149 10081 10183 10115
rect 10977 10081 11011 10115
rect 11161 10081 11195 10115
rect 11897 10081 11931 10115
rect 12725 10081 12759 10115
rect 13001 10081 13035 10115
rect 17509 10081 17543 10115
rect 17601 10081 17635 10115
rect 1501 10013 1535 10047
rect 1869 10013 1903 10047
rect 2329 10013 2363 10047
rect 2421 10013 2455 10047
rect 3157 10013 3191 10047
rect 4077 10013 4111 10047
rect 6009 10013 6043 10047
rect 7389 10013 7423 10047
rect 7656 10013 7690 10047
rect 9965 10013 9999 10047
rect 10057 10013 10091 10047
rect 11713 10013 11747 10047
rect 12541 10013 12575 10047
rect 13277 10013 13311 10047
rect 15485 10013 15519 10047
rect 15577 10013 15611 10047
rect 15844 10013 15878 10047
rect 18429 10013 18463 10047
rect 1685 9945 1719 9979
rect 3893 9945 3927 9979
rect 4261 9945 4295 9979
rect 5181 9945 5215 9979
rect 10885 9945 10919 9979
rect 11805 9945 11839 9979
rect 15240 9945 15274 9979
rect 18245 9945 18279 9979
rect 2145 9877 2179 9911
rect 2605 9877 2639 9911
rect 3249 9877 3283 9911
rect 5641 9877 5675 9911
rect 6101 9877 6135 9911
rect 6837 9877 6871 9911
rect 8769 9877 8803 9911
rect 12633 9877 12667 9911
rect 14105 9877 14139 9911
rect 16957 9877 16991 9911
rect 17417 9877 17451 9911
rect 17877 9877 17911 9911
rect 5825 9673 5859 9707
rect 6377 9673 6411 9707
rect 6745 9673 6779 9707
rect 12541 9673 12575 9707
rect 12909 9673 12943 9707
rect 15577 9673 15611 9707
rect 16313 9673 16347 9707
rect 16681 9673 16715 9707
rect 4445 9605 4479 9639
rect 7205 9605 7239 9639
rect 8686 9605 8720 9639
rect 10333 9605 10367 9639
rect 1501 9537 1535 9571
rect 2044 9537 2078 9571
rect 3617 9537 3651 9571
rect 4537 9537 4571 9571
rect 5089 9537 5123 9571
rect 5273 9537 5307 9571
rect 6837 9537 6871 9571
rect 7481 9537 7515 9571
rect 14197 9537 14231 9571
rect 14464 9537 14498 9571
rect 15669 9537 15703 9571
rect 17049 9537 17083 9571
rect 17969 9537 18003 9571
rect 1777 9469 1811 9503
rect 3709 9469 3743 9503
rect 3893 9469 3927 9503
rect 4629 9469 4663 9503
rect 5641 9469 5675 9503
rect 5733 9469 5767 9503
rect 7021 9469 7055 9503
rect 8953 9469 8987 9503
rect 11529 9469 11563 9503
rect 12265 9469 12299 9503
rect 12449 9469 12483 9503
rect 13001 9469 13035 9503
rect 13277 9469 13311 9503
rect 17141 9469 17175 9503
rect 17233 9469 17267 9503
rect 17693 9469 17727 9503
rect 3249 9401 3283 9435
rect 4077 9401 4111 9435
rect 6193 9401 6227 9435
rect 1593 9333 1627 9367
rect 3157 9333 3191 9367
rect 4905 9333 4939 9367
rect 7573 9333 7607 9367
rect 13921 9333 13955 9367
rect 16405 9333 16439 9367
rect 17601 9333 17635 9367
rect 1501 9129 1535 9163
rect 9045 9129 9079 9163
rect 12909 9129 12943 9163
rect 14289 9129 14323 9163
rect 15945 9129 15979 9163
rect 17233 9129 17267 9163
rect 17325 9129 17359 9163
rect 3249 9061 3283 9095
rect 2973 8993 3007 9027
rect 8585 8993 8619 9027
rect 9873 8993 9907 9027
rect 10609 8993 10643 9027
rect 13461 8993 13495 9027
rect 13829 8993 13863 9027
rect 16589 8993 16623 9027
rect 17877 8993 17911 9027
rect 3065 8925 3099 8959
rect 3525 8925 3559 8959
rect 5181 8925 5215 8959
rect 5273 8925 5307 8959
rect 8401 8925 8435 8959
rect 12817 8925 12851 8959
rect 14565 8925 14599 8959
rect 16405 8925 16439 8959
rect 17693 8925 17727 8959
rect 17785 8925 17819 8959
rect 18245 8925 18279 8959
rect 2706 8857 2740 8891
rect 3433 8857 3467 8891
rect 4914 8857 4948 8891
rect 7021 8857 7055 8891
rect 8493 8857 8527 8891
rect 9689 8857 9723 8891
rect 12572 8857 12606 8891
rect 13277 8857 13311 8891
rect 14832 8857 14866 8891
rect 16773 8857 16807 8891
rect 1593 8789 1627 8823
rect 3801 8789 3835 8823
rect 8033 8789 8067 8823
rect 9229 8789 9263 8823
rect 9597 8789 9631 8823
rect 10057 8789 10091 8823
rect 10425 8789 10459 8823
rect 10517 8789 10551 8823
rect 11437 8789 11471 8823
rect 13369 8789 13403 8823
rect 14105 8789 14139 8823
rect 16037 8789 16071 8823
rect 16221 8789 16255 8823
rect 16865 8789 16899 8823
rect 18429 8789 18463 8823
rect 1777 8585 1811 8619
rect 2237 8585 2271 8619
rect 2605 8585 2639 8619
rect 3433 8585 3467 8619
rect 5365 8585 5399 8619
rect 5825 8585 5859 8619
rect 6745 8585 6779 8619
rect 7481 8585 7515 8619
rect 7941 8585 7975 8619
rect 13001 8585 13035 8619
rect 13369 8585 13403 8619
rect 14289 8585 14323 8619
rect 14749 8585 14783 8619
rect 16497 8585 16531 8619
rect 17417 8585 17451 8619
rect 17509 8585 17543 8619
rect 17969 8585 18003 8619
rect 6193 8517 6227 8551
rect 6653 8517 6687 8551
rect 7205 8517 7239 8551
rect 8309 8517 8343 8551
rect 8769 8517 8803 8551
rect 12081 8517 12115 8551
rect 13737 8517 13771 8551
rect 13829 8517 13863 8551
rect 4353 8449 4387 8483
rect 5273 8449 5307 8483
rect 6009 8449 6043 8483
rect 10701 8449 10735 8483
rect 11989 8449 12023 8483
rect 12909 8449 12943 8483
rect 14540 8449 14574 8483
rect 15862 8449 15896 8483
rect 16129 8449 16163 8483
rect 16313 8449 16347 8483
rect 17049 8449 17083 8483
rect 17877 8449 17911 8483
rect 18521 8449 18555 8483
rect 1593 8381 1627 8415
rect 1685 8381 1719 8415
rect 2697 8381 2731 8415
rect 2881 8381 2915 8415
rect 3157 8381 3191 8415
rect 3709 8381 3743 8415
rect 4445 8381 4479 8415
rect 4537 8381 4571 8415
rect 5457 8381 5491 8415
rect 6469 8381 6503 8415
rect 8401 8381 8435 8415
rect 8493 8381 8527 8415
rect 11897 8381 11931 8415
rect 13185 8381 13219 8415
rect 14013 8381 14047 8415
rect 16773 8381 16807 8415
rect 16957 8381 16991 8415
rect 18061 8381 18095 8415
rect 3985 8313 4019 8347
rect 10057 8313 10091 8347
rect 11529 8313 11563 8347
rect 12541 8313 12575 8347
rect 14611 8313 14645 8347
rect 18337 8313 18371 8347
rect 2145 8245 2179 8279
rect 3893 8245 3927 8279
rect 4905 8245 4939 8279
rect 7113 8245 7147 8279
rect 7849 8245 7883 8279
rect 11345 8245 11379 8279
rect 12449 8245 12483 8279
rect 1501 8041 1535 8075
rect 2329 8041 2363 8075
rect 2697 8041 2731 8075
rect 4169 8041 4203 8075
rect 11713 8041 11747 8075
rect 15853 8041 15887 8075
rect 16773 8041 16807 8075
rect 17601 8041 17635 8075
rect 8033 7973 8067 8007
rect 9045 7973 9079 8007
rect 10241 7973 10275 8007
rect 14105 7973 14139 8007
rect 15117 7973 15151 8007
rect 16129 7973 16163 8007
rect 3341 7905 3375 7939
rect 4629 7905 4663 7939
rect 7297 7905 7331 7939
rect 7481 7905 7515 7939
rect 8677 7905 8711 7939
rect 9597 7905 9631 7939
rect 9965 7905 9999 7939
rect 10149 7905 10183 7939
rect 14657 7905 14691 7939
rect 17325 7905 17359 7939
rect 18153 7905 18187 7939
rect 1685 7837 1719 7871
rect 2605 7837 2639 7871
rect 3065 7837 3099 7871
rect 3157 7837 3191 7871
rect 3525 7837 3559 7871
rect 4353 7837 4387 7871
rect 4813 7837 4847 7871
rect 7021 7837 7055 7871
rect 7573 7837 7607 7871
rect 9413 7837 9447 7871
rect 10425 7837 10459 7871
rect 12265 7837 12299 7871
rect 13737 7837 13771 7871
rect 14933 7837 14967 7871
rect 15209 7837 15243 7871
rect 15945 7837 15979 7871
rect 16405 7837 16439 7871
rect 16681 7837 16715 7871
rect 17969 7837 18003 7871
rect 4721 7769 4755 7803
rect 8493 7769 8527 7803
rect 9505 7769 9539 7803
rect 12510 7769 12544 7803
rect 2421 7701 2455 7735
rect 3985 7701 4019 7735
rect 5181 7701 5215 7735
rect 5733 7701 5767 7735
rect 7941 7701 7975 7735
rect 8401 7701 8435 7735
rect 13645 7701 13679 7735
rect 13921 7701 13955 7735
rect 14473 7701 14507 7735
rect 14565 7701 14599 7735
rect 16221 7701 16255 7735
rect 16497 7701 16531 7735
rect 17141 7701 17175 7735
rect 17233 7701 17267 7735
rect 18061 7701 18095 7735
rect 18429 7701 18463 7735
rect 1593 7497 1627 7531
rect 1869 7497 1903 7531
rect 2697 7497 2731 7531
rect 3065 7497 3099 7531
rect 4077 7497 4111 7531
rect 4629 7497 4663 7531
rect 5089 7497 5123 7531
rect 5457 7497 5491 7531
rect 5917 7497 5951 7531
rect 9505 7497 9539 7531
rect 9597 7497 9631 7531
rect 11069 7497 11103 7531
rect 11621 7497 11655 7531
rect 12357 7497 12391 7531
rect 12817 7497 12851 7531
rect 16405 7497 16439 7531
rect 17693 7497 17727 7531
rect 17969 7497 18003 7531
rect 18429 7497 18463 7531
rect 4997 7429 5031 7463
rect 7849 7429 7883 7463
rect 8392 7429 8426 7463
rect 10710 7429 10744 7463
rect 13277 7429 13311 7463
rect 14096 7429 14130 7463
rect 17325 7429 17359 7463
rect 1409 7361 1443 7395
rect 2053 7361 2087 7395
rect 2421 7361 2455 7395
rect 2605 7361 2639 7395
rect 3157 7361 3191 7395
rect 3709 7361 3743 7395
rect 4169 7361 4203 7395
rect 5825 7361 5859 7395
rect 7490 7361 7524 7395
rect 7757 7361 7791 7395
rect 8125 7361 8159 7395
rect 12265 7361 12299 7395
rect 13185 7361 13219 7395
rect 13829 7361 13863 7395
rect 15301 7361 15335 7395
rect 15577 7361 15611 7395
rect 15853 7361 15887 7395
rect 16129 7361 16163 7395
rect 16681 7361 16715 7395
rect 17417 7361 17451 7395
rect 18153 7361 18187 7395
rect 18245 7361 18279 7395
rect 3341 7293 3375 7327
rect 3985 7293 4019 7327
rect 5181 7293 5215 7327
rect 6101 7293 6135 7327
rect 10977 7293 11011 7327
rect 12081 7293 12115 7327
rect 13461 7293 13495 7327
rect 2237 7225 2271 7259
rect 3525 7225 3559 7259
rect 4537 7225 4571 7259
rect 11345 7225 11379 7259
rect 16313 7225 16347 7259
rect 17601 7225 17635 7259
rect 6377 7157 6411 7191
rect 11805 7157 11839 7191
rect 12725 7157 12759 7191
rect 13737 7157 13771 7191
rect 15209 7157 15243 7191
rect 15485 7157 15519 7191
rect 15761 7157 15795 7191
rect 16037 7157 16071 7191
rect 1501 6953 1535 6987
rect 2605 6953 2639 6987
rect 5181 6953 5215 6987
rect 7665 6953 7699 6987
rect 8585 6953 8619 6987
rect 10425 6953 10459 6987
rect 11989 6953 12023 6987
rect 18429 6953 18463 6987
rect 2329 6885 2363 6919
rect 8953 6885 8987 6919
rect 3341 6817 3375 6851
rect 6837 6817 6871 6851
rect 7113 6817 7147 6851
rect 7941 6817 7975 6851
rect 9505 6817 9539 6851
rect 12173 6817 12207 6851
rect 13553 6817 13587 6851
rect 16865 6817 16899 6851
rect 17693 6817 17727 6851
rect 1685 6749 1719 6783
rect 2053 6749 2087 6783
rect 2145 6749 2179 6783
rect 2697 6749 2731 6783
rect 3617 6749 3651 6783
rect 3801 6749 3835 6783
rect 5273 6749 5307 6783
rect 7757 6749 7791 6783
rect 9781 6749 9815 6783
rect 10609 6749 10643 6783
rect 14105 6749 14139 6783
rect 14841 6749 14875 6783
rect 18245 6749 18279 6783
rect 4046 6681 4080 6715
rect 8217 6681 8251 6715
rect 9413 6681 9447 6715
rect 10876 6681 10910 6715
rect 12357 6681 12391 6715
rect 13277 6681 13311 6715
rect 13369 6681 13403 6715
rect 15108 6681 15142 6715
rect 17509 6681 17543 6715
rect 1869 6613 1903 6647
rect 3433 6613 3467 6647
rect 7297 6613 7331 6647
rect 8125 6613 8159 6647
rect 8769 6613 8803 6647
rect 9321 6613 9355 6647
rect 12449 6613 12483 6647
rect 12817 6613 12851 6647
rect 12909 6613 12943 6647
rect 13737 6613 13771 6647
rect 14749 6613 14783 6647
rect 16221 6613 16255 6647
rect 16313 6613 16347 6647
rect 16681 6613 16715 6647
rect 16773 6613 16807 6647
rect 17141 6613 17175 6647
rect 17601 6613 17635 6647
rect 17969 6613 18003 6647
rect 2053 6409 2087 6443
rect 2513 6409 2547 6443
rect 4353 6409 4387 6443
rect 6745 6409 6779 6443
rect 7665 6409 7699 6443
rect 8033 6409 8067 6443
rect 8401 6409 8435 6443
rect 12909 6409 12943 6443
rect 14565 6409 14599 6443
rect 15209 6409 15243 6443
rect 15577 6409 15611 6443
rect 16681 6409 16715 6443
rect 17049 6409 17083 6443
rect 18337 6409 18371 6443
rect 6837 6341 6871 6375
rect 10342 6341 10376 6375
rect 15117 6341 15151 6375
rect 1685 6273 1719 6307
rect 1869 6273 1903 6307
rect 2329 6273 2363 6307
rect 3729 6273 3763 6307
rect 3985 6273 4019 6307
rect 4261 6273 4295 6307
rect 4537 6273 4571 6307
rect 5834 6273 5868 6307
rect 9137 6273 9171 6307
rect 10701 6273 10735 6307
rect 11796 6273 11830 6307
rect 13093 6273 13127 6307
rect 13360 6273 13394 6307
rect 15945 6273 15979 6307
rect 17877 6273 17911 6307
rect 18521 6273 18555 6307
rect 6101 6205 6135 6239
rect 6929 6205 6963 6239
rect 7481 6205 7515 6239
rect 7573 6205 7607 6239
rect 10609 6205 10643 6239
rect 11529 6205 11563 6239
rect 15301 6205 15335 6239
rect 16037 6205 16071 6239
rect 16129 6205 16163 6239
rect 16497 6205 16531 6239
rect 17141 6205 17175 6239
rect 17233 6205 17267 6239
rect 17969 6205 18003 6239
rect 18061 6205 18095 6239
rect 9229 6137 9263 6171
rect 14749 6137 14783 6171
rect 1501 6069 1535 6103
rect 2145 6069 2179 6103
rect 2605 6069 2639 6103
rect 4077 6069 4111 6103
rect 4721 6069 4755 6103
rect 6377 6069 6411 6103
rect 8493 6069 8527 6103
rect 11345 6069 11379 6103
rect 14473 6069 14507 6103
rect 17509 6069 17543 6103
rect 13093 5865 13127 5899
rect 15669 5865 15703 5899
rect 16221 5865 16255 5899
rect 17049 5865 17083 5899
rect 18061 5865 18095 5899
rect 18429 5865 18463 5899
rect 4353 5797 4387 5831
rect 2237 5729 2271 5763
rect 3433 5729 3467 5763
rect 3985 5729 4019 5763
rect 5089 5729 5123 5763
rect 7665 5729 7699 5763
rect 8769 5729 8803 5763
rect 10333 5729 10367 5763
rect 12725 5729 12759 5763
rect 12909 5729 12943 5763
rect 13645 5729 13679 5763
rect 16773 5729 16807 5763
rect 17601 5729 17635 5763
rect 1685 5661 1719 5695
rect 1777 5661 1811 5695
rect 2329 5661 2363 5695
rect 7021 5661 7055 5695
rect 7941 5661 7975 5695
rect 10077 5661 10111 5695
rect 10425 5661 10459 5695
rect 12173 5661 12207 5695
rect 14289 5661 14323 5695
rect 14556 5661 14590 5695
rect 16129 5661 16163 5695
rect 17417 5661 17451 5695
rect 17877 5661 17911 5695
rect 18245 5661 18279 5695
rect 3341 5593 3375 5627
rect 4169 5593 4203 5627
rect 8585 5593 8619 5627
rect 12633 5593 12667 5627
rect 13461 5593 13495 5627
rect 13553 5593 13587 5627
rect 1501 5525 1535 5559
rect 1961 5525 1995 5559
rect 2421 5525 2455 5559
rect 2789 5525 2823 5559
rect 2881 5525 2915 5559
rect 3249 5525 3283 5559
rect 4445 5525 4479 5559
rect 4813 5525 4847 5559
rect 4905 5525 4939 5559
rect 5733 5525 5767 5559
rect 7113 5525 7147 5559
rect 7481 5525 7515 5559
rect 7573 5525 7607 5559
rect 8953 5525 8987 5559
rect 12265 5525 12299 5559
rect 14105 5525 14139 5559
rect 15945 5525 15979 5559
rect 16589 5525 16623 5559
rect 16681 5525 16715 5559
rect 17509 5525 17543 5559
rect 2145 5321 2179 5355
rect 2421 5321 2455 5355
rect 5457 5321 5491 5355
rect 5825 5321 5859 5355
rect 8033 5321 8067 5355
rect 13093 5321 13127 5355
rect 16773 5321 16807 5355
rect 17141 5321 17175 5355
rect 17601 5321 17635 5355
rect 17969 5321 18003 5355
rect 4353 5253 4387 5287
rect 5089 5253 5123 5287
rect 12955 5253 12989 5287
rect 13461 5253 13495 5287
rect 15117 5253 15151 5287
rect 1685 5185 1719 5219
rect 2053 5185 2087 5219
rect 2329 5185 2363 5219
rect 4537 5185 4571 5219
rect 4997 5185 5031 5219
rect 6469 5185 6503 5219
rect 6736 5185 6770 5219
rect 8309 5185 8343 5219
rect 8576 5185 8610 5219
rect 10241 5185 10275 5219
rect 10333 5185 10367 5219
rect 11161 5185 11195 5219
rect 11529 5185 11563 5219
rect 11805 5185 11839 5219
rect 12265 5185 12299 5219
rect 12852 5185 12886 5219
rect 15209 5185 15243 5219
rect 15634 5185 15668 5219
rect 15945 5185 15979 5219
rect 16037 5185 16071 5219
rect 16313 5185 16347 5219
rect 17233 5185 17267 5219
rect 18521 5185 18555 5219
rect 2605 5117 2639 5151
rect 5273 5117 5307 5151
rect 5917 5117 5951 5151
rect 6009 5117 6043 5151
rect 12081 5117 12115 5151
rect 13277 5117 13311 5151
rect 17325 5117 17359 5151
rect 18061 5117 18095 5151
rect 18153 5117 18187 5151
rect 1501 5049 1535 5083
rect 8125 5049 8159 5083
rect 9689 5049 9723 5083
rect 11713 5049 11747 5083
rect 15761 5049 15795 5083
rect 16221 5049 16255 5083
rect 1869 4981 1903 5015
rect 4629 4981 4663 5015
rect 7849 4981 7883 5015
rect 9781 4981 9815 5015
rect 10149 4981 10183 5015
rect 10977 4981 11011 5015
rect 11345 4981 11379 5015
rect 11989 4981 12023 5015
rect 12725 4981 12759 5015
rect 15393 4981 15427 5015
rect 15531 4981 15565 5015
rect 16497 4981 16531 5015
rect 1777 4777 1811 4811
rect 2053 4777 2087 4811
rect 3617 4777 3651 4811
rect 4077 4777 4111 4811
rect 4445 4777 4479 4811
rect 4537 4777 4571 4811
rect 8953 4777 8987 4811
rect 9689 4777 9723 4811
rect 11529 4777 11563 4811
rect 13553 4777 13587 4811
rect 18429 4777 18463 4811
rect 6929 4709 6963 4743
rect 13829 4709 13863 4743
rect 4997 4641 5031 4675
rect 5181 4641 5215 4675
rect 12357 4641 12391 4675
rect 14197 4641 14231 4675
rect 16129 4641 16163 4675
rect 16313 4641 16347 4675
rect 16865 4641 16899 4675
rect 18061 4641 18095 4675
rect 1685 4573 1719 4607
rect 1961 4573 1995 4607
rect 2237 4573 2271 4607
rect 2513 4573 2547 4607
rect 2881 4573 2915 4607
rect 3157 4573 3191 4607
rect 3409 4573 3443 4607
rect 4905 4573 4939 4607
rect 5365 4573 5399 4607
rect 7205 4573 7239 4607
rect 7389 4573 7423 4607
rect 9597 4573 9631 4607
rect 9873 4573 9907 4607
rect 10149 4573 10183 4607
rect 11621 4573 11655 4607
rect 12541 4573 12575 4607
rect 13093 4573 13127 4607
rect 13369 4573 13403 4607
rect 13645 4573 13679 4607
rect 16037 4573 16071 4607
rect 18245 4573 18279 4607
rect 3893 4505 3927 4539
rect 5610 4505 5644 4539
rect 7656 4505 7690 4539
rect 10416 4505 10450 4539
rect 14381 4505 14415 4539
rect 1501 4437 1535 4471
rect 2329 4437 2363 4471
rect 2697 4437 2731 4471
rect 2973 4437 3007 4471
rect 3249 4437 3283 4471
rect 4169 4437 4203 4471
rect 6745 4437 6779 4471
rect 7021 4437 7055 4471
rect 8769 4437 8803 4471
rect 10057 4437 10091 4471
rect 12265 4437 12299 4471
rect 13001 4437 13035 4471
rect 13277 4437 13311 4471
rect 3525 4233 3559 4267
rect 4261 4233 4295 4267
rect 4997 4233 5031 4267
rect 5457 4233 5491 4267
rect 9413 4233 9447 4267
rect 12449 4233 12483 4267
rect 17325 4233 17359 4267
rect 15393 4165 15427 4199
rect 1685 4097 1719 4131
rect 2053 4097 2087 4131
rect 2329 4097 2363 4131
rect 2605 4097 2639 4131
rect 2881 4097 2915 4131
rect 3157 4097 3191 4131
rect 3433 4097 3467 4131
rect 3709 4097 3743 4131
rect 4169 4097 4203 4131
rect 5089 4097 5123 4131
rect 5733 4097 5767 4131
rect 6469 4097 6503 4131
rect 6736 4097 6770 4131
rect 7941 4097 7975 4131
rect 8585 4097 8619 4131
rect 8677 4097 8711 4131
rect 8953 4097 8987 4131
rect 9597 4097 9631 4131
rect 10241 4097 10275 4131
rect 10517 4097 10551 4131
rect 11161 4097 11195 4131
rect 11713 4097 11747 4131
rect 11989 4097 12023 4131
rect 12265 4097 12299 4131
rect 12541 4097 12575 4131
rect 14657 4097 14691 4131
rect 15531 4097 15565 4131
rect 15634 4097 15668 4131
rect 15853 4097 15887 4131
rect 16497 4097 16531 4131
rect 17509 4097 17543 4131
rect 17877 4097 17911 4131
rect 18245 4097 18279 4131
rect 4445 4029 4479 4063
rect 5273 4029 5307 4063
rect 10977 4029 11011 4063
rect 12817 4029 12851 4063
rect 13001 4029 13035 4063
rect 14749 4029 14783 4063
rect 14933 4029 14967 4063
rect 16681 4029 16715 4063
rect 16865 4029 16899 4063
rect 3249 3961 3283 3995
rect 3801 3961 3835 3995
rect 4629 3961 4663 3995
rect 6193 3961 6227 3995
rect 7849 3961 7883 3995
rect 8861 3961 8895 3995
rect 10425 3961 10459 3995
rect 11345 3961 11379 3995
rect 11897 3961 11931 3995
rect 18061 3961 18095 3995
rect 1501 3893 1535 3927
rect 1869 3893 1903 3927
rect 2145 3893 2179 3927
rect 2421 3893 2455 3927
rect 2697 3893 2731 3927
rect 2973 3893 3007 3927
rect 5917 3893 5951 3927
rect 9137 3893 9171 3927
rect 9873 3893 9907 3927
rect 10057 3893 10091 3927
rect 10793 3893 10827 3927
rect 11621 3893 11655 3927
rect 12173 3893 12207 3927
rect 12725 3893 12759 3927
rect 16037 3893 16071 3927
rect 16313 3893 16347 3927
rect 17693 3893 17727 3927
rect 18429 3893 18463 3927
rect 3341 3689 3375 3723
rect 3893 3689 3927 3723
rect 5365 3689 5399 3723
rect 6929 3689 6963 3723
rect 7941 3689 7975 3723
rect 9597 3689 9631 3723
rect 12679 3689 12713 3723
rect 18429 3689 18463 3723
rect 3065 3621 3099 3655
rect 6837 3621 6871 3655
rect 8125 3621 8159 3655
rect 9965 3621 9999 3655
rect 14473 3621 14507 3655
rect 8953 3553 8987 3587
rect 14289 3553 14323 3587
rect 15301 3553 15335 3587
rect 15485 3553 15519 3587
rect 1685 3485 1719 3519
rect 2053 3485 2087 3519
rect 2605 3485 2639 3519
rect 2973 3485 3007 3519
rect 3249 3485 3283 3519
rect 3525 3485 3559 3519
rect 3985 3485 4019 3519
rect 5457 3485 5491 3519
rect 7573 3485 7607 3519
rect 7665 3485 7699 3519
rect 8217 3485 8251 3519
rect 8620 3485 8654 3519
rect 9137 3485 9171 3519
rect 9740 3485 9774 3519
rect 10149 3485 10183 3519
rect 10425 3485 10459 3519
rect 12173 3485 12207 3519
rect 12300 3485 12334 3519
rect 12576 3485 12610 3519
rect 12817 3485 12851 3519
rect 13093 3485 13127 3519
rect 13461 3485 13495 3519
rect 13737 3485 13771 3519
rect 14105 3485 14139 3519
rect 15209 3485 15243 3519
rect 17233 3485 17267 3519
rect 17509 3485 17543 3519
rect 17877 3485 17911 3519
rect 18245 3485 18279 3519
rect 2329 3417 2363 3451
rect 4252 3417 4286 3451
rect 5724 3417 5758 3451
rect 9827 3417 9861 3451
rect 11906 3417 11940 3451
rect 17141 3417 17175 3451
rect 1501 3349 1535 3383
rect 1869 3349 1903 3383
rect 2789 3349 2823 3383
rect 8401 3349 8435 3383
rect 8723 3349 8757 3383
rect 10241 3349 10275 3383
rect 10609 3349 10643 3383
rect 10793 3349 10827 3383
rect 12403 3349 12437 3383
rect 13001 3349 13035 3383
rect 13277 3349 13311 3383
rect 13645 3349 13679 3383
rect 13921 3349 13955 3383
rect 15025 3349 15059 3383
rect 17417 3349 17451 3383
rect 17693 3349 17727 3383
rect 18061 3349 18095 3383
rect 2237 3145 2271 3179
rect 3617 3145 3651 3179
rect 4629 3145 4663 3179
rect 5089 3145 5123 3179
rect 5273 3145 5307 3179
rect 6561 3145 6595 3179
rect 7389 3145 7423 3179
rect 15393 3145 15427 3179
rect 16497 3145 16531 3179
rect 13645 3077 13679 3111
rect 1685 3009 1719 3043
rect 2053 3009 2087 3043
rect 2421 3009 2455 3043
rect 2789 3009 2823 3043
rect 3157 3009 3191 3043
rect 3249 3009 3283 3043
rect 3801 3009 3835 3043
rect 4169 3009 4203 3043
rect 4445 3009 4479 3043
rect 6009 3009 6043 3043
rect 6377 3009 6411 3043
rect 6653 3009 6687 3043
rect 6929 3009 6963 3043
rect 7481 3009 7515 3043
rect 8217 3009 8251 3043
rect 8493 3009 8527 3043
rect 10701 3009 10735 3043
rect 11253 3009 11287 3043
rect 11529 3009 11563 3043
rect 13461 3009 13495 3043
rect 15577 3009 15611 3043
rect 15761 3009 15795 3043
rect 16313 3009 16347 3043
rect 16773 3009 16807 3043
rect 17141 3009 17175 3043
rect 17509 3009 17543 3043
rect 17877 3009 17911 3043
rect 18245 3009 18279 3043
rect 4905 2941 4939 2975
rect 5917 2941 5951 2975
rect 7941 2941 7975 2975
rect 9229 2941 9263 2975
rect 10425 2941 10459 2975
rect 10609 2941 10643 2975
rect 11713 2941 11747 2975
rect 12449 2941 12483 2975
rect 15117 2941 15151 2975
rect 1869 2873 1903 2907
rect 2605 2873 2639 2907
rect 6193 2873 6227 2907
rect 6837 2873 6871 2907
rect 8033 2873 8067 2907
rect 11161 2873 11195 2907
rect 15945 2873 15979 2907
rect 1501 2805 1535 2839
rect 2973 2805 3007 2839
rect 3433 2805 3467 2839
rect 3985 2805 4019 2839
rect 4261 2805 4295 2839
rect 4721 2805 4755 2839
rect 5641 2805 5675 2839
rect 7113 2805 7147 2839
rect 7573 2805 7607 2839
rect 8401 2805 8435 2839
rect 8677 2805 8711 2839
rect 10885 2805 10919 2839
rect 16957 2805 16991 2839
rect 17325 2805 17359 2839
rect 17693 2805 17727 2839
rect 18061 2805 18095 2839
rect 18429 2805 18463 2839
rect 2605 2601 2639 2635
rect 4721 2601 4755 2635
rect 5917 2601 5951 2635
rect 11805 2601 11839 2635
rect 12541 2601 12575 2635
rect 13277 2601 13311 2635
rect 16405 2601 16439 2635
rect 4997 2533 5031 2567
rect 11253 2533 11287 2567
rect 11529 2533 11563 2567
rect 16865 2533 16899 2567
rect 17601 2533 17635 2567
rect 9781 2465 9815 2499
rect 9965 2465 9999 2499
rect 12357 2465 12391 2499
rect 14105 2465 14139 2499
rect 15945 2465 15979 2499
rect 1685 2397 1719 2431
rect 2053 2397 2087 2431
rect 2513 2397 2547 2431
rect 2789 2397 2823 2431
rect 3525 2397 3559 2431
rect 4077 2397 4111 2431
rect 4537 2397 4571 2431
rect 4905 2397 4939 2431
rect 5181 2397 5215 2431
rect 5549 2397 5583 2431
rect 5733 2397 5767 2431
rect 6653 2397 6687 2431
rect 6745 2397 6779 2431
rect 7205 2397 7239 2431
rect 7757 2397 7791 2431
rect 8401 2397 8435 2431
rect 8493 2397 8527 2431
rect 9045 2397 9079 2431
rect 9689 2397 9723 2431
rect 10977 2397 11011 2431
rect 11069 2397 11103 2431
rect 11713 2397 11747 2431
rect 11989 2397 12023 2431
rect 12173 2397 12207 2431
rect 13036 2397 13070 2431
rect 13461 2397 13495 2431
rect 13645 2397 13679 2431
rect 16037 2397 16071 2431
rect 16681 2397 16715 2431
rect 17049 2397 17083 2431
rect 17417 2397 17451 2431
rect 17785 2397 17819 2431
rect 18245 2397 18279 2431
rect 10425 2329 10459 2363
rect 13139 2329 13173 2363
rect 14289 2329 14323 2363
rect 1501 2261 1535 2295
rect 1869 2261 1903 2295
rect 2329 2261 2363 2295
rect 2973 2261 3007 2295
rect 3341 2261 3375 2295
rect 3893 2261 3927 2295
rect 4353 2261 4387 2295
rect 5365 2261 5399 2295
rect 6101 2261 6135 2295
rect 6469 2261 6503 2295
rect 6929 2261 6963 2295
rect 7389 2261 7423 2295
rect 7573 2261 7607 2295
rect 7941 2261 7975 2295
rect 8217 2261 8251 2295
rect 8677 2261 8711 2295
rect 9229 2261 9263 2295
rect 9505 2261 9539 2295
rect 10517 2261 10551 2295
rect 10793 2261 10827 2295
rect 13829 2261 13863 2295
rect 16221 2261 16255 2295
rect 17233 2261 17267 2295
rect 17969 2261 18003 2295
rect 18429 2261 18463 2295
<< metal1 >>
rect 15930 16056 15936 16108
rect 15988 16096 15994 16108
rect 16390 16096 16396 16108
rect 15988 16068 16396 16096
rect 15988 16056 15994 16068
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 3786 15172 3792 15224
rect 3844 15212 3850 15224
rect 5534 15212 5540 15224
rect 3844 15184 5540 15212
rect 3844 15172 3850 15184
rect 5534 15172 5540 15184
rect 5592 15172 5598 15224
rect 4430 15036 4436 15088
rect 4488 15076 4494 15088
rect 4488 15048 12434 15076
rect 4488 15036 4494 15048
rect 3602 14968 3608 15020
rect 3660 15008 3666 15020
rect 7282 15008 7288 15020
rect 3660 14980 7288 15008
rect 3660 14968 3666 14980
rect 7282 14968 7288 14980
rect 7340 14968 7346 15020
rect 12406 15008 12434 15048
rect 14182 15008 14188 15020
rect 12406 14980 14188 15008
rect 14182 14968 14188 14980
rect 14240 14968 14246 15020
rect 3878 14900 3884 14952
rect 3936 14940 3942 14952
rect 5074 14940 5080 14952
rect 3936 14912 5080 14940
rect 3936 14900 3942 14912
rect 5074 14900 5080 14912
rect 5132 14900 5138 14952
rect 5166 14900 5172 14952
rect 5224 14940 5230 14952
rect 15194 14940 15200 14952
rect 5224 14912 15200 14940
rect 5224 14900 5230 14912
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 3694 14832 3700 14884
rect 3752 14872 3758 14884
rect 6638 14872 6644 14884
rect 3752 14844 6644 14872
rect 3752 14832 3758 14844
rect 6638 14832 6644 14844
rect 6696 14832 6702 14884
rect 9122 14832 9128 14884
rect 9180 14872 9186 14884
rect 17034 14872 17040 14884
rect 9180 14844 17040 14872
rect 9180 14832 9186 14844
rect 17034 14832 17040 14844
rect 17092 14832 17098 14884
rect 1210 14764 1216 14816
rect 1268 14804 1274 14816
rect 4062 14804 4068 14816
rect 1268 14776 4068 14804
rect 1268 14764 1274 14776
rect 4062 14764 4068 14776
rect 4120 14764 4126 14816
rect 4154 14764 4160 14816
rect 4212 14804 4218 14816
rect 7466 14804 7472 14816
rect 4212 14776 7472 14804
rect 4212 14764 4218 14776
rect 7466 14764 7472 14776
rect 7524 14764 7530 14816
rect 8110 14764 8116 14816
rect 8168 14804 8174 14816
rect 17954 14804 17960 14816
rect 8168 14776 17960 14804
rect 8168 14764 8174 14776
rect 17954 14764 17960 14776
rect 18012 14764 18018 14816
rect 1104 14714 18860 14736
rect 1104 14662 3174 14714
rect 3226 14662 3238 14714
rect 3290 14662 3302 14714
rect 3354 14662 3366 14714
rect 3418 14662 3430 14714
rect 3482 14662 7622 14714
rect 7674 14662 7686 14714
rect 7738 14662 7750 14714
rect 7802 14662 7814 14714
rect 7866 14662 7878 14714
rect 7930 14662 12070 14714
rect 12122 14662 12134 14714
rect 12186 14662 12198 14714
rect 12250 14662 12262 14714
rect 12314 14662 12326 14714
rect 12378 14662 16518 14714
rect 16570 14662 16582 14714
rect 16634 14662 16646 14714
rect 16698 14662 16710 14714
rect 16762 14662 16774 14714
rect 16826 14662 18860 14714
rect 1104 14640 18860 14662
rect 3421 14603 3479 14609
rect 3421 14569 3433 14603
rect 3467 14600 3479 14603
rect 3510 14600 3516 14612
rect 3467 14572 3516 14600
rect 3467 14569 3479 14572
rect 3421 14563 3479 14569
rect 3510 14560 3516 14572
rect 3568 14560 3574 14612
rect 5442 14560 5448 14612
rect 5500 14600 5506 14612
rect 5721 14603 5779 14609
rect 5721 14600 5733 14603
rect 5500 14572 5733 14600
rect 5500 14560 5506 14572
rect 5721 14569 5733 14572
rect 5767 14569 5779 14603
rect 5721 14563 5779 14569
rect 5810 14560 5816 14612
rect 5868 14600 5874 14612
rect 5868 14572 6684 14600
rect 5868 14560 5874 14572
rect 4062 14492 4068 14544
rect 4120 14532 4126 14544
rect 6549 14535 6607 14541
rect 6549 14532 6561 14535
rect 4120 14504 6561 14532
rect 4120 14492 4126 14504
rect 6549 14501 6561 14504
rect 6595 14501 6607 14535
rect 6656 14532 6684 14572
rect 6914 14560 6920 14612
rect 6972 14600 6978 14612
rect 7009 14603 7067 14609
rect 7009 14600 7021 14603
rect 6972 14572 7021 14600
rect 6972 14560 6978 14572
rect 7009 14569 7021 14572
rect 7055 14569 7067 14603
rect 7374 14600 7380 14612
rect 7335 14572 7380 14600
rect 7009 14563 7067 14569
rect 7374 14560 7380 14572
rect 7432 14560 7438 14612
rect 7466 14560 7472 14612
rect 7524 14600 7530 14612
rect 8021 14603 8079 14609
rect 8021 14600 8033 14603
rect 7524 14572 8033 14600
rect 7524 14560 7530 14572
rect 8021 14569 8033 14572
rect 8067 14569 8079 14603
rect 8662 14600 8668 14612
rect 8623 14572 8668 14600
rect 8021 14563 8079 14569
rect 8662 14560 8668 14572
rect 8720 14560 8726 14612
rect 9306 14600 9312 14612
rect 9267 14572 9312 14600
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 9950 14600 9956 14612
rect 9911 14572 9956 14600
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 10594 14600 10600 14612
rect 10555 14572 10600 14600
rect 10594 14560 10600 14572
rect 10652 14560 10658 14612
rect 11882 14560 11888 14612
rect 11940 14600 11946 14612
rect 12253 14603 12311 14609
rect 12253 14600 12265 14603
rect 11940 14572 12265 14600
rect 11940 14560 11946 14572
rect 7837 14535 7895 14541
rect 7837 14532 7849 14535
rect 6656 14504 7849 14532
rect 6549 14495 6607 14501
rect 7837 14501 7849 14504
rect 7883 14501 7895 14535
rect 8202 14532 8208 14544
rect 8163 14504 8208 14532
rect 7837 14495 7895 14501
rect 8202 14492 8208 14504
rect 8260 14492 8266 14544
rect 11701 14535 11759 14541
rect 11701 14501 11713 14535
rect 11747 14532 11759 14535
rect 11974 14532 11980 14544
rect 11747 14504 11980 14532
rect 11747 14501 11759 14504
rect 11701 14495 11759 14501
rect 11974 14492 11980 14504
rect 12032 14492 12038 14544
rect 1949 14467 2007 14473
rect 1949 14433 1961 14467
rect 1995 14464 2007 14467
rect 2682 14464 2688 14476
rect 1995 14436 2688 14464
rect 1995 14433 2007 14436
rect 1949 14427 2007 14433
rect 2682 14424 2688 14436
rect 2740 14424 2746 14476
rect 2958 14424 2964 14476
rect 3016 14464 3022 14476
rect 3145 14467 3203 14473
rect 3145 14464 3157 14467
rect 3016 14436 3157 14464
rect 3016 14424 3022 14436
rect 3145 14433 3157 14436
rect 3191 14464 3203 14467
rect 3694 14464 3700 14476
rect 3191 14436 3700 14464
rect 3191 14433 3203 14436
rect 3145 14427 3203 14433
rect 3694 14424 3700 14436
rect 3752 14424 3758 14476
rect 4154 14424 4160 14476
rect 4212 14464 4218 14476
rect 4617 14467 4675 14473
rect 4617 14464 4629 14467
rect 4212 14436 4629 14464
rect 4212 14424 4218 14436
rect 4617 14433 4629 14436
rect 4663 14433 4675 14467
rect 4617 14427 4675 14433
rect 5261 14467 5319 14473
rect 5261 14433 5273 14467
rect 5307 14464 5319 14467
rect 5718 14464 5724 14476
rect 5307 14436 5724 14464
rect 5307 14433 5319 14436
rect 5261 14427 5319 14433
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 2222 14396 2228 14408
rect 2183 14368 2228 14396
rect 2222 14356 2228 14368
rect 2280 14356 2286 14408
rect 2869 14399 2927 14405
rect 2869 14365 2881 14399
rect 2915 14365 2927 14399
rect 2869 14359 2927 14365
rect 3605 14399 3663 14405
rect 3605 14365 3617 14399
rect 3651 14365 3663 14399
rect 3605 14359 3663 14365
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14396 4399 14399
rect 4522 14396 4528 14408
rect 4387 14368 4528 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 2884 14328 2912 14359
rect 3418 14328 3424 14340
rect 2884 14300 3424 14328
rect 3418 14288 3424 14300
rect 3476 14288 3482 14340
rect 3620 14260 3648 14359
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 5534 14396 5540 14408
rect 5495 14368 5540 14396
rect 5534 14356 5540 14368
rect 5592 14356 5598 14408
rect 5905 14399 5963 14405
rect 5905 14365 5917 14399
rect 5951 14365 5963 14399
rect 5905 14359 5963 14365
rect 5920 14328 5948 14359
rect 5994 14356 6000 14408
rect 6052 14396 6058 14408
rect 6052 14368 6097 14396
rect 6052 14356 6058 14368
rect 6178 14356 6184 14408
rect 6236 14396 6242 14408
rect 6365 14399 6423 14405
rect 6365 14396 6377 14399
rect 6236 14368 6377 14396
rect 6236 14356 6242 14368
rect 6365 14365 6377 14368
rect 6411 14365 6423 14399
rect 6365 14359 6423 14365
rect 6546 14356 6552 14408
rect 6604 14396 6610 14408
rect 6825 14399 6883 14405
rect 6825 14396 6837 14399
rect 6604 14368 6837 14396
rect 6604 14356 6610 14368
rect 6825 14365 6837 14368
rect 6871 14365 6883 14399
rect 6825 14359 6883 14365
rect 7374 14356 7380 14408
rect 7432 14396 7438 14408
rect 7561 14399 7619 14405
rect 7561 14396 7573 14399
rect 7432 14368 7573 14396
rect 7432 14356 7438 14368
rect 7561 14365 7573 14368
rect 7607 14365 7619 14399
rect 7561 14359 7619 14365
rect 8662 14356 8668 14408
rect 8720 14396 8726 14408
rect 9125 14399 9183 14405
rect 9125 14396 9137 14399
rect 8720 14368 9137 14396
rect 8720 14356 8726 14368
rect 9125 14365 9137 14368
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 9306 14356 9312 14408
rect 9364 14396 9370 14408
rect 9401 14399 9459 14405
rect 9401 14396 9413 14399
rect 9364 14368 9413 14396
rect 9364 14356 9370 14368
rect 9401 14365 9413 14368
rect 9447 14365 9459 14399
rect 9401 14359 9459 14365
rect 9950 14356 9956 14408
rect 10008 14396 10014 14408
rect 10045 14399 10103 14405
rect 10045 14396 10057 14399
rect 10008 14368 10057 14396
rect 10008 14356 10014 14368
rect 10045 14365 10057 14368
rect 10091 14365 10103 14399
rect 10045 14359 10103 14365
rect 10594 14356 10600 14408
rect 10652 14396 10658 14408
rect 10689 14399 10747 14405
rect 10689 14396 10701 14399
rect 10652 14368 10701 14396
rect 10652 14356 10658 14368
rect 10689 14365 10701 14368
rect 10735 14365 10747 14399
rect 11514 14396 11520 14408
rect 11475 14368 11520 14396
rect 10689 14359 10747 14365
rect 11514 14356 11520 14368
rect 11572 14396 11578 14408
rect 12176 14405 12204 14572
rect 12253 14569 12265 14572
rect 12299 14569 12311 14603
rect 12526 14600 12532 14612
rect 12487 14572 12532 14600
rect 12253 14563 12311 14569
rect 12526 14560 12532 14572
rect 12584 14560 12590 14612
rect 13170 14600 13176 14612
rect 13131 14572 13176 14600
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 13262 14560 13268 14612
rect 13320 14600 13326 14612
rect 13320 14572 16528 14600
rect 13320 14560 13326 14572
rect 16500 14544 16528 14572
rect 12342 14492 12348 14544
rect 12400 14532 12406 14544
rect 15838 14532 15844 14544
rect 12400 14504 15844 14532
rect 12400 14492 12406 14504
rect 15838 14492 15844 14504
rect 15896 14492 15902 14544
rect 16482 14492 16488 14544
rect 16540 14492 16546 14544
rect 14645 14467 14703 14473
rect 14645 14433 14657 14467
rect 14691 14464 14703 14467
rect 16761 14467 16819 14473
rect 16761 14464 16773 14467
rect 14691 14436 16773 14464
rect 14691 14433 14703 14436
rect 14645 14427 14703 14433
rect 16761 14433 16773 14436
rect 16807 14464 16819 14467
rect 17402 14464 17408 14476
rect 16807 14436 17408 14464
rect 16807 14433 16819 14436
rect 16761 14427 16819 14433
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 17954 14464 17960 14476
rect 17915 14436 17960 14464
rect 17954 14424 17960 14436
rect 18012 14424 18018 14476
rect 11793 14399 11851 14405
rect 11793 14396 11805 14399
rect 11572 14368 11805 14396
rect 11572 14356 11578 14368
rect 11793 14365 11805 14368
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14365 12219 14399
rect 12161 14359 12219 14365
rect 12526 14356 12532 14408
rect 12584 14396 12590 14408
rect 12621 14399 12679 14405
rect 12621 14396 12633 14399
rect 12584 14368 12633 14396
rect 12584 14356 12590 14368
rect 12621 14365 12633 14368
rect 12667 14365 12679 14399
rect 12621 14359 12679 14365
rect 13170 14356 13176 14408
rect 13228 14396 13234 14408
rect 13265 14399 13323 14405
rect 13265 14396 13277 14399
rect 13228 14368 13277 14396
rect 13228 14356 13234 14368
rect 13265 14365 13277 14368
rect 13311 14365 13323 14399
rect 13265 14359 13323 14365
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13872 14368 14105 14396
rect 13872 14356 13878 14368
rect 14093 14365 14105 14368
rect 14139 14396 14151 14399
rect 14369 14399 14427 14405
rect 14369 14396 14381 14399
rect 14139 14368 14381 14396
rect 14139 14365 14151 14368
rect 14093 14359 14151 14365
rect 14369 14365 14381 14368
rect 14415 14365 14427 14399
rect 14369 14359 14427 14365
rect 14826 14356 14832 14408
rect 14884 14396 14890 14408
rect 15289 14399 15347 14405
rect 15289 14396 15301 14399
rect 14884 14368 15301 14396
rect 14884 14356 14890 14368
rect 15289 14365 15301 14368
rect 15335 14365 15347 14399
rect 15562 14396 15568 14408
rect 15475 14368 15568 14396
rect 15289 14359 15347 14365
rect 15562 14356 15568 14368
rect 15620 14396 15626 14408
rect 16022 14396 16028 14408
rect 15620 14368 16028 14396
rect 15620 14356 15626 14368
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16485 14399 16543 14405
rect 16485 14396 16497 14399
rect 16408 14368 16497 14396
rect 15654 14328 15660 14340
rect 5920 14300 15660 14328
rect 15654 14288 15660 14300
rect 15712 14288 15718 14340
rect 16114 14288 16120 14340
rect 16172 14328 16178 14340
rect 16408 14328 16436 14368
rect 16485 14365 16497 14368
rect 16531 14365 16543 14399
rect 16485 14359 16543 14365
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14365 17095 14399
rect 17678 14396 17684 14408
rect 17639 14368 17684 14396
rect 17037 14359 17095 14365
rect 17052 14328 17080 14359
rect 17678 14356 17684 14368
rect 17736 14356 17742 14408
rect 16172 14300 16436 14328
rect 16546 14300 17080 14328
rect 16172 14288 16178 14300
rect 16546 14272 16574 14300
rect 5718 14260 5724 14272
rect 3620 14232 5724 14260
rect 5718 14220 5724 14232
rect 5776 14220 5782 14272
rect 6181 14263 6239 14269
rect 6181 14229 6193 14263
rect 6227 14260 6239 14263
rect 6454 14260 6460 14272
rect 6227 14232 6460 14260
rect 6227 14229 6239 14232
rect 6181 14223 6239 14229
rect 6454 14220 6460 14232
rect 6512 14220 6518 14272
rect 7190 14220 7196 14272
rect 7248 14260 7254 14272
rect 7653 14263 7711 14269
rect 7653 14260 7665 14263
rect 7248 14232 7665 14260
rect 7248 14220 7254 14232
rect 7653 14229 7665 14232
rect 7699 14229 7711 14263
rect 7653 14223 7711 14229
rect 8846 14220 8852 14272
rect 8904 14260 8910 14272
rect 8941 14263 8999 14269
rect 8941 14260 8953 14263
rect 8904 14232 8953 14260
rect 8904 14220 8910 14232
rect 8941 14229 8953 14232
rect 8987 14229 8999 14263
rect 8941 14223 8999 14229
rect 9585 14263 9643 14269
rect 9585 14229 9597 14263
rect 9631 14260 9643 14263
rect 9766 14260 9772 14272
rect 9631 14232 9772 14260
rect 9631 14229 9643 14232
rect 9585 14223 9643 14229
rect 9766 14220 9772 14232
rect 9824 14220 9830 14272
rect 10229 14263 10287 14269
rect 10229 14229 10241 14263
rect 10275 14260 10287 14263
rect 10686 14260 10692 14272
rect 10275 14232 10692 14260
rect 10275 14229 10287 14232
rect 10229 14223 10287 14229
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 10870 14260 10876 14272
rect 10831 14232 10876 14260
rect 10870 14220 10876 14232
rect 10928 14220 10934 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 11977 14263 12035 14269
rect 11977 14260 11989 14263
rect 11940 14232 11989 14260
rect 11940 14220 11946 14232
rect 11977 14229 11989 14232
rect 12023 14229 12035 14263
rect 12802 14260 12808 14272
rect 12763 14232 12808 14260
rect 11977 14223 12035 14229
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 13446 14260 13452 14272
rect 13407 14232 13452 14260
rect 13446 14220 13452 14232
rect 13504 14220 13510 14272
rect 14277 14263 14335 14269
rect 14277 14229 14289 14263
rect 14323 14260 14335 14263
rect 15102 14260 15108 14272
rect 14323 14232 15108 14260
rect 14323 14229 14335 14232
rect 14277 14223 14335 14229
rect 15102 14220 15108 14232
rect 15160 14220 15166 14272
rect 15746 14220 15752 14272
rect 15804 14260 15810 14272
rect 16255 14263 16313 14269
rect 16255 14260 16267 14263
rect 15804 14232 16267 14260
rect 15804 14220 15810 14232
rect 16255 14229 16267 14232
rect 16301 14229 16313 14263
rect 16255 14223 16313 14229
rect 16482 14220 16488 14272
rect 16540 14232 16574 14272
rect 16540 14220 16546 14232
rect 1104 14170 18860 14192
rect 1104 14118 5398 14170
rect 5450 14118 5462 14170
rect 5514 14118 5526 14170
rect 5578 14118 5590 14170
rect 5642 14118 5654 14170
rect 5706 14118 9846 14170
rect 9898 14118 9910 14170
rect 9962 14118 9974 14170
rect 10026 14118 10038 14170
rect 10090 14118 10102 14170
rect 10154 14118 14294 14170
rect 14346 14118 14358 14170
rect 14410 14118 14422 14170
rect 14474 14118 14486 14170
rect 14538 14118 14550 14170
rect 14602 14118 18860 14170
rect 1104 14096 18860 14118
rect 2915 14059 2973 14065
rect 2915 14025 2927 14059
rect 2961 14056 2973 14059
rect 4154 14056 4160 14068
rect 2961 14028 4160 14056
rect 2961 14025 2973 14028
rect 2915 14019 2973 14025
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 4338 14056 4344 14068
rect 4299 14028 4344 14056
rect 4338 14016 4344 14028
rect 4396 14016 4402 14068
rect 4798 14016 4804 14068
rect 4856 14056 4862 14068
rect 4985 14059 5043 14065
rect 4985 14056 4997 14059
rect 4856 14028 4997 14056
rect 4856 14016 4862 14028
rect 4985 14025 4997 14028
rect 5031 14025 5043 14059
rect 4985 14019 5043 14025
rect 5353 14059 5411 14065
rect 5353 14025 5365 14059
rect 5399 14025 5411 14059
rect 5997 14059 6055 14065
rect 5997 14056 6009 14059
rect 5353 14019 5411 14025
rect 5644 14028 6009 14056
rect 4062 13988 4068 14000
rect 2746 13960 4068 13988
rect 2225 13923 2283 13929
rect 2225 13889 2237 13923
rect 2271 13920 2283 13923
rect 2746 13920 2774 13960
rect 4062 13948 4068 13960
rect 4120 13948 4126 14000
rect 5368 13988 5396 14019
rect 4172 13960 5396 13988
rect 3145 13923 3203 13929
rect 2271 13892 2820 13920
rect 2271 13889 2283 13892
rect 2225 13883 2283 13889
rect 2792 13864 2820 13892
rect 3145 13889 3157 13923
rect 3191 13920 3203 13923
rect 3602 13920 3608 13932
rect 3191 13892 3608 13920
rect 3191 13889 3203 13892
rect 3145 13883 3203 13889
rect 3602 13880 3608 13892
rect 3660 13880 3666 13932
rect 3970 13880 3976 13932
rect 4028 13920 4034 13932
rect 4172 13920 4200 13960
rect 4028 13892 4200 13920
rect 4028 13880 4034 13892
rect 4430 13880 4436 13932
rect 4488 13920 4494 13932
rect 4525 13923 4583 13929
rect 4525 13920 4537 13923
rect 4488 13892 4537 13920
rect 4488 13880 4494 13892
rect 4525 13889 4537 13892
rect 4571 13889 4583 13923
rect 4798 13920 4804 13932
rect 4759 13892 4804 13920
rect 4525 13883 4583 13889
rect 4798 13880 4804 13892
rect 4856 13880 4862 13932
rect 5166 13920 5172 13932
rect 5127 13892 5172 13920
rect 5166 13880 5172 13892
rect 5224 13880 5230 13932
rect 5534 13920 5540 13932
rect 5495 13892 5540 13920
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 5644 13920 5672 14028
rect 5997 14025 6009 14028
rect 6043 14025 6055 14059
rect 6546 14056 6552 14068
rect 6507 14028 6552 14056
rect 5997 14019 6055 14025
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 6638 14016 6644 14068
rect 6696 14056 6702 14068
rect 7469 14059 7527 14065
rect 7469 14056 7481 14059
rect 6696 14028 7481 14056
rect 6696 14016 6702 14028
rect 7469 14025 7481 14028
rect 7515 14025 7527 14059
rect 7469 14019 7527 14025
rect 9306 14016 9312 14068
rect 9364 14056 9370 14068
rect 13262 14056 13268 14068
rect 9364 14028 13268 14056
rect 9364 14016 9370 14028
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 13633 14059 13691 14065
rect 13633 14025 13645 14059
rect 13679 14025 13691 14059
rect 13633 14019 13691 14025
rect 5718 13948 5724 14000
rect 5776 13988 5782 14000
rect 13648 13988 13676 14019
rect 14182 14016 14188 14068
rect 14240 14056 14246 14068
rect 14461 14059 14519 14065
rect 14461 14056 14473 14059
rect 14240 14028 14473 14056
rect 14240 14016 14246 14028
rect 14461 14025 14473 14028
rect 14507 14025 14519 14059
rect 14461 14019 14519 14025
rect 15197 14059 15255 14065
rect 15197 14025 15209 14059
rect 15243 14056 15255 14059
rect 15562 14056 15568 14068
rect 15243 14028 15568 14056
rect 15243 14025 15255 14028
rect 15197 14019 15255 14025
rect 15562 14016 15568 14028
rect 15620 14016 15626 14068
rect 14826 13988 14832 14000
rect 5776 13960 13676 13988
rect 13740 13960 14832 13988
rect 5776 13948 5782 13960
rect 5905 13923 5963 13929
rect 5905 13920 5917 13923
rect 5644 13892 5917 13920
rect 5905 13889 5917 13892
rect 5951 13889 5963 13923
rect 6178 13920 6184 13932
rect 6139 13892 6184 13920
rect 5905 13883 5963 13889
rect 6178 13880 6184 13892
rect 6236 13880 6242 13932
rect 6270 13880 6276 13932
rect 6328 13920 6334 13932
rect 6365 13923 6423 13929
rect 6365 13920 6377 13923
rect 6328 13892 6377 13920
rect 6328 13880 6334 13892
rect 6365 13889 6377 13892
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 6454 13880 6460 13932
rect 6512 13920 6518 13932
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 6512 13892 6837 13920
rect 6512 13880 6518 13892
rect 6825 13889 6837 13892
rect 6871 13889 6883 13923
rect 6825 13883 6883 13889
rect 7006 13880 7012 13932
rect 7064 13920 7070 13932
rect 7374 13920 7380 13932
rect 7064 13892 7236 13920
rect 7335 13892 7380 13920
rect 7064 13880 7070 13892
rect 1949 13855 2007 13861
rect 1949 13821 1961 13855
rect 1995 13852 2007 13855
rect 2038 13852 2044 13864
rect 1995 13824 2044 13852
rect 1995 13821 2007 13824
rect 1949 13815 2007 13821
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2774 13812 2780 13864
rect 2832 13812 2838 13864
rect 3694 13812 3700 13864
rect 3752 13852 3758 13864
rect 3789 13855 3847 13861
rect 3789 13852 3801 13855
rect 3752 13824 3801 13852
rect 3752 13812 3758 13824
rect 3789 13821 3801 13824
rect 3835 13821 3847 13855
rect 3789 13815 3847 13821
rect 3878 13812 3884 13864
rect 3936 13852 3942 13864
rect 4065 13855 4123 13861
rect 4065 13852 4077 13855
rect 3936 13824 4077 13852
rect 3936 13812 3942 13824
rect 4065 13821 4077 13824
rect 4111 13821 4123 13855
rect 4065 13815 4123 13821
rect 4172 13824 5764 13852
rect 1578 13744 1584 13796
rect 1636 13784 1642 13796
rect 3970 13784 3976 13796
rect 1636 13756 3976 13784
rect 1636 13744 1642 13756
rect 3970 13744 3976 13756
rect 4028 13744 4034 13796
rect 4172 13784 4200 13824
rect 5736 13793 5764 13824
rect 5994 13812 6000 13864
rect 6052 13852 6058 13864
rect 7101 13855 7159 13861
rect 7101 13852 7113 13855
rect 6052 13824 7113 13852
rect 6052 13812 6058 13824
rect 7101 13821 7113 13824
rect 7147 13821 7159 13855
rect 7208 13852 7236 13892
rect 7374 13880 7380 13892
rect 7432 13880 7438 13932
rect 8202 13880 8208 13932
rect 8260 13920 8266 13932
rect 13740 13920 13768 13960
rect 14826 13948 14832 13960
rect 14884 13948 14890 14000
rect 15013 13991 15071 13997
rect 15013 13957 15025 13991
rect 15059 13988 15071 13991
rect 15059 13960 17724 13988
rect 15059 13957 15071 13960
rect 15013 13951 15071 13957
rect 8260 13892 13768 13920
rect 13817 13923 13875 13929
rect 8260 13880 8266 13892
rect 13817 13889 13829 13923
rect 13863 13889 13875 13923
rect 13817 13883 13875 13889
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13920 14703 13923
rect 14918 13920 14924 13932
rect 14691 13892 14924 13920
rect 14691 13889 14703 13892
rect 14645 13883 14703 13889
rect 9122 13852 9128 13864
rect 7208 13824 9128 13852
rect 7101 13815 7159 13821
rect 9122 13812 9128 13824
rect 9180 13812 9186 13864
rect 11606 13812 11612 13864
rect 11664 13852 11670 13864
rect 12342 13852 12348 13864
rect 11664 13824 12348 13852
rect 11664 13812 11670 13824
rect 12342 13812 12348 13824
rect 12400 13812 12406 13864
rect 13832 13852 13860 13883
rect 14918 13880 14924 13892
rect 14976 13920 14982 13932
rect 14976 13892 15148 13920
rect 14976 13880 14982 13892
rect 14734 13852 14740 13864
rect 13832 13824 14740 13852
rect 14734 13812 14740 13824
rect 14792 13852 14798 13864
rect 15010 13852 15016 13864
rect 14792 13824 15016 13852
rect 14792 13812 14798 13824
rect 15010 13812 15016 13824
rect 15068 13812 15074 13864
rect 4080 13756 4200 13784
rect 5721 13787 5779 13793
rect 290 13676 296 13728
rect 348 13716 354 13728
rect 4080 13716 4108 13756
rect 5721 13753 5733 13787
rect 5767 13753 5779 13787
rect 5721 13747 5779 13753
rect 6730 13744 6736 13796
rect 6788 13784 6794 13796
rect 8110 13784 8116 13796
rect 6788 13756 8116 13784
rect 6788 13744 6794 13756
rect 8110 13744 8116 13756
rect 8168 13744 8174 13796
rect 348 13688 4108 13716
rect 348 13676 354 13688
rect 4430 13676 4436 13728
rect 4488 13716 4494 13728
rect 4617 13719 4675 13725
rect 4617 13716 4629 13719
rect 4488 13688 4629 13716
rect 4488 13676 4494 13688
rect 4617 13685 4629 13688
rect 4663 13685 4675 13719
rect 4617 13679 4675 13685
rect 5074 13676 5080 13728
rect 5132 13716 5138 13728
rect 6546 13716 6552 13728
rect 5132 13688 6552 13716
rect 5132 13676 5138 13688
rect 6546 13676 6552 13688
rect 6604 13676 6610 13728
rect 6638 13676 6644 13728
rect 6696 13716 6702 13728
rect 15120 13716 15148 13892
rect 15378 13880 15384 13932
rect 15436 13920 15442 13932
rect 15473 13923 15531 13929
rect 15473 13920 15485 13923
rect 15436 13892 15485 13920
rect 15436 13880 15442 13892
rect 15473 13889 15485 13892
rect 15519 13889 15531 13923
rect 15473 13883 15531 13889
rect 15838 13880 15844 13932
rect 15896 13920 15902 13932
rect 16209 13923 16267 13929
rect 16209 13920 16221 13923
rect 15896 13892 16221 13920
rect 15896 13880 15902 13892
rect 16209 13889 16221 13892
rect 16255 13889 16267 13923
rect 16209 13883 16267 13889
rect 16298 13880 16304 13932
rect 16356 13920 16362 13932
rect 16485 13923 16543 13929
rect 16485 13920 16497 13923
rect 16356 13892 16497 13920
rect 16356 13880 16362 13892
rect 16485 13889 16497 13892
rect 16531 13920 16543 13923
rect 16850 13920 16856 13932
rect 16531 13892 16856 13920
rect 16531 13889 16543 13892
rect 16485 13883 16543 13889
rect 16850 13880 16856 13892
rect 16908 13880 16914 13932
rect 17696 13864 17724 13960
rect 15194 13812 15200 13864
rect 15252 13852 15258 13864
rect 16761 13855 16819 13861
rect 16761 13852 16773 13855
rect 15252 13824 15332 13852
rect 15252 13812 15258 13824
rect 15304 13793 15332 13824
rect 16546 13824 16773 13852
rect 15289 13787 15347 13793
rect 15289 13753 15301 13787
rect 15335 13753 15347 13787
rect 15289 13747 15347 13753
rect 16298 13744 16304 13796
rect 16356 13784 16362 13796
rect 16546 13784 16574 13824
rect 16761 13821 16773 13824
rect 16807 13821 16819 13855
rect 17034 13852 17040 13864
rect 16995 13824 17040 13852
rect 16761 13815 16819 13821
rect 17034 13812 17040 13824
rect 17092 13812 17098 13864
rect 17678 13852 17684 13864
rect 17639 13824 17684 13852
rect 17678 13812 17684 13824
rect 17736 13812 17742 13864
rect 17957 13855 18015 13861
rect 17957 13821 17969 13855
rect 18003 13852 18015 13855
rect 18046 13852 18052 13864
rect 18003 13824 18052 13852
rect 18003 13821 18015 13824
rect 17957 13815 18015 13821
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 16356 13756 16574 13784
rect 16356 13744 16362 13756
rect 16022 13716 16028 13728
rect 6696 13688 6741 13716
rect 15120 13688 16028 13716
rect 6696 13676 6702 13688
rect 16022 13676 16028 13688
rect 16080 13676 16086 13728
rect 1104 13626 18860 13648
rect 1104 13574 3174 13626
rect 3226 13574 3238 13626
rect 3290 13574 3302 13626
rect 3354 13574 3366 13626
rect 3418 13574 3430 13626
rect 3482 13574 7622 13626
rect 7674 13574 7686 13626
rect 7738 13574 7750 13626
rect 7802 13574 7814 13626
rect 7866 13574 7878 13626
rect 7930 13574 12070 13626
rect 12122 13574 12134 13626
rect 12186 13574 12198 13626
rect 12250 13574 12262 13626
rect 12314 13574 12326 13626
rect 12378 13574 16518 13626
rect 16570 13574 16582 13626
rect 16634 13574 16646 13626
rect 16698 13574 16710 13626
rect 16762 13574 16774 13626
rect 16826 13574 18860 13626
rect 1104 13552 18860 13574
rect 2866 13472 2872 13524
rect 2924 13512 2930 13524
rect 3329 13515 3387 13521
rect 3329 13512 3341 13515
rect 2924 13484 3341 13512
rect 2924 13472 2930 13484
rect 3329 13481 3341 13484
rect 3375 13481 3387 13515
rect 5445 13515 5503 13521
rect 5445 13512 5457 13515
rect 3329 13475 3387 13481
rect 3436 13484 5457 13512
rect 3436 13444 3464 13484
rect 5445 13481 5457 13484
rect 5491 13481 5503 13515
rect 5445 13475 5503 13481
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 5721 13515 5779 13521
rect 5721 13512 5733 13515
rect 5592 13484 5733 13512
rect 5592 13472 5598 13484
rect 5721 13481 5733 13484
rect 5767 13481 5779 13515
rect 6825 13515 6883 13521
rect 6825 13512 6837 13515
rect 5721 13475 5779 13481
rect 5828 13484 6837 13512
rect 5828 13444 5856 13484
rect 6825 13481 6837 13484
rect 6871 13481 6883 13515
rect 6825 13475 6883 13481
rect 15654 13472 15660 13524
rect 15712 13512 15718 13524
rect 15749 13515 15807 13521
rect 15749 13512 15761 13515
rect 15712 13484 15761 13512
rect 15712 13472 15718 13484
rect 15749 13481 15761 13484
rect 15795 13481 15807 13515
rect 15749 13475 15807 13481
rect 16114 13472 16120 13524
rect 16172 13512 16178 13524
rect 16393 13515 16451 13521
rect 16393 13512 16405 13515
rect 16172 13484 16405 13512
rect 16172 13472 16178 13484
rect 16393 13481 16405 13484
rect 16439 13481 16451 13515
rect 16393 13475 16451 13481
rect 16669 13515 16727 13521
rect 16669 13481 16681 13515
rect 16715 13512 16727 13515
rect 16850 13512 16856 13524
rect 16715 13484 16856 13512
rect 16715 13481 16727 13484
rect 16669 13475 16727 13481
rect 16850 13472 16856 13484
rect 16908 13472 16914 13524
rect 3344 13416 3464 13444
rect 3528 13416 5856 13444
rect 5997 13447 6055 13453
rect 2498 13336 2504 13388
rect 2556 13376 2562 13388
rect 2556 13348 2774 13376
rect 2556 13336 2562 13348
rect 1946 13308 1952 13320
rect 1907 13280 1952 13308
rect 1946 13268 1952 13280
rect 2004 13268 2010 13320
rect 2222 13308 2228 13320
rect 2183 13280 2228 13308
rect 2222 13268 2228 13280
rect 2280 13268 2286 13320
rect 2746 13240 2774 13348
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13308 2927 13311
rect 2958 13308 2964 13320
rect 2915 13280 2964 13308
rect 2915 13277 2927 13280
rect 2869 13271 2927 13277
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13308 3203 13311
rect 3234 13308 3240 13320
rect 3191 13280 3240 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 3344 13240 3372 13416
rect 3528 13376 3556 13416
rect 5997 13413 6009 13447
rect 6043 13413 6055 13447
rect 5997 13407 6055 13413
rect 2746 13212 3372 13240
rect 3436 13348 3556 13376
rect 2222 13132 2228 13184
rect 2280 13172 2286 13184
rect 3436 13172 3464 13348
rect 3602 13336 3608 13388
rect 3660 13376 3666 13388
rect 3881 13379 3939 13385
rect 3881 13376 3893 13379
rect 3660 13348 3893 13376
rect 3660 13336 3666 13348
rect 3881 13345 3893 13348
rect 3927 13345 3939 13379
rect 3881 13339 3939 13345
rect 4154 13336 4160 13388
rect 4212 13376 4218 13388
rect 6012 13376 6040 13407
rect 6546 13404 6552 13456
rect 6604 13444 6610 13456
rect 6641 13447 6699 13453
rect 6641 13444 6653 13447
rect 6604 13416 6653 13444
rect 6604 13404 6610 13416
rect 6641 13413 6653 13416
rect 6687 13413 6699 13447
rect 16298 13444 16304 13456
rect 16259 13416 16304 13444
rect 6641 13407 6699 13413
rect 16298 13404 16304 13416
rect 16356 13404 16362 13456
rect 4212 13348 4660 13376
rect 4212 13336 4218 13348
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13308 3571 13311
rect 4430 13308 4436 13320
rect 3559 13280 4436 13308
rect 3559 13277 3571 13280
rect 3513 13271 3571 13277
rect 4430 13268 4436 13280
rect 4488 13268 4494 13320
rect 4632 13317 4660 13348
rect 5644 13348 6040 13376
rect 5644 13317 5672 13348
rect 16390 13336 16396 13388
rect 16448 13376 16454 13388
rect 17589 13379 17647 13385
rect 17589 13376 17601 13379
rect 16448 13348 17601 13376
rect 16448 13336 16454 13348
rect 17589 13345 17601 13348
rect 17635 13345 17647 13379
rect 17589 13339 17647 13345
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13277 4675 13311
rect 4617 13271 4675 13277
rect 5629 13311 5687 13317
rect 5629 13277 5641 13311
rect 5675 13277 5687 13311
rect 5629 13271 5687 13277
rect 5905 13311 5963 13317
rect 5905 13277 5917 13311
rect 5951 13277 5963 13311
rect 5905 13271 5963 13277
rect 6181 13311 6239 13317
rect 6181 13277 6193 13311
rect 6227 13308 6239 13311
rect 15930 13308 15936 13320
rect 6227 13280 6408 13308
rect 15891 13280 15936 13308
rect 6227 13277 6239 13280
rect 6181 13271 6239 13277
rect 3786 13200 3792 13252
rect 3844 13240 3850 13252
rect 4157 13243 4215 13249
rect 4157 13240 4169 13243
rect 3844 13212 4169 13240
rect 3844 13200 3850 13212
rect 4157 13209 4169 13212
rect 4203 13209 4215 13243
rect 4157 13203 4215 13209
rect 4338 13200 4344 13252
rect 4396 13240 4402 13252
rect 5074 13240 5080 13252
rect 4396 13212 5080 13240
rect 4396 13200 4402 13212
rect 5074 13200 5080 13212
rect 5132 13200 5138 13252
rect 2280 13144 3464 13172
rect 2280 13132 2286 13144
rect 3510 13132 3516 13184
rect 3568 13172 3574 13184
rect 3878 13172 3884 13184
rect 3568 13144 3884 13172
rect 3568 13132 3574 13144
rect 3878 13132 3884 13144
rect 3936 13132 3942 13184
rect 4065 13175 4123 13181
rect 4065 13141 4077 13175
rect 4111 13172 4123 13175
rect 4246 13172 4252 13184
rect 4111 13144 4252 13172
rect 4111 13141 4123 13144
rect 4065 13135 4123 13141
rect 4246 13132 4252 13144
rect 4304 13132 4310 13184
rect 4525 13175 4583 13181
rect 4525 13141 4537 13175
rect 4571 13172 4583 13175
rect 5166 13172 5172 13184
rect 4571 13144 5172 13172
rect 4571 13141 4583 13144
rect 4525 13135 4583 13141
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 5258 13132 5264 13184
rect 5316 13172 5322 13184
rect 5920 13172 5948 13271
rect 6380 13252 6408 13280
rect 15930 13268 15936 13280
rect 15988 13268 15994 13320
rect 17218 13268 17224 13320
rect 17276 13308 17282 13320
rect 17313 13311 17371 13317
rect 17313 13308 17325 13311
rect 17276 13280 17325 13308
rect 17276 13268 17282 13280
rect 17313 13277 17325 13280
rect 17359 13277 17371 13311
rect 17678 13308 17684 13320
rect 17639 13280 17684 13308
rect 17313 13271 17371 13277
rect 17678 13268 17684 13280
rect 17736 13268 17742 13320
rect 17957 13311 18015 13317
rect 17957 13308 17969 13311
rect 17788 13280 17969 13308
rect 6362 13240 6368 13252
rect 6323 13212 6368 13240
rect 6362 13200 6368 13212
rect 6420 13200 6426 13252
rect 6549 13243 6607 13249
rect 6549 13209 6561 13243
rect 6595 13240 6607 13243
rect 15194 13240 15200 13252
rect 6595 13212 15200 13240
rect 6595 13209 6607 13212
rect 6549 13203 6607 13209
rect 6564 13172 6592 13203
rect 15194 13200 15200 13212
rect 15252 13200 15258 13252
rect 16117 13243 16175 13249
rect 16117 13209 16129 13243
rect 16163 13240 16175 13243
rect 17696 13240 17724 13268
rect 16163 13212 17724 13240
rect 16163 13209 16175 13212
rect 16117 13203 16175 13209
rect 5316 13144 5361 13172
rect 5920 13144 6592 13172
rect 5316 13132 5322 13144
rect 17402 13132 17408 13184
rect 17460 13172 17466 13184
rect 17788 13172 17816 13280
rect 17957 13277 17969 13280
rect 18003 13277 18015 13311
rect 17957 13271 18015 13277
rect 17460 13144 17816 13172
rect 17460 13132 17466 13144
rect 1104 13082 18860 13104
rect 1104 13030 5398 13082
rect 5450 13030 5462 13082
rect 5514 13030 5526 13082
rect 5578 13030 5590 13082
rect 5642 13030 5654 13082
rect 5706 13030 9846 13082
rect 9898 13030 9910 13082
rect 9962 13030 9974 13082
rect 10026 13030 10038 13082
rect 10090 13030 10102 13082
rect 10154 13030 14294 13082
rect 14346 13030 14358 13082
rect 14410 13030 14422 13082
rect 14474 13030 14486 13082
rect 14538 13030 14550 13082
rect 14602 13030 18860 13082
rect 1104 13008 18860 13030
rect 2746 12940 4016 12968
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12764 2007 12767
rect 2130 12764 2136 12776
rect 1995 12736 2136 12764
rect 1995 12733 2007 12736
rect 1949 12727 2007 12733
rect 2130 12724 2136 12736
rect 2188 12724 2194 12776
rect 2222 12724 2228 12776
rect 2280 12764 2286 12776
rect 2746 12764 2774 12940
rect 3418 12900 3424 12912
rect 3344 12872 3424 12900
rect 3142 12832 3148 12844
rect 3103 12804 3148 12832
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3344 12841 3372 12872
rect 3418 12860 3424 12872
rect 3476 12860 3482 12912
rect 3602 12909 3608 12912
rect 3596 12863 3608 12909
rect 3660 12900 3666 12912
rect 3988 12900 4016 12940
rect 4062 12928 4068 12980
rect 4120 12968 4126 12980
rect 4982 12968 4988 12980
rect 4120 12940 4988 12968
rect 4120 12928 4126 12940
rect 4982 12928 4988 12940
rect 5040 12928 5046 12980
rect 5166 12968 5172 12980
rect 5127 12940 5172 12968
rect 5166 12928 5172 12940
rect 5224 12928 5230 12980
rect 5902 12968 5908 12980
rect 5863 12940 5908 12968
rect 5902 12928 5908 12940
rect 5960 12928 5966 12980
rect 16390 12928 16396 12980
rect 16448 12968 16454 12980
rect 16945 12971 17003 12977
rect 16945 12968 16957 12971
rect 16448 12940 16957 12968
rect 16448 12928 16454 12940
rect 16945 12937 16957 12940
rect 16991 12937 17003 12971
rect 16945 12931 17003 12937
rect 5997 12903 6055 12909
rect 5997 12900 6009 12903
rect 3660 12872 3696 12900
rect 3988 12872 6009 12900
rect 3602 12860 3608 12863
rect 3660 12860 3666 12872
rect 5997 12869 6009 12872
rect 6043 12869 6055 12903
rect 5997 12863 6055 12869
rect 17221 12903 17279 12909
rect 17221 12869 17233 12903
rect 17267 12900 17279 12903
rect 17494 12900 17500 12912
rect 17267 12872 17500 12900
rect 17267 12869 17279 12872
rect 17221 12863 17279 12869
rect 17494 12860 17500 12872
rect 17552 12860 17558 12912
rect 3329 12835 3387 12841
rect 3329 12801 3341 12835
rect 3375 12801 3387 12835
rect 4890 12832 4896 12844
rect 3329 12795 3387 12801
rect 3436 12804 4896 12832
rect 2280 12736 2774 12764
rect 2869 12767 2927 12773
rect 2280 12724 2286 12736
rect 2869 12733 2881 12767
rect 2915 12764 2927 12767
rect 2958 12764 2964 12776
rect 2915 12736 2964 12764
rect 2915 12733 2927 12736
rect 2869 12727 2927 12733
rect 2958 12724 2964 12736
rect 3016 12724 3022 12776
rect 3160 12764 3188 12792
rect 3436 12764 3464 12804
rect 4890 12792 4896 12804
rect 4948 12792 4954 12844
rect 4982 12792 4988 12844
rect 5040 12832 5046 12844
rect 6365 12835 6423 12841
rect 6365 12832 6377 12835
rect 5040 12804 6377 12832
rect 5040 12792 5046 12804
rect 6365 12801 6377 12804
rect 6411 12801 6423 12835
rect 14550 12832 14556 12844
rect 6365 12795 6423 12801
rect 9646 12804 14556 12832
rect 3160 12736 3464 12764
rect 4522 12724 4528 12776
rect 4580 12764 4586 12776
rect 5261 12767 5319 12773
rect 5261 12764 5273 12767
rect 4580 12736 5273 12764
rect 4580 12724 4586 12736
rect 5261 12733 5273 12736
rect 5307 12733 5319 12767
rect 5261 12727 5319 12733
rect 5353 12767 5411 12773
rect 5353 12733 5365 12767
rect 5399 12733 5411 12767
rect 5718 12764 5724 12776
rect 5631 12736 5724 12764
rect 5353 12727 5411 12733
rect 4706 12696 4712 12708
rect 4619 12668 4712 12696
rect 4706 12656 4712 12668
rect 4764 12696 4770 12708
rect 5368 12696 5396 12727
rect 5718 12724 5724 12736
rect 5776 12764 5782 12776
rect 9646 12764 9674 12804
rect 14550 12792 14556 12804
rect 14608 12832 14614 12844
rect 19610 12832 19616 12844
rect 14608 12804 19616 12832
rect 14608 12792 14614 12804
rect 19610 12792 19616 12804
rect 19668 12792 19674 12844
rect 5776 12736 9674 12764
rect 16853 12767 16911 12773
rect 5776 12724 5782 12736
rect 16853 12733 16865 12767
rect 16899 12764 16911 12767
rect 17678 12764 17684 12776
rect 16899 12736 17684 12764
rect 16899 12733 16911 12736
rect 16853 12727 16911 12733
rect 17678 12724 17684 12736
rect 17736 12724 17742 12776
rect 17954 12764 17960 12776
rect 17915 12736 17960 12764
rect 17954 12724 17960 12736
rect 18012 12724 18018 12776
rect 4764 12668 5396 12696
rect 4764 12656 4770 12668
rect 10962 12656 10968 12708
rect 11020 12696 11026 12708
rect 17313 12699 17371 12705
rect 17313 12696 17325 12699
rect 11020 12668 17325 12696
rect 11020 12656 11026 12668
rect 17313 12665 17325 12668
rect 17359 12665 17371 12699
rect 17313 12659 17371 12665
rect 4798 12588 4804 12640
rect 4856 12628 4862 12640
rect 4856 12600 4901 12628
rect 4856 12588 4862 12600
rect 5074 12588 5080 12640
rect 5132 12628 5138 12640
rect 11054 12628 11060 12640
rect 5132 12600 11060 12628
rect 5132 12588 5138 12600
rect 11054 12588 11060 12600
rect 11112 12588 11118 12640
rect 15194 12588 15200 12640
rect 15252 12628 15258 12640
rect 18322 12628 18328 12640
rect 15252 12600 18328 12628
rect 15252 12588 15258 12600
rect 18322 12588 18328 12600
rect 18380 12588 18386 12640
rect 1104 12538 18860 12560
rect 1104 12486 3174 12538
rect 3226 12486 3238 12538
rect 3290 12486 3302 12538
rect 3354 12486 3366 12538
rect 3418 12486 3430 12538
rect 3482 12486 7622 12538
rect 7674 12486 7686 12538
rect 7738 12486 7750 12538
rect 7802 12486 7814 12538
rect 7866 12486 7878 12538
rect 7930 12486 12070 12538
rect 12122 12486 12134 12538
rect 12186 12486 12198 12538
rect 12250 12486 12262 12538
rect 12314 12486 12326 12538
rect 12378 12486 16518 12538
rect 16570 12486 16582 12538
rect 16634 12486 16646 12538
rect 16698 12486 16710 12538
rect 16762 12486 16774 12538
rect 16826 12486 18860 12538
rect 1104 12464 18860 12486
rect 2774 12424 2780 12436
rect 2332 12396 2780 12424
rect 2225 12291 2283 12297
rect 2225 12257 2237 12291
rect 2271 12288 2283 12291
rect 2332 12288 2360 12396
rect 2774 12384 2780 12396
rect 2832 12424 2838 12436
rect 4062 12424 4068 12436
rect 2832 12396 4068 12424
rect 2832 12384 2838 12396
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4522 12424 4528 12436
rect 4483 12396 4528 12424
rect 4522 12384 4528 12396
rect 4580 12384 4586 12436
rect 4890 12424 4896 12436
rect 4851 12396 4896 12424
rect 4890 12384 4896 12396
rect 4948 12384 4954 12436
rect 17221 12427 17279 12433
rect 17221 12393 17233 12427
rect 17267 12424 17279 12427
rect 17586 12424 17592 12436
rect 17267 12396 17592 12424
rect 17267 12393 17279 12396
rect 17221 12387 17279 12393
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 4706 12356 4712 12368
rect 2976 12328 4712 12356
rect 2976 12297 3004 12328
rect 4706 12316 4712 12328
rect 4764 12316 4770 12368
rect 2271 12260 2360 12288
rect 2961 12291 3019 12297
rect 2271 12257 2283 12260
rect 2225 12251 2283 12257
rect 2961 12257 2973 12291
rect 3007 12257 3019 12291
rect 2961 12251 3019 12257
rect 3602 12248 3608 12300
rect 3660 12288 3666 12300
rect 3881 12291 3939 12297
rect 3881 12288 3893 12291
rect 3660 12260 3893 12288
rect 3660 12248 3666 12260
rect 3881 12257 3893 12260
rect 3927 12257 3939 12291
rect 3881 12251 3939 12257
rect 15838 12248 15844 12300
rect 15896 12288 15902 12300
rect 17957 12291 18015 12297
rect 17957 12288 17969 12291
rect 15896 12260 17969 12288
rect 15896 12248 15902 12260
rect 17957 12257 17969 12260
rect 18003 12288 18015 12291
rect 18138 12288 18144 12300
rect 18003 12260 18144 12288
rect 18003 12257 18015 12260
rect 17957 12251 18015 12257
rect 18138 12248 18144 12260
rect 18196 12248 18202 12300
rect 1949 12223 2007 12229
rect 1949 12189 1961 12223
rect 1995 12220 2007 12223
rect 2590 12220 2596 12232
rect 1995 12192 2596 12220
rect 1995 12189 2007 12192
rect 1949 12183 2007 12189
rect 2590 12180 2596 12192
rect 2648 12180 2654 12232
rect 3234 12220 3240 12232
rect 3195 12192 3240 12220
rect 3234 12180 3240 12192
rect 3292 12220 3298 12232
rect 3510 12220 3516 12232
rect 3292 12192 3516 12220
rect 3292 12180 3298 12192
rect 3510 12180 3516 12192
rect 3568 12180 3574 12232
rect 3970 12180 3976 12232
rect 4028 12220 4034 12232
rect 5350 12229 5356 12232
rect 5077 12223 5135 12229
rect 5077 12220 5089 12223
rect 4028 12192 5089 12220
rect 4028 12180 4034 12192
rect 5077 12189 5089 12192
rect 5123 12189 5135 12223
rect 5344 12220 5356 12229
rect 5311 12192 5356 12220
rect 5077 12183 5135 12189
rect 5344 12183 5356 12192
rect 5350 12180 5356 12183
rect 5408 12180 5414 12232
rect 6914 12180 6920 12232
rect 6972 12220 6978 12232
rect 7745 12223 7803 12229
rect 7745 12220 7757 12223
rect 6972 12192 7757 12220
rect 6972 12180 6978 12192
rect 7745 12189 7757 12192
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 16853 12223 16911 12229
rect 16853 12189 16865 12223
rect 16899 12220 16911 12223
rect 17310 12220 17316 12232
rect 16899 12192 17316 12220
rect 16899 12189 16911 12192
rect 16853 12183 16911 12189
rect 17310 12180 17316 12192
rect 17368 12180 17374 12232
rect 17589 12223 17647 12229
rect 17589 12189 17601 12223
rect 17635 12220 17647 12223
rect 17678 12220 17684 12232
rect 17635 12192 17684 12220
rect 17635 12189 17647 12192
rect 17589 12183 17647 12189
rect 17678 12180 17684 12192
rect 17736 12180 17742 12232
rect 2498 12112 2504 12164
rect 2556 12152 2562 12164
rect 2777 12155 2835 12161
rect 2777 12152 2789 12155
rect 2556 12124 2789 12152
rect 2556 12112 2562 12124
rect 2777 12121 2789 12124
rect 2823 12121 2835 12155
rect 2777 12115 2835 12121
rect 3605 12155 3663 12161
rect 3605 12121 3617 12155
rect 3651 12152 3663 12155
rect 3694 12152 3700 12164
rect 3651 12124 3700 12152
rect 3651 12121 3663 12124
rect 3605 12115 3663 12121
rect 3694 12112 3700 12124
rect 3752 12152 3758 12164
rect 4157 12155 4215 12161
rect 4157 12152 4169 12155
rect 3752 12124 4169 12152
rect 3752 12112 3758 12124
rect 4157 12121 4169 12124
rect 4203 12152 4215 12155
rect 4203 12124 8524 12152
rect 4203 12121 4215 12124
rect 4157 12115 4215 12121
rect 2314 12084 2320 12096
rect 2275 12056 2320 12084
rect 2314 12044 2320 12056
rect 2372 12044 2378 12096
rect 2406 12044 2412 12096
rect 2464 12084 2470 12096
rect 2685 12087 2743 12093
rect 2685 12084 2697 12087
rect 2464 12056 2697 12084
rect 2464 12044 2470 12056
rect 2685 12053 2697 12056
rect 2731 12053 2743 12087
rect 2685 12047 2743 12053
rect 3329 12087 3387 12093
rect 3329 12053 3341 12087
rect 3375 12084 3387 12087
rect 3970 12084 3976 12096
rect 3375 12056 3976 12084
rect 3375 12053 3387 12056
rect 3329 12047 3387 12053
rect 3970 12044 3976 12056
rect 4028 12044 4034 12096
rect 4065 12087 4123 12093
rect 4065 12053 4077 12087
rect 4111 12084 4123 12087
rect 4338 12084 4344 12096
rect 4111 12056 4344 12084
rect 4111 12053 4123 12056
rect 4065 12047 4123 12053
rect 4338 12044 4344 12056
rect 4396 12084 4402 12096
rect 4617 12087 4675 12093
rect 4617 12084 4629 12087
rect 4396 12056 4629 12084
rect 4396 12044 4402 12056
rect 4617 12053 4629 12056
rect 4663 12053 4675 12087
rect 6454 12084 6460 12096
rect 6415 12056 6460 12084
rect 4617 12047 4675 12053
rect 6454 12044 6460 12056
rect 6512 12044 6518 12096
rect 8496 12084 8524 12124
rect 8570 12112 8576 12164
rect 8628 12152 8634 12164
rect 8628 12124 8673 12152
rect 8628 12112 8634 12124
rect 14918 12112 14924 12164
rect 14976 12152 14982 12164
rect 17954 12152 17960 12164
rect 14976 12124 17960 12152
rect 14976 12112 14982 12124
rect 17954 12112 17960 12124
rect 18012 12112 18018 12164
rect 10226 12084 10232 12096
rect 8496 12056 10232 12084
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 16945 12087 17003 12093
rect 16945 12084 16957 12087
rect 13872 12056 16957 12084
rect 13872 12044 13878 12056
rect 16945 12053 16957 12056
rect 16991 12053 17003 12087
rect 17402 12084 17408 12096
rect 17315 12056 17408 12084
rect 16945 12047 17003 12053
rect 17402 12044 17408 12056
rect 17460 12084 17466 12096
rect 17862 12084 17868 12096
rect 17460 12056 17868 12084
rect 17460 12044 17466 12056
rect 17862 12044 17868 12056
rect 17920 12044 17926 12096
rect 1104 11994 18860 12016
rect 1104 11942 5398 11994
rect 5450 11942 5462 11994
rect 5514 11942 5526 11994
rect 5578 11942 5590 11994
rect 5642 11942 5654 11994
rect 5706 11942 9846 11994
rect 9898 11942 9910 11994
rect 9962 11942 9974 11994
rect 10026 11942 10038 11994
rect 10090 11942 10102 11994
rect 10154 11942 14294 11994
rect 14346 11942 14358 11994
rect 14410 11942 14422 11994
rect 14474 11942 14486 11994
rect 14538 11942 14550 11994
rect 14602 11942 18860 11994
rect 1104 11920 18860 11942
rect 2406 11880 2412 11892
rect 2367 11852 2412 11880
rect 2406 11840 2412 11852
rect 2464 11840 2470 11892
rect 2958 11880 2964 11892
rect 2746 11852 2964 11880
rect 2746 11812 2774 11852
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 3421 11883 3479 11889
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 3786 11880 3792 11892
rect 3467 11852 3792 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 3786 11840 3792 11852
rect 3844 11840 3850 11892
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 8294 11880 8300 11892
rect 4028 11852 8300 11880
rect 4028 11840 4034 11852
rect 8294 11840 8300 11852
rect 8352 11880 8358 11892
rect 13630 11880 13636 11892
rect 8352 11852 13636 11880
rect 8352 11840 8358 11852
rect 13630 11840 13636 11852
rect 13688 11840 13694 11892
rect 17126 11840 17132 11892
rect 17184 11880 17190 11892
rect 18046 11880 18052 11892
rect 17184 11852 18052 11880
rect 17184 11840 17190 11852
rect 18046 11840 18052 11852
rect 18104 11840 18110 11892
rect 1964 11784 2774 11812
rect 1964 11753 1992 11784
rect 2866 11772 2872 11824
rect 2924 11772 2930 11824
rect 3436 11784 3832 11812
rect 1949 11747 2007 11753
rect 1949 11713 1961 11747
rect 1995 11713 2007 11747
rect 1949 11707 2007 11713
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11744 2835 11747
rect 2884 11744 2912 11772
rect 3436 11744 3464 11784
rect 2823 11716 3464 11744
rect 3513 11747 3571 11753
rect 2823 11713 2835 11716
rect 2777 11707 2835 11713
rect 3513 11713 3525 11747
rect 3559 11744 3571 11747
rect 3694 11744 3700 11756
rect 3559 11716 3700 11744
rect 3559 11713 3571 11716
rect 3513 11707 3571 11713
rect 3694 11704 3700 11716
rect 3752 11704 3758 11756
rect 3804 11744 3832 11784
rect 3878 11772 3884 11824
rect 3936 11812 3942 11824
rect 3936 11784 5304 11812
rect 3936 11772 3942 11784
rect 3970 11744 3976 11756
rect 3804 11716 3976 11744
rect 3970 11704 3976 11716
rect 4028 11704 4034 11756
rect 4706 11704 4712 11756
rect 4764 11744 4770 11756
rect 5276 11753 5304 11784
rect 6454 11772 6460 11824
rect 6512 11812 6518 11824
rect 6610 11815 6668 11821
rect 6610 11812 6622 11815
rect 6512 11784 6622 11812
rect 6512 11772 6518 11784
rect 6610 11781 6622 11784
rect 6656 11781 6668 11815
rect 6610 11775 6668 11781
rect 7006 11772 7012 11824
rect 7064 11812 7070 11824
rect 7064 11784 9674 11812
rect 7064 11772 7070 11784
rect 4994 11747 5052 11753
rect 4994 11744 5006 11747
rect 4764 11716 5006 11744
rect 4764 11704 4770 11716
rect 4994 11713 5006 11716
rect 5040 11713 5052 11747
rect 4994 11707 5052 11713
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11744 5319 11747
rect 6362 11744 6368 11756
rect 5307 11716 6368 11744
rect 5307 11713 5319 11716
rect 5261 11707 5319 11713
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 8386 11744 8392 11756
rect 8347 11716 8392 11744
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 9646 11744 9674 11784
rect 12802 11772 12808 11824
rect 12860 11812 12866 11824
rect 13998 11812 14004 11824
rect 12860 11784 14004 11812
rect 12860 11772 12866 11784
rect 13998 11772 14004 11784
rect 14056 11772 14062 11824
rect 17037 11815 17095 11821
rect 17037 11781 17049 11815
rect 17083 11812 17095 11815
rect 17083 11784 17724 11812
rect 17083 11781 17095 11784
rect 17037 11775 17095 11781
rect 15838 11744 15844 11756
rect 9646 11716 15844 11744
rect 15838 11704 15844 11716
rect 15896 11704 15902 11756
rect 17221 11747 17279 11753
rect 17221 11713 17233 11747
rect 17267 11744 17279 11747
rect 17494 11744 17500 11756
rect 17267 11716 17500 11744
rect 17267 11713 17279 11716
rect 17221 11707 17279 11713
rect 17494 11704 17500 11716
rect 17552 11704 17558 11756
rect 17696 11753 17724 11784
rect 17681 11747 17739 11753
rect 17681 11713 17693 11747
rect 17727 11744 17739 11747
rect 17770 11744 17776 11756
rect 17727 11716 17776 11744
rect 17727 11713 17739 11716
rect 17681 11707 17739 11713
rect 17770 11704 17776 11716
rect 17828 11704 17834 11756
rect 2222 11676 2228 11688
rect 2183 11648 2228 11676
rect 2222 11636 2228 11648
rect 2280 11636 2286 11688
rect 2866 11676 2872 11688
rect 2827 11648 2872 11676
rect 2866 11636 2872 11648
rect 2924 11636 2930 11688
rect 3050 11636 3056 11688
rect 3108 11676 3114 11688
rect 3602 11676 3608 11688
rect 3108 11648 3608 11676
rect 3108 11636 3114 11648
rect 3602 11636 3608 11648
rect 3660 11636 3666 11688
rect 15746 11636 15752 11688
rect 15804 11676 15810 11688
rect 17310 11676 17316 11688
rect 15804 11648 17316 11676
rect 15804 11636 15810 11648
rect 17310 11636 17316 11648
rect 17368 11636 17374 11688
rect 17954 11676 17960 11688
rect 17915 11648 17960 11676
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 3697 11611 3755 11617
rect 3697 11577 3709 11611
rect 3743 11608 3755 11611
rect 3743 11580 4384 11608
rect 3743 11577 3755 11580
rect 3697 11571 3755 11577
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3602 11540 3608 11552
rect 3016 11512 3608 11540
rect 3016 11500 3022 11512
rect 3602 11500 3608 11512
rect 3660 11500 3666 11552
rect 3881 11543 3939 11549
rect 3881 11509 3893 11543
rect 3927 11540 3939 11543
rect 4154 11540 4160 11552
rect 3927 11512 4160 11540
rect 3927 11509 3939 11512
rect 3881 11503 3939 11509
rect 4154 11500 4160 11512
rect 4212 11500 4218 11552
rect 4356 11540 4384 11580
rect 15102 11568 15108 11620
rect 15160 11608 15166 11620
rect 16393 11611 16451 11617
rect 16393 11608 16405 11611
rect 15160 11580 16405 11608
rect 15160 11568 15166 11580
rect 16393 11577 16405 11580
rect 16439 11577 16451 11611
rect 16393 11571 16451 11577
rect 16853 11611 16911 11617
rect 16853 11577 16865 11611
rect 16899 11608 16911 11611
rect 17770 11608 17776 11620
rect 16899 11580 17776 11608
rect 16899 11577 16911 11580
rect 16853 11571 16911 11577
rect 17770 11568 17776 11580
rect 17828 11568 17834 11620
rect 6086 11540 6092 11552
rect 4356 11512 6092 11540
rect 6086 11500 6092 11512
rect 6144 11500 6150 11552
rect 7466 11500 7472 11552
rect 7524 11540 7530 11552
rect 7745 11543 7803 11549
rect 7745 11540 7757 11543
rect 7524 11512 7757 11540
rect 7524 11500 7530 11512
rect 7745 11509 7757 11512
rect 7791 11509 7803 11543
rect 7745 11503 7803 11509
rect 8110 11500 8116 11552
rect 8168 11540 8174 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8168 11512 9045 11540
rect 8168 11500 8174 11512
rect 9033 11509 9045 11512
rect 9079 11509 9091 11543
rect 9033 11503 9091 11509
rect 10226 11500 10232 11552
rect 10284 11540 10290 11552
rect 15654 11540 15660 11552
rect 10284 11512 15660 11540
rect 10284 11500 10290 11512
rect 15654 11500 15660 11512
rect 15712 11540 15718 11552
rect 16117 11543 16175 11549
rect 16117 11540 16129 11543
rect 15712 11512 16129 11540
rect 15712 11500 15718 11512
rect 16117 11509 16129 11512
rect 16163 11509 16175 11543
rect 17402 11540 17408 11552
rect 17363 11512 17408 11540
rect 16117 11503 16175 11509
rect 17402 11500 17408 11512
rect 17460 11500 17466 11552
rect 1104 11450 18860 11472
rect 1104 11398 3174 11450
rect 3226 11398 3238 11450
rect 3290 11398 3302 11450
rect 3354 11398 3366 11450
rect 3418 11398 3430 11450
rect 3482 11398 7622 11450
rect 7674 11398 7686 11450
rect 7738 11398 7750 11450
rect 7802 11398 7814 11450
rect 7866 11398 7878 11450
rect 7930 11398 12070 11450
rect 12122 11398 12134 11450
rect 12186 11398 12198 11450
rect 12250 11398 12262 11450
rect 12314 11398 12326 11450
rect 12378 11398 16518 11450
rect 16570 11398 16582 11450
rect 16634 11398 16646 11450
rect 16698 11398 16710 11450
rect 16762 11398 16774 11450
rect 16826 11398 18860 11450
rect 1104 11376 18860 11398
rect 2498 11336 2504 11348
rect 2459 11308 2504 11336
rect 2498 11296 2504 11308
rect 2556 11296 2562 11348
rect 3421 11339 3479 11345
rect 3421 11305 3433 11339
rect 3467 11336 3479 11339
rect 3510 11336 3516 11348
rect 3467 11308 3516 11336
rect 3467 11305 3479 11308
rect 3421 11299 3479 11305
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 3694 11296 3700 11348
rect 3752 11336 3758 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 3752 11308 3801 11336
rect 3752 11296 3758 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 3789 11299 3847 11305
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4341 11339 4399 11345
rect 4341 11336 4353 11339
rect 4120 11308 4353 11336
rect 4120 11296 4126 11308
rect 4341 11305 4353 11308
rect 4387 11305 4399 11339
rect 8386 11336 8392 11348
rect 4341 11299 4399 11305
rect 5184 11308 8392 11336
rect 3605 11271 3663 11277
rect 3605 11237 3617 11271
rect 3651 11268 3663 11271
rect 3970 11268 3976 11280
rect 3651 11240 3976 11268
rect 3651 11237 3663 11240
rect 3605 11231 3663 11237
rect 3970 11228 3976 11240
rect 4028 11228 4034 11280
rect 4246 11228 4252 11280
rect 4304 11268 4310 11280
rect 4525 11271 4583 11277
rect 4525 11268 4537 11271
rect 4304 11240 4537 11268
rect 4304 11228 4310 11240
rect 4525 11237 4537 11240
rect 4571 11237 4583 11271
rect 4525 11231 4583 11237
rect 2958 11200 2964 11212
rect 2919 11172 2964 11200
rect 2958 11160 2964 11172
rect 3016 11160 3022 11212
rect 3050 11160 3056 11212
rect 3108 11200 3114 11212
rect 3108 11172 3153 11200
rect 3108 11160 3114 11172
rect 3418 11160 3424 11212
rect 3476 11200 3482 11212
rect 5184 11209 5212 11308
rect 8386 11296 8392 11308
rect 8444 11296 8450 11348
rect 11146 11296 11152 11348
rect 11204 11336 11210 11348
rect 12253 11339 12311 11345
rect 12253 11336 12265 11339
rect 11204 11308 12265 11336
rect 11204 11296 11210 11308
rect 12253 11305 12265 11308
rect 12299 11336 12311 11339
rect 12710 11336 12716 11348
rect 12299 11308 12716 11336
rect 12299 11305 12311 11308
rect 12253 11299 12311 11305
rect 12710 11296 12716 11308
rect 12768 11336 12774 11348
rect 17221 11339 17279 11345
rect 17221 11336 17233 11339
rect 12768 11308 17233 11336
rect 12768 11296 12774 11308
rect 17221 11305 17233 11308
rect 17267 11336 17279 11339
rect 17586 11336 17592 11348
rect 17267 11308 17592 11336
rect 17267 11305 17279 11308
rect 17221 11299 17279 11305
rect 17586 11296 17592 11308
rect 17644 11296 17650 11348
rect 6549 11271 6607 11277
rect 6549 11268 6561 11271
rect 5920 11240 6561 11268
rect 4157 11203 4215 11209
rect 4157 11200 4169 11203
rect 3476 11172 4169 11200
rect 3476 11160 3482 11172
rect 4157 11169 4169 11172
rect 4203 11169 4215 11203
rect 4157 11163 4215 11169
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 1946 11132 1952 11144
rect 1907 11104 1952 11132
rect 1946 11092 1952 11104
rect 2004 11092 2010 11144
rect 2222 11132 2228 11144
rect 2183 11104 2228 11132
rect 2222 11092 2228 11104
rect 2280 11132 2286 11144
rect 3973 11135 4031 11141
rect 3973 11132 3985 11135
rect 2280 11104 3985 11132
rect 2280 11092 2286 11104
rect 3973 11101 3985 11104
rect 4019 11101 4031 11135
rect 4890 11132 4896 11144
rect 4851 11104 4896 11132
rect 3973 11095 4031 11101
rect 4890 11092 4896 11104
rect 4948 11092 4954 11144
rect 5810 11132 5816 11144
rect 5771 11104 5816 11132
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 2869 11067 2927 11073
rect 2869 11033 2881 11067
rect 2915 11064 2927 11067
rect 3050 11064 3056 11076
rect 2915 11036 3056 11064
rect 2915 11033 2927 11036
rect 2869 11027 2927 11033
rect 3050 11024 3056 11036
rect 3108 11024 3114 11076
rect 5718 11024 5724 11076
rect 5776 11064 5782 11076
rect 5920 11073 5948 11240
rect 6549 11237 6561 11240
rect 6595 11268 6607 11271
rect 6730 11268 6736 11280
rect 6595 11240 6736 11268
rect 6595 11237 6607 11240
rect 6549 11231 6607 11237
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 15746 11268 15752 11280
rect 15707 11240 15752 11268
rect 15746 11228 15752 11240
rect 15804 11228 15810 11280
rect 15838 11228 15844 11280
rect 15896 11268 15902 11280
rect 16025 11271 16083 11277
rect 16025 11268 16037 11271
rect 15896 11240 16037 11268
rect 15896 11228 15902 11240
rect 16025 11237 16037 11240
rect 16071 11237 16083 11271
rect 16025 11231 16083 11237
rect 6089 11203 6147 11209
rect 6089 11169 6101 11203
rect 6135 11169 6147 11203
rect 6089 11163 6147 11169
rect 5905 11067 5963 11073
rect 5905 11064 5917 11067
rect 5776 11036 5917 11064
rect 5776 11024 5782 11036
rect 5905 11033 5917 11036
rect 5951 11033 5963 11067
rect 6104 11064 6132 11163
rect 14642 11160 14648 11212
rect 14700 11200 14706 11212
rect 17957 11203 18015 11209
rect 17957 11200 17969 11203
rect 14700 11172 17969 11200
rect 14700 11160 14706 11172
rect 17957 11169 17969 11172
rect 18003 11169 18015 11203
rect 17957 11163 18015 11169
rect 6362 11092 6368 11144
rect 6420 11132 6426 11144
rect 8113 11135 8171 11141
rect 8113 11132 8125 11135
rect 6420 11104 8125 11132
rect 6420 11092 6426 11104
rect 8113 11101 8125 11104
rect 8159 11101 8171 11135
rect 8113 11095 8171 11101
rect 10321 11135 10379 11141
rect 10321 11101 10333 11135
rect 10367 11132 10379 11135
rect 11885 11135 11943 11141
rect 11885 11132 11897 11135
rect 10367 11104 11897 11132
rect 10367 11101 10379 11104
rect 10321 11095 10379 11101
rect 11885 11101 11897 11104
rect 11931 11132 11943 11135
rect 13909 11135 13967 11141
rect 13909 11132 13921 11135
rect 11931 11104 13921 11132
rect 11931 11101 11943 11104
rect 11885 11095 11943 11101
rect 13909 11101 13921 11104
rect 13955 11132 13967 11135
rect 14182 11132 14188 11144
rect 13955 11104 14188 11132
rect 13955 11101 13967 11104
rect 13909 11095 13967 11101
rect 14182 11092 14188 11104
rect 14240 11092 14246 11144
rect 15470 11132 15476 11144
rect 15431 11104 15476 11132
rect 15470 11092 15476 11104
rect 15528 11092 15534 11144
rect 15933 11135 15991 11141
rect 15933 11101 15945 11135
rect 15979 11132 15991 11135
rect 16390 11132 16396 11144
rect 15979 11104 16396 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 17218 11092 17224 11144
rect 17276 11132 17282 11144
rect 17402 11132 17408 11144
rect 17276 11104 17408 11132
rect 17276 11092 17282 11104
rect 17402 11092 17408 11104
rect 17460 11092 17466 11144
rect 17586 11132 17592 11144
rect 17547 11104 17592 11132
rect 17586 11092 17592 11104
rect 17644 11092 17650 11144
rect 17678 11092 17684 11144
rect 17736 11132 17742 11144
rect 17736 11104 17781 11132
rect 17736 11092 17742 11104
rect 6822 11064 6828 11076
rect 6104 11036 6828 11064
rect 5905 11027 5963 11033
rect 6822 11024 6828 11036
rect 6880 11064 6886 11076
rect 7466 11064 7472 11076
rect 6880 11036 7472 11064
rect 6880 11024 6886 11036
rect 7466 11024 7472 11036
rect 7524 11064 7530 11076
rect 7846 11067 7904 11073
rect 7846 11064 7858 11067
rect 7524 11036 7858 11064
rect 7524 11024 7530 11036
rect 7846 11033 7858 11036
rect 7892 11033 7904 11067
rect 7846 11027 7904 11033
rect 10076 11067 10134 11073
rect 10076 11033 10088 11067
rect 10122 11064 10134 11067
rect 11640 11067 11698 11073
rect 10122 11036 10548 11064
rect 10122 11033 10134 11036
rect 10076 11027 10134 11033
rect 2406 10996 2412 11008
rect 2367 10968 2412 10996
rect 2406 10956 2412 10968
rect 2464 10956 2470 11008
rect 4982 10996 4988 11008
rect 4943 10968 4988 10996
rect 4982 10956 4988 10968
rect 5040 10956 5046 11008
rect 5074 10956 5080 11008
rect 5132 10996 5138 11008
rect 5445 10999 5503 11005
rect 5445 10996 5457 10999
rect 5132 10968 5457 10996
rect 5132 10956 5138 10968
rect 5445 10965 5457 10968
rect 5491 10965 5503 10999
rect 6270 10996 6276 11008
rect 6231 10968 6276 10996
rect 5445 10959 5503 10965
rect 6270 10956 6276 10968
rect 6328 10956 6334 11008
rect 6733 10999 6791 11005
rect 6733 10965 6745 10999
rect 6779 10996 6791 10999
rect 7282 10996 7288 11008
rect 6779 10968 7288 10996
rect 6779 10965 6791 10968
rect 6733 10959 6791 10965
rect 7282 10956 7288 10968
rect 7340 10956 7346 11008
rect 8941 10999 8999 11005
rect 8941 10965 8953 10999
rect 8987 10996 8999 10999
rect 9030 10996 9036 11008
rect 8987 10968 9036 10996
rect 8987 10965 8999 10968
rect 8941 10959 8999 10965
rect 9030 10956 9036 10968
rect 9088 10956 9094 11008
rect 10520 11005 10548 11036
rect 11640 11033 11652 11067
rect 11686 11064 11698 11067
rect 11686 11036 12434 11064
rect 11686 11033 11698 11036
rect 11640 11027 11698 11033
rect 10505 10999 10563 11005
rect 10505 10965 10517 10999
rect 10551 10996 10563 10999
rect 10686 10996 10692 11008
rect 10551 10968 10692 10996
rect 10551 10965 10563 10968
rect 10505 10959 10563 10965
rect 10686 10956 10692 10968
rect 10744 10956 10750 11008
rect 12406 10996 12434 11036
rect 13446 11024 13452 11076
rect 13504 11064 13510 11076
rect 13642 11067 13700 11073
rect 13642 11064 13654 11067
rect 13504 11036 13654 11064
rect 13504 11024 13510 11036
rect 13642 11033 13654 11036
rect 13688 11033 13700 11067
rect 13642 11027 13700 11033
rect 15286 11024 15292 11076
rect 15344 11064 15350 11076
rect 15344 11036 15792 11064
rect 15344 11024 15350 11036
rect 12529 10999 12587 11005
rect 12529 10996 12541 10999
rect 12406 10968 12541 10996
rect 12529 10965 12541 10968
rect 12575 10996 12587 10999
rect 12894 10996 12900 11008
rect 12575 10968 12900 10996
rect 12575 10965 12587 10968
rect 12529 10959 12587 10965
rect 12894 10956 12900 10968
rect 12952 10956 12958 11008
rect 15764 10996 15792 11036
rect 15838 11024 15844 11076
rect 15896 11064 15902 11076
rect 16485 11067 16543 11073
rect 16485 11064 16497 11067
rect 15896 11036 16497 11064
rect 15896 11024 15902 11036
rect 16485 11033 16497 11036
rect 16531 11033 16543 11067
rect 16485 11027 16543 11033
rect 16945 11067 17003 11073
rect 16945 11033 16957 11067
rect 16991 11064 17003 11067
rect 17696 11064 17724 11092
rect 16991 11036 17724 11064
rect 16991 11033 17003 11036
rect 16945 11027 17003 11033
rect 16209 10999 16267 11005
rect 16209 10996 16221 10999
rect 15764 10968 16221 10996
rect 16209 10965 16221 10968
rect 16255 10965 16267 10999
rect 16666 10996 16672 11008
rect 16627 10968 16672 10996
rect 16209 10959 16267 10965
rect 16666 10956 16672 10968
rect 16724 10956 16730 11008
rect 17126 10996 17132 11008
rect 17087 10968 17132 10996
rect 17126 10956 17132 10968
rect 17184 10956 17190 11008
rect 17218 10956 17224 11008
rect 17276 10996 17282 11008
rect 17405 10999 17463 11005
rect 17405 10996 17417 10999
rect 17276 10968 17417 10996
rect 17276 10956 17282 10968
rect 17405 10965 17417 10968
rect 17451 10965 17463 10999
rect 17405 10959 17463 10965
rect 1104 10906 18860 10928
rect 1104 10854 5398 10906
rect 5450 10854 5462 10906
rect 5514 10854 5526 10906
rect 5578 10854 5590 10906
rect 5642 10854 5654 10906
rect 5706 10854 9846 10906
rect 9898 10854 9910 10906
rect 9962 10854 9974 10906
rect 10026 10854 10038 10906
rect 10090 10854 10102 10906
rect 10154 10854 14294 10906
rect 14346 10854 14358 10906
rect 14410 10854 14422 10906
rect 14474 10854 14486 10906
rect 14538 10854 14550 10906
rect 14602 10854 18860 10906
rect 1104 10832 18860 10854
rect 1949 10795 2007 10801
rect 1949 10761 1961 10795
rect 1995 10792 2007 10795
rect 2314 10792 2320 10804
rect 1995 10764 2320 10792
rect 1995 10761 2007 10764
rect 1949 10755 2007 10761
rect 2314 10752 2320 10764
rect 2372 10752 2378 10804
rect 2501 10795 2559 10801
rect 2501 10761 2513 10795
rect 2547 10792 2559 10795
rect 3142 10792 3148 10804
rect 2547 10764 3148 10792
rect 2547 10761 2559 10764
rect 2501 10755 2559 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 4154 10792 4160 10804
rect 3436 10764 4160 10792
rect 3436 10724 3464 10764
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4617 10795 4675 10801
rect 4617 10761 4629 10795
rect 4663 10792 4675 10795
rect 4890 10792 4896 10804
rect 4663 10764 4896 10792
rect 4663 10761 4675 10764
rect 4617 10755 4675 10761
rect 4890 10752 4896 10764
rect 4948 10752 4954 10804
rect 5074 10792 5080 10804
rect 5035 10764 5080 10792
rect 5074 10752 5080 10764
rect 5132 10752 5138 10804
rect 5445 10795 5503 10801
rect 5445 10761 5457 10795
rect 5491 10761 5503 10795
rect 5445 10755 5503 10761
rect 5813 10795 5871 10801
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 6270 10792 6276 10804
rect 5859 10764 6276 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 1872 10696 3464 10724
rect 1578 10656 1584 10668
rect 1539 10628 1584 10656
rect 1578 10616 1584 10628
rect 1636 10616 1642 10668
rect 1872 10597 1900 10696
rect 3510 10684 3516 10736
rect 3568 10724 3574 10736
rect 3614 10727 3672 10733
rect 3614 10724 3626 10727
rect 3568 10696 3626 10724
rect 3568 10684 3574 10696
rect 3614 10693 3626 10696
rect 3660 10693 3672 10727
rect 3614 10687 3672 10693
rect 4985 10727 5043 10733
rect 4985 10693 4997 10727
rect 5031 10724 5043 10727
rect 5460 10724 5488 10755
rect 6270 10752 6276 10764
rect 6328 10752 6334 10804
rect 8386 10792 8392 10804
rect 8347 10764 8392 10792
rect 8386 10752 8392 10764
rect 8444 10752 8450 10804
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 12345 10795 12403 10801
rect 12345 10792 12357 10795
rect 11931 10764 12357 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 12345 10761 12357 10764
rect 12391 10761 12403 10795
rect 12710 10792 12716 10804
rect 12671 10764 12716 10792
rect 12345 10755 12403 10761
rect 12710 10752 12716 10764
rect 12768 10752 12774 10804
rect 12805 10795 12863 10801
rect 12805 10761 12817 10795
rect 12851 10792 12863 10795
rect 13173 10795 13231 10801
rect 13173 10792 13185 10795
rect 12851 10764 13185 10792
rect 12851 10761 12863 10764
rect 12805 10755 12863 10761
rect 13173 10761 13185 10764
rect 13219 10761 13231 10795
rect 13538 10792 13544 10804
rect 13451 10764 13544 10792
rect 13173 10755 13231 10761
rect 13538 10752 13544 10764
rect 13596 10792 13602 10804
rect 14277 10795 14335 10801
rect 14277 10792 14289 10795
rect 13596 10764 14289 10792
rect 13596 10752 13602 10764
rect 14277 10761 14289 10764
rect 14323 10792 14335 10795
rect 17954 10792 17960 10804
rect 14323 10764 17960 10792
rect 14323 10761 14335 10764
rect 14277 10755 14335 10761
rect 17954 10752 17960 10764
rect 18012 10752 18018 10804
rect 7282 10733 7288 10736
rect 7276 10724 7288 10733
rect 5031 10696 5488 10724
rect 5828 10696 7288 10724
rect 5031 10693 5043 10696
rect 4985 10687 5043 10693
rect 2041 10659 2099 10665
rect 2041 10625 2053 10659
rect 2087 10656 2099 10659
rect 4798 10656 4804 10668
rect 2087 10628 4804 10656
rect 2087 10625 2099 10628
rect 2041 10619 2099 10625
rect 4798 10616 4804 10628
rect 4856 10616 4862 10668
rect 1857 10591 1915 10597
rect 1857 10557 1869 10591
rect 1903 10557 1915 10591
rect 3878 10588 3884 10600
rect 3839 10560 3884 10588
rect 1857 10551 1915 10557
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 5261 10591 5319 10597
rect 5261 10557 5273 10591
rect 5307 10588 5319 10591
rect 5442 10588 5448 10600
rect 5307 10560 5448 10588
rect 5307 10557 5319 10560
rect 5261 10551 5319 10557
rect 5442 10548 5448 10560
rect 5500 10588 5506 10600
rect 5828 10588 5856 10696
rect 7276 10687 7288 10696
rect 7282 10684 7288 10687
rect 7340 10684 7346 10736
rect 14090 10684 14096 10736
rect 14148 10724 14154 10736
rect 14645 10727 14703 10733
rect 14645 10724 14657 10727
rect 14148 10696 14657 10724
rect 14148 10684 14154 10696
rect 14645 10693 14657 10696
rect 14691 10724 14703 10727
rect 16669 10727 16727 10733
rect 16669 10724 16681 10727
rect 14691 10696 16681 10724
rect 14691 10693 14703 10696
rect 14645 10687 14703 10693
rect 16669 10693 16681 10696
rect 16715 10724 16727 10727
rect 17126 10724 17132 10736
rect 16715 10696 16988 10724
rect 17087 10696 17132 10724
rect 16715 10693 16727 10696
rect 16669 10687 16727 10693
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 5960 10628 6005 10656
rect 5960 10616 5966 10628
rect 6362 10616 6368 10668
rect 6420 10656 6426 10668
rect 6822 10656 6828 10668
rect 6420 10628 6828 10656
rect 6420 10616 6426 10628
rect 6822 10616 6828 10628
rect 6880 10656 6886 10668
rect 7009 10659 7067 10665
rect 7009 10656 7021 10659
rect 6880 10628 7021 10656
rect 6880 10616 6886 10628
rect 7009 10625 7021 10628
rect 7055 10625 7067 10659
rect 8478 10656 8484 10668
rect 7009 10619 7067 10625
rect 7116 10628 8484 10656
rect 5500 10560 5856 10588
rect 6089 10591 6147 10597
rect 5500 10548 5506 10560
rect 6089 10557 6101 10591
rect 6135 10588 6147 10591
rect 6730 10588 6736 10600
rect 6135 10560 6736 10588
rect 6135 10557 6147 10560
rect 6089 10551 6147 10557
rect 6730 10548 6736 10560
rect 6788 10548 6794 10600
rect 7116 10588 7144 10628
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 9030 10656 9036 10668
rect 8991 10628 9036 10656
rect 9030 10616 9036 10628
rect 9088 10616 9094 10668
rect 10413 10659 10471 10665
rect 10413 10625 10425 10659
rect 10459 10656 10471 10659
rect 11330 10656 11336 10668
rect 10459 10628 11336 10656
rect 10459 10625 10471 10628
rect 10413 10619 10471 10625
rect 11330 10616 11336 10628
rect 11388 10616 11394 10668
rect 13630 10656 13636 10668
rect 13543 10628 13636 10656
rect 13630 10616 13636 10628
rect 13688 10656 13694 10668
rect 14001 10659 14059 10665
rect 14001 10656 14013 10659
rect 13688 10628 14013 10656
rect 13688 10616 13694 10628
rect 14001 10625 14013 10628
rect 14047 10625 14059 10659
rect 15562 10656 15568 10668
rect 15523 10628 15568 10656
rect 14001 10619 14059 10625
rect 15562 10616 15568 10628
rect 15620 10616 15626 10668
rect 15657 10659 15715 10665
rect 15657 10625 15669 10659
rect 15703 10656 15715 10659
rect 16850 10656 16856 10668
rect 15703 10628 16856 10656
rect 15703 10625 15715 10628
rect 15657 10619 15715 10625
rect 16850 10616 16856 10628
rect 16908 10616 16914 10668
rect 16960 10656 16988 10696
rect 17126 10684 17132 10696
rect 17184 10684 17190 10736
rect 17221 10659 17279 10665
rect 17221 10656 17233 10659
rect 16960 10628 17233 10656
rect 17221 10625 17233 10628
rect 17267 10656 17279 10659
rect 18598 10656 18604 10668
rect 17267 10628 18604 10656
rect 17267 10625 17279 10628
rect 17221 10619 17279 10625
rect 18598 10616 18604 10628
rect 18656 10616 18662 10668
rect 10502 10588 10508 10600
rect 6840 10560 7144 10588
rect 10463 10560 10508 10588
rect 4065 10523 4123 10529
rect 4065 10489 4077 10523
rect 4111 10520 4123 10523
rect 6840 10520 6868 10560
rect 10502 10548 10508 10560
rect 10560 10548 10566 10600
rect 10686 10548 10692 10600
rect 10744 10588 10750 10600
rect 11149 10591 11207 10597
rect 10744 10560 10837 10588
rect 10744 10548 10750 10560
rect 11149 10557 11161 10591
rect 11195 10588 11207 10591
rect 11698 10588 11704 10600
rect 11195 10560 11704 10588
rect 11195 10557 11207 10560
rect 11149 10551 11207 10557
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 11974 10588 11980 10600
rect 11935 10560 11980 10588
rect 11974 10548 11980 10560
rect 12032 10548 12038 10600
rect 12069 10591 12127 10597
rect 12069 10557 12081 10591
rect 12115 10557 12127 10591
rect 12894 10588 12900 10600
rect 12855 10560 12900 10588
rect 12069 10551 12127 10557
rect 4111 10492 6868 10520
rect 9677 10523 9735 10529
rect 4111 10489 4123 10492
rect 4065 10483 4123 10489
rect 9677 10489 9689 10523
rect 9723 10520 9735 10523
rect 10318 10520 10324 10532
rect 9723 10492 10324 10520
rect 9723 10489 9735 10492
rect 9677 10483 9735 10489
rect 1394 10452 1400 10464
rect 1355 10424 1400 10452
rect 1394 10412 1400 10424
rect 1452 10412 1458 10464
rect 2409 10455 2467 10461
rect 2409 10421 2421 10455
rect 2455 10452 2467 10455
rect 2682 10452 2688 10464
rect 2455 10424 2688 10452
rect 2455 10421 2467 10424
rect 2409 10415 2467 10421
rect 2682 10412 2688 10424
rect 2740 10412 2746 10464
rect 3694 10412 3700 10464
rect 3752 10452 3758 10464
rect 4080 10452 4108 10483
rect 10318 10480 10324 10492
rect 10376 10480 10382 10532
rect 10704 10520 10732 10548
rect 12084 10520 12112 10551
rect 12894 10548 12900 10560
rect 12952 10548 12958 10600
rect 13446 10548 13452 10600
rect 13504 10588 13510 10600
rect 13725 10591 13783 10597
rect 13725 10588 13737 10591
rect 13504 10560 13737 10588
rect 13504 10548 13510 10560
rect 13725 10557 13737 10560
rect 13771 10557 13783 10591
rect 13725 10551 13783 10557
rect 15746 10548 15752 10600
rect 15804 10588 15810 10600
rect 15804 10560 15849 10588
rect 15804 10548 15810 10560
rect 16114 10548 16120 10600
rect 16172 10588 16178 10600
rect 16945 10591 17003 10597
rect 16945 10588 16957 10591
rect 16172 10560 16957 10588
rect 16172 10548 16178 10560
rect 16945 10557 16957 10560
rect 16991 10557 17003 10591
rect 17678 10588 17684 10600
rect 17639 10560 17684 10588
rect 16945 10551 17003 10557
rect 17678 10548 17684 10560
rect 17736 10548 17742 10600
rect 17954 10588 17960 10600
rect 17915 10560 17960 10588
rect 17954 10548 17960 10560
rect 18012 10548 18018 10600
rect 10704 10492 12112 10520
rect 14090 10480 14096 10532
rect 14148 10520 14154 10532
rect 14829 10523 14887 10529
rect 14829 10520 14841 10523
rect 14148 10492 14841 10520
rect 14148 10480 14154 10492
rect 14829 10489 14841 10492
rect 14875 10489 14887 10523
rect 15194 10520 15200 10532
rect 15155 10492 15200 10520
rect 14829 10483 14887 10489
rect 15194 10480 15200 10492
rect 15252 10480 15258 10532
rect 16025 10523 16083 10529
rect 16025 10489 16037 10523
rect 16071 10520 16083 10523
rect 16206 10520 16212 10532
rect 16071 10492 16212 10520
rect 16071 10489 16083 10492
rect 16025 10483 16083 10489
rect 16206 10480 16212 10492
rect 16264 10480 16270 10532
rect 16485 10523 16543 10529
rect 16485 10489 16497 10523
rect 16531 10520 16543 10523
rect 17696 10520 17724 10548
rect 16531 10492 17724 10520
rect 16531 10489 16543 10492
rect 16485 10483 16543 10489
rect 3752 10424 4108 10452
rect 3752 10412 3758 10424
rect 4522 10412 4528 10464
rect 4580 10452 4586 10464
rect 5810 10452 5816 10464
rect 4580 10424 5816 10452
rect 4580 10412 4586 10424
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 5902 10412 5908 10464
rect 5960 10452 5966 10464
rect 8202 10452 8208 10464
rect 5960 10424 8208 10452
rect 5960 10412 5966 10424
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 9950 10412 9956 10464
rect 10008 10452 10014 10464
rect 10045 10455 10103 10461
rect 10045 10452 10057 10455
rect 10008 10424 10057 10452
rect 10008 10412 10014 10424
rect 10045 10421 10057 10424
rect 10091 10421 10103 10455
rect 11514 10452 11520 10464
rect 11475 10424 11520 10452
rect 10045 10415 10103 10421
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 13078 10412 13084 10464
rect 13136 10452 13142 10464
rect 15013 10455 15071 10461
rect 15013 10452 15025 10455
rect 13136 10424 15025 10452
rect 13136 10412 13142 10424
rect 15013 10421 15025 10424
rect 15059 10421 15071 10455
rect 16298 10452 16304 10464
rect 16259 10424 16304 10452
rect 15013 10415 15071 10421
rect 16298 10412 16304 10424
rect 16356 10412 16362 10464
rect 17494 10412 17500 10464
rect 17552 10452 17558 10464
rect 17589 10455 17647 10461
rect 17589 10452 17601 10455
rect 17552 10424 17601 10452
rect 17552 10412 17558 10424
rect 17589 10421 17601 10424
rect 17635 10421 17647 10455
rect 17589 10415 17647 10421
rect 1104 10362 18860 10384
rect 1104 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 3430 10362
rect 3482 10310 7622 10362
rect 7674 10310 7686 10362
rect 7738 10310 7750 10362
rect 7802 10310 7814 10362
rect 7866 10310 7878 10362
rect 7930 10310 12070 10362
rect 12122 10310 12134 10362
rect 12186 10310 12198 10362
rect 12250 10310 12262 10362
rect 12314 10310 12326 10362
rect 12378 10310 16518 10362
rect 16570 10310 16582 10362
rect 16634 10310 16646 10362
rect 16698 10310 16710 10362
rect 16762 10310 16774 10362
rect 16826 10310 18860 10362
rect 1104 10288 18860 10310
rect 2038 10208 2044 10260
rect 2096 10208 2102 10260
rect 2777 10251 2835 10257
rect 2777 10217 2789 10251
rect 2823 10248 2835 10251
rect 2866 10248 2872 10260
rect 2823 10220 2872 10248
rect 2823 10217 2835 10220
rect 2777 10211 2835 10217
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 4522 10208 4528 10260
rect 4580 10248 4586 10260
rect 4617 10251 4675 10257
rect 4617 10248 4629 10251
rect 4580 10220 4629 10248
rect 4580 10208 4586 10220
rect 4617 10217 4629 10220
rect 4663 10217 4675 10251
rect 4617 10211 4675 10217
rect 4801 10251 4859 10257
rect 4801 10217 4813 10251
rect 4847 10248 4859 10251
rect 4982 10248 4988 10260
rect 4847 10220 4988 10248
rect 4847 10217 4859 10220
rect 4801 10211 4859 10217
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 8570 10248 8576 10260
rect 5184 10220 8576 10248
rect 2056 10180 2084 10208
rect 3970 10180 3976 10192
rect 2056 10152 3976 10180
rect 3970 10140 3976 10152
rect 4028 10140 4034 10192
rect 4433 10183 4491 10189
rect 4433 10149 4445 10183
rect 4479 10180 4491 10183
rect 5184 10180 5212 10220
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 10502 10248 10508 10260
rect 10463 10220 10508 10248
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 11330 10248 11336 10260
rect 11291 10220 11336 10248
rect 11330 10208 11336 10220
rect 11388 10208 11394 10260
rect 11974 10208 11980 10260
rect 12032 10248 12038 10260
rect 12161 10251 12219 10257
rect 12161 10248 12173 10251
rect 12032 10220 12173 10248
rect 12032 10208 12038 10220
rect 12161 10217 12173 10220
rect 12207 10217 12219 10251
rect 12161 10211 12219 10217
rect 15562 10208 15568 10260
rect 15620 10248 15626 10260
rect 17037 10251 17095 10257
rect 17037 10248 17049 10251
rect 15620 10220 17049 10248
rect 15620 10208 15626 10220
rect 17037 10217 17049 10220
rect 17083 10217 17095 10251
rect 17037 10211 17095 10217
rect 6457 10183 6515 10189
rect 6457 10180 6469 10183
rect 4479 10152 5212 10180
rect 5276 10152 5580 10180
rect 4479 10149 4491 10152
rect 4433 10143 4491 10149
rect 2041 10115 2099 10121
rect 2041 10081 2053 10115
rect 2087 10112 2099 10115
rect 2498 10112 2504 10124
rect 2087 10084 2504 10112
rect 2087 10081 2099 10084
rect 2041 10075 2099 10081
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 3421 10115 3479 10121
rect 3421 10081 3433 10115
rect 3467 10112 3479 10115
rect 3510 10112 3516 10124
rect 3467 10084 3516 10112
rect 3467 10081 3479 10084
rect 3421 10075 3479 10081
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 5276 10121 5304 10152
rect 5261 10115 5319 10121
rect 5261 10081 5273 10115
rect 5307 10081 5319 10115
rect 5442 10112 5448 10124
rect 5403 10084 5448 10112
rect 5261 10075 5319 10081
rect 5442 10072 5448 10084
rect 5500 10072 5506 10124
rect 5552 10112 5580 10152
rect 5828 10152 6469 10180
rect 5828 10112 5856 10152
rect 6457 10149 6469 10152
rect 6503 10149 6515 10183
rect 6457 10143 6515 10149
rect 6730 10140 6736 10192
rect 6788 10180 6794 10192
rect 6788 10152 7052 10180
rect 6788 10140 6794 10152
rect 5552 10084 5856 10112
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10081 6239 10115
rect 6181 10075 6239 10081
rect 1486 10044 1492 10056
rect 1447 10016 1492 10044
rect 1486 10004 1492 10016
rect 1544 10004 1550 10056
rect 1854 10044 1860 10056
rect 1815 10016 1860 10044
rect 1854 10004 1860 10016
rect 1912 10004 1918 10056
rect 2314 10044 2320 10056
rect 2275 10016 2320 10044
rect 2314 10004 2320 10016
rect 2372 10004 2378 10056
rect 2406 10004 2412 10056
rect 2464 10044 2470 10056
rect 3145 10047 3203 10053
rect 2464 10016 2509 10044
rect 2464 10004 2470 10016
rect 3145 10013 3157 10047
rect 3191 10044 3203 10047
rect 3694 10044 3700 10056
rect 3191 10016 3700 10044
rect 3191 10013 3203 10016
rect 3145 10007 3203 10013
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 4065 10047 4123 10053
rect 4065 10013 4077 10047
rect 4111 10044 4123 10047
rect 4111 10040 5580 10044
rect 4111 10016 5764 10040
rect 4111 10013 4123 10016
rect 4065 10007 4123 10013
rect 5552 10012 5764 10016
rect 1673 9979 1731 9985
rect 1673 9945 1685 9979
rect 1719 9976 1731 9979
rect 2222 9976 2228 9988
rect 1719 9948 2228 9976
rect 1719 9945 1731 9948
rect 1673 9939 1731 9945
rect 2222 9936 2228 9948
rect 2280 9936 2286 9988
rect 3786 9976 3792 9988
rect 2608 9948 3792 9976
rect 2038 9868 2044 9920
rect 2096 9908 2102 9920
rect 2608 9917 2636 9948
rect 3786 9936 3792 9948
rect 3844 9976 3850 9988
rect 3881 9979 3939 9985
rect 3881 9976 3893 9979
rect 3844 9948 3893 9976
rect 3844 9936 3850 9948
rect 3881 9945 3893 9948
rect 3927 9945 3939 9979
rect 3881 9939 3939 9945
rect 4249 9979 4307 9985
rect 4249 9945 4261 9979
rect 4295 9976 4307 9979
rect 4522 9976 4528 9988
rect 4295 9948 4528 9976
rect 4295 9945 4307 9948
rect 4249 9939 4307 9945
rect 4522 9936 4528 9948
rect 4580 9936 4586 9988
rect 5169 9979 5227 9985
rect 5169 9945 5181 9979
rect 5215 9976 5227 9979
rect 5736 9976 5764 10012
rect 5810 10004 5816 10056
rect 5868 10044 5874 10056
rect 5994 10044 6000 10056
rect 5868 10016 6000 10044
rect 5868 10004 5874 10016
rect 5994 10004 6000 10016
rect 6052 10004 6058 10056
rect 6196 10044 6224 10075
rect 6270 10072 6276 10124
rect 6328 10112 6334 10124
rect 7024 10121 7052 10152
rect 8478 10140 8484 10192
rect 8536 10180 8542 10192
rect 9585 10183 9643 10189
rect 9585 10180 9597 10183
rect 8536 10152 9597 10180
rect 8536 10140 8542 10152
rect 9585 10149 9597 10152
rect 9631 10149 9643 10183
rect 9585 10143 9643 10149
rect 10686 10140 10692 10192
rect 10744 10180 10750 10192
rect 13538 10180 13544 10192
rect 10744 10152 13544 10180
rect 10744 10140 10750 10152
rect 13538 10140 13544 10152
rect 13596 10140 13602 10192
rect 16942 10140 16948 10192
rect 17000 10180 17006 10192
rect 17000 10152 17632 10180
rect 17000 10140 17006 10152
rect 6917 10115 6975 10121
rect 6917 10112 6929 10115
rect 6328 10084 6929 10112
rect 6328 10072 6334 10084
rect 6917 10081 6929 10084
rect 6963 10081 6975 10115
rect 6917 10075 6975 10081
rect 7009 10115 7067 10121
rect 7009 10081 7021 10115
rect 7055 10081 7067 10115
rect 7009 10075 7067 10081
rect 9030 10072 9036 10124
rect 9088 10112 9094 10124
rect 10137 10115 10195 10121
rect 10137 10112 10149 10115
rect 9088 10084 10149 10112
rect 9088 10072 9094 10084
rect 10137 10081 10149 10084
rect 10183 10081 10195 10115
rect 10137 10075 10195 10081
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 10962 10112 10968 10124
rect 10468 10084 10968 10112
rect 10468 10072 10474 10084
rect 10962 10072 10968 10084
rect 11020 10072 11026 10124
rect 11149 10115 11207 10121
rect 11149 10081 11161 10115
rect 11195 10112 11207 10115
rect 11885 10115 11943 10121
rect 11885 10112 11897 10115
rect 11195 10084 11897 10112
rect 11195 10081 11207 10084
rect 11149 10075 11207 10081
rect 11885 10081 11897 10084
rect 11931 10112 11943 10115
rect 12713 10115 12771 10121
rect 12713 10112 12725 10115
rect 11931 10084 12725 10112
rect 11931 10081 11943 10084
rect 11885 10075 11943 10081
rect 12713 10081 12725 10084
rect 12759 10112 12771 10115
rect 12894 10112 12900 10124
rect 12759 10084 12900 10112
rect 12759 10081 12771 10084
rect 12713 10075 12771 10081
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 12989 10115 13047 10121
rect 12989 10081 13001 10115
rect 13035 10112 13047 10115
rect 13630 10112 13636 10124
rect 13035 10084 13636 10112
rect 13035 10081 13047 10084
rect 12989 10075 13047 10081
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 17494 10112 17500 10124
rect 17455 10084 17500 10112
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 17604 10121 17632 10152
rect 17589 10115 17647 10121
rect 17589 10081 17601 10115
rect 17635 10081 17647 10115
rect 17589 10075 17647 10081
rect 6730 10044 6736 10056
rect 6196 10016 6736 10044
rect 6730 10004 6736 10016
rect 6788 10004 6794 10056
rect 6822 10004 6828 10056
rect 6880 10044 6886 10056
rect 7377 10047 7435 10053
rect 7377 10044 7389 10047
rect 6880 10016 7389 10044
rect 6880 10004 6886 10016
rect 7377 10013 7389 10016
rect 7423 10013 7435 10047
rect 7377 10007 7435 10013
rect 7644 10047 7702 10053
rect 7644 10013 7656 10047
rect 7690 10044 7702 10047
rect 8110 10044 8116 10056
rect 7690 10016 8116 10044
rect 7690 10013 7702 10016
rect 7644 10007 7702 10013
rect 8110 10004 8116 10016
rect 8168 10004 8174 10056
rect 9950 10044 9956 10056
rect 9911 10016 9956 10044
rect 9950 10004 9956 10016
rect 10008 10004 10014 10056
rect 10045 10047 10103 10053
rect 10045 10013 10057 10047
rect 10091 10044 10103 10047
rect 11514 10044 11520 10056
rect 10091 10016 11520 10044
rect 10091 10013 10103 10016
rect 10045 10007 10103 10013
rect 11514 10004 11520 10016
rect 11572 10004 11578 10056
rect 11698 10044 11704 10056
rect 11659 10016 11704 10044
rect 11698 10004 11704 10016
rect 11756 10004 11762 10056
rect 12529 10047 12587 10053
rect 12529 10013 12541 10047
rect 12575 10044 12587 10047
rect 12802 10044 12808 10056
rect 12575 10016 12808 10044
rect 12575 10013 12587 10016
rect 12529 10007 12587 10013
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 9674 9976 9680 9988
rect 5215 9948 5672 9976
rect 5736 9948 9680 9976
rect 5215 9945 5227 9948
rect 5169 9939 5227 9945
rect 2133 9911 2191 9917
rect 2133 9908 2145 9911
rect 2096 9880 2145 9908
rect 2096 9868 2102 9880
rect 2133 9877 2145 9880
rect 2179 9877 2191 9911
rect 2133 9871 2191 9877
rect 2593 9911 2651 9917
rect 2593 9877 2605 9911
rect 2639 9877 2651 9911
rect 2593 9871 2651 9877
rect 3237 9911 3295 9917
rect 3237 9877 3249 9911
rect 3283 9908 3295 9911
rect 3694 9908 3700 9920
rect 3283 9880 3700 9908
rect 3283 9877 3295 9880
rect 3237 9871 3295 9877
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 5644 9917 5672 9948
rect 9674 9936 9680 9948
rect 9732 9936 9738 9988
rect 10226 9936 10232 9988
rect 10284 9976 10290 9988
rect 10873 9979 10931 9985
rect 10873 9976 10885 9979
rect 10284 9948 10885 9976
rect 10284 9936 10290 9948
rect 10873 9945 10885 9948
rect 10919 9945 10931 9979
rect 10873 9939 10931 9945
rect 11606 9936 11612 9988
rect 11664 9976 11670 9988
rect 11793 9979 11851 9985
rect 11793 9976 11805 9979
rect 11664 9948 11805 9976
rect 11664 9936 11670 9948
rect 11793 9945 11805 9948
rect 11839 9945 11851 9979
rect 13280 9976 13308 10007
rect 14182 10004 14188 10056
rect 14240 10044 14246 10056
rect 15473 10047 15531 10053
rect 15473 10044 15485 10047
rect 14240 10016 15485 10044
rect 14240 10004 14246 10016
rect 15473 10013 15485 10016
rect 15519 10044 15531 10047
rect 15565 10047 15623 10053
rect 15565 10044 15577 10047
rect 15519 10016 15577 10044
rect 15519 10013 15531 10016
rect 15473 10007 15531 10013
rect 15565 10013 15577 10016
rect 15611 10013 15623 10047
rect 15565 10007 15623 10013
rect 15832 10047 15890 10053
rect 15832 10013 15844 10047
rect 15878 10044 15890 10047
rect 16114 10044 16120 10056
rect 15878 10016 16120 10044
rect 15878 10013 15890 10016
rect 15832 10007 15890 10013
rect 16114 10004 16120 10016
rect 16172 10004 16178 10056
rect 16298 10004 16304 10056
rect 16356 10044 16362 10056
rect 18414 10044 18420 10056
rect 16356 10016 18420 10044
rect 16356 10004 16362 10016
rect 18414 10004 18420 10016
rect 18472 10004 18478 10056
rect 11793 9939 11851 9945
rect 12406 9948 13308 9976
rect 15228 9979 15286 9985
rect 5629 9911 5687 9917
rect 5629 9877 5641 9911
rect 5675 9877 5687 9911
rect 5629 9871 5687 9877
rect 6086 9868 6092 9920
rect 6144 9908 6150 9920
rect 6825 9911 6883 9917
rect 6144 9880 6189 9908
rect 6144 9868 6150 9880
rect 6825 9877 6837 9911
rect 6871 9908 6883 9911
rect 7190 9908 7196 9920
rect 6871 9880 7196 9908
rect 6871 9877 6883 9880
rect 6825 9871 6883 9877
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 8662 9868 8668 9920
rect 8720 9908 8726 9920
rect 8757 9911 8815 9917
rect 8757 9908 8769 9911
rect 8720 9880 8769 9908
rect 8720 9868 8726 9880
rect 8757 9877 8769 9880
rect 8803 9877 8815 9911
rect 8757 9871 8815 9877
rect 10410 9868 10416 9920
rect 10468 9908 10474 9920
rect 12406 9908 12434 9948
rect 15228 9945 15240 9979
rect 15274 9976 15286 9979
rect 18230 9976 18236 9988
rect 15274 9948 15792 9976
rect 18191 9948 18236 9976
rect 15274 9945 15286 9948
rect 15228 9939 15286 9945
rect 10468 9880 12434 9908
rect 10468 9868 10474 9880
rect 12618 9868 12624 9920
rect 12676 9908 12682 9920
rect 12676 9880 12721 9908
rect 12676 9868 12682 9880
rect 13446 9868 13452 9920
rect 13504 9908 13510 9920
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 13504 9880 14105 9908
rect 13504 9868 13510 9880
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 15764 9908 15792 9948
rect 18230 9936 18236 9948
rect 18288 9936 18294 9988
rect 16298 9908 16304 9920
rect 15764 9880 16304 9908
rect 14093 9871 14151 9877
rect 16298 9868 16304 9880
rect 16356 9868 16362 9920
rect 16942 9908 16948 9920
rect 16903 9880 16948 9908
rect 16942 9868 16948 9880
rect 17000 9868 17006 9920
rect 17402 9908 17408 9920
rect 17363 9880 17408 9908
rect 17402 9868 17408 9880
rect 17460 9868 17466 9920
rect 17678 9868 17684 9920
rect 17736 9908 17742 9920
rect 17865 9911 17923 9917
rect 17865 9908 17877 9911
rect 17736 9880 17877 9908
rect 17736 9868 17742 9880
rect 17865 9877 17877 9880
rect 17911 9877 17923 9911
rect 17865 9871 17923 9877
rect 1104 9818 18860 9840
rect 1104 9766 5398 9818
rect 5450 9766 5462 9818
rect 5514 9766 5526 9818
rect 5578 9766 5590 9818
rect 5642 9766 5654 9818
rect 5706 9766 9846 9818
rect 9898 9766 9910 9818
rect 9962 9766 9974 9818
rect 10026 9766 10038 9818
rect 10090 9766 10102 9818
rect 10154 9766 14294 9818
rect 14346 9766 14358 9818
rect 14410 9766 14422 9818
rect 14474 9766 14486 9818
rect 14538 9766 14550 9818
rect 14602 9766 18860 9818
rect 1104 9744 18860 9766
rect 3878 9704 3884 9716
rect 2746 9676 3884 9704
rect 2746 9636 2774 9676
rect 3878 9664 3884 9676
rect 3936 9664 3942 9716
rect 5810 9704 5816 9716
rect 5771 9676 5816 9704
rect 5810 9664 5816 9676
rect 5868 9664 5874 9716
rect 6086 9664 6092 9716
rect 6144 9704 6150 9716
rect 6365 9707 6423 9713
rect 6365 9704 6377 9707
rect 6144 9676 6377 9704
rect 6144 9664 6150 9676
rect 6365 9673 6377 9676
rect 6411 9673 6423 9707
rect 6733 9707 6791 9713
rect 6733 9704 6745 9707
rect 6365 9667 6423 9673
rect 6656 9676 6745 9704
rect 1780 9608 2774 9636
rect 4433 9639 4491 9645
rect 1489 9571 1547 9577
rect 1489 9537 1501 9571
rect 1535 9537 1547 9571
rect 1489 9531 1547 9537
rect 1302 9392 1308 9444
rect 1360 9432 1366 9444
rect 1504 9432 1532 9531
rect 1780 9512 1808 9608
rect 4433 9605 4445 9639
rect 4479 9636 4491 9639
rect 4614 9636 4620 9648
rect 4479 9608 4620 9636
rect 4479 9605 4491 9608
rect 4433 9599 4491 9605
rect 4614 9596 4620 9608
rect 4672 9636 4678 9648
rect 5442 9636 5448 9648
rect 4672 9608 5448 9636
rect 4672 9596 4678 9608
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 6546 9596 6552 9648
rect 6604 9636 6610 9648
rect 6656 9636 6684 9676
rect 6733 9673 6745 9676
rect 6779 9704 6791 9707
rect 12529 9707 12587 9713
rect 6779 9676 6868 9704
rect 6779 9673 6791 9676
rect 6733 9667 6791 9673
rect 6604 9608 6684 9636
rect 6840 9636 6868 9676
rect 12529 9673 12541 9707
rect 12575 9704 12587 9707
rect 12710 9704 12716 9716
rect 12575 9676 12716 9704
rect 12575 9673 12587 9676
rect 12529 9667 12587 9673
rect 12710 9664 12716 9676
rect 12768 9664 12774 9716
rect 12802 9664 12808 9716
rect 12860 9704 12866 9716
rect 12897 9707 12955 9713
rect 12897 9704 12909 9707
rect 12860 9676 12909 9704
rect 12860 9664 12866 9676
rect 12897 9673 12909 9676
rect 12943 9673 12955 9707
rect 12897 9667 12955 9673
rect 15565 9707 15623 9713
rect 15565 9673 15577 9707
rect 15611 9704 15623 9707
rect 15746 9704 15752 9716
rect 15611 9676 15752 9704
rect 15611 9673 15623 9676
rect 15565 9667 15623 9673
rect 7006 9636 7012 9648
rect 6840 9608 7012 9636
rect 6604 9596 6610 9608
rect 7006 9596 7012 9608
rect 7064 9636 7070 9648
rect 7193 9639 7251 9645
rect 7193 9636 7205 9639
rect 7064 9608 7205 9636
rect 7064 9596 7070 9608
rect 7193 9605 7205 9608
rect 7239 9605 7251 9639
rect 7193 9599 7251 9605
rect 8662 9596 8668 9648
rect 8720 9645 8726 9648
rect 8720 9636 8732 9645
rect 9582 9636 9588 9648
rect 8720 9608 9588 9636
rect 8720 9599 8732 9608
rect 8720 9596 8726 9599
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 10226 9596 10232 9648
rect 10284 9636 10290 9648
rect 10321 9639 10379 9645
rect 10321 9636 10333 9639
rect 10284 9608 10333 9636
rect 10284 9596 10290 9608
rect 10321 9605 10333 9608
rect 10367 9605 10379 9639
rect 10321 9599 10379 9605
rect 2032 9571 2090 9577
rect 2032 9537 2044 9571
rect 2078 9568 2090 9571
rect 2314 9568 2320 9580
rect 2078 9540 2320 9568
rect 2078 9537 2090 9540
rect 2032 9531 2090 9537
rect 2314 9528 2320 9540
rect 2372 9528 2378 9580
rect 2866 9528 2872 9580
rect 2924 9568 2930 9580
rect 3602 9568 3608 9580
rect 2924 9540 3608 9568
rect 2924 9528 2930 9540
rect 3602 9528 3608 9540
rect 3660 9528 3666 9580
rect 4522 9528 4528 9580
rect 4580 9568 4586 9580
rect 4982 9568 4988 9580
rect 4580 9540 4988 9568
rect 4580 9528 4586 9540
rect 4982 9528 4988 9540
rect 5040 9528 5046 9580
rect 5077 9571 5135 9577
rect 5077 9537 5089 9571
rect 5123 9537 5135 9571
rect 5077 9531 5135 9537
rect 1762 9500 1768 9512
rect 1723 9472 1768 9500
rect 1762 9460 1768 9472
rect 1820 9460 1826 9512
rect 2958 9460 2964 9512
rect 3016 9500 3022 9512
rect 3697 9503 3755 9509
rect 3016 9472 3556 9500
rect 3016 9460 3022 9472
rect 1360 9404 1716 9432
rect 1360 9392 1366 9404
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 1688 9364 1716 9404
rect 3050 9392 3056 9444
rect 3108 9432 3114 9444
rect 3237 9435 3295 9441
rect 3237 9432 3249 9435
rect 3108 9404 3249 9432
rect 3108 9392 3114 9404
rect 3237 9401 3249 9404
rect 3283 9401 3295 9435
rect 3528 9432 3556 9472
rect 3697 9469 3709 9503
rect 3743 9500 3755 9503
rect 3786 9500 3792 9512
rect 3743 9472 3792 9500
rect 3743 9469 3755 9472
rect 3697 9463 3755 9469
rect 3786 9460 3792 9472
rect 3844 9460 3850 9512
rect 3881 9503 3939 9509
rect 3881 9469 3893 9503
rect 3927 9500 3939 9503
rect 4617 9503 4675 9509
rect 3927 9472 4200 9500
rect 3927 9469 3939 9472
rect 3881 9463 3939 9469
rect 4065 9435 4123 9441
rect 4065 9432 4077 9435
rect 3528 9404 4077 9432
rect 3237 9395 3295 9401
rect 4065 9401 4077 9404
rect 4111 9401 4123 9435
rect 4065 9395 4123 9401
rect 4172 9432 4200 9472
rect 4617 9469 4629 9503
rect 4663 9469 4675 9503
rect 5092 9500 5120 9531
rect 5166 9528 5172 9580
rect 5224 9568 5230 9580
rect 5261 9571 5319 9577
rect 5261 9568 5273 9571
rect 5224 9540 5273 9568
rect 5224 9528 5230 9540
rect 5261 9537 5273 9540
rect 5307 9568 5319 9571
rect 6822 9568 6828 9580
rect 5307 9540 6828 9568
rect 5307 9537 5319 9540
rect 5261 9531 5319 9537
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 7469 9571 7527 9577
rect 7469 9537 7481 9571
rect 7515 9568 7527 9571
rect 11974 9568 11980 9580
rect 7515 9540 11980 9568
rect 7515 9537 7527 9540
rect 7469 9531 7527 9537
rect 5350 9500 5356 9512
rect 5092 9472 5356 9500
rect 4617 9463 4675 9469
rect 4632 9432 4660 9463
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 5629 9503 5687 9509
rect 5629 9469 5641 9503
rect 5675 9469 5687 9503
rect 5629 9463 5687 9469
rect 5721 9503 5779 9509
rect 5721 9469 5733 9503
rect 5767 9469 5779 9503
rect 5721 9463 5779 9469
rect 4172 9404 4660 9432
rect 2958 9364 2964 9376
rect 1688 9336 2964 9364
rect 2958 9324 2964 9336
rect 3016 9324 3022 9376
rect 3145 9367 3203 9373
rect 3145 9333 3157 9367
rect 3191 9364 3203 9367
rect 3510 9364 3516 9376
rect 3191 9336 3516 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 3510 9324 3516 9336
rect 3568 9364 3574 9376
rect 4172 9364 4200 9404
rect 3568 9336 4200 9364
rect 3568 9324 3574 9336
rect 4798 9324 4804 9376
rect 4856 9364 4862 9376
rect 4893 9367 4951 9373
rect 4893 9364 4905 9367
rect 4856 9336 4905 9364
rect 4856 9324 4862 9336
rect 4893 9333 4905 9336
rect 4939 9333 4951 9367
rect 5644 9364 5672 9463
rect 5736 9432 5764 9463
rect 5810 9460 5816 9512
rect 5868 9500 5874 9512
rect 6730 9500 6736 9512
rect 5868 9472 6736 9500
rect 5868 9460 5874 9472
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 7009 9503 7067 9509
rect 7009 9469 7021 9503
rect 7055 9469 7067 9503
rect 7009 9463 7067 9469
rect 5994 9432 6000 9444
rect 5736 9404 6000 9432
rect 5994 9392 6000 9404
rect 6052 9392 6058 9444
rect 6181 9435 6239 9441
rect 6181 9401 6193 9435
rect 6227 9432 6239 9435
rect 6270 9432 6276 9444
rect 6227 9404 6276 9432
rect 6227 9401 6239 9404
rect 6181 9395 6239 9401
rect 6270 9392 6276 9404
rect 6328 9392 6334 9444
rect 7024 9432 7052 9463
rect 6472 9404 7052 9432
rect 6472 9376 6500 9404
rect 6454 9364 6460 9376
rect 5644 9336 6460 9364
rect 4893 9327 4951 9333
rect 6454 9324 6460 9336
rect 6512 9324 6518 9376
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 7484 9364 7512 9531
rect 11974 9528 11980 9540
rect 12032 9528 12038 9580
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 13630 9568 13636 9580
rect 12768 9540 13636 9568
rect 12768 9528 12774 9540
rect 13630 9528 13636 9540
rect 13688 9528 13694 9580
rect 14182 9568 14188 9580
rect 14143 9540 14188 9568
rect 14182 9528 14188 9540
rect 14240 9528 14246 9580
rect 15672 9577 15700 9676
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 16298 9704 16304 9716
rect 16259 9676 16304 9704
rect 16298 9664 16304 9676
rect 16356 9664 16362 9716
rect 16669 9707 16727 9713
rect 16669 9673 16681 9707
rect 16715 9704 16727 9707
rect 16850 9704 16856 9716
rect 16715 9676 16856 9704
rect 16715 9673 16727 9676
rect 16669 9667 16727 9673
rect 16850 9664 16856 9676
rect 16908 9664 16914 9716
rect 16868 9608 18000 9636
rect 16868 9580 16896 9608
rect 14452 9571 14510 9577
rect 14452 9537 14464 9571
rect 14498 9568 14510 9571
rect 15657 9571 15715 9577
rect 14498 9540 15608 9568
rect 14498 9537 14510 9540
rect 14452 9531 14510 9537
rect 8938 9500 8944 9512
rect 8899 9472 8944 9500
rect 8938 9460 8944 9472
rect 8996 9460 9002 9512
rect 10962 9460 10968 9512
rect 11020 9500 11026 9512
rect 11517 9503 11575 9509
rect 11517 9500 11529 9503
rect 11020 9472 11529 9500
rect 11020 9460 11026 9472
rect 11517 9469 11529 9472
rect 11563 9469 11575 9503
rect 11517 9463 11575 9469
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9469 12311 9503
rect 12253 9463 12311 9469
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9500 12495 9503
rect 12986 9500 12992 9512
rect 12483 9472 12848 9500
rect 12947 9472 12992 9500
rect 12483 9469 12495 9472
rect 12437 9463 12495 9469
rect 9674 9392 9680 9444
rect 9732 9432 9738 9444
rect 11146 9432 11152 9444
rect 9732 9404 11152 9432
rect 9732 9392 9738 9404
rect 11146 9392 11152 9404
rect 11204 9392 11210 9444
rect 12268 9432 12296 9463
rect 12710 9432 12716 9444
rect 12268 9404 12716 9432
rect 12710 9392 12716 9404
rect 12768 9392 12774 9444
rect 12820 9376 12848 9472
rect 12986 9460 12992 9472
rect 13044 9460 13050 9512
rect 13262 9500 13268 9512
rect 13223 9472 13268 9500
rect 13262 9460 13268 9472
rect 13320 9460 13326 9512
rect 15580 9500 15608 9540
rect 15657 9537 15669 9571
rect 15703 9537 15715 9571
rect 15657 9531 15715 9537
rect 16850 9528 16856 9580
rect 16908 9528 16914 9580
rect 17034 9568 17040 9580
rect 16995 9540 17040 9568
rect 17034 9528 17040 9540
rect 17092 9528 17098 9580
rect 17972 9577 18000 9608
rect 17957 9571 18015 9577
rect 17957 9537 17969 9571
rect 18003 9537 18015 9571
rect 17957 9531 18015 9537
rect 16942 9500 16948 9512
rect 15580 9472 16948 9500
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17126 9500 17132 9512
rect 17087 9472 17132 9500
rect 17126 9460 17132 9472
rect 17184 9460 17190 9512
rect 17221 9503 17279 9509
rect 17221 9469 17233 9503
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 17681 9503 17739 9509
rect 17681 9469 17693 9503
rect 17727 9500 17739 9503
rect 17770 9500 17776 9512
rect 17727 9472 17776 9500
rect 17727 9469 17739 9472
rect 17681 9463 17739 9469
rect 12894 9392 12900 9444
rect 12952 9432 12958 9444
rect 13446 9432 13452 9444
rect 12952 9404 13452 9432
rect 12952 9392 12958 9404
rect 13446 9392 13452 9404
rect 13504 9392 13510 9444
rect 13630 9392 13636 9444
rect 13688 9432 13694 9444
rect 16960 9432 16988 9460
rect 17236 9432 17264 9463
rect 17770 9460 17776 9472
rect 17828 9460 17834 9512
rect 18322 9432 18328 9444
rect 13688 9404 14044 9432
rect 13688 9392 13694 9404
rect 6788 9336 7512 9364
rect 7561 9367 7619 9373
rect 6788 9324 6794 9336
rect 7561 9333 7573 9367
rect 7607 9364 7619 9367
rect 8662 9364 8668 9376
rect 7607 9336 8668 9364
rect 7607 9333 7619 9336
rect 7561 9327 7619 9333
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 8754 9324 8760 9376
rect 8812 9364 8818 9376
rect 10226 9364 10232 9376
rect 8812 9336 10232 9364
rect 8812 9324 8818 9336
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 10778 9324 10784 9376
rect 10836 9364 10842 9376
rect 12434 9364 12440 9376
rect 10836 9336 12440 9364
rect 10836 9324 10842 9336
rect 12434 9324 12440 9336
rect 12492 9324 12498 9376
rect 12802 9324 12808 9376
rect 12860 9324 12866 9376
rect 13906 9364 13912 9376
rect 13867 9336 13912 9364
rect 13906 9324 13912 9336
rect 13964 9324 13970 9376
rect 14016 9364 14044 9404
rect 15120 9404 16528 9432
rect 16960 9404 17264 9432
rect 17328 9404 18328 9432
rect 15120 9364 15148 9404
rect 14016 9336 15148 9364
rect 15562 9324 15568 9376
rect 15620 9364 15626 9376
rect 15930 9364 15936 9376
rect 15620 9336 15936 9364
rect 15620 9324 15626 9336
rect 15930 9324 15936 9336
rect 15988 9364 15994 9376
rect 16393 9367 16451 9373
rect 16393 9364 16405 9367
rect 15988 9336 16405 9364
rect 15988 9324 15994 9336
rect 16393 9333 16405 9336
rect 16439 9333 16451 9367
rect 16500 9364 16528 9404
rect 17328 9364 17356 9404
rect 18322 9392 18328 9404
rect 18380 9392 18386 9444
rect 17586 9364 17592 9376
rect 16500 9336 17356 9364
rect 17547 9336 17592 9364
rect 16393 9327 16451 9333
rect 17586 9324 17592 9336
rect 17644 9324 17650 9376
rect 1104 9274 18860 9296
rect 1104 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 3430 9274
rect 3482 9222 7622 9274
rect 7674 9222 7686 9274
rect 7738 9222 7750 9274
rect 7802 9222 7814 9274
rect 7866 9222 7878 9274
rect 7930 9222 12070 9274
rect 12122 9222 12134 9274
rect 12186 9222 12198 9274
rect 12250 9222 12262 9274
rect 12314 9222 12326 9274
rect 12378 9222 16518 9274
rect 16570 9222 16582 9274
rect 16634 9222 16646 9274
rect 16698 9222 16710 9274
rect 16762 9222 16774 9274
rect 16826 9222 18860 9274
rect 1104 9200 18860 9222
rect 1489 9163 1547 9169
rect 1489 9129 1501 9163
rect 1535 9160 1547 9163
rect 1854 9160 1860 9172
rect 1535 9132 1860 9160
rect 1535 9129 1547 9132
rect 1489 9123 1547 9129
rect 1854 9120 1860 9132
rect 1912 9120 1918 9172
rect 2682 9120 2688 9172
rect 2740 9160 2746 9172
rect 3602 9160 3608 9172
rect 2740 9132 3608 9160
rect 2740 9120 2746 9132
rect 3602 9120 3608 9132
rect 3660 9120 3666 9172
rect 4522 9160 4528 9172
rect 4264 9132 4528 9160
rect 3237 9095 3295 9101
rect 3237 9061 3249 9095
rect 3283 9092 3295 9095
rect 4264 9092 4292 9132
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 8478 9160 8484 9172
rect 5408 9132 8484 9160
rect 5408 9120 5414 9132
rect 8478 9120 8484 9132
rect 8536 9120 8542 9172
rect 8570 9120 8576 9172
rect 8628 9160 8634 9172
rect 9033 9163 9091 9169
rect 9033 9160 9045 9163
rect 8628 9132 9045 9160
rect 8628 9120 8634 9132
rect 9033 9129 9045 9132
rect 9079 9160 9091 9163
rect 9490 9160 9496 9172
rect 9079 9132 9496 9160
rect 9079 9129 9091 9132
rect 9033 9123 9091 9129
rect 9490 9120 9496 9132
rect 9548 9160 9554 9172
rect 12526 9160 12532 9172
rect 9548 9132 12532 9160
rect 9548 9120 9554 9132
rect 12526 9120 12532 9132
rect 12584 9120 12590 9172
rect 12618 9120 12624 9172
rect 12676 9160 12682 9172
rect 12897 9163 12955 9169
rect 12897 9160 12909 9163
rect 12676 9132 12909 9160
rect 12676 9120 12682 9132
rect 12897 9129 12909 9132
rect 12943 9129 12955 9163
rect 12897 9123 12955 9129
rect 13722 9120 13728 9172
rect 13780 9160 13786 9172
rect 14277 9163 14335 9169
rect 14277 9160 14289 9163
rect 13780 9132 14289 9160
rect 13780 9120 13786 9132
rect 14277 9129 14289 9132
rect 14323 9160 14335 9163
rect 15286 9160 15292 9172
rect 14323 9132 15292 9160
rect 14323 9129 14335 9132
rect 14277 9123 14335 9129
rect 15286 9120 15292 9132
rect 15344 9160 15350 9172
rect 15933 9163 15991 9169
rect 15344 9132 15893 9160
rect 15344 9120 15350 9132
rect 3283 9064 4292 9092
rect 3283 9061 3295 9064
rect 3237 9055 3295 9061
rect 5994 9052 6000 9104
rect 6052 9092 6058 9104
rect 11514 9092 11520 9104
rect 6052 9064 9168 9092
rect 6052 9052 6058 9064
rect 2961 9027 3019 9033
rect 2961 8993 2973 9027
rect 3007 9024 3019 9027
rect 3007 8996 4108 9024
rect 3007 8993 3019 8996
rect 2961 8987 3019 8993
rect 1578 8916 1584 8968
rect 1636 8916 1642 8968
rect 1762 8916 1768 8968
rect 1820 8956 1826 8968
rect 2976 8956 3004 8987
rect 1820 8928 3004 8956
rect 1820 8916 1826 8928
rect 3050 8916 3056 8968
rect 3108 8956 3114 8968
rect 3513 8959 3571 8965
rect 3513 8956 3525 8959
rect 3108 8928 3525 8956
rect 3108 8916 3114 8928
rect 3513 8925 3525 8928
rect 3559 8925 3571 8959
rect 4080 8956 4108 8996
rect 5442 8984 5448 9036
rect 5500 9024 5506 9036
rect 8570 9024 8576 9036
rect 5500 8996 8156 9024
rect 8531 8996 8576 9024
rect 5500 8984 5506 8996
rect 5169 8959 5227 8965
rect 5169 8956 5181 8959
rect 4080 8928 5181 8956
rect 3513 8919 3571 8925
rect 5169 8925 5181 8928
rect 5215 8956 5227 8959
rect 5261 8959 5319 8965
rect 5261 8956 5273 8959
rect 5215 8928 5273 8956
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5261 8925 5273 8928
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 8018 8916 8024 8968
rect 8076 8916 8082 8968
rect 1596 8888 1624 8916
rect 1596 8860 2636 8888
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 2608 8820 2636 8860
rect 2682 8848 2688 8900
rect 2740 8897 2746 8900
rect 2740 8888 2752 8897
rect 3418 8888 3424 8900
rect 2740 8860 2785 8888
rect 3379 8860 3424 8888
rect 2740 8851 2752 8860
rect 2740 8848 2746 8851
rect 3418 8848 3424 8860
rect 3476 8848 3482 8900
rect 3712 8860 4660 8888
rect 3712 8820 3740 8860
rect 2608 8792 3740 8820
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8820 3847 8823
rect 3878 8820 3884 8832
rect 3835 8792 3884 8820
rect 3835 8789 3847 8792
rect 3789 8783 3847 8789
rect 3878 8780 3884 8792
rect 3936 8820 3942 8832
rect 4522 8820 4528 8832
rect 3936 8792 4528 8820
rect 3936 8780 3942 8792
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 4632 8820 4660 8860
rect 4890 8848 4896 8900
rect 4948 8897 4954 8900
rect 4948 8888 4960 8897
rect 7009 8891 7067 8897
rect 4948 8860 4993 8888
rect 4948 8851 4960 8860
rect 7009 8857 7021 8891
rect 7055 8888 7067 8891
rect 7098 8888 7104 8900
rect 7055 8860 7104 8888
rect 7055 8857 7067 8860
rect 7009 8851 7067 8857
rect 4948 8848 4954 8851
rect 7098 8848 7104 8860
rect 7156 8848 7162 8900
rect 7558 8848 7564 8900
rect 7616 8888 7622 8900
rect 8036 8888 8064 8916
rect 7616 8860 8064 8888
rect 7616 8848 7622 8860
rect 5994 8820 6000 8832
rect 4632 8792 6000 8820
rect 5994 8780 6000 8792
rect 6052 8780 6058 8832
rect 7466 8780 7472 8832
rect 7524 8820 7530 8832
rect 8021 8823 8079 8829
rect 8021 8820 8033 8823
rect 7524 8792 8033 8820
rect 7524 8780 7530 8792
rect 8021 8789 8033 8792
rect 8067 8789 8079 8823
rect 8128 8820 8156 8996
rect 8570 8984 8576 8996
rect 8628 8984 8634 9036
rect 9140 9024 9168 9064
rect 9508 9064 11520 9092
rect 9508 9024 9536 9064
rect 11514 9052 11520 9064
rect 11572 9052 11578 9104
rect 12802 9052 12808 9104
rect 12860 9092 12866 9104
rect 13906 9092 13912 9104
rect 12860 9064 13912 9092
rect 12860 9052 12866 9064
rect 13906 9052 13912 9064
rect 13964 9052 13970 9104
rect 15865 9092 15893 9132
rect 15933 9129 15945 9163
rect 15979 9160 15991 9163
rect 16114 9160 16120 9172
rect 15979 9132 16120 9160
rect 15979 9129 15991 9132
rect 15933 9123 15991 9129
rect 16114 9120 16120 9132
rect 16172 9120 16178 9172
rect 16850 9160 16856 9172
rect 16500 9132 16856 9160
rect 16500 9092 16528 9132
rect 16850 9120 16856 9132
rect 16908 9120 16914 9172
rect 17034 9120 17040 9172
rect 17092 9160 17098 9172
rect 17221 9163 17279 9169
rect 17221 9160 17233 9163
rect 17092 9132 17233 9160
rect 17092 9120 17098 9132
rect 17221 9129 17233 9132
rect 17267 9129 17279 9163
rect 17221 9123 17279 9129
rect 17313 9163 17371 9169
rect 17313 9129 17325 9163
rect 17359 9160 17371 9163
rect 17402 9160 17408 9172
rect 17359 9132 17408 9160
rect 17359 9129 17371 9132
rect 17313 9123 17371 9129
rect 17402 9120 17408 9132
rect 17460 9120 17466 9172
rect 17494 9120 17500 9172
rect 17552 9160 17558 9172
rect 17552 9132 18000 9160
rect 17552 9120 17558 9132
rect 15865 9064 16528 9092
rect 16592 9064 17908 9092
rect 9140 8996 9536 9024
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 9861 9027 9919 9033
rect 9861 9024 9873 9027
rect 9640 8996 9873 9024
rect 9640 8984 9646 8996
rect 9861 8993 9873 8996
rect 9907 9024 9919 9027
rect 10597 9027 10655 9033
rect 10597 9024 10609 9027
rect 9907 8996 10609 9024
rect 9907 8993 9919 8996
rect 9861 8987 9919 8993
rect 10597 8993 10609 8996
rect 10643 8993 10655 9027
rect 13262 9024 13268 9036
rect 10597 8987 10655 8993
rect 12728 8996 13268 9024
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 8754 8956 8760 8968
rect 8435 8928 8760 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 12728 8956 12756 8996
rect 13262 8984 13268 8996
rect 13320 8984 13326 9036
rect 13446 9024 13452 9036
rect 13407 8996 13452 9024
rect 13446 8984 13452 8996
rect 13504 8984 13510 9036
rect 13538 8984 13544 9036
rect 13596 9024 13602 9036
rect 13814 9024 13820 9036
rect 13596 8996 13820 9024
rect 13596 8984 13602 8996
rect 13814 8984 13820 8996
rect 13872 8984 13878 9036
rect 16114 8984 16120 9036
rect 16172 9024 16178 9036
rect 16482 9024 16488 9036
rect 16172 8996 16488 9024
rect 16172 8984 16178 8996
rect 16482 8984 16488 8996
rect 16540 9024 16546 9036
rect 16592 9033 16620 9064
rect 16577 9027 16635 9033
rect 16577 9024 16589 9027
rect 16540 8996 16589 9024
rect 16540 8984 16546 8996
rect 16577 8993 16589 8996
rect 16623 8993 16635 9027
rect 17586 9024 17592 9036
rect 16577 8987 16635 8993
rect 17512 8996 17592 9024
rect 9784 8928 12756 8956
rect 12805 8959 12863 8965
rect 8481 8891 8539 8897
rect 8481 8857 8493 8891
rect 8527 8888 8539 8891
rect 8527 8860 9260 8888
rect 8527 8857 8539 8860
rect 8481 8851 8539 8857
rect 8754 8820 8760 8832
rect 8128 8792 8760 8820
rect 8021 8783 8079 8789
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9232 8829 9260 8860
rect 9490 8848 9496 8900
rect 9548 8888 9554 8900
rect 9677 8891 9735 8897
rect 9677 8888 9689 8891
rect 9548 8860 9689 8888
rect 9548 8848 9554 8860
rect 9677 8857 9689 8860
rect 9723 8857 9735 8891
rect 9677 8851 9735 8857
rect 9217 8823 9275 8829
rect 9217 8789 9229 8823
rect 9263 8789 9275 8823
rect 9217 8783 9275 8789
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 9585 8823 9643 8829
rect 9585 8820 9597 8823
rect 9364 8792 9597 8820
rect 9364 8780 9370 8792
rect 9585 8789 9597 8792
rect 9631 8820 9643 8823
rect 9784 8820 9812 8928
rect 12805 8925 12817 8959
rect 12851 8956 12863 8959
rect 14182 8956 14188 8968
rect 12851 8928 14188 8956
rect 12851 8925 12863 8928
rect 12805 8919 12863 8925
rect 14182 8916 14188 8928
rect 14240 8956 14246 8968
rect 14553 8959 14611 8965
rect 14553 8956 14565 8959
rect 14240 8928 14565 8956
rect 14240 8916 14246 8928
rect 14553 8925 14565 8928
rect 14599 8925 14611 8959
rect 16393 8959 16451 8965
rect 14553 8919 14611 8925
rect 14752 8928 16160 8956
rect 12560 8891 12618 8897
rect 12560 8857 12572 8891
rect 12606 8888 12618 8891
rect 12710 8888 12716 8900
rect 12606 8860 12716 8888
rect 12606 8857 12618 8860
rect 12560 8851 12618 8857
rect 12710 8848 12716 8860
rect 12768 8848 12774 8900
rect 12986 8848 12992 8900
rect 13044 8888 13050 8900
rect 13265 8891 13323 8897
rect 13265 8888 13277 8891
rect 13044 8860 13277 8888
rect 13044 8848 13050 8860
rect 13265 8857 13277 8860
rect 13311 8888 13323 8891
rect 14752 8888 14780 8928
rect 14826 8897 14832 8900
rect 13311 8860 14780 8888
rect 13311 8857 13323 8860
rect 13265 8851 13323 8857
rect 14820 8851 14832 8897
rect 14884 8888 14890 8900
rect 14884 8860 14920 8888
rect 14826 8848 14832 8851
rect 14884 8848 14890 8860
rect 16132 8832 16160 8928
rect 16393 8925 16405 8959
rect 16439 8956 16451 8959
rect 17512 8956 17540 8996
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 17880 9033 17908 9064
rect 17865 9027 17923 9033
rect 17865 8993 17877 9027
rect 17911 8993 17923 9027
rect 17865 8987 17923 8993
rect 17972 9024 18000 9132
rect 18782 9024 18788 9036
rect 17972 8996 18788 9024
rect 17678 8956 17684 8968
rect 16439 8928 17540 8956
rect 17639 8928 17684 8956
rect 16439 8925 16451 8928
rect 16393 8919 16451 8925
rect 17678 8916 17684 8928
rect 17736 8916 17742 8968
rect 17773 8959 17831 8965
rect 17773 8925 17785 8959
rect 17819 8956 17831 8959
rect 17972 8956 18000 8996
rect 18782 8984 18788 8996
rect 18840 8984 18846 9036
rect 17819 8928 18000 8956
rect 18233 8959 18291 8965
rect 17819 8925 17831 8928
rect 17773 8919 17831 8925
rect 18233 8925 18245 8959
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 16761 8891 16819 8897
rect 16761 8857 16773 8891
rect 16807 8888 16819 8891
rect 17494 8888 17500 8900
rect 16807 8860 17500 8888
rect 16807 8857 16819 8860
rect 16761 8851 16819 8857
rect 17494 8848 17500 8860
rect 17552 8848 17558 8900
rect 18248 8888 18276 8919
rect 17604 8860 18276 8888
rect 9631 8792 9812 8820
rect 10045 8823 10103 8829
rect 9631 8789 9643 8792
rect 9585 8783 9643 8789
rect 10045 8789 10057 8823
rect 10091 8820 10103 8823
rect 10226 8820 10232 8832
rect 10091 8792 10232 8820
rect 10091 8789 10103 8792
rect 10045 8783 10103 8789
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 10410 8820 10416 8832
rect 10371 8792 10416 8820
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 10505 8823 10563 8829
rect 10505 8789 10517 8823
rect 10551 8820 10563 8823
rect 11146 8820 11152 8832
rect 10551 8792 11152 8820
rect 10551 8789 10563 8792
rect 10505 8783 10563 8789
rect 11146 8780 11152 8792
rect 11204 8780 11210 8832
rect 11425 8823 11483 8829
rect 11425 8789 11437 8823
rect 11471 8820 11483 8823
rect 13170 8820 13176 8832
rect 11471 8792 13176 8820
rect 11471 8789 11483 8792
rect 11425 8783 11483 8789
rect 13170 8780 13176 8792
rect 13228 8780 13234 8832
rect 13357 8823 13415 8829
rect 13357 8789 13369 8823
rect 13403 8820 13415 8823
rect 13538 8820 13544 8832
rect 13403 8792 13544 8820
rect 13403 8789 13415 8792
rect 13357 8783 13415 8789
rect 13538 8780 13544 8792
rect 13596 8780 13602 8832
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 14093 8823 14151 8829
rect 14093 8820 14105 8823
rect 13872 8792 14105 8820
rect 13872 8780 13878 8792
rect 14093 8789 14105 8792
rect 14139 8789 14151 8823
rect 14093 8783 14151 8789
rect 15746 8780 15752 8832
rect 15804 8820 15810 8832
rect 16025 8823 16083 8829
rect 16025 8820 16037 8823
rect 15804 8792 16037 8820
rect 15804 8780 15810 8792
rect 16025 8789 16037 8792
rect 16071 8789 16083 8823
rect 16025 8783 16083 8789
rect 16114 8780 16120 8832
rect 16172 8820 16178 8832
rect 16209 8823 16267 8829
rect 16209 8820 16221 8823
rect 16172 8792 16221 8820
rect 16172 8780 16178 8792
rect 16209 8789 16221 8792
rect 16255 8789 16267 8823
rect 16209 8783 16267 8789
rect 16666 8780 16672 8832
rect 16724 8820 16730 8832
rect 16853 8823 16911 8829
rect 16853 8820 16865 8823
rect 16724 8792 16865 8820
rect 16724 8780 16730 8792
rect 16853 8789 16865 8792
rect 16899 8789 16911 8823
rect 16853 8783 16911 8789
rect 16942 8780 16948 8832
rect 17000 8820 17006 8832
rect 17604 8820 17632 8860
rect 18414 8820 18420 8832
rect 17000 8792 17632 8820
rect 18375 8792 18420 8820
rect 17000 8780 17006 8792
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 1104 8730 18860 8752
rect 1104 8678 5398 8730
rect 5450 8678 5462 8730
rect 5514 8678 5526 8730
rect 5578 8678 5590 8730
rect 5642 8678 5654 8730
rect 5706 8678 9846 8730
rect 9898 8678 9910 8730
rect 9962 8678 9974 8730
rect 10026 8678 10038 8730
rect 10090 8678 10102 8730
rect 10154 8678 14294 8730
rect 14346 8678 14358 8730
rect 14410 8678 14422 8730
rect 14474 8678 14486 8730
rect 14538 8678 14550 8730
rect 14602 8678 18860 8730
rect 1104 8656 18860 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 2225 8619 2283 8625
rect 2225 8616 2237 8619
rect 1811 8588 2237 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 2225 8585 2237 8588
rect 2271 8585 2283 8619
rect 2590 8616 2596 8628
rect 2551 8588 2596 8616
rect 2225 8579 2283 8585
rect 2590 8576 2596 8588
rect 2648 8576 2654 8628
rect 2958 8576 2964 8628
rect 3016 8616 3022 8628
rect 3421 8619 3479 8625
rect 3421 8616 3433 8619
rect 3016 8588 3433 8616
rect 3016 8576 3022 8588
rect 3421 8585 3433 8588
rect 3467 8585 3479 8619
rect 3421 8579 3479 8585
rect 3694 8576 3700 8628
rect 3752 8616 3758 8628
rect 4062 8616 4068 8628
rect 3752 8588 4068 8616
rect 3752 8576 3758 8588
rect 4062 8576 4068 8588
rect 4120 8576 4126 8628
rect 5258 8576 5264 8628
rect 5316 8616 5322 8628
rect 5353 8619 5411 8625
rect 5353 8616 5365 8619
rect 5316 8588 5365 8616
rect 5316 8576 5322 8588
rect 5353 8585 5365 8588
rect 5399 8585 5411 8619
rect 5353 8579 5411 8585
rect 5813 8619 5871 8625
rect 5813 8585 5825 8619
rect 5859 8616 5871 8619
rect 5994 8616 6000 8628
rect 5859 8588 6000 8616
rect 5859 8585 5871 8588
rect 5813 8579 5871 8585
rect 2682 8508 2688 8560
rect 2740 8548 2746 8560
rect 3878 8548 3884 8560
rect 2740 8520 3884 8548
rect 2740 8508 2746 8520
rect 1578 8412 1584 8424
rect 1539 8384 1584 8412
rect 1578 8372 1584 8384
rect 1636 8372 1642 8424
rect 1673 8415 1731 8421
rect 1673 8381 1685 8415
rect 1719 8381 1731 8415
rect 2682 8412 2688 8424
rect 2643 8384 2688 8412
rect 1673 8375 1731 8381
rect 1688 8344 1716 8375
rect 2682 8372 2688 8384
rect 2740 8372 2746 8424
rect 2884 8421 2912 8520
rect 3878 8508 3884 8520
rect 3936 8508 3942 8560
rect 5534 8508 5540 8560
rect 5592 8548 5598 8560
rect 5828 8548 5856 8579
rect 5994 8576 6000 8588
rect 6052 8576 6058 8628
rect 6730 8616 6736 8628
rect 6691 8588 6736 8616
rect 6730 8576 6736 8588
rect 6788 8616 6794 8628
rect 6788 8588 6960 8616
rect 6788 8576 6794 8588
rect 5592 8520 5856 8548
rect 5592 8508 5598 8520
rect 5902 8508 5908 8560
rect 5960 8548 5966 8560
rect 6181 8551 6239 8557
rect 6181 8548 6193 8551
rect 5960 8520 6193 8548
rect 5960 8508 5966 8520
rect 6181 8517 6193 8520
rect 6227 8548 6239 8551
rect 6641 8551 6699 8557
rect 6641 8548 6653 8551
rect 6227 8520 6653 8548
rect 6227 8517 6239 8520
rect 6181 8511 6239 8517
rect 6641 8517 6653 8520
rect 6687 8548 6699 8551
rect 6822 8548 6828 8560
rect 6687 8520 6828 8548
rect 6687 8517 6699 8520
rect 6641 8511 6699 8517
rect 6822 8508 6828 8520
rect 6880 8508 6886 8560
rect 6932 8548 6960 8588
rect 7006 8576 7012 8628
rect 7064 8616 7070 8628
rect 7469 8619 7527 8625
rect 7469 8616 7481 8619
rect 7064 8588 7481 8616
rect 7064 8576 7070 8588
rect 7469 8585 7481 8588
rect 7515 8616 7527 8619
rect 7558 8616 7564 8628
rect 7515 8588 7564 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 7929 8619 7987 8625
rect 7929 8616 7941 8619
rect 7861 8588 7941 8616
rect 7193 8551 7251 8557
rect 7193 8548 7205 8551
rect 6932 8520 7205 8548
rect 7193 8517 7205 8520
rect 7239 8517 7251 8551
rect 7193 8511 7251 8517
rect 7650 8508 7656 8560
rect 7708 8548 7714 8560
rect 7861 8548 7889 8588
rect 7929 8585 7941 8588
rect 7975 8585 7987 8619
rect 7929 8579 7987 8585
rect 8110 8576 8116 8628
rect 8168 8616 8174 8628
rect 10778 8616 10784 8628
rect 8168 8588 10784 8616
rect 8168 8576 8174 8588
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 12989 8619 13047 8625
rect 12989 8585 13001 8619
rect 13035 8616 13047 8619
rect 13357 8619 13415 8625
rect 13357 8616 13369 8619
rect 13035 8588 13369 8616
rect 13035 8585 13047 8588
rect 12989 8579 13047 8585
rect 13357 8585 13369 8588
rect 13403 8585 13415 8619
rect 14277 8619 14335 8625
rect 14277 8616 14289 8619
rect 13357 8579 13415 8585
rect 13464 8588 14289 8616
rect 7708 8520 7889 8548
rect 7708 8508 7714 8520
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 8352 8520 8397 8548
rect 8352 8508 8358 8520
rect 8478 8508 8484 8560
rect 8536 8548 8542 8560
rect 8757 8551 8815 8557
rect 8757 8548 8769 8551
rect 8536 8520 8769 8548
rect 8536 8508 8542 8520
rect 8757 8517 8769 8520
rect 8803 8517 8815 8551
rect 12069 8551 12127 8557
rect 12069 8548 12081 8551
rect 8757 8511 8815 8517
rect 9048 8520 12081 8548
rect 4338 8480 4344 8492
rect 4299 8452 4344 8480
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 5166 8440 5172 8492
rect 5224 8480 5230 8492
rect 5261 8483 5319 8489
rect 5261 8480 5273 8483
rect 5224 8452 5273 8480
rect 5224 8440 5230 8452
rect 5261 8449 5273 8452
rect 5307 8480 5319 8483
rect 5997 8483 6055 8489
rect 5997 8480 6009 8483
rect 5307 8452 6009 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5997 8449 6009 8452
rect 6043 8480 6055 8483
rect 8018 8480 8024 8492
rect 6043 8452 8024 8480
rect 6043 8449 6055 8452
rect 5997 8443 6055 8449
rect 8018 8440 8024 8452
rect 8076 8440 8082 8492
rect 8110 8440 8116 8492
rect 8168 8480 8174 8492
rect 9048 8480 9076 8520
rect 12069 8517 12081 8520
rect 12115 8548 12127 8551
rect 13464 8548 13492 8588
rect 14277 8585 14289 8588
rect 14323 8616 14335 8619
rect 14642 8616 14648 8628
rect 14323 8588 14648 8616
rect 14323 8585 14335 8588
rect 14277 8579 14335 8585
rect 14642 8576 14648 8588
rect 14700 8576 14706 8628
rect 14737 8619 14795 8625
rect 14737 8585 14749 8619
rect 14783 8616 14795 8619
rect 14826 8616 14832 8628
rect 14783 8588 14832 8616
rect 14783 8585 14795 8588
rect 14737 8579 14795 8585
rect 14826 8576 14832 8588
rect 14884 8616 14890 8628
rect 16485 8619 16543 8625
rect 14884 8588 16436 8616
rect 14884 8576 14890 8588
rect 13722 8548 13728 8560
rect 12115 8520 13492 8548
rect 13683 8520 13728 8548
rect 12115 8517 12127 8520
rect 12069 8511 12127 8517
rect 13722 8508 13728 8520
rect 13780 8508 13786 8560
rect 13814 8508 13820 8560
rect 13872 8548 13878 8560
rect 13872 8520 13917 8548
rect 13872 8508 13878 8520
rect 14182 8508 14188 8560
rect 14240 8548 14246 8560
rect 16408 8548 16436 8588
rect 16485 8585 16497 8619
rect 16531 8616 16543 8619
rect 16942 8616 16948 8628
rect 16531 8588 16948 8616
rect 16531 8585 16543 8588
rect 16485 8579 16543 8585
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17405 8619 17463 8625
rect 17405 8616 17417 8619
rect 17184 8588 17417 8616
rect 17184 8576 17190 8588
rect 17405 8585 17417 8588
rect 17451 8585 17463 8619
rect 17405 8579 17463 8585
rect 17494 8576 17500 8628
rect 17552 8616 17558 8628
rect 17552 8588 17597 8616
rect 17552 8576 17558 8588
rect 17862 8576 17868 8628
rect 17920 8616 17926 8628
rect 17957 8619 18015 8625
rect 17957 8616 17969 8619
rect 17920 8588 17969 8616
rect 17920 8576 17926 8588
rect 17957 8585 17969 8588
rect 18003 8585 18015 8619
rect 17957 8579 18015 8585
rect 17310 8548 17316 8560
rect 14240 8520 16160 8548
rect 16408 8520 17316 8548
rect 14240 8508 14246 8520
rect 8168 8479 8717 8480
rect 8772 8479 9076 8480
rect 8168 8452 9076 8479
rect 8168 8440 8174 8452
rect 8689 8451 8800 8452
rect 9766 8440 9772 8492
rect 9824 8480 9830 8492
rect 10689 8483 10747 8489
rect 10689 8480 10701 8483
rect 9824 8452 10701 8480
rect 9824 8440 9830 8452
rect 10689 8449 10701 8452
rect 10735 8449 10747 8483
rect 11974 8480 11980 8492
rect 11935 8452 11980 8480
rect 10689 8443 10747 8449
rect 11974 8440 11980 8452
rect 12032 8440 12038 8492
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8480 12955 8483
rect 13630 8480 13636 8492
rect 12943 8452 13636 8480
rect 12943 8449 12955 8452
rect 12897 8443 12955 8449
rect 13630 8440 13636 8452
rect 13688 8440 13694 8492
rect 14528 8483 14586 8489
rect 14528 8449 14540 8483
rect 14574 8480 14586 8483
rect 14826 8480 14832 8492
rect 14574 8452 14832 8480
rect 14574 8449 14586 8452
rect 14528 8443 14586 8449
rect 14826 8440 14832 8452
rect 14884 8440 14890 8492
rect 15838 8480 15844 8492
rect 15896 8489 15902 8492
rect 16132 8489 16160 8520
rect 17310 8508 17316 8520
rect 17368 8548 17374 8560
rect 17368 8520 18092 8548
rect 17368 8508 17374 8520
rect 15808 8452 15844 8480
rect 15838 8440 15844 8452
rect 15896 8443 15908 8489
rect 16117 8483 16175 8489
rect 16117 8449 16129 8483
rect 16163 8449 16175 8483
rect 16298 8480 16304 8492
rect 16259 8452 16304 8480
rect 16117 8443 16175 8449
rect 15896 8440 15902 8443
rect 16298 8440 16304 8452
rect 16356 8440 16362 8492
rect 17034 8480 17040 8492
rect 16995 8452 17040 8480
rect 17034 8440 17040 8452
rect 17092 8440 17098 8492
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8480 17923 8483
rect 17954 8480 17960 8492
rect 17911 8452 17960 8480
rect 17911 8449 17923 8452
rect 17865 8443 17923 8449
rect 17954 8440 17960 8452
rect 18012 8440 18018 8492
rect 2869 8415 2927 8421
rect 2869 8381 2881 8415
rect 2915 8381 2927 8415
rect 2869 8375 2927 8381
rect 3050 8372 3056 8424
rect 3108 8412 3114 8424
rect 3145 8415 3203 8421
rect 3145 8412 3157 8415
rect 3108 8384 3157 8412
rect 3108 8372 3114 8384
rect 3145 8381 3157 8384
rect 3191 8381 3203 8415
rect 3145 8375 3203 8381
rect 3697 8415 3755 8421
rect 3697 8381 3709 8415
rect 3743 8412 3755 8415
rect 3878 8412 3884 8424
rect 3743 8384 3884 8412
rect 3743 8381 3755 8384
rect 3697 8375 3755 8381
rect 3878 8372 3884 8384
rect 3936 8372 3942 8424
rect 4430 8412 4436 8424
rect 4391 8384 4436 8412
rect 4430 8372 4436 8384
rect 4488 8372 4494 8424
rect 4522 8372 4528 8424
rect 4580 8412 4586 8424
rect 5445 8415 5503 8421
rect 4580 8384 4625 8412
rect 4580 8372 4586 8384
rect 5445 8381 5457 8415
rect 5491 8381 5503 8415
rect 6454 8412 6460 8424
rect 6415 8384 6460 8412
rect 5445 8375 5503 8381
rect 3973 8347 4031 8353
rect 3973 8344 3985 8347
rect 1688 8316 3985 8344
rect 3973 8313 3985 8316
rect 4019 8313 4031 8347
rect 3973 8307 4031 8313
rect 5074 8304 5080 8356
rect 5132 8344 5138 8356
rect 5132 8316 5212 8344
rect 5132 8304 5138 8316
rect 2133 8279 2191 8285
rect 2133 8245 2145 8279
rect 2179 8276 2191 8279
rect 2958 8276 2964 8288
rect 2179 8248 2964 8276
rect 2179 8245 2191 8248
rect 2133 8239 2191 8245
rect 2958 8236 2964 8248
rect 3016 8236 3022 8288
rect 3881 8279 3939 8285
rect 3881 8245 3893 8279
rect 3927 8276 3939 8279
rect 4062 8276 4068 8288
rect 3927 8248 4068 8276
rect 3927 8245 3939 8248
rect 3881 8239 3939 8245
rect 4062 8236 4068 8248
rect 4120 8236 4126 8288
rect 4154 8236 4160 8288
rect 4212 8276 4218 8288
rect 4893 8279 4951 8285
rect 4893 8276 4905 8279
rect 4212 8248 4905 8276
rect 4212 8236 4218 8248
rect 4893 8245 4905 8248
rect 4939 8245 4951 8279
rect 5184 8276 5212 8316
rect 5258 8304 5264 8356
rect 5316 8344 5322 8356
rect 5460 8344 5488 8375
rect 6454 8372 6460 8384
rect 6512 8372 6518 8424
rect 7098 8372 7104 8424
rect 7156 8412 7162 8424
rect 8386 8412 8392 8424
rect 7156 8384 7512 8412
rect 8347 8384 8392 8412
rect 7156 8372 7162 8384
rect 6822 8344 6828 8356
rect 5316 8316 5488 8344
rect 6012 8316 6828 8344
rect 5316 8304 5322 8316
rect 6012 8276 6040 8316
rect 6822 8304 6828 8316
rect 6880 8304 6886 8356
rect 7190 8304 7196 8356
rect 7248 8304 7254 8356
rect 7484 8344 7512 8384
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 8478 8372 8484 8424
rect 8536 8412 8542 8424
rect 11885 8415 11943 8421
rect 8536 8384 8581 8412
rect 8536 8372 8542 8384
rect 11885 8381 11897 8415
rect 11931 8412 11943 8415
rect 13170 8412 13176 8424
rect 11931 8384 12756 8412
rect 13083 8384 13176 8412
rect 11931 8381 11943 8384
rect 11885 8375 11943 8381
rect 12728 8356 12756 8384
rect 13170 8372 13176 8384
rect 13228 8412 13234 8424
rect 13446 8412 13452 8424
rect 13228 8384 13452 8412
rect 13228 8372 13234 8384
rect 13446 8372 13452 8384
rect 13504 8372 13510 8424
rect 14001 8415 14059 8421
rect 14001 8381 14013 8415
rect 14047 8412 14059 8415
rect 14274 8412 14280 8424
rect 14047 8384 14280 8412
rect 14047 8381 14059 8384
rect 14001 8375 14059 8381
rect 10045 8347 10103 8353
rect 10045 8344 10057 8347
rect 7484 8316 10057 8344
rect 10045 8313 10057 8316
rect 10091 8344 10103 8347
rect 10410 8344 10416 8356
rect 10091 8316 10416 8344
rect 10091 8313 10103 8316
rect 10045 8307 10103 8313
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 11514 8344 11520 8356
rect 11475 8316 11520 8344
rect 11514 8304 11520 8316
rect 11572 8304 11578 8356
rect 12526 8304 12532 8356
rect 12584 8344 12590 8356
rect 12584 8316 12629 8344
rect 12584 8304 12590 8316
rect 12710 8304 12716 8356
rect 12768 8344 12774 8356
rect 14016 8344 14044 8375
rect 14274 8372 14280 8384
rect 14332 8372 14338 8424
rect 16482 8372 16488 8424
rect 16540 8412 16546 8424
rect 16761 8415 16819 8421
rect 16761 8412 16773 8415
rect 16540 8384 16773 8412
rect 16540 8372 16546 8384
rect 16761 8381 16773 8384
rect 16807 8381 16819 8415
rect 16942 8412 16948 8424
rect 16903 8384 16948 8412
rect 16761 8375 16819 8381
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 18064 8421 18092 8520
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 18156 8452 18521 8480
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 12768 8316 14044 8344
rect 12768 8304 12774 8316
rect 14550 8304 14556 8356
rect 14608 8353 14614 8356
rect 14608 8347 14657 8353
rect 14608 8313 14611 8347
rect 14645 8313 14657 8347
rect 14608 8307 14657 8313
rect 14608 8304 14614 8307
rect 16390 8304 16396 8356
rect 16448 8344 16454 8356
rect 18156 8344 18184 8452
rect 18509 8449 18521 8452
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 18322 8344 18328 8356
rect 16448 8316 18184 8344
rect 18283 8316 18328 8344
rect 16448 8304 16454 8316
rect 18322 8304 18328 8316
rect 18380 8304 18386 8356
rect 5184 8248 6040 8276
rect 4893 8239 4951 8245
rect 6086 8236 6092 8288
rect 6144 8276 6150 8288
rect 6454 8276 6460 8288
rect 6144 8248 6460 8276
rect 6144 8236 6150 8248
rect 6454 8236 6460 8248
rect 6512 8236 6518 8288
rect 7101 8279 7159 8285
rect 7101 8245 7113 8279
rect 7147 8276 7159 8279
rect 7208 8276 7236 8304
rect 7147 8248 7236 8276
rect 7837 8279 7895 8285
rect 7147 8245 7159 8248
rect 7101 8239 7159 8245
rect 7837 8245 7849 8279
rect 7883 8276 7895 8279
rect 8110 8276 8116 8288
rect 7883 8248 8116 8276
rect 7883 8245 7895 8248
rect 7837 8239 7895 8245
rect 8110 8236 8116 8248
rect 8168 8236 8174 8288
rect 8202 8236 8208 8288
rect 8260 8276 8266 8288
rect 10226 8276 10232 8288
rect 8260 8248 10232 8276
rect 8260 8236 8266 8248
rect 10226 8236 10232 8248
rect 10284 8236 10290 8288
rect 11330 8276 11336 8288
rect 11291 8248 11336 8276
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 12434 8236 12440 8288
rect 12492 8276 12498 8288
rect 12492 8248 12537 8276
rect 12492 8236 12498 8248
rect 13906 8236 13912 8288
rect 13964 8276 13970 8288
rect 15930 8276 15936 8288
rect 13964 8248 15936 8276
rect 13964 8236 13970 8248
rect 15930 8236 15936 8248
rect 15988 8276 15994 8288
rect 18046 8276 18052 8288
rect 15988 8248 18052 8276
rect 15988 8236 15994 8248
rect 18046 8236 18052 8248
rect 18104 8236 18110 8288
rect 1104 8186 18860 8208
rect 1104 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 3430 8186
rect 3482 8134 7622 8186
rect 7674 8134 7686 8186
rect 7738 8134 7750 8186
rect 7802 8134 7814 8186
rect 7866 8134 7878 8186
rect 7930 8134 12070 8186
rect 12122 8134 12134 8186
rect 12186 8134 12198 8186
rect 12250 8134 12262 8186
rect 12314 8134 12326 8186
rect 12378 8134 16518 8186
rect 16570 8134 16582 8186
rect 16634 8134 16646 8186
rect 16698 8134 16710 8186
rect 16762 8134 16774 8186
rect 16826 8134 18860 8186
rect 1104 8112 18860 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 2314 8072 2320 8084
rect 2275 8044 2320 8072
rect 2314 8032 2320 8044
rect 2372 8032 2378 8084
rect 2682 8072 2688 8084
rect 2643 8044 2688 8072
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 4157 8075 4215 8081
rect 4157 8072 4169 8075
rect 3344 8044 4169 8072
rect 2498 7964 2504 8016
rect 2556 8004 2562 8016
rect 3344 8004 3372 8044
rect 4157 8041 4169 8044
rect 4203 8072 4215 8075
rect 5902 8072 5908 8084
rect 4203 8044 5908 8072
rect 4203 8041 4215 8044
rect 4157 8035 4215 8041
rect 5902 8032 5908 8044
rect 5960 8032 5966 8084
rect 5994 8032 6000 8084
rect 6052 8072 6058 8084
rect 8754 8072 8760 8084
rect 6052 8044 8760 8072
rect 6052 8032 6058 8044
rect 8754 8032 8760 8044
rect 8812 8032 8818 8084
rect 8938 8032 8944 8084
rect 8996 8072 9002 8084
rect 11701 8075 11759 8081
rect 11701 8072 11713 8075
rect 8996 8044 11713 8072
rect 8996 8032 9002 8044
rect 11701 8041 11713 8044
rect 11747 8072 11759 8075
rect 13814 8072 13820 8084
rect 11747 8044 13820 8072
rect 11747 8041 11759 8044
rect 11701 8035 11759 8041
rect 13814 8032 13820 8044
rect 13872 8072 13878 8084
rect 14182 8072 14188 8084
rect 13872 8044 14188 8072
rect 13872 8032 13878 8044
rect 14182 8032 14188 8044
rect 14240 8032 14246 8084
rect 15838 8072 15844 8084
rect 15799 8044 15844 8072
rect 15838 8032 15844 8044
rect 15896 8032 15902 8084
rect 16761 8075 16819 8081
rect 16040 8044 16712 8072
rect 2556 7976 3372 8004
rect 2556 7964 2562 7976
rect 3970 7964 3976 8016
rect 4028 8004 4034 8016
rect 8021 8007 8079 8013
rect 8021 8004 8033 8007
rect 4028 7976 8033 8004
rect 4028 7964 4034 7976
rect 8021 7973 8033 7976
rect 8067 7973 8079 8007
rect 8021 7967 8079 7973
rect 8386 7964 8392 8016
rect 8444 8004 8450 8016
rect 9033 8007 9091 8013
rect 9033 8004 9045 8007
rect 8444 7976 9045 8004
rect 8444 7964 8450 7976
rect 9033 7973 9045 7976
rect 9079 7973 9091 8007
rect 9766 8004 9772 8016
rect 9033 7967 9091 7973
rect 9324 7976 9772 8004
rect 3326 7936 3332 7948
rect 3287 7908 3332 7936
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 4617 7939 4675 7945
rect 4617 7905 4629 7939
rect 4663 7936 4675 7939
rect 5258 7936 5264 7948
rect 4663 7908 5264 7936
rect 4663 7905 4675 7908
rect 4617 7899 4675 7905
rect 5258 7896 5264 7908
rect 5316 7896 5322 7948
rect 7282 7936 7288 7948
rect 7243 7908 7288 7936
rect 7282 7896 7288 7908
rect 7340 7896 7346 7948
rect 7466 7936 7472 7948
rect 7427 7908 7472 7936
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 8665 7939 8723 7945
rect 8665 7905 8677 7939
rect 8711 7936 8723 7939
rect 9324 7936 9352 7976
rect 9766 7964 9772 7976
rect 9824 7964 9830 8016
rect 10042 8004 10048 8016
rect 9968 7976 10048 8004
rect 9582 7936 9588 7948
rect 8711 7908 9352 7936
rect 9543 7908 9588 7936
rect 8711 7905 8723 7908
rect 8665 7899 8723 7905
rect 9582 7896 9588 7908
rect 9640 7896 9646 7948
rect 9968 7945 9996 7976
rect 10042 7964 10048 7976
rect 10100 7964 10106 8016
rect 10226 8004 10232 8016
rect 10187 7976 10232 8004
rect 10226 7964 10232 7976
rect 10284 8004 10290 8016
rect 12250 8004 12256 8016
rect 10284 7976 12256 8004
rect 10284 7964 10290 7976
rect 12250 7964 12256 7976
rect 12308 7964 12314 8016
rect 13630 7964 13636 8016
rect 13688 8004 13694 8016
rect 14093 8007 14151 8013
rect 14093 8004 14105 8007
rect 13688 7976 14105 8004
rect 13688 7964 13694 7976
rect 14093 7973 14105 7976
rect 14139 7973 14151 8007
rect 15105 8007 15163 8013
rect 14093 7967 14151 7973
rect 14200 7976 14964 8004
rect 9953 7939 10011 7945
rect 9953 7905 9965 7939
rect 9999 7905 10011 7939
rect 9953 7899 10011 7905
rect 10137 7939 10195 7945
rect 10137 7905 10149 7939
rect 10183 7936 10195 7939
rect 14200 7936 14228 7976
rect 10183 7908 12388 7936
rect 10183 7905 10195 7908
rect 10137 7899 10195 7905
rect 1578 7828 1584 7880
rect 1636 7868 1642 7880
rect 1673 7871 1731 7877
rect 1673 7868 1685 7871
rect 1636 7840 1685 7868
rect 1636 7828 1642 7840
rect 1673 7837 1685 7840
rect 1719 7837 1731 7871
rect 1673 7831 1731 7837
rect 2593 7871 2651 7877
rect 2593 7837 2605 7871
rect 2639 7868 2651 7871
rect 2682 7868 2688 7880
rect 2639 7840 2688 7868
rect 2639 7837 2651 7840
rect 2593 7831 2651 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 3053 7871 3111 7877
rect 3053 7868 3065 7871
rect 2832 7840 3065 7868
rect 2832 7828 2838 7840
rect 3053 7837 3065 7840
rect 3099 7837 3111 7871
rect 3053 7831 3111 7837
rect 3142 7828 3148 7880
rect 3200 7868 3206 7880
rect 3513 7871 3571 7877
rect 3513 7868 3525 7871
rect 3200 7840 3525 7868
rect 3200 7828 3206 7840
rect 3513 7837 3525 7840
rect 3559 7837 3571 7871
rect 3513 7831 3571 7837
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7868 4399 7871
rect 4801 7871 4859 7877
rect 4801 7868 4813 7871
rect 4387 7840 4813 7868
rect 4387 7837 4399 7840
rect 4341 7831 4399 7837
rect 4801 7837 4813 7840
rect 4847 7868 4859 7871
rect 5810 7868 5816 7880
rect 4847 7840 5816 7868
rect 4847 7837 4859 7840
rect 4801 7831 4859 7837
rect 2314 7760 2320 7812
rect 2372 7800 2378 7812
rect 4356 7800 4384 7831
rect 5810 7828 5816 7840
rect 5868 7828 5874 7880
rect 7006 7868 7012 7880
rect 6967 7840 7012 7868
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 7561 7871 7619 7877
rect 7561 7837 7573 7871
rect 7607 7868 7619 7871
rect 8018 7868 8024 7880
rect 7607 7840 8024 7868
rect 7607 7837 7619 7840
rect 7561 7831 7619 7837
rect 8018 7828 8024 7840
rect 8076 7828 8082 7880
rect 8202 7828 8208 7880
rect 8260 7868 8266 7880
rect 8260 7840 8708 7868
rect 8260 7828 8266 7840
rect 2372 7772 4384 7800
rect 4709 7803 4767 7809
rect 2372 7760 2378 7772
rect 4709 7769 4721 7803
rect 4755 7800 4767 7803
rect 5534 7800 5540 7812
rect 4755 7772 5540 7800
rect 4755 7769 4767 7772
rect 4709 7763 4767 7769
rect 1762 7692 1768 7744
rect 1820 7732 1826 7744
rect 2409 7735 2467 7741
rect 2409 7732 2421 7735
rect 1820 7704 2421 7732
rect 1820 7692 1826 7704
rect 2409 7701 2421 7704
rect 2455 7701 2467 7735
rect 2409 7695 2467 7701
rect 3973 7735 4031 7741
rect 3973 7701 3985 7735
rect 4019 7732 4031 7735
rect 4724 7732 4752 7763
rect 5534 7760 5540 7772
rect 5592 7800 5598 7812
rect 6270 7800 6276 7812
rect 5592 7772 6276 7800
rect 5592 7760 5598 7772
rect 6270 7760 6276 7772
rect 6328 7760 6334 7812
rect 8481 7803 8539 7809
rect 8481 7800 8493 7803
rect 7944 7772 8493 7800
rect 4019 7704 4752 7732
rect 4019 7701 4031 7704
rect 3973 7695 4031 7701
rect 5074 7692 5080 7744
rect 5132 7732 5138 7744
rect 5169 7735 5227 7741
rect 5169 7732 5181 7735
rect 5132 7704 5181 7732
rect 5132 7692 5138 7704
rect 5169 7701 5181 7704
rect 5215 7701 5227 7735
rect 5718 7732 5724 7744
rect 5679 7704 5724 7732
rect 5169 7695 5227 7701
rect 5718 7692 5724 7704
rect 5776 7692 5782 7744
rect 7944 7741 7972 7772
rect 8481 7769 8493 7772
rect 8527 7769 8539 7803
rect 8680 7800 8708 7840
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 9401 7871 9459 7877
rect 9401 7868 9413 7871
rect 8812 7840 9413 7868
rect 8812 7828 8818 7840
rect 9401 7837 9413 7840
rect 9447 7868 9459 7871
rect 9674 7868 9680 7880
rect 9447 7840 9680 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 10152 7868 10180 7899
rect 10410 7868 10416 7880
rect 9968 7844 10180 7868
rect 9784 7840 10180 7844
rect 10371 7840 10416 7868
rect 9784 7816 9996 7840
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 11146 7828 11152 7880
rect 11204 7868 11210 7880
rect 12253 7871 12311 7877
rect 12253 7868 12265 7871
rect 11204 7840 12265 7868
rect 11204 7828 11210 7840
rect 12253 7837 12265 7840
rect 12299 7837 12311 7871
rect 12360 7868 12388 7908
rect 13280 7908 14228 7936
rect 14645 7939 14703 7945
rect 13280 7868 13308 7908
rect 14645 7905 14657 7939
rect 14691 7905 14703 7939
rect 14645 7899 14703 7905
rect 12360 7840 13308 7868
rect 12253 7831 12311 7837
rect 13630 7828 13636 7880
rect 13688 7868 13694 7880
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13688 7840 13737 7868
rect 13688 7828 13694 7840
rect 13725 7837 13737 7840
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 9493 7803 9551 7809
rect 9493 7800 9505 7803
rect 8680 7772 9505 7800
rect 8481 7763 8539 7769
rect 9493 7769 9505 7772
rect 9539 7800 9551 7803
rect 9784 7800 9812 7816
rect 9539 7772 9812 7800
rect 9539 7769 9551 7772
rect 9493 7763 9551 7769
rect 11330 7760 11336 7812
rect 11388 7800 11394 7812
rect 12498 7803 12556 7809
rect 12498 7800 12510 7803
rect 11388 7772 12510 7800
rect 11388 7760 11394 7772
rect 12498 7769 12510 7772
rect 12544 7769 12556 7803
rect 14274 7800 14280 7812
rect 12498 7763 12556 7769
rect 13648 7772 14280 7800
rect 7929 7735 7987 7741
rect 7929 7701 7941 7735
rect 7975 7701 7987 7735
rect 8386 7732 8392 7744
rect 8347 7704 8392 7732
rect 7929 7695 7987 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 13648 7741 13676 7772
rect 14274 7760 14280 7772
rect 14332 7800 14338 7812
rect 14660 7800 14688 7899
rect 14936 7880 14964 7976
rect 15105 7973 15117 8007
rect 15151 8004 15163 8007
rect 16040 8004 16068 8044
rect 15151 7976 16068 8004
rect 16117 8007 16175 8013
rect 15151 7973 15163 7976
rect 15105 7967 15163 7973
rect 16117 7973 16129 8007
rect 16163 7973 16175 8007
rect 16684 8004 16712 8044
rect 16761 8041 16773 8075
rect 16807 8072 16819 8075
rect 16942 8072 16948 8084
rect 16807 8044 16948 8072
rect 16807 8041 16819 8044
rect 16761 8035 16819 8041
rect 16942 8032 16948 8044
rect 17000 8032 17006 8084
rect 17034 8032 17040 8084
rect 17092 8072 17098 8084
rect 17589 8075 17647 8081
rect 17589 8072 17601 8075
rect 17092 8044 17601 8072
rect 17092 8032 17098 8044
rect 17589 8041 17601 8044
rect 17635 8041 17647 8075
rect 17589 8035 17647 8041
rect 17494 8004 17500 8016
rect 16684 7976 17500 8004
rect 16117 7967 16175 7973
rect 15654 7896 15660 7948
rect 15712 7936 15718 7948
rect 16132 7936 16160 7967
rect 17494 7964 17500 7976
rect 17552 7964 17558 8016
rect 16942 7936 16948 7948
rect 15712 7908 16068 7936
rect 16132 7908 16948 7936
rect 15712 7896 15718 7908
rect 14918 7868 14924 7880
rect 14879 7840 14924 7868
rect 14918 7828 14924 7840
rect 14976 7828 14982 7880
rect 15102 7828 15108 7880
rect 15160 7868 15166 7880
rect 15197 7871 15255 7877
rect 15197 7868 15209 7871
rect 15160 7840 15209 7868
rect 15160 7828 15166 7840
rect 15197 7837 15209 7840
rect 15243 7837 15255 7871
rect 15930 7868 15936 7880
rect 15197 7831 15255 7837
rect 15764 7840 15936 7868
rect 15764 7800 15792 7840
rect 15930 7828 15936 7840
rect 15988 7828 15994 7880
rect 16040 7868 16068 7908
rect 16942 7896 16948 7908
rect 17000 7896 17006 7948
rect 17310 7936 17316 7948
rect 17271 7908 17316 7936
rect 17310 7896 17316 7908
rect 17368 7936 17374 7948
rect 18141 7939 18199 7945
rect 18141 7936 18153 7939
rect 17368 7908 18153 7936
rect 17368 7896 17374 7908
rect 18141 7905 18153 7908
rect 18187 7905 18199 7939
rect 18141 7899 18199 7905
rect 16206 7868 16212 7880
rect 16040 7840 16212 7868
rect 16206 7828 16212 7840
rect 16264 7828 16270 7880
rect 16393 7871 16451 7877
rect 16393 7837 16405 7871
rect 16439 7837 16451 7871
rect 16393 7831 16451 7837
rect 16669 7871 16727 7877
rect 16669 7837 16681 7871
rect 16715 7868 16727 7871
rect 17126 7868 17132 7880
rect 16715 7840 17132 7868
rect 16715 7837 16727 7840
rect 16669 7831 16727 7837
rect 14332 7772 14688 7800
rect 15120 7772 15792 7800
rect 14332 7760 14338 7772
rect 13633 7735 13691 7741
rect 13633 7701 13645 7735
rect 13679 7701 13691 7735
rect 13906 7732 13912 7744
rect 13867 7704 13912 7732
rect 13633 7695 13691 7701
rect 13906 7692 13912 7704
rect 13964 7692 13970 7744
rect 14182 7692 14188 7744
rect 14240 7732 14246 7744
rect 14461 7735 14519 7741
rect 14461 7732 14473 7735
rect 14240 7704 14473 7732
rect 14240 7692 14246 7704
rect 14461 7701 14473 7704
rect 14507 7701 14519 7735
rect 14461 7695 14519 7701
rect 14553 7735 14611 7741
rect 14553 7701 14565 7735
rect 14599 7732 14611 7735
rect 15120 7732 15148 7772
rect 15838 7760 15844 7812
rect 15896 7800 15902 7812
rect 16408 7800 16436 7831
rect 17126 7828 17132 7840
rect 17184 7828 17190 7880
rect 17954 7868 17960 7880
rect 17915 7840 17960 7868
rect 17954 7828 17960 7840
rect 18012 7868 18018 7880
rect 18230 7868 18236 7880
rect 18012 7840 18236 7868
rect 18012 7828 18018 7840
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 15896 7772 16436 7800
rect 15896 7760 15902 7772
rect 14599 7704 15148 7732
rect 14599 7701 14611 7704
rect 14553 7695 14611 7701
rect 15194 7692 15200 7744
rect 15252 7732 15258 7744
rect 16209 7735 16267 7741
rect 16209 7732 16221 7735
rect 15252 7704 16221 7732
rect 15252 7692 15258 7704
rect 16209 7701 16221 7704
rect 16255 7701 16267 7735
rect 16209 7695 16267 7701
rect 16390 7692 16396 7744
rect 16448 7732 16454 7744
rect 16485 7735 16543 7741
rect 16485 7732 16497 7735
rect 16448 7704 16497 7732
rect 16448 7692 16454 7704
rect 16485 7701 16497 7704
rect 16531 7701 16543 7735
rect 16485 7695 16543 7701
rect 16850 7692 16856 7744
rect 16908 7732 16914 7744
rect 17129 7735 17187 7741
rect 17129 7732 17141 7735
rect 16908 7704 17141 7732
rect 16908 7692 16914 7704
rect 17129 7701 17141 7704
rect 17175 7701 17187 7735
rect 17129 7695 17187 7701
rect 17218 7692 17224 7744
rect 17276 7732 17282 7744
rect 18046 7732 18052 7744
rect 17276 7704 17321 7732
rect 17959 7704 18052 7732
rect 17276 7692 17282 7704
rect 18046 7692 18052 7704
rect 18104 7732 18110 7744
rect 18417 7735 18475 7741
rect 18417 7732 18429 7735
rect 18104 7704 18429 7732
rect 18104 7692 18110 7704
rect 18417 7701 18429 7704
rect 18463 7732 18475 7735
rect 18690 7732 18696 7744
rect 18463 7704 18696 7732
rect 18463 7701 18475 7704
rect 18417 7695 18475 7701
rect 18690 7692 18696 7704
rect 18748 7692 18754 7744
rect 1104 7642 18860 7664
rect 1104 7590 5398 7642
rect 5450 7590 5462 7642
rect 5514 7590 5526 7642
rect 5578 7590 5590 7642
rect 5642 7590 5654 7642
rect 5706 7590 9846 7642
rect 9898 7590 9910 7642
rect 9962 7590 9974 7642
rect 10026 7590 10038 7642
rect 10090 7590 10102 7642
rect 10154 7590 14294 7642
rect 14346 7590 14358 7642
rect 14410 7590 14422 7642
rect 14474 7590 14486 7642
rect 14538 7590 14550 7642
rect 14602 7590 18860 7642
rect 1104 7568 18860 7590
rect 1581 7531 1639 7537
rect 1581 7497 1593 7531
rect 1627 7528 1639 7531
rect 1670 7528 1676 7540
rect 1627 7500 1676 7528
rect 1627 7497 1639 7500
rect 1581 7491 1639 7497
rect 1670 7488 1676 7500
rect 1728 7488 1734 7540
rect 1854 7528 1860 7540
rect 1815 7500 1860 7528
rect 1854 7488 1860 7500
rect 1912 7488 1918 7540
rect 2590 7488 2596 7540
rect 2648 7528 2654 7540
rect 2685 7531 2743 7537
rect 2685 7528 2697 7531
rect 2648 7500 2697 7528
rect 2648 7488 2654 7500
rect 2685 7497 2697 7500
rect 2731 7497 2743 7531
rect 3050 7528 3056 7540
rect 3011 7500 3056 7528
rect 2685 7491 2743 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 4065 7531 4123 7537
rect 4065 7497 4077 7531
rect 4111 7528 4123 7531
rect 4154 7528 4160 7540
rect 4111 7500 4160 7528
rect 4111 7497 4123 7500
rect 4065 7491 4123 7497
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4430 7488 4436 7540
rect 4488 7528 4494 7540
rect 4617 7531 4675 7537
rect 4617 7528 4629 7531
rect 4488 7500 4629 7528
rect 4488 7488 4494 7500
rect 4617 7497 4629 7500
rect 4663 7497 4675 7531
rect 5074 7528 5080 7540
rect 5035 7500 5080 7528
rect 4617 7491 4675 7497
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5445 7531 5503 7537
rect 5445 7497 5457 7531
rect 5491 7497 5503 7531
rect 5902 7528 5908 7540
rect 5863 7500 5908 7528
rect 5445 7491 5503 7497
rect 3878 7420 3884 7472
rect 3936 7460 3942 7472
rect 4985 7463 5043 7469
rect 3936 7432 4200 7460
rect 3936 7420 3942 7432
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 2038 7392 2044 7404
rect 1999 7364 2044 7392
rect 2038 7352 2044 7364
rect 2096 7352 2102 7404
rect 2409 7395 2467 7401
rect 2409 7361 2421 7395
rect 2455 7361 2467 7395
rect 2409 7355 2467 7361
rect 2222 7256 2228 7268
rect 2183 7228 2228 7256
rect 2222 7216 2228 7228
rect 2280 7216 2286 7268
rect 2424 7256 2452 7355
rect 2590 7352 2596 7404
rect 2648 7392 2654 7404
rect 3142 7392 3148 7404
rect 2648 7364 3148 7392
rect 2648 7352 2654 7364
rect 3142 7352 3148 7364
rect 3200 7352 3206 7404
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7392 3755 7395
rect 4062 7392 4068 7404
rect 3743 7364 4068 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4172 7401 4200 7432
rect 4985 7429 4997 7463
rect 5031 7460 5043 7463
rect 5460 7460 5488 7491
rect 5902 7488 5908 7500
rect 5960 7488 5966 7540
rect 7282 7488 7288 7540
rect 7340 7528 7346 7540
rect 9493 7531 9551 7537
rect 9493 7528 9505 7531
rect 7340 7500 9505 7528
rect 7340 7488 7346 7500
rect 9493 7497 9505 7500
rect 9539 7497 9551 7531
rect 9493 7491 9551 7497
rect 9585 7531 9643 7537
rect 9585 7497 9597 7531
rect 9631 7528 9643 7531
rect 9766 7528 9772 7540
rect 9631 7500 9772 7528
rect 9631 7497 9643 7500
rect 9585 7491 9643 7497
rect 5031 7432 5488 7460
rect 5031 7429 5043 7432
rect 4985 7423 5043 7429
rect 7006 7420 7012 7472
rect 7064 7460 7070 7472
rect 7837 7463 7895 7469
rect 7837 7460 7849 7463
rect 7064 7432 7849 7460
rect 7064 7420 7070 7432
rect 7837 7429 7849 7432
rect 7883 7429 7895 7463
rect 7837 7423 7895 7429
rect 8380 7463 8438 7469
rect 8380 7429 8392 7463
rect 8426 7460 8438 7463
rect 8478 7460 8484 7472
rect 8426 7432 8484 7460
rect 8426 7429 8438 7432
rect 8380 7423 8438 7429
rect 8478 7420 8484 7432
rect 8536 7420 8542 7472
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 5813 7395 5871 7401
rect 5813 7361 5825 7395
rect 5859 7392 5871 7395
rect 5902 7392 5908 7404
rect 5859 7364 5908 7392
rect 5859 7361 5871 7364
rect 5813 7355 5871 7361
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 7478 7395 7536 7401
rect 7478 7392 7490 7395
rect 6104 7364 7490 7392
rect 3326 7324 3332 7336
rect 3239 7296 3332 7324
rect 3326 7284 3332 7296
rect 3384 7324 3390 7336
rect 3973 7327 4031 7333
rect 3973 7324 3985 7327
rect 3384 7296 3985 7324
rect 3384 7284 3390 7296
rect 3973 7293 3985 7296
rect 4019 7324 4031 7327
rect 4890 7324 4896 7336
rect 4019 7296 4896 7324
rect 4019 7293 4031 7296
rect 3973 7287 4031 7293
rect 4890 7284 4896 7296
rect 4948 7324 4954 7336
rect 6104 7333 6132 7364
rect 7478 7361 7490 7364
rect 7524 7361 7536 7395
rect 7478 7355 7536 7361
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7392 7803 7395
rect 8110 7392 8116 7404
rect 7791 7364 8116 7392
rect 7791 7361 7803 7364
rect 7745 7355 7803 7361
rect 8110 7352 8116 7364
rect 8168 7352 8174 7404
rect 9508 7392 9536 7491
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 11054 7528 11060 7540
rect 11015 7500 11060 7528
rect 11054 7488 11060 7500
rect 11112 7528 11118 7540
rect 11609 7531 11667 7537
rect 11609 7528 11621 7531
rect 11112 7500 11621 7528
rect 11112 7488 11118 7500
rect 11609 7497 11621 7500
rect 11655 7528 11667 7531
rect 11790 7528 11796 7540
rect 11655 7500 11796 7528
rect 11655 7497 11667 7500
rect 11609 7491 11667 7497
rect 11790 7488 11796 7500
rect 11848 7488 11854 7540
rect 12345 7531 12403 7537
rect 12345 7497 12357 7531
rect 12391 7528 12403 7531
rect 12805 7531 12863 7537
rect 12805 7528 12817 7531
rect 12391 7500 12817 7528
rect 12391 7497 12403 7500
rect 12345 7491 12403 7497
rect 12805 7497 12817 7500
rect 12851 7497 12863 7531
rect 14182 7528 14188 7540
rect 12805 7491 12863 7497
rect 13924 7500 14188 7528
rect 10502 7420 10508 7472
rect 10560 7460 10566 7472
rect 10698 7463 10756 7469
rect 10698 7460 10710 7463
rect 10560 7432 10710 7460
rect 10560 7420 10566 7432
rect 10698 7429 10710 7432
rect 10744 7429 10756 7463
rect 10698 7423 10756 7429
rect 12434 7420 12440 7472
rect 12492 7460 12498 7472
rect 13265 7463 13323 7469
rect 13265 7460 13277 7463
rect 12492 7432 13277 7460
rect 12492 7420 12498 7432
rect 13265 7429 13277 7432
rect 13311 7429 13323 7463
rect 13265 7423 13323 7429
rect 9674 7392 9680 7404
rect 9508 7364 9680 7392
rect 9674 7352 9680 7364
rect 9732 7352 9738 7404
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7392 12311 7395
rect 12526 7392 12532 7404
rect 12299 7364 12532 7392
rect 12299 7361 12311 7364
rect 12253 7355 12311 7361
rect 12526 7352 12532 7364
rect 12584 7352 12590 7404
rect 13173 7395 13231 7401
rect 13173 7361 13185 7395
rect 13219 7392 13231 7395
rect 13538 7392 13544 7404
rect 13219 7364 13544 7392
rect 13219 7361 13231 7364
rect 13173 7355 13231 7361
rect 5169 7327 5227 7333
rect 5169 7324 5181 7327
rect 4948 7296 5181 7324
rect 4948 7284 4954 7296
rect 5169 7293 5181 7296
rect 5215 7293 5227 7327
rect 5169 7287 5227 7293
rect 6089 7327 6147 7333
rect 6089 7293 6101 7327
rect 6135 7293 6147 7327
rect 6089 7287 6147 7293
rect 10965 7327 11023 7333
rect 10965 7293 10977 7327
rect 11011 7324 11023 7327
rect 11146 7324 11152 7336
rect 11011 7296 11152 7324
rect 11011 7293 11023 7296
rect 10965 7287 11023 7293
rect 3513 7259 3571 7265
rect 3513 7256 3525 7259
rect 2424 7228 3525 7256
rect 3513 7225 3525 7228
rect 3559 7225 3571 7259
rect 3513 7219 3571 7225
rect 4338 7216 4344 7268
rect 4396 7256 4402 7268
rect 4525 7259 4583 7265
rect 4525 7256 4537 7259
rect 4396 7228 4537 7256
rect 4396 7216 4402 7228
rect 4525 7225 4537 7228
rect 4571 7225 4583 7259
rect 4525 7219 4583 7225
rect 5184 7188 5212 7287
rect 5258 7216 5264 7268
rect 5316 7256 5322 7268
rect 6104 7256 6132 7287
rect 11146 7284 11152 7296
rect 11204 7284 11210 7336
rect 11974 7284 11980 7336
rect 12032 7324 12038 7336
rect 12069 7327 12127 7333
rect 12069 7324 12081 7327
rect 12032 7296 12081 7324
rect 12032 7284 12038 7296
rect 12069 7293 12081 7296
rect 12115 7293 12127 7327
rect 13188 7324 13216 7355
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 13814 7392 13820 7404
rect 13775 7364 13820 7392
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 13924 7392 13952 7500
rect 14182 7488 14188 7500
rect 14240 7488 14246 7540
rect 14918 7488 14924 7540
rect 14976 7528 14982 7540
rect 16393 7531 16451 7537
rect 16393 7528 16405 7531
rect 14976 7500 16405 7528
rect 14976 7488 14982 7500
rect 16393 7497 16405 7500
rect 16439 7497 16451 7531
rect 16393 7491 16451 7497
rect 16758 7488 16764 7540
rect 16816 7528 16822 7540
rect 17681 7531 17739 7537
rect 17681 7528 17693 7531
rect 16816 7500 17693 7528
rect 16816 7488 16822 7500
rect 17681 7497 17693 7500
rect 17727 7528 17739 7531
rect 17954 7528 17960 7540
rect 17727 7500 17816 7528
rect 17915 7500 17960 7528
rect 17727 7497 17739 7500
rect 17681 7491 17739 7497
rect 14084 7463 14142 7469
rect 14084 7429 14096 7463
rect 14130 7460 14142 7463
rect 17313 7463 17371 7469
rect 17313 7460 17325 7463
rect 14130 7432 17325 7460
rect 14130 7429 14142 7432
rect 14084 7423 14142 7429
rect 17313 7429 17325 7432
rect 17359 7429 17371 7463
rect 17788 7460 17816 7500
rect 17954 7488 17960 7500
rect 18012 7488 18018 7540
rect 18414 7528 18420 7540
rect 18375 7500 18420 7528
rect 18414 7488 18420 7500
rect 18472 7488 18478 7540
rect 17862 7460 17868 7472
rect 17788 7432 17868 7460
rect 17313 7423 17371 7429
rect 17862 7420 17868 7432
rect 17920 7420 17926 7472
rect 15286 7392 15292 7404
rect 13924 7364 15148 7392
rect 15247 7364 15292 7392
rect 13446 7324 13452 7336
rect 12069 7287 12127 7293
rect 12176 7296 13216 7324
rect 13359 7296 13452 7324
rect 5316 7228 6132 7256
rect 11333 7259 11391 7265
rect 5316 7216 5322 7228
rect 11333 7225 11345 7259
rect 11379 7256 11391 7259
rect 11698 7256 11704 7268
rect 11379 7228 11704 7256
rect 11379 7225 11391 7228
rect 11333 7219 11391 7225
rect 11698 7216 11704 7228
rect 11756 7216 11762 7268
rect 12176 7256 12204 7296
rect 13446 7284 13452 7296
rect 13504 7324 13510 7336
rect 13630 7324 13636 7336
rect 13504 7296 13636 7324
rect 13504 7284 13510 7296
rect 13630 7284 13636 7296
rect 13688 7284 13694 7336
rect 13924 7324 13952 7364
rect 13832 7296 13952 7324
rect 15120 7324 15148 7364
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 15565 7395 15623 7401
rect 15565 7392 15577 7395
rect 15528 7364 15577 7392
rect 15528 7352 15534 7364
rect 15565 7361 15577 7364
rect 15611 7361 15623 7395
rect 15565 7355 15623 7361
rect 15654 7352 15660 7404
rect 15712 7392 15718 7404
rect 15841 7395 15899 7401
rect 15841 7392 15853 7395
rect 15712 7364 15853 7392
rect 15712 7352 15718 7364
rect 15841 7361 15853 7364
rect 15887 7361 15899 7395
rect 16114 7392 16120 7404
rect 16075 7364 16120 7392
rect 15841 7355 15899 7361
rect 15746 7324 15752 7336
rect 15120 7296 15752 7324
rect 11808 7228 12204 7256
rect 6365 7191 6423 7197
rect 6365 7188 6377 7191
rect 5184 7160 6377 7188
rect 6365 7157 6377 7160
rect 6411 7157 6423 7191
rect 6365 7151 6423 7157
rect 6822 7148 6828 7200
rect 6880 7188 6886 7200
rect 11808 7197 11836 7228
rect 12250 7216 12256 7268
rect 12308 7256 12314 7268
rect 13832 7256 13860 7296
rect 15746 7284 15752 7296
rect 15804 7284 15810 7336
rect 15856 7324 15884 7355
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 16669 7395 16727 7401
rect 16669 7361 16681 7395
rect 16715 7392 16727 7395
rect 16850 7392 16856 7404
rect 16715 7364 16856 7392
rect 16715 7361 16727 7364
rect 16669 7355 16727 7361
rect 16850 7352 16856 7364
rect 16908 7352 16914 7404
rect 17402 7392 17408 7404
rect 17363 7364 17408 7392
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 18138 7392 18144 7404
rect 18099 7364 18144 7392
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 18230 7352 18236 7404
rect 18288 7392 18294 7404
rect 18288 7364 18333 7392
rect 18288 7352 18294 7364
rect 16758 7324 16764 7336
rect 15856 7296 16764 7324
rect 16758 7284 16764 7296
rect 16816 7284 16822 7336
rect 18046 7324 18052 7336
rect 17512 7296 18052 7324
rect 12308 7228 13860 7256
rect 12308 7216 12314 7228
rect 15930 7216 15936 7268
rect 15988 7256 15994 7268
rect 16301 7259 16359 7265
rect 16301 7256 16313 7259
rect 15988 7228 16313 7256
rect 15988 7216 15994 7228
rect 16301 7225 16313 7228
rect 16347 7225 16359 7259
rect 16301 7219 16359 7225
rect 11793 7191 11851 7197
rect 11793 7188 11805 7191
rect 6880 7160 11805 7188
rect 6880 7148 6886 7160
rect 11793 7157 11805 7160
rect 11839 7157 11851 7191
rect 12710 7188 12716 7200
rect 12671 7160 12716 7188
rect 11793 7151 11851 7157
rect 12710 7148 12716 7160
rect 12768 7148 12774 7200
rect 13722 7188 13728 7200
rect 13683 7160 13728 7188
rect 13722 7148 13728 7160
rect 13780 7148 13786 7200
rect 15102 7148 15108 7200
rect 15160 7188 15166 7200
rect 15197 7191 15255 7197
rect 15197 7188 15209 7191
rect 15160 7160 15209 7188
rect 15160 7148 15166 7160
rect 15197 7157 15209 7160
rect 15243 7157 15255 7191
rect 15197 7151 15255 7157
rect 15473 7191 15531 7197
rect 15473 7157 15485 7191
rect 15519 7188 15531 7191
rect 15562 7188 15568 7200
rect 15519 7160 15568 7188
rect 15519 7157 15531 7160
rect 15473 7151 15531 7157
rect 15562 7148 15568 7160
rect 15620 7148 15626 7200
rect 15746 7188 15752 7200
rect 15707 7160 15752 7188
rect 15746 7148 15752 7160
rect 15804 7148 15810 7200
rect 16025 7191 16083 7197
rect 16025 7157 16037 7191
rect 16071 7188 16083 7191
rect 17512 7188 17540 7296
rect 18046 7284 18052 7296
rect 18104 7284 18110 7336
rect 17589 7259 17647 7265
rect 17589 7225 17601 7259
rect 17635 7256 17647 7259
rect 17770 7256 17776 7268
rect 17635 7228 17776 7256
rect 17635 7225 17647 7228
rect 17589 7219 17647 7225
rect 17770 7216 17776 7228
rect 17828 7216 17834 7268
rect 16071 7160 17540 7188
rect 16071 7157 16083 7160
rect 16025 7151 16083 7157
rect 1104 7098 18860 7120
rect 1104 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 3430 7098
rect 3482 7046 7622 7098
rect 7674 7046 7686 7098
rect 7738 7046 7750 7098
rect 7802 7046 7814 7098
rect 7866 7046 7878 7098
rect 7930 7046 12070 7098
rect 12122 7046 12134 7098
rect 12186 7046 12198 7098
rect 12250 7046 12262 7098
rect 12314 7046 12326 7098
rect 12378 7046 16518 7098
rect 16570 7046 16582 7098
rect 16634 7046 16646 7098
rect 16698 7046 16710 7098
rect 16762 7046 16774 7098
rect 16826 7046 18860 7098
rect 1104 7024 18860 7046
rect 1486 6984 1492 6996
rect 1447 6956 1492 6984
rect 1486 6944 1492 6956
rect 1544 6944 1550 6996
rect 2590 6984 2596 6996
rect 2551 6956 2596 6984
rect 2590 6944 2596 6956
rect 2648 6944 2654 6996
rect 5169 6987 5227 6993
rect 5169 6953 5181 6987
rect 5215 6984 5227 6987
rect 5258 6984 5264 6996
rect 5215 6956 5264 6984
rect 5215 6953 5227 6956
rect 5169 6947 5227 6953
rect 5258 6944 5264 6956
rect 5316 6944 5322 6996
rect 7653 6987 7711 6993
rect 7653 6953 7665 6987
rect 7699 6984 7711 6987
rect 8294 6984 8300 6996
rect 7699 6956 8300 6984
rect 7699 6953 7711 6956
rect 7653 6947 7711 6953
rect 8294 6944 8300 6956
rect 8352 6944 8358 6996
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 8573 6987 8631 6993
rect 8573 6984 8585 6987
rect 8444 6956 8585 6984
rect 8444 6944 8450 6956
rect 8573 6953 8585 6956
rect 8619 6953 8631 6987
rect 8573 6947 8631 6953
rect 10413 6987 10471 6993
rect 10413 6953 10425 6987
rect 10459 6984 10471 6987
rect 10502 6984 10508 6996
rect 10459 6956 10508 6984
rect 10459 6953 10471 6956
rect 10413 6947 10471 6953
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 11974 6984 11980 6996
rect 11935 6956 11980 6984
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 12492 6956 13584 6984
rect 12492 6944 12498 6956
rect 2314 6916 2320 6928
rect 2275 6888 2320 6916
rect 2314 6876 2320 6888
rect 2372 6876 2378 6928
rect 5902 6876 5908 6928
rect 5960 6916 5966 6928
rect 6730 6916 6736 6928
rect 5960 6888 6736 6916
rect 5960 6876 5966 6888
rect 6730 6876 6736 6888
rect 6788 6916 6794 6928
rect 6788 6888 7144 6916
rect 6788 6876 6794 6888
rect 3329 6851 3387 6857
rect 3329 6817 3341 6851
rect 3375 6848 3387 6851
rect 6825 6851 6883 6857
rect 3375 6820 3740 6848
rect 3375 6817 3387 6820
rect 3329 6811 3387 6817
rect 1673 6783 1731 6789
rect 1673 6749 1685 6783
rect 1719 6780 1731 6783
rect 1762 6780 1768 6792
rect 1719 6752 1768 6780
rect 1719 6749 1731 6752
rect 1673 6743 1731 6749
rect 1762 6740 1768 6752
rect 1820 6740 1826 6792
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6749 2099 6783
rect 2041 6743 2099 6749
rect 2056 6712 2084 6743
rect 2130 6740 2136 6792
rect 2188 6780 2194 6792
rect 2188 6752 2233 6780
rect 2188 6740 2194 6752
rect 2590 6740 2596 6792
rect 2648 6780 2654 6792
rect 2685 6783 2743 6789
rect 2685 6780 2697 6783
rect 2648 6752 2697 6780
rect 2648 6740 2654 6752
rect 2685 6749 2697 6752
rect 2731 6749 2743 6783
rect 2685 6743 2743 6749
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6749 3663 6783
rect 3605 6743 3663 6749
rect 3234 6712 3240 6724
rect 2056 6684 3240 6712
rect 3234 6672 3240 6684
rect 3292 6672 3298 6724
rect 1854 6644 1860 6656
rect 1815 6616 1860 6644
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 3421 6647 3479 6653
rect 3421 6613 3433 6647
rect 3467 6644 3479 6647
rect 3510 6644 3516 6656
rect 3467 6616 3516 6644
rect 3467 6613 3479 6616
rect 3421 6607 3479 6613
rect 3510 6604 3516 6616
rect 3568 6604 3574 6656
rect 3620 6644 3648 6743
rect 3712 6712 3740 6820
rect 6825 6817 6837 6851
rect 6871 6848 6883 6851
rect 6914 6848 6920 6860
rect 6871 6820 6920 6848
rect 6871 6817 6883 6820
rect 6825 6811 6883 6817
rect 6914 6808 6920 6820
rect 6972 6808 6978 6860
rect 7116 6857 7144 6888
rect 7282 6876 7288 6928
rect 7340 6916 7346 6928
rect 8938 6916 8944 6928
rect 7340 6888 7972 6916
rect 8899 6888 8944 6916
rect 7340 6876 7346 6888
rect 7101 6851 7159 6857
rect 7101 6817 7113 6851
rect 7147 6817 7159 6851
rect 7101 6811 7159 6817
rect 7190 6808 7196 6860
rect 7248 6848 7254 6860
rect 7650 6848 7656 6860
rect 7248 6820 7656 6848
rect 7248 6808 7254 6820
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 7944 6857 7972 6888
rect 8938 6876 8944 6888
rect 8996 6876 9002 6928
rect 11790 6876 11796 6928
rect 11848 6916 11854 6928
rect 11848 6888 12572 6916
rect 11848 6876 11854 6888
rect 7929 6851 7987 6857
rect 7929 6817 7941 6851
rect 7975 6817 7987 6851
rect 7929 6811 7987 6817
rect 8478 6808 8484 6860
rect 8536 6848 8542 6860
rect 9493 6851 9551 6857
rect 9493 6848 9505 6851
rect 8536 6820 9505 6848
rect 8536 6808 8542 6820
rect 9493 6817 9505 6820
rect 9539 6817 9551 6851
rect 9493 6811 9551 6817
rect 11974 6808 11980 6860
rect 12032 6848 12038 6860
rect 12161 6851 12219 6857
rect 12161 6848 12173 6851
rect 12032 6820 12173 6848
rect 12032 6808 12038 6820
rect 12161 6817 12173 6820
rect 12207 6817 12219 6851
rect 12434 6848 12440 6860
rect 12161 6811 12219 6817
rect 12268 6820 12440 6848
rect 3789 6783 3847 6789
rect 3789 6749 3801 6783
rect 3835 6780 3847 6783
rect 3878 6780 3884 6792
rect 3835 6752 3884 6780
rect 3835 6749 3847 6752
rect 3789 6743 3847 6749
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 4338 6740 4344 6792
rect 4396 6780 4402 6792
rect 5261 6783 5319 6789
rect 5261 6780 5273 6783
rect 4396 6752 5273 6780
rect 4396 6740 4402 6752
rect 5261 6749 5273 6752
rect 5307 6780 5319 6783
rect 5718 6780 5724 6792
rect 5307 6752 5724 6780
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 7374 6740 7380 6792
rect 7432 6780 7438 6792
rect 7745 6783 7803 6789
rect 7745 6780 7757 6783
rect 7432 6752 7757 6780
rect 7432 6740 7438 6752
rect 7745 6749 7757 6752
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 8128 6752 9628 6780
rect 4034 6715 4092 6721
rect 4034 6712 4046 6715
rect 3712 6684 4046 6712
rect 4034 6681 4046 6684
rect 4080 6681 4092 6715
rect 4034 6675 4092 6681
rect 4154 6672 4160 6724
rect 4212 6712 4218 6724
rect 6914 6712 6920 6724
rect 4212 6684 6920 6712
rect 4212 6672 4218 6684
rect 6914 6672 6920 6684
rect 6972 6672 6978 6724
rect 8128 6712 8156 6752
rect 7024 6684 8156 6712
rect 8205 6715 8263 6721
rect 7024 6644 7052 6684
rect 8205 6681 8217 6715
rect 8251 6712 8263 6715
rect 8938 6712 8944 6724
rect 8251 6684 8944 6712
rect 8251 6681 8263 6684
rect 8205 6675 8263 6681
rect 8938 6672 8944 6684
rect 8996 6672 9002 6724
rect 9398 6712 9404 6724
rect 9048 6684 9404 6712
rect 3620 6616 7052 6644
rect 7285 6647 7343 6653
rect 7285 6613 7297 6647
rect 7331 6644 7343 6647
rect 7926 6644 7932 6656
rect 7331 6616 7932 6644
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 8018 6604 8024 6656
rect 8076 6644 8082 6656
rect 8113 6647 8171 6653
rect 8113 6644 8125 6647
rect 8076 6616 8125 6644
rect 8076 6604 8082 6616
rect 8113 6613 8125 6616
rect 8159 6613 8171 6647
rect 8754 6644 8760 6656
rect 8667 6616 8760 6644
rect 8113 6607 8171 6613
rect 8754 6604 8760 6616
rect 8812 6644 8818 6656
rect 9048 6644 9076 6684
rect 9398 6672 9404 6684
rect 9456 6672 9462 6724
rect 9306 6644 9312 6656
rect 8812 6616 9076 6644
rect 9267 6616 9312 6644
rect 8812 6604 8818 6616
rect 9306 6604 9312 6616
rect 9364 6604 9370 6656
rect 9600 6644 9628 6752
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 9769 6783 9827 6789
rect 9769 6780 9781 6783
rect 9732 6752 9781 6780
rect 9732 6740 9738 6752
rect 9769 6749 9781 6752
rect 9815 6749 9827 6783
rect 9769 6743 9827 6749
rect 10597 6783 10655 6789
rect 10597 6749 10609 6783
rect 10643 6780 10655 6783
rect 11146 6780 11152 6792
rect 10643 6752 11152 6780
rect 10643 6749 10655 6752
rect 10597 6743 10655 6749
rect 11146 6740 11152 6752
rect 11204 6740 11210 6792
rect 10864 6715 10922 6721
rect 10864 6681 10876 6715
rect 10910 6712 10922 6715
rect 12268 6712 12296 6820
rect 12434 6808 12440 6820
rect 12492 6808 12498 6860
rect 12544 6848 12572 6888
rect 13262 6848 13268 6860
rect 12544 6820 13268 6848
rect 13262 6808 13268 6820
rect 13320 6808 13326 6860
rect 13556 6857 13584 6956
rect 15470 6944 15476 6996
rect 15528 6984 15534 6996
rect 15528 6956 16528 6984
rect 15528 6944 15534 6956
rect 16500 6928 16528 6956
rect 16592 6956 17172 6984
rect 13814 6876 13820 6928
rect 13872 6916 13878 6928
rect 14734 6916 14740 6928
rect 13872 6888 14740 6916
rect 13872 6876 13878 6888
rect 14734 6876 14740 6888
rect 14792 6876 14798 6928
rect 16482 6876 16488 6928
rect 16540 6876 16546 6928
rect 13541 6851 13599 6857
rect 13541 6817 13553 6851
rect 13587 6848 13599 6851
rect 13630 6848 13636 6860
rect 13587 6820 13636 6848
rect 13587 6817 13599 6820
rect 13541 6811 13599 6817
rect 13630 6808 13636 6820
rect 13688 6808 13694 6860
rect 13906 6808 13912 6860
rect 13964 6848 13970 6860
rect 13964 6820 14964 6848
rect 13964 6808 13970 6820
rect 12894 6740 12900 6792
rect 12952 6780 12958 6792
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 12952 6752 14105 6780
rect 12952 6740 12958 6752
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14826 6780 14832 6792
rect 14787 6752 14832 6780
rect 14093 6743 14151 6749
rect 14826 6740 14832 6752
rect 14884 6740 14890 6792
rect 14936 6780 14964 6820
rect 16592 6780 16620 6956
rect 16684 6888 16988 6916
rect 16684 6860 16712 6888
rect 16666 6808 16672 6860
rect 16724 6808 16730 6860
rect 16850 6848 16856 6860
rect 16811 6820 16856 6848
rect 16850 6808 16856 6820
rect 16908 6808 16914 6860
rect 16960 6848 16988 6888
rect 16960 6820 17080 6848
rect 14936 6752 16620 6780
rect 10910 6684 12296 6712
rect 12345 6715 12403 6721
rect 10910 6681 10922 6684
rect 10864 6675 10922 6681
rect 12345 6681 12357 6715
rect 12391 6712 12403 6715
rect 13262 6712 13268 6724
rect 12391 6684 12940 6712
rect 13223 6684 13268 6712
rect 12391 6681 12403 6684
rect 12345 6675 12403 6681
rect 11422 6644 11428 6656
rect 9600 6616 11428 6644
rect 11422 6604 11428 6616
rect 11480 6604 11486 6656
rect 12434 6604 12440 6656
rect 12492 6644 12498 6656
rect 12492 6616 12537 6644
rect 12492 6604 12498 6616
rect 12618 6604 12624 6656
rect 12676 6644 12682 6656
rect 12912 6653 12940 6684
rect 13262 6672 13268 6684
rect 13320 6672 13326 6724
rect 13357 6715 13415 6721
rect 13357 6681 13369 6715
rect 13403 6712 13415 6715
rect 13814 6712 13820 6724
rect 13403 6684 13820 6712
rect 13403 6681 13415 6684
rect 13357 6675 13415 6681
rect 13814 6672 13820 6684
rect 13872 6672 13878 6724
rect 15096 6715 15154 6721
rect 15096 6681 15108 6715
rect 15142 6712 15154 6715
rect 15654 6712 15660 6724
rect 15142 6684 15660 6712
rect 15142 6681 15154 6684
rect 15096 6675 15154 6681
rect 15654 6672 15660 6684
rect 15712 6672 15718 6724
rect 16850 6712 16856 6724
rect 16224 6684 16856 6712
rect 12805 6647 12863 6653
rect 12805 6644 12817 6647
rect 12676 6616 12817 6644
rect 12676 6604 12682 6616
rect 12805 6613 12817 6616
rect 12851 6613 12863 6647
rect 12805 6607 12863 6613
rect 12897 6647 12955 6653
rect 12897 6613 12909 6647
rect 12943 6613 12955 6647
rect 12897 6607 12955 6613
rect 13446 6604 13452 6656
rect 13504 6644 13510 6656
rect 13725 6647 13783 6653
rect 13725 6644 13737 6647
rect 13504 6616 13737 6644
rect 13504 6604 13510 6616
rect 13725 6613 13737 6616
rect 13771 6613 13783 6647
rect 14734 6644 14740 6656
rect 14695 6616 14740 6644
rect 13725 6607 13783 6613
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 16114 6604 16120 6656
rect 16172 6644 16178 6656
rect 16224 6653 16252 6684
rect 16850 6672 16856 6684
rect 16908 6672 16914 6724
rect 17052 6712 17080 6820
rect 17144 6780 17172 6956
rect 17218 6944 17224 6996
rect 17276 6984 17282 6996
rect 18414 6984 18420 6996
rect 17276 6956 17448 6984
rect 18375 6956 18420 6984
rect 17276 6944 17282 6956
rect 17420 6928 17448 6956
rect 18414 6944 18420 6956
rect 18472 6944 18478 6996
rect 17402 6876 17408 6928
rect 17460 6876 17466 6928
rect 17218 6808 17224 6860
rect 17276 6848 17282 6860
rect 17681 6851 17739 6857
rect 17681 6848 17693 6851
rect 17276 6820 17693 6848
rect 17276 6808 17282 6820
rect 17681 6817 17693 6820
rect 17727 6817 17739 6851
rect 17681 6811 17739 6817
rect 18233 6783 18291 6789
rect 18233 6780 18245 6783
rect 17144 6752 18245 6780
rect 18233 6749 18245 6752
rect 18279 6749 18291 6783
rect 18233 6743 18291 6749
rect 17497 6715 17555 6721
rect 17497 6712 17509 6715
rect 17052 6684 17509 6712
rect 17497 6681 17509 6684
rect 17543 6681 17555 6715
rect 17497 6675 17555 6681
rect 16209 6647 16267 6653
rect 16209 6644 16221 6647
rect 16172 6616 16221 6644
rect 16172 6604 16178 6616
rect 16209 6613 16221 6616
rect 16255 6613 16267 6647
rect 16209 6607 16267 6613
rect 16298 6604 16304 6656
rect 16356 6644 16362 6656
rect 16666 6644 16672 6656
rect 16356 6616 16401 6644
rect 16627 6616 16672 6644
rect 16356 6604 16362 6616
rect 16666 6604 16672 6616
rect 16724 6604 16730 6656
rect 16761 6647 16819 6653
rect 16761 6613 16773 6647
rect 16807 6644 16819 6647
rect 17129 6647 17187 6653
rect 17129 6644 17141 6647
rect 16807 6616 17141 6644
rect 16807 6613 16819 6616
rect 16761 6607 16819 6613
rect 17129 6613 17141 6616
rect 17175 6613 17187 6647
rect 17129 6607 17187 6613
rect 17402 6604 17408 6656
rect 17460 6644 17466 6656
rect 17589 6647 17647 6653
rect 17589 6644 17601 6647
rect 17460 6616 17601 6644
rect 17460 6604 17466 6616
rect 17589 6613 17601 6616
rect 17635 6644 17647 6647
rect 17678 6644 17684 6656
rect 17635 6616 17684 6644
rect 17635 6613 17647 6616
rect 17589 6607 17647 6613
rect 17678 6604 17684 6616
rect 17736 6604 17742 6656
rect 17954 6644 17960 6656
rect 17915 6616 17960 6644
rect 17954 6604 17960 6616
rect 18012 6604 18018 6656
rect 1104 6554 18860 6576
rect 1104 6502 5398 6554
rect 5450 6502 5462 6554
rect 5514 6502 5526 6554
rect 5578 6502 5590 6554
rect 5642 6502 5654 6554
rect 5706 6502 9846 6554
rect 9898 6502 9910 6554
rect 9962 6502 9974 6554
rect 10026 6502 10038 6554
rect 10090 6502 10102 6554
rect 10154 6502 14294 6554
rect 14346 6502 14358 6554
rect 14410 6502 14422 6554
rect 14474 6502 14486 6554
rect 14538 6502 14550 6554
rect 14602 6502 18860 6554
rect 1104 6480 18860 6502
rect 2041 6443 2099 6449
rect 2041 6409 2053 6443
rect 2087 6440 2099 6443
rect 2130 6440 2136 6452
rect 2087 6412 2136 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 2130 6400 2136 6412
rect 2188 6400 2194 6452
rect 2501 6443 2559 6449
rect 2501 6409 2513 6443
rect 2547 6440 2559 6443
rect 2682 6440 2688 6452
rect 2547 6412 2688 6440
rect 2547 6409 2559 6412
rect 2501 6403 2559 6409
rect 2682 6400 2688 6412
rect 2740 6400 2746 6452
rect 3234 6400 3240 6452
rect 3292 6440 3298 6452
rect 4341 6443 4399 6449
rect 4341 6440 4353 6443
rect 3292 6412 4353 6440
rect 3292 6400 3298 6412
rect 4341 6409 4353 6412
rect 4387 6409 4399 6443
rect 4341 6403 4399 6409
rect 6733 6443 6791 6449
rect 6733 6409 6745 6443
rect 6779 6440 6791 6443
rect 7006 6440 7012 6452
rect 6779 6412 7012 6440
rect 6779 6409 6791 6412
rect 6733 6403 6791 6409
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 7466 6440 7472 6452
rect 7116 6412 7472 6440
rect 3878 6332 3884 6384
rect 3936 6372 3942 6384
rect 5534 6372 5540 6384
rect 3936 6344 5540 6372
rect 3936 6332 3942 6344
rect 1670 6304 1676 6316
rect 1631 6276 1676 6304
rect 1670 6264 1676 6276
rect 1728 6264 1734 6316
rect 1854 6304 1860 6316
rect 1815 6276 1860 6304
rect 1854 6264 1860 6276
rect 1912 6264 1918 6316
rect 2314 6304 2320 6316
rect 2275 6276 2320 6304
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 2498 6264 2504 6316
rect 2556 6304 2562 6316
rect 3988 6313 4016 6344
rect 5534 6332 5540 6344
rect 5592 6332 5598 6384
rect 6825 6375 6883 6381
rect 6825 6341 6837 6375
rect 6871 6372 6883 6375
rect 6914 6372 6920 6384
rect 6871 6344 6920 6372
rect 6871 6341 6883 6344
rect 6825 6335 6883 6341
rect 6914 6332 6920 6344
rect 6972 6372 6978 6384
rect 7116 6372 7144 6412
rect 7466 6400 7472 6412
rect 7524 6400 7530 6452
rect 7650 6440 7656 6452
rect 7611 6412 7656 6440
rect 7650 6400 7656 6412
rect 7708 6400 7714 6452
rect 8018 6440 8024 6452
rect 7979 6412 8024 6440
rect 8018 6400 8024 6412
rect 8076 6400 8082 6452
rect 8389 6443 8447 6449
rect 8389 6409 8401 6443
rect 8435 6440 8447 6443
rect 9306 6440 9312 6452
rect 8435 6412 9312 6440
rect 8435 6409 8447 6412
rect 8389 6403 8447 6409
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 10686 6440 10692 6452
rect 9416 6412 10692 6440
rect 8478 6372 8484 6384
rect 6972 6344 7144 6372
rect 7484 6344 8484 6372
rect 6972 6332 6978 6344
rect 3717 6307 3775 6313
rect 3717 6304 3729 6307
rect 2556 6276 3729 6304
rect 2556 6264 2562 6276
rect 3717 6273 3729 6276
rect 3763 6304 3775 6307
rect 3973 6307 4031 6313
rect 3763 6276 3924 6304
rect 3763 6273 3775 6276
rect 3717 6267 3775 6273
rect 3896 6236 3924 6276
rect 3973 6273 3985 6307
rect 4019 6273 4031 6307
rect 3973 6267 4031 6273
rect 4154 6264 4160 6316
rect 4212 6304 4218 6316
rect 4249 6307 4307 6313
rect 4249 6304 4261 6307
rect 4212 6276 4261 6304
rect 4212 6264 4218 6276
rect 4249 6273 4261 6276
rect 4295 6273 4307 6307
rect 4522 6304 4528 6316
rect 4483 6276 4528 6304
rect 4249 6267 4307 6273
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 5810 6264 5816 6316
rect 5868 6313 5874 6316
rect 5868 6304 5880 6313
rect 5868 6276 5913 6304
rect 5868 6267 5880 6276
rect 5868 6264 5874 6267
rect 6086 6236 6092 6248
rect 3896 6208 4752 6236
rect 6047 6208 6092 6236
rect 1486 6100 1492 6112
rect 1447 6072 1492 6100
rect 1486 6060 1492 6072
rect 1544 6060 1550 6112
rect 2130 6100 2136 6112
rect 2091 6072 2136 6100
rect 2130 6060 2136 6072
rect 2188 6060 2194 6112
rect 2590 6100 2596 6112
rect 2551 6072 2596 6100
rect 2590 6060 2596 6072
rect 2648 6060 2654 6112
rect 4062 6100 4068 6112
rect 4023 6072 4068 6100
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4724 6109 4752 6208
rect 6086 6196 6092 6208
rect 6144 6196 6150 6248
rect 7484 6245 7512 6344
rect 8478 6332 8484 6344
rect 8536 6332 8542 6384
rect 8938 6332 8944 6384
rect 8996 6372 9002 6384
rect 9416 6372 9444 6412
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 12894 6440 12900 6452
rect 12855 6412 12900 6440
rect 12894 6400 12900 6412
rect 12952 6400 12958 6452
rect 13814 6400 13820 6452
rect 13872 6440 13878 6452
rect 14553 6443 14611 6449
rect 14553 6440 14565 6443
rect 13872 6412 14565 6440
rect 13872 6400 13878 6412
rect 14553 6409 14565 6412
rect 14599 6409 14611 6443
rect 14553 6403 14611 6409
rect 15197 6443 15255 6449
rect 15197 6409 15209 6443
rect 15243 6440 15255 6443
rect 15565 6443 15623 6449
rect 15565 6440 15577 6443
rect 15243 6412 15577 6440
rect 15243 6409 15255 6412
rect 15197 6403 15255 6409
rect 15565 6409 15577 6412
rect 15611 6409 15623 6443
rect 15565 6403 15623 6409
rect 16298 6400 16304 6452
rect 16356 6400 16362 6452
rect 16666 6440 16672 6452
rect 16627 6412 16672 6440
rect 16666 6400 16672 6412
rect 16724 6400 16730 6452
rect 17037 6443 17095 6449
rect 17037 6409 17049 6443
rect 17083 6440 17095 6443
rect 17954 6440 17960 6452
rect 17083 6412 17960 6440
rect 17083 6409 17095 6412
rect 17037 6403 17095 6409
rect 17954 6400 17960 6412
rect 18012 6400 18018 6452
rect 18138 6400 18144 6452
rect 18196 6440 18202 6452
rect 18325 6443 18383 6449
rect 18325 6440 18337 6443
rect 18196 6412 18337 6440
rect 18196 6400 18202 6412
rect 18325 6409 18337 6412
rect 18371 6409 18383 6443
rect 18325 6403 18383 6409
rect 8996 6344 9444 6372
rect 8996 6332 9002 6344
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 10226 6372 10232 6384
rect 9824 6344 10232 6372
rect 9824 6332 9830 6344
rect 10226 6332 10232 6344
rect 10284 6332 10290 6384
rect 10318 6332 10324 6384
rect 10376 6381 10382 6384
rect 10376 6372 10388 6381
rect 14274 6372 14280 6384
rect 10376 6344 10421 6372
rect 11532 6344 14280 6372
rect 10376 6335 10388 6344
rect 10376 6332 10382 6335
rect 8294 6264 8300 6316
rect 8352 6304 8358 6316
rect 9125 6307 9183 6313
rect 9125 6304 9137 6307
rect 8352 6276 9137 6304
rect 8352 6264 8358 6276
rect 9125 6273 9137 6276
rect 9171 6273 9183 6307
rect 10686 6304 10692 6316
rect 10647 6276 10692 6304
rect 9125 6267 9183 6273
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6205 6975 6239
rect 6917 6199 6975 6205
rect 7469 6239 7527 6245
rect 7469 6205 7481 6239
rect 7515 6205 7527 6239
rect 7469 6199 7527 6205
rect 7561 6239 7619 6245
rect 7561 6205 7573 6239
rect 7607 6236 7619 6239
rect 8938 6236 8944 6248
rect 7607 6208 8944 6236
rect 7607 6205 7619 6208
rect 7561 6199 7619 6205
rect 6932 6168 6960 6199
rect 6196 6140 6960 6168
rect 4709 6103 4767 6109
rect 4709 6069 4721 6103
rect 4755 6100 4767 6103
rect 5718 6100 5724 6112
rect 4755 6072 5724 6100
rect 4755 6069 4767 6072
rect 4709 6063 4767 6069
rect 5718 6060 5724 6072
rect 5776 6060 5782 6112
rect 5810 6060 5816 6112
rect 5868 6100 5874 6112
rect 6196 6100 6224 6140
rect 6362 6100 6368 6112
rect 5868 6072 6224 6100
rect 6323 6072 6368 6100
rect 5868 6060 5874 6072
rect 6362 6060 6368 6072
rect 6420 6060 6426 6112
rect 6914 6060 6920 6112
rect 6972 6100 6978 6112
rect 7659 6100 7687 6208
rect 8938 6196 8944 6208
rect 8996 6196 9002 6248
rect 7742 6128 7748 6180
rect 7800 6168 7806 6180
rect 8754 6168 8760 6180
rect 7800 6140 8760 6168
rect 7800 6128 7806 6140
rect 8754 6128 8760 6140
rect 8812 6128 8818 6180
rect 9140 6168 9168 6267
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 10597 6239 10655 6245
rect 10597 6205 10609 6239
rect 10643 6236 10655 6239
rect 11146 6236 11152 6248
rect 10643 6208 11152 6236
rect 10643 6205 10655 6208
rect 10597 6199 10655 6205
rect 11146 6196 11152 6208
rect 11204 6236 11210 6248
rect 11532 6245 11560 6344
rect 11784 6307 11842 6313
rect 11784 6273 11796 6307
rect 11830 6304 11842 6307
rect 12066 6304 12072 6316
rect 11830 6276 12072 6304
rect 11830 6273 11842 6276
rect 11784 6267 11842 6273
rect 12066 6264 12072 6276
rect 12124 6264 12130 6316
rect 13096 6313 13124 6344
rect 14274 6332 14280 6344
rect 14332 6372 14338 6384
rect 14826 6372 14832 6384
rect 14332 6344 14832 6372
rect 14332 6332 14338 6344
rect 14826 6332 14832 6344
rect 14884 6332 14890 6384
rect 15105 6375 15163 6381
rect 15105 6341 15117 6375
rect 15151 6372 15163 6375
rect 16316 6372 16344 6400
rect 15151 6344 16344 6372
rect 15151 6341 15163 6344
rect 15105 6335 15163 6341
rect 16482 6332 16488 6384
rect 16540 6372 16546 6384
rect 16540 6344 17448 6372
rect 16540 6332 16546 6344
rect 13081 6307 13139 6313
rect 13081 6273 13093 6307
rect 13127 6273 13139 6307
rect 13081 6267 13139 6273
rect 13348 6307 13406 6313
rect 13348 6273 13360 6307
rect 13394 6304 13406 6307
rect 14734 6304 14740 6316
rect 13394 6276 14740 6304
rect 13394 6273 13406 6276
rect 13348 6267 13406 6273
rect 14734 6264 14740 6276
rect 14792 6264 14798 6316
rect 15933 6307 15991 6313
rect 15933 6273 15945 6307
rect 15979 6273 15991 6307
rect 15933 6267 15991 6273
rect 11517 6239 11575 6245
rect 11517 6236 11529 6239
rect 11204 6208 11529 6236
rect 11204 6196 11210 6208
rect 11517 6205 11529 6208
rect 11563 6205 11575 6239
rect 11517 6199 11575 6205
rect 15102 6196 15108 6248
rect 15160 6236 15166 6248
rect 15289 6239 15347 6245
rect 15289 6236 15301 6239
rect 15160 6208 15301 6236
rect 15160 6196 15166 6208
rect 15289 6205 15301 6208
rect 15335 6205 15347 6239
rect 15289 6199 15347 6205
rect 9217 6171 9275 6177
rect 9217 6168 9229 6171
rect 9140 6140 9229 6168
rect 9217 6137 9229 6140
rect 9263 6137 9275 6171
rect 14737 6171 14795 6177
rect 14737 6168 14749 6171
rect 9217 6131 9275 6137
rect 12820 6140 13032 6168
rect 6972 6072 7687 6100
rect 6972 6060 6978 6072
rect 8386 6060 8392 6112
rect 8444 6100 8450 6112
rect 8481 6103 8539 6109
rect 8481 6100 8493 6103
rect 8444 6072 8493 6100
rect 8444 6060 8450 6072
rect 8481 6069 8493 6072
rect 8527 6069 8539 6103
rect 8481 6063 8539 6069
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 11333 6103 11391 6109
rect 11333 6100 11345 6103
rect 10284 6072 11345 6100
rect 10284 6060 10290 6072
rect 11333 6069 11345 6072
rect 11379 6069 11391 6103
rect 11333 6063 11391 6069
rect 11422 6060 11428 6112
rect 11480 6100 11486 6112
rect 12820 6100 12848 6140
rect 11480 6072 12848 6100
rect 13004 6100 13032 6140
rect 14016 6140 14749 6168
rect 14016 6100 14044 6140
rect 14737 6137 14749 6140
rect 14783 6137 14795 6171
rect 14737 6131 14795 6137
rect 14458 6100 14464 6112
rect 13004 6072 14044 6100
rect 14419 6072 14464 6100
rect 11480 6060 11486 6072
rect 14458 6060 14464 6072
rect 14516 6060 14522 6112
rect 15948 6100 15976 6267
rect 16850 6264 16856 6316
rect 16908 6304 16914 6316
rect 17034 6304 17040 6316
rect 16908 6276 17040 6304
rect 16908 6264 16914 6276
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 17310 6304 17316 6316
rect 17144 6276 17316 6304
rect 16025 6239 16083 6245
rect 16025 6205 16037 6239
rect 16071 6205 16083 6239
rect 16025 6199 16083 6205
rect 16040 6168 16068 6199
rect 16114 6196 16120 6248
rect 16172 6236 16178 6248
rect 16482 6236 16488 6248
rect 16172 6208 16217 6236
rect 16443 6208 16488 6236
rect 16172 6196 16178 6208
rect 16482 6196 16488 6208
rect 16540 6196 16546 6248
rect 16758 6196 16764 6248
rect 16816 6236 16822 6248
rect 17144 6245 17172 6276
rect 17310 6264 17316 6276
rect 17368 6264 17374 6316
rect 17129 6239 17187 6245
rect 17129 6236 17141 6239
rect 16816 6208 17141 6236
rect 16816 6196 16822 6208
rect 17129 6205 17141 6208
rect 17175 6205 17187 6239
rect 17129 6199 17187 6205
rect 17218 6196 17224 6248
rect 17276 6236 17282 6248
rect 17420 6236 17448 6344
rect 17865 6307 17923 6313
rect 17865 6273 17877 6307
rect 17911 6304 17923 6307
rect 18322 6304 18328 6316
rect 17911 6276 18328 6304
rect 17911 6273 17923 6276
rect 17865 6267 17923 6273
rect 18322 6264 18328 6276
rect 18380 6264 18386 6316
rect 18509 6307 18567 6313
rect 18509 6273 18521 6307
rect 18555 6304 18567 6307
rect 18598 6304 18604 6316
rect 18555 6276 18604 6304
rect 18555 6273 18567 6276
rect 18509 6267 18567 6273
rect 18598 6264 18604 6276
rect 18656 6264 18662 6316
rect 17957 6239 18015 6245
rect 17957 6236 17969 6239
rect 17276 6208 17321 6236
rect 17420 6208 17969 6236
rect 17276 6196 17282 6208
rect 17957 6205 17969 6208
rect 18003 6205 18015 6239
rect 17957 6199 18015 6205
rect 18049 6239 18107 6245
rect 18049 6205 18061 6239
rect 18095 6205 18107 6239
rect 18049 6199 18107 6205
rect 17034 6168 17040 6180
rect 16040 6140 17040 6168
rect 17034 6128 17040 6140
rect 17092 6128 17098 6180
rect 17310 6128 17316 6180
rect 17368 6168 17374 6180
rect 18064 6168 18092 6199
rect 17368 6140 18092 6168
rect 17368 6128 17374 6140
rect 16206 6100 16212 6112
rect 15948 6072 16212 6100
rect 16206 6060 16212 6072
rect 16264 6060 16270 6112
rect 17497 6103 17555 6109
rect 17497 6069 17509 6103
rect 17543 6100 17555 6103
rect 17678 6100 17684 6112
rect 17543 6072 17684 6100
rect 17543 6069 17555 6072
rect 17497 6063 17555 6069
rect 17678 6060 17684 6072
rect 17736 6060 17742 6112
rect 1104 6010 18860 6032
rect 1104 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 3430 6010
rect 3482 5958 7622 6010
rect 7674 5958 7686 6010
rect 7738 5958 7750 6010
rect 7802 5958 7814 6010
rect 7866 5958 7878 6010
rect 7930 5958 12070 6010
rect 12122 5958 12134 6010
rect 12186 5958 12198 6010
rect 12250 5958 12262 6010
rect 12314 5958 12326 6010
rect 12378 5958 16518 6010
rect 16570 5958 16582 6010
rect 16634 5958 16646 6010
rect 16698 5958 16710 6010
rect 16762 5958 16774 6010
rect 16826 5958 18860 6010
rect 1104 5936 18860 5958
rect 3878 5856 3884 5908
rect 3936 5896 3942 5908
rect 3936 5868 12388 5896
rect 3936 5856 3942 5868
rect 4062 5828 4068 5840
rect 1688 5800 4068 5828
rect 1688 5701 1716 5800
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 4341 5831 4399 5837
rect 4341 5797 4353 5831
rect 4387 5828 4399 5831
rect 4706 5828 4712 5840
rect 4387 5800 4712 5828
rect 4387 5797 4399 5800
rect 4341 5791 4399 5797
rect 4706 5788 4712 5800
rect 4764 5788 4770 5840
rect 5534 5788 5540 5840
rect 5592 5828 5598 5840
rect 6086 5828 6092 5840
rect 5592 5800 6092 5828
rect 5592 5788 5598 5800
rect 6086 5788 6092 5800
rect 6144 5788 6150 5840
rect 6822 5788 6828 5840
rect 6880 5828 6886 5840
rect 12360 5828 12388 5868
rect 12434 5856 12440 5908
rect 12492 5896 12498 5908
rect 13081 5899 13139 5905
rect 13081 5896 13093 5899
rect 12492 5868 13093 5896
rect 12492 5856 12498 5868
rect 13081 5865 13093 5868
rect 13127 5865 13139 5899
rect 15654 5896 15660 5908
rect 15615 5868 15660 5896
rect 13081 5859 13139 5865
rect 15654 5856 15660 5868
rect 15712 5856 15718 5908
rect 16206 5896 16212 5908
rect 16167 5868 16212 5896
rect 16206 5856 16212 5868
rect 16264 5856 16270 5908
rect 17034 5896 17040 5908
rect 16995 5868 17040 5896
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 18046 5896 18052 5908
rect 18007 5868 18052 5896
rect 18046 5856 18052 5868
rect 18104 5856 18110 5908
rect 18414 5896 18420 5908
rect 18375 5868 18420 5896
rect 18414 5856 18420 5868
rect 18472 5856 18478 5908
rect 13814 5828 13820 5840
rect 6880 5800 9352 5828
rect 12360 5800 13820 5828
rect 6880 5788 6886 5800
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5760 2283 5763
rect 2498 5760 2504 5772
rect 2271 5732 2504 5760
rect 2271 5729 2283 5732
rect 2225 5723 2283 5729
rect 2498 5720 2504 5732
rect 2556 5720 2562 5772
rect 2590 5720 2596 5772
rect 2648 5760 2654 5772
rect 3421 5763 3479 5769
rect 3421 5760 3433 5763
rect 2648 5732 3433 5760
rect 2648 5720 2654 5732
rect 3421 5729 3433 5732
rect 3467 5729 3479 5763
rect 3421 5723 3479 5729
rect 3694 5720 3700 5772
rect 3752 5760 3758 5772
rect 3973 5763 4031 5769
rect 3973 5760 3985 5763
rect 3752 5732 3985 5760
rect 3752 5720 3758 5732
rect 3973 5729 3985 5732
rect 4019 5760 4031 5763
rect 4154 5760 4160 5772
rect 4019 5732 4160 5760
rect 4019 5729 4031 5732
rect 3973 5723 4031 5729
rect 4154 5720 4160 5732
rect 4212 5720 4218 5772
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5661 1731 5695
rect 1673 5655 1731 5661
rect 1762 5652 1768 5704
rect 1820 5692 1826 5704
rect 2317 5695 2375 5701
rect 1820 5664 1865 5692
rect 1820 5652 1826 5664
rect 2317 5661 2329 5695
rect 2363 5692 2375 5695
rect 2363 5664 3648 5692
rect 2363 5661 2375 5664
rect 2317 5655 2375 5661
rect 3329 5627 3387 5633
rect 3329 5624 3341 5627
rect 2792 5596 3341 5624
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 1946 5556 1952 5568
rect 1907 5528 1952 5556
rect 1946 5516 1952 5528
rect 2004 5516 2010 5568
rect 2409 5559 2467 5565
rect 2409 5525 2421 5559
rect 2455 5556 2467 5559
rect 2498 5556 2504 5568
rect 2455 5528 2504 5556
rect 2455 5525 2467 5528
rect 2409 5519 2467 5525
rect 2498 5516 2504 5528
rect 2556 5516 2562 5568
rect 2792 5565 2820 5596
rect 3329 5593 3341 5596
rect 3375 5593 3387 5627
rect 3329 5587 3387 5593
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5525 2835 5559
rect 2777 5519 2835 5525
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 3234 5556 3240 5568
rect 2924 5528 2969 5556
rect 3195 5528 3240 5556
rect 2924 5516 2930 5528
rect 3234 5516 3240 5528
rect 3292 5516 3298 5568
rect 3620 5556 3648 5664
rect 4157 5627 4215 5633
rect 4157 5593 4169 5627
rect 4203 5624 4215 5627
rect 4522 5624 4528 5636
rect 4203 5596 4528 5624
rect 4203 5593 4215 5596
rect 4157 5587 4215 5593
rect 4522 5584 4528 5596
rect 4580 5584 4586 5636
rect 4724 5624 4752 5788
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5760 5135 5763
rect 5810 5760 5816 5772
rect 5123 5732 5816 5760
rect 5123 5729 5135 5732
rect 5077 5723 5135 5729
rect 5810 5720 5816 5732
rect 5868 5760 5874 5772
rect 7653 5763 7711 5769
rect 7653 5760 7665 5763
rect 5868 5732 7665 5760
rect 5868 5720 5874 5732
rect 7653 5729 7665 5732
rect 7699 5729 7711 5763
rect 7653 5723 7711 5729
rect 8757 5763 8815 5769
rect 8757 5729 8769 5763
rect 8803 5760 8815 5763
rect 8938 5760 8944 5772
rect 8803 5732 8944 5760
rect 8803 5729 8815 5732
rect 8757 5723 8815 5729
rect 8938 5720 8944 5732
rect 8996 5720 9002 5772
rect 7009 5695 7067 5701
rect 7009 5661 7021 5695
rect 7055 5692 7067 5695
rect 7098 5692 7104 5704
rect 7055 5664 7104 5692
rect 7055 5661 7067 5664
rect 7009 5655 7067 5661
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 7466 5652 7472 5704
rect 7524 5692 7530 5704
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 7524 5664 7941 5692
rect 7524 5652 7530 5664
rect 7929 5661 7941 5664
rect 7975 5661 7987 5695
rect 7929 5655 7987 5661
rect 6822 5624 6828 5636
rect 4724 5596 6828 5624
rect 6822 5584 6828 5596
rect 6880 5624 6886 5636
rect 6880 5596 7236 5624
rect 6880 5584 6886 5596
rect 4433 5559 4491 5565
rect 4433 5556 4445 5559
rect 3620 5528 4445 5556
rect 4433 5525 4445 5528
rect 4479 5525 4491 5559
rect 4433 5519 4491 5525
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 4801 5559 4859 5565
rect 4801 5556 4813 5559
rect 4672 5528 4813 5556
rect 4672 5516 4678 5528
rect 4801 5525 4813 5528
rect 4847 5525 4859 5559
rect 4801 5519 4859 5525
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 5721 5559 5779 5565
rect 4948 5528 4993 5556
rect 4948 5516 4954 5528
rect 5721 5525 5733 5559
rect 5767 5556 5779 5559
rect 6086 5556 6092 5568
rect 5767 5528 6092 5556
rect 5767 5525 5779 5528
rect 5721 5519 5779 5525
rect 6086 5516 6092 5528
rect 6144 5516 6150 5568
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 6730 5556 6736 5568
rect 6604 5528 6736 5556
rect 6604 5516 6610 5528
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 7098 5556 7104 5568
rect 7059 5528 7104 5556
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 7208 5556 7236 5596
rect 7650 5584 7656 5636
rect 7708 5624 7714 5636
rect 8573 5627 8631 5633
rect 8573 5624 8585 5627
rect 7708 5596 8585 5624
rect 7708 5584 7714 5596
rect 8573 5593 8585 5596
rect 8619 5593 8631 5627
rect 9324 5624 9352 5800
rect 13814 5788 13820 5800
rect 13872 5788 13878 5840
rect 10321 5763 10379 5769
rect 10321 5729 10333 5763
rect 10367 5760 10379 5763
rect 11146 5760 11152 5772
rect 10367 5732 11152 5760
rect 10367 5729 10379 5732
rect 10321 5723 10379 5729
rect 11146 5720 11152 5732
rect 11204 5720 11210 5772
rect 12710 5760 12716 5772
rect 12671 5732 12716 5760
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 12894 5760 12900 5772
rect 12855 5732 12900 5760
rect 12894 5720 12900 5732
rect 12952 5720 12958 5772
rect 13630 5760 13636 5772
rect 13591 5732 13636 5760
rect 13630 5720 13636 5732
rect 13688 5720 13694 5772
rect 15672 5760 15700 5856
rect 15930 5788 15936 5840
rect 15988 5828 15994 5840
rect 15988 5800 17724 5828
rect 15988 5788 15994 5800
rect 16761 5763 16819 5769
rect 16761 5760 16773 5763
rect 15672 5732 16773 5760
rect 16761 5729 16773 5732
rect 16807 5760 16819 5763
rect 17218 5760 17224 5772
rect 16807 5732 17224 5760
rect 16807 5729 16819 5732
rect 16761 5723 16819 5729
rect 17218 5720 17224 5732
rect 17276 5760 17282 5772
rect 17589 5763 17647 5769
rect 17589 5760 17601 5763
rect 17276 5732 17601 5760
rect 17276 5720 17282 5732
rect 17589 5729 17601 5732
rect 17635 5729 17647 5763
rect 17589 5723 17647 5729
rect 10065 5695 10123 5701
rect 10065 5661 10077 5695
rect 10111 5692 10123 5695
rect 10226 5692 10232 5704
rect 10111 5664 10232 5692
rect 10111 5661 10123 5664
rect 10065 5655 10123 5661
rect 10226 5652 10232 5664
rect 10284 5652 10290 5704
rect 10410 5692 10416 5704
rect 10371 5664 10416 5692
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 12161 5695 12219 5701
rect 12161 5661 12173 5695
rect 12207 5692 12219 5695
rect 14274 5692 14280 5704
rect 12207 5664 14280 5692
rect 12207 5661 12219 5664
rect 12161 5655 12219 5661
rect 14274 5652 14280 5664
rect 14332 5652 14338 5704
rect 14544 5695 14602 5701
rect 14544 5661 14556 5695
rect 14590 5661 14602 5695
rect 14544 5655 14602 5661
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5692 16175 5695
rect 16850 5692 16856 5704
rect 16163 5664 16856 5692
rect 16163 5661 16175 5664
rect 16117 5655 16175 5661
rect 11514 5624 11520 5636
rect 9324 5596 11520 5624
rect 8573 5587 8631 5593
rect 11514 5584 11520 5596
rect 11572 5584 11578 5636
rect 12618 5624 12624 5636
rect 12579 5596 12624 5624
rect 12618 5584 12624 5596
rect 12676 5584 12682 5636
rect 13446 5624 13452 5636
rect 13407 5596 13452 5624
rect 13446 5584 13452 5596
rect 13504 5584 13510 5636
rect 13541 5627 13599 5633
rect 13541 5593 13553 5627
rect 13587 5624 13599 5627
rect 13722 5624 13728 5636
rect 13587 5596 13728 5624
rect 13587 5593 13599 5596
rect 13541 5587 13599 5593
rect 13722 5584 13728 5596
rect 13780 5624 13786 5636
rect 13780 5596 14412 5624
rect 13780 5584 13786 5596
rect 7469 5559 7527 5565
rect 7469 5556 7481 5559
rect 7208 5528 7481 5556
rect 7469 5525 7481 5528
rect 7515 5525 7527 5559
rect 7469 5519 7527 5525
rect 7561 5559 7619 5565
rect 7561 5525 7573 5559
rect 7607 5556 7619 5559
rect 8202 5556 8208 5568
rect 7607 5528 8208 5556
rect 7607 5525 7619 5528
rect 7561 5519 7619 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 8941 5559 8999 5565
rect 8941 5525 8953 5559
rect 8987 5556 8999 5559
rect 10318 5556 10324 5568
rect 8987 5528 10324 5556
rect 8987 5525 8999 5528
rect 8941 5519 8999 5525
rect 10318 5516 10324 5528
rect 10376 5516 10382 5568
rect 11054 5516 11060 5568
rect 11112 5556 11118 5568
rect 12253 5559 12311 5565
rect 12253 5556 12265 5559
rect 11112 5528 12265 5556
rect 11112 5516 11118 5528
rect 12253 5525 12265 5528
rect 12299 5525 12311 5559
rect 12253 5519 12311 5525
rect 13998 5516 14004 5568
rect 14056 5556 14062 5568
rect 14093 5559 14151 5565
rect 14093 5556 14105 5559
rect 14056 5528 14105 5556
rect 14056 5516 14062 5528
rect 14093 5525 14105 5528
rect 14139 5525 14151 5559
rect 14384 5556 14412 5596
rect 14458 5584 14464 5636
rect 14516 5624 14522 5636
rect 14568 5624 14596 5655
rect 16850 5652 16856 5664
rect 16908 5652 16914 5704
rect 17405 5695 17463 5701
rect 17405 5661 17417 5695
rect 17451 5661 17463 5695
rect 17696 5692 17724 5800
rect 17770 5720 17776 5772
rect 17828 5760 17834 5772
rect 17828 5732 18276 5760
rect 17828 5720 17834 5732
rect 18248 5701 18276 5732
rect 17865 5695 17923 5701
rect 17865 5692 17877 5695
rect 17696 5664 17877 5692
rect 17405 5655 17463 5661
rect 17865 5661 17877 5664
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5661 18291 5695
rect 18233 5655 18291 5661
rect 17310 5624 17316 5636
rect 14516 5596 17316 5624
rect 14516 5584 14522 5596
rect 17310 5584 17316 5596
rect 17368 5584 17374 5636
rect 17420 5624 17448 5655
rect 17678 5624 17684 5636
rect 17420 5596 17684 5624
rect 17678 5584 17684 5596
rect 17736 5584 17742 5636
rect 15286 5556 15292 5568
rect 14384 5528 15292 5556
rect 14093 5519 14151 5525
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 15930 5556 15936 5568
rect 15891 5528 15936 5556
rect 15930 5516 15936 5528
rect 15988 5516 15994 5568
rect 16574 5556 16580 5568
rect 16535 5528 16580 5556
rect 16574 5516 16580 5528
rect 16632 5516 16638 5568
rect 16666 5516 16672 5568
rect 16724 5556 16730 5568
rect 16724 5528 16769 5556
rect 16724 5516 16730 5528
rect 17494 5516 17500 5568
rect 17552 5556 17558 5568
rect 17552 5528 17597 5556
rect 17552 5516 17558 5528
rect 1104 5466 18860 5488
rect 1104 5414 5398 5466
rect 5450 5414 5462 5466
rect 5514 5414 5526 5466
rect 5578 5414 5590 5466
rect 5642 5414 5654 5466
rect 5706 5414 9846 5466
rect 9898 5414 9910 5466
rect 9962 5414 9974 5466
rect 10026 5414 10038 5466
rect 10090 5414 10102 5466
rect 10154 5414 14294 5466
rect 14346 5414 14358 5466
rect 14410 5414 14422 5466
rect 14474 5414 14486 5466
rect 14538 5414 14550 5466
rect 14602 5414 18860 5466
rect 1104 5392 18860 5414
rect 1670 5312 1676 5364
rect 1728 5352 1734 5364
rect 2133 5355 2191 5361
rect 2133 5352 2145 5355
rect 1728 5324 2145 5352
rect 1728 5312 1734 5324
rect 2133 5321 2145 5324
rect 2179 5321 2191 5355
rect 2133 5315 2191 5321
rect 2314 5312 2320 5364
rect 2372 5352 2378 5364
rect 2409 5355 2467 5361
rect 2409 5352 2421 5355
rect 2372 5324 2421 5352
rect 2372 5312 2378 5324
rect 2409 5321 2421 5324
rect 2455 5321 2467 5355
rect 2409 5315 2467 5321
rect 3234 5312 3240 5364
rect 3292 5352 3298 5364
rect 5445 5355 5503 5361
rect 5445 5352 5457 5355
rect 3292 5324 5457 5352
rect 3292 5312 3298 5324
rect 5445 5321 5457 5324
rect 5491 5321 5503 5355
rect 5445 5315 5503 5321
rect 5813 5355 5871 5361
rect 5813 5321 5825 5355
rect 5859 5352 5871 5355
rect 6362 5352 6368 5364
rect 5859 5324 6368 5352
rect 5859 5321 5871 5324
rect 5813 5315 5871 5321
rect 6362 5312 6368 5324
rect 6420 5312 6426 5364
rect 6546 5312 6552 5364
rect 6604 5352 6610 5364
rect 8021 5355 8079 5361
rect 8021 5352 8033 5355
rect 6604 5324 8033 5352
rect 6604 5312 6610 5324
rect 8021 5321 8033 5324
rect 8067 5352 8079 5355
rect 8202 5352 8208 5364
rect 8067 5324 8208 5352
rect 8067 5321 8079 5324
rect 8021 5315 8079 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 9582 5312 9588 5364
rect 9640 5352 9646 5364
rect 9640 5324 11376 5352
rect 9640 5312 9646 5324
rect 4338 5284 4344 5296
rect 4299 5256 4344 5284
rect 4338 5244 4344 5256
rect 4396 5244 4402 5296
rect 4430 5244 4436 5296
rect 4488 5284 4494 5296
rect 5077 5287 5135 5293
rect 5077 5284 5089 5287
rect 4488 5256 5089 5284
rect 4488 5244 4494 5256
rect 5077 5253 5089 5256
rect 5123 5253 5135 5287
rect 5994 5284 6000 5296
rect 5077 5247 5135 5253
rect 5644 5256 6000 5284
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 1762 5216 1768 5228
rect 1719 5188 1768 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 1762 5176 1768 5188
rect 1820 5176 1826 5228
rect 2038 5216 2044 5228
rect 1999 5188 2044 5216
rect 2038 5176 2044 5188
rect 2096 5176 2102 5228
rect 2314 5216 2320 5228
rect 2275 5188 2320 5216
rect 2314 5176 2320 5188
rect 2372 5176 2378 5228
rect 4525 5219 4583 5225
rect 4525 5185 4537 5219
rect 4571 5216 4583 5219
rect 4985 5219 5043 5225
rect 4985 5216 4997 5219
rect 4571 5188 4997 5216
rect 4571 5185 4583 5188
rect 4525 5179 4583 5185
rect 4985 5185 4997 5188
rect 5031 5216 5043 5219
rect 5644 5216 5672 5256
rect 5994 5244 6000 5256
rect 6052 5244 6058 5296
rect 6086 5244 6092 5296
rect 6144 5284 6150 5296
rect 6144 5256 8156 5284
rect 6144 5244 6150 5256
rect 5031 5188 5672 5216
rect 5031 5185 5043 5188
rect 4985 5179 5043 5185
rect 5718 5176 5724 5228
rect 5776 5216 5782 5228
rect 6472 5225 6500 5256
rect 8128 5228 8156 5256
rect 8478 5244 8484 5296
rect 8536 5284 8542 5296
rect 11054 5284 11060 5296
rect 8536 5256 11060 5284
rect 8536 5244 8542 5256
rect 11054 5244 11060 5256
rect 11112 5244 11118 5296
rect 11348 5284 11376 5324
rect 11422 5312 11428 5364
rect 11480 5352 11486 5364
rect 13081 5355 13139 5361
rect 13081 5352 13093 5355
rect 11480 5324 13093 5352
rect 11480 5312 11486 5324
rect 13081 5321 13093 5324
rect 13127 5321 13139 5355
rect 13081 5315 13139 5321
rect 14090 5312 14096 5364
rect 14148 5352 14154 5364
rect 14826 5352 14832 5364
rect 14148 5324 14832 5352
rect 14148 5312 14154 5324
rect 14826 5312 14832 5324
rect 14884 5352 14890 5364
rect 14884 5324 15875 5352
rect 14884 5312 14890 5324
rect 12943 5287 13001 5293
rect 11348 5256 12388 5284
rect 6457 5219 6515 5225
rect 5776 5188 6040 5216
rect 5776 5176 5782 5188
rect 1854 5108 1860 5160
rect 1912 5148 1918 5160
rect 2406 5148 2412 5160
rect 1912 5120 2412 5148
rect 1912 5108 1918 5120
rect 2406 5108 2412 5120
rect 2464 5108 2470 5160
rect 2590 5148 2596 5160
rect 2551 5120 2596 5148
rect 2590 5108 2596 5120
rect 2648 5108 2654 5160
rect 5258 5148 5264 5160
rect 5219 5120 5264 5148
rect 5258 5108 5264 5120
rect 5316 5108 5322 5160
rect 6012 5157 6040 5188
rect 6457 5185 6469 5219
rect 6503 5185 6515 5219
rect 6457 5179 6515 5185
rect 6724 5219 6782 5225
rect 6724 5185 6736 5219
rect 6770 5216 6782 5219
rect 6770 5188 7604 5216
rect 6770 5185 6782 5188
rect 6724 5179 6782 5185
rect 5905 5151 5963 5157
rect 5905 5117 5917 5151
rect 5951 5117 5963 5151
rect 5905 5111 5963 5117
rect 5997 5151 6055 5157
rect 5997 5117 6009 5151
rect 6043 5117 6055 5151
rect 7576 5148 7604 5188
rect 8110 5176 8116 5228
rect 8168 5216 8174 5228
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 8168 5188 8309 5216
rect 8168 5176 8174 5188
rect 8297 5185 8309 5188
rect 8343 5185 8355 5219
rect 8297 5179 8355 5185
rect 8386 5176 8392 5228
rect 8444 5176 8450 5228
rect 8564 5219 8622 5225
rect 8564 5185 8576 5219
rect 8610 5216 8622 5219
rect 8938 5216 8944 5228
rect 8610 5188 8944 5216
rect 8610 5185 8622 5188
rect 8564 5179 8622 5185
rect 8938 5176 8944 5188
rect 8996 5176 9002 5228
rect 10229 5219 10287 5225
rect 10229 5185 10241 5219
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 8404 5148 8432 5176
rect 7576 5120 8432 5148
rect 10244 5148 10272 5179
rect 10318 5176 10324 5228
rect 10376 5216 10382 5228
rect 11149 5219 11207 5225
rect 10376 5188 10421 5216
rect 10376 5176 10382 5188
rect 11149 5185 11161 5219
rect 11195 5216 11207 5219
rect 11422 5216 11428 5228
rect 11195 5188 11428 5216
rect 11195 5185 11207 5188
rect 11149 5179 11207 5185
rect 11422 5176 11428 5188
rect 11480 5176 11486 5228
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5216 11575 5219
rect 11698 5216 11704 5228
rect 11563 5188 11704 5216
rect 11563 5185 11575 5188
rect 11517 5179 11575 5185
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 11793 5219 11851 5225
rect 11793 5185 11805 5219
rect 11839 5216 11851 5219
rect 12253 5219 12311 5225
rect 11839 5188 12204 5216
rect 11839 5185 11851 5188
rect 11793 5179 11851 5185
rect 10502 5148 10508 5160
rect 10244 5120 10508 5148
rect 5997 5111 6055 5117
rect 1486 5080 1492 5092
rect 1447 5052 1492 5080
rect 1486 5040 1492 5052
rect 1544 5040 1550 5092
rect 2774 5040 2780 5092
rect 2832 5080 2838 5092
rect 4154 5080 4160 5092
rect 2832 5052 4160 5080
rect 2832 5040 2838 5052
rect 4154 5040 4160 5052
rect 4212 5080 4218 5092
rect 5166 5080 5172 5092
rect 4212 5052 5172 5080
rect 4212 5040 4218 5052
rect 5166 5040 5172 5052
rect 5224 5040 5230 5092
rect 1854 5012 1860 5024
rect 1815 4984 1860 5012
rect 1854 4972 1860 4984
rect 1912 4972 1918 5024
rect 3050 4972 3056 5024
rect 3108 5012 3114 5024
rect 4062 5012 4068 5024
rect 3108 4984 4068 5012
rect 3108 4972 3114 4984
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4522 4972 4528 5024
rect 4580 5012 4586 5024
rect 4617 5015 4675 5021
rect 4617 5012 4629 5015
rect 4580 4984 4629 5012
rect 4580 4972 4586 4984
rect 4617 4981 4629 4984
rect 4663 4981 4675 5015
rect 5920 5012 5948 5111
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 11606 5108 11612 5160
rect 11664 5148 11670 5160
rect 12069 5151 12127 5157
rect 12069 5148 12081 5151
rect 11664 5120 12081 5148
rect 11664 5108 11670 5120
rect 12069 5117 12081 5120
rect 12115 5117 12127 5151
rect 12176 5148 12204 5188
rect 12253 5185 12265 5219
rect 12299 5216 12311 5219
rect 12360 5216 12388 5256
rect 12943 5253 12955 5287
rect 12989 5284 13001 5287
rect 13449 5287 13507 5293
rect 13449 5284 13461 5287
rect 12989 5256 13461 5284
rect 12989 5253 13001 5256
rect 12943 5247 13001 5253
rect 13449 5253 13461 5256
rect 13495 5253 13507 5287
rect 13449 5247 13507 5253
rect 15010 5244 15016 5296
rect 15068 5284 15074 5296
rect 15105 5287 15163 5293
rect 15105 5284 15117 5287
rect 15068 5256 15117 5284
rect 15068 5244 15074 5256
rect 15105 5253 15117 5256
rect 15151 5253 15163 5287
rect 15105 5247 15163 5253
rect 12840 5219 12898 5225
rect 12840 5216 12852 5219
rect 12299 5188 12852 5216
rect 12299 5185 12311 5188
rect 12253 5179 12311 5185
rect 12840 5185 12852 5188
rect 12886 5185 12898 5219
rect 14734 5216 14740 5228
rect 12840 5179 12898 5185
rect 14660 5188 14740 5216
rect 12176 5120 13170 5148
rect 12069 5111 12127 5117
rect 7558 5040 7564 5092
rect 7616 5080 7622 5092
rect 8113 5083 8171 5089
rect 8113 5080 8125 5083
rect 7616 5052 8125 5080
rect 7616 5040 7622 5052
rect 8113 5049 8125 5052
rect 8159 5049 8171 5083
rect 8113 5043 8171 5049
rect 9677 5083 9735 5089
rect 9677 5049 9689 5083
rect 9723 5080 9735 5083
rect 11701 5083 11759 5089
rect 9723 5052 10180 5080
rect 9723 5049 9735 5052
rect 9677 5043 9735 5049
rect 7098 5012 7104 5024
rect 5920 4984 7104 5012
rect 4617 4975 4675 4981
rect 7098 4972 7104 4984
rect 7156 4972 7162 5024
rect 7466 4972 7472 5024
rect 7524 5012 7530 5024
rect 7837 5015 7895 5021
rect 7837 5012 7849 5015
rect 7524 4984 7849 5012
rect 7524 4972 7530 4984
rect 7837 4981 7849 4984
rect 7883 4981 7895 5015
rect 7837 4975 7895 4981
rect 9030 4972 9036 5024
rect 9088 5012 9094 5024
rect 9582 5012 9588 5024
rect 9088 4984 9588 5012
rect 9088 4972 9094 4984
rect 9582 4972 9588 4984
rect 9640 5012 9646 5024
rect 10152 5021 10180 5052
rect 11701 5049 11713 5083
rect 11747 5080 11759 5083
rect 12618 5080 12624 5092
rect 11747 5052 12624 5080
rect 11747 5049 11759 5052
rect 11701 5043 11759 5049
rect 12618 5040 12624 5052
rect 12676 5040 12682 5092
rect 9769 5015 9827 5021
rect 9769 5012 9781 5015
rect 9640 4984 9781 5012
rect 9640 4972 9646 4984
rect 9769 4981 9781 4984
rect 9815 4981 9827 5015
rect 9769 4975 9827 4981
rect 10137 5015 10195 5021
rect 10137 4981 10149 5015
rect 10183 5012 10195 5015
rect 10686 5012 10692 5024
rect 10183 4984 10692 5012
rect 10183 4981 10195 4984
rect 10137 4975 10195 4981
rect 10686 4972 10692 4984
rect 10744 4972 10750 5024
rect 10962 5012 10968 5024
rect 10923 4984 10968 5012
rect 10962 4972 10968 4984
rect 11020 4972 11026 5024
rect 11330 5012 11336 5024
rect 11291 4984 11336 5012
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 11977 5015 12035 5021
rect 11977 4981 11989 5015
rect 12023 5012 12035 5015
rect 12434 5012 12440 5024
rect 12023 4984 12440 5012
rect 12023 4981 12035 4984
rect 11977 4975 12035 4981
rect 12434 4972 12440 4984
rect 12492 4972 12498 5024
rect 12710 5012 12716 5024
rect 12671 4984 12716 5012
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 13142 5012 13170 5120
rect 13262 5108 13268 5160
rect 13320 5148 13326 5160
rect 13320 5120 13365 5148
rect 13320 5108 13326 5120
rect 13814 5108 13820 5160
rect 13872 5148 13878 5160
rect 14660 5148 14688 5188
rect 14734 5176 14740 5188
rect 14792 5216 14798 5228
rect 15654 5225 15660 5228
rect 15197 5219 15255 5225
rect 15197 5216 15209 5219
rect 14792 5188 15209 5216
rect 14792 5176 14798 5188
rect 15197 5185 15209 5188
rect 15243 5185 15255 5219
rect 15197 5179 15255 5185
rect 15622 5219 15660 5225
rect 15622 5185 15634 5219
rect 15622 5179 15660 5185
rect 15654 5176 15660 5179
rect 15712 5176 15718 5228
rect 15847 5216 15875 5324
rect 16298 5312 16304 5364
rect 16356 5312 16362 5364
rect 16666 5312 16672 5364
rect 16724 5352 16730 5364
rect 16761 5355 16819 5361
rect 16761 5352 16773 5355
rect 16724 5324 16773 5352
rect 16724 5312 16730 5324
rect 16761 5321 16773 5324
rect 16807 5321 16819 5355
rect 17126 5352 17132 5364
rect 17087 5324 17132 5352
rect 16761 5315 16819 5321
rect 17126 5312 17132 5324
rect 17184 5312 17190 5364
rect 17494 5312 17500 5364
rect 17552 5352 17558 5364
rect 17589 5355 17647 5361
rect 17589 5352 17601 5355
rect 17552 5324 17601 5352
rect 17552 5312 17558 5324
rect 17589 5321 17601 5324
rect 17635 5321 17647 5355
rect 17589 5315 17647 5321
rect 17957 5355 18015 5361
rect 17957 5321 17969 5355
rect 18003 5352 18015 5355
rect 18506 5352 18512 5364
rect 18003 5324 18512 5352
rect 18003 5321 18015 5324
rect 17957 5315 18015 5321
rect 18506 5312 18512 5324
rect 18564 5312 18570 5364
rect 15933 5219 15991 5225
rect 15933 5216 15945 5219
rect 15847 5188 15945 5216
rect 15933 5185 15945 5188
rect 15979 5185 15991 5219
rect 15933 5179 15991 5185
rect 16025 5219 16083 5225
rect 16025 5185 16037 5219
rect 16071 5216 16083 5219
rect 16206 5216 16212 5228
rect 16071 5188 16212 5216
rect 16071 5185 16083 5188
rect 16025 5179 16083 5185
rect 16206 5176 16212 5188
rect 16264 5176 16270 5228
rect 16316 5225 16344 5312
rect 17310 5244 17316 5296
rect 17368 5284 17374 5296
rect 17368 5256 18184 5284
rect 17368 5244 17374 5256
rect 16301 5219 16359 5225
rect 16301 5185 16313 5219
rect 16347 5185 16359 5219
rect 16301 5179 16359 5185
rect 17221 5219 17279 5225
rect 17221 5185 17233 5219
rect 17267 5216 17279 5219
rect 17862 5216 17868 5228
rect 17267 5188 17868 5216
rect 17267 5185 17279 5188
rect 17221 5179 17279 5185
rect 17862 5176 17868 5188
rect 17920 5176 17926 5228
rect 13872 5120 14688 5148
rect 13872 5108 13878 5120
rect 14918 5108 14924 5160
rect 14976 5148 14982 5160
rect 14976 5120 16160 5148
rect 14976 5108 14982 5120
rect 15286 5040 15292 5092
rect 15344 5080 15350 5092
rect 15749 5083 15807 5089
rect 15749 5080 15761 5083
rect 15344 5052 15761 5080
rect 15344 5040 15350 5052
rect 15749 5049 15761 5052
rect 15795 5049 15807 5083
rect 15749 5043 15807 5049
rect 13998 5012 14004 5024
rect 13142 4984 14004 5012
rect 13998 4972 14004 4984
rect 14056 4972 14062 5024
rect 15378 5012 15384 5024
rect 15339 4984 15384 5012
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 15470 4972 15476 5024
rect 15528 5021 15534 5024
rect 15528 5015 15577 5021
rect 15528 4981 15531 5015
rect 15565 4981 15577 5015
rect 16132 5012 16160 5120
rect 17310 5108 17316 5160
rect 17368 5148 17374 5160
rect 18046 5148 18052 5160
rect 17368 5120 17413 5148
rect 18007 5120 18052 5148
rect 17368 5108 17374 5120
rect 18046 5108 18052 5120
rect 18104 5108 18110 5160
rect 18156 5157 18184 5256
rect 18509 5219 18567 5225
rect 18509 5185 18521 5219
rect 18555 5216 18567 5219
rect 18782 5216 18788 5228
rect 18555 5188 18788 5216
rect 18555 5185 18567 5188
rect 18509 5179 18567 5185
rect 18782 5176 18788 5188
rect 18840 5176 18846 5228
rect 18141 5151 18199 5157
rect 18141 5117 18153 5151
rect 18187 5117 18199 5151
rect 18141 5111 18199 5117
rect 16209 5083 16267 5089
rect 16209 5049 16221 5083
rect 16255 5080 16267 5083
rect 18230 5080 18236 5092
rect 16255 5052 18236 5080
rect 16255 5049 16267 5052
rect 16209 5043 16267 5049
rect 18230 5040 18236 5052
rect 18288 5040 18294 5092
rect 16298 5012 16304 5024
rect 16132 4984 16304 5012
rect 15528 4975 15577 4981
rect 15528 4972 15534 4975
rect 16298 4972 16304 4984
rect 16356 4972 16362 5024
rect 16485 5015 16543 5021
rect 16485 4981 16497 5015
rect 16531 5012 16543 5015
rect 18138 5012 18144 5024
rect 16531 4984 18144 5012
rect 16531 4981 16543 4984
rect 16485 4975 16543 4981
rect 18138 4972 18144 4984
rect 18196 4972 18202 5024
rect 1104 4922 18860 4944
rect 1104 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 3430 4922
rect 3482 4870 7622 4922
rect 7674 4870 7686 4922
rect 7738 4870 7750 4922
rect 7802 4870 7814 4922
rect 7866 4870 7878 4922
rect 7930 4870 12070 4922
rect 12122 4870 12134 4922
rect 12186 4870 12198 4922
rect 12250 4870 12262 4922
rect 12314 4870 12326 4922
rect 12378 4870 16518 4922
rect 16570 4870 16582 4922
rect 16634 4870 16646 4922
rect 16698 4870 16710 4922
rect 16762 4870 16774 4922
rect 16826 4870 18860 4922
rect 1104 4848 18860 4870
rect 1762 4808 1768 4820
rect 1723 4780 1768 4808
rect 1762 4768 1768 4780
rect 1820 4768 1826 4820
rect 2038 4808 2044 4820
rect 1999 4780 2044 4808
rect 2038 4768 2044 4780
rect 2096 4768 2102 4820
rect 3605 4811 3663 4817
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 3694 4808 3700 4820
rect 3651 4780 3700 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 3694 4768 3700 4780
rect 3752 4768 3758 4820
rect 4062 4808 4068 4820
rect 4023 4780 4068 4808
rect 4062 4768 4068 4780
rect 4120 4768 4126 4820
rect 4430 4808 4436 4820
rect 4391 4780 4436 4808
rect 4430 4768 4436 4780
rect 4488 4768 4494 4820
rect 4525 4811 4583 4817
rect 4525 4777 4537 4811
rect 4571 4808 4583 4811
rect 4890 4808 4896 4820
rect 4571 4780 4896 4808
rect 4571 4777 4583 4780
rect 4525 4771 4583 4777
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 8478 4808 8484 4820
rect 5000 4780 8484 4808
rect 5000 4740 5028 4780
rect 8478 4768 8484 4780
rect 8536 4768 8542 4820
rect 8938 4808 8944 4820
rect 8899 4780 8944 4808
rect 8938 4768 8944 4780
rect 8996 4768 9002 4820
rect 9674 4808 9680 4820
rect 9635 4780 9680 4808
rect 9674 4768 9680 4780
rect 9732 4768 9738 4820
rect 10778 4768 10784 4820
rect 10836 4808 10842 4820
rect 11517 4811 11575 4817
rect 11517 4808 11529 4811
rect 10836 4780 11529 4808
rect 10836 4768 10842 4780
rect 11517 4777 11529 4780
rect 11563 4777 11575 4811
rect 11517 4771 11575 4777
rect 2884 4712 5028 4740
rect 6917 4743 6975 4749
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4573 1731 4607
rect 1673 4567 1731 4573
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4604 2007 4607
rect 2038 4604 2044 4616
rect 1995 4576 2044 4604
rect 1995 4573 2007 4576
rect 1949 4567 2007 4573
rect 1688 4536 1716 4567
rect 2038 4564 2044 4576
rect 2096 4564 2102 4616
rect 2222 4604 2228 4616
rect 2183 4576 2228 4604
rect 2222 4564 2228 4576
rect 2280 4564 2286 4616
rect 2501 4607 2559 4613
rect 2501 4573 2513 4607
rect 2547 4604 2559 4607
rect 2774 4604 2780 4616
rect 2547 4576 2780 4604
rect 2547 4573 2559 4576
rect 2501 4567 2559 4573
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 2884 4613 2912 4712
rect 6917 4709 6929 4743
rect 6963 4740 6975 4743
rect 7282 4740 7288 4752
rect 6963 4712 7288 4740
rect 6963 4709 6975 4712
rect 6917 4703 6975 4709
rect 7282 4700 7288 4712
rect 7340 4700 7346 4752
rect 2958 4632 2964 4684
rect 3016 4672 3022 4684
rect 4982 4672 4988 4684
rect 3016 4644 3280 4672
rect 4943 4644 4988 4672
rect 3016 4632 3022 4644
rect 2869 4607 2927 4613
rect 2869 4573 2881 4607
rect 2915 4573 2927 4607
rect 2869 4567 2927 4573
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4573 3203 4607
rect 3252 4604 3280 4644
rect 4982 4632 4988 4644
rect 5040 4632 5046 4684
rect 5169 4675 5227 4681
rect 5169 4641 5181 4675
rect 5215 4672 5227 4675
rect 5258 4672 5264 4684
rect 5215 4644 5264 4672
rect 5215 4641 5227 4644
rect 5169 4635 5227 4641
rect 5258 4632 5264 4644
rect 5316 4632 5322 4684
rect 3397 4607 3455 4613
rect 3397 4604 3409 4607
rect 3252 4576 3409 4604
rect 3145 4567 3203 4573
rect 3397 4573 3409 4576
rect 3443 4573 3455 4607
rect 3397 4567 3455 4573
rect 3160 4536 3188 4567
rect 4706 4564 4712 4616
rect 4764 4604 4770 4616
rect 4893 4607 4951 4613
rect 4893 4604 4905 4607
rect 4764 4576 4905 4604
rect 4764 4564 4770 4576
rect 4893 4573 4905 4576
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 5353 4607 5411 4613
rect 5353 4573 5365 4607
rect 5399 4604 5411 4607
rect 6086 4604 6092 4616
rect 5399 4576 6092 4604
rect 5399 4573 5411 4576
rect 5353 4567 5411 4573
rect 6086 4564 6092 4576
rect 6144 4564 6150 4616
rect 6914 4564 6920 4616
rect 6972 4564 6978 4616
rect 7193 4607 7251 4613
rect 7193 4573 7205 4607
rect 7239 4604 7251 4607
rect 7282 4604 7288 4616
rect 7239 4576 7288 4604
rect 7239 4573 7251 4576
rect 7193 4567 7251 4573
rect 7282 4564 7288 4576
rect 7340 4564 7346 4616
rect 7377 4607 7435 4613
rect 7377 4573 7389 4607
rect 7423 4604 7435 4607
rect 8110 4604 8116 4616
rect 7423 4576 8116 4604
rect 7423 4573 7435 4576
rect 7377 4567 7435 4573
rect 8110 4564 8116 4576
rect 8168 4564 8174 4616
rect 9122 4604 9128 4616
rect 8772 4576 9128 4604
rect 3881 4539 3939 4545
rect 3881 4536 3893 4539
rect 1688 4508 2820 4536
rect 3160 4508 3893 4536
rect 2792 4480 2820 4508
rect 3881 4505 3893 4508
rect 3927 4536 3939 4539
rect 3927 4508 5212 4536
rect 3927 4505 3939 4508
rect 3881 4499 3939 4505
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 2317 4471 2375 4477
rect 2317 4437 2329 4471
rect 2363 4468 2375 4471
rect 2406 4468 2412 4480
rect 2363 4440 2412 4468
rect 2363 4437 2375 4440
rect 2317 4431 2375 4437
rect 2406 4428 2412 4440
rect 2464 4428 2470 4480
rect 2682 4468 2688 4480
rect 2643 4440 2688 4468
rect 2682 4428 2688 4440
rect 2740 4428 2746 4480
rect 2774 4428 2780 4480
rect 2832 4428 2838 4480
rect 2958 4468 2964 4480
rect 2919 4440 2964 4468
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 3050 4428 3056 4480
rect 3108 4468 3114 4480
rect 3237 4471 3295 4477
rect 3237 4468 3249 4471
rect 3108 4440 3249 4468
rect 3108 4428 3114 4440
rect 3237 4437 3249 4440
rect 3283 4437 3295 4471
rect 4154 4468 4160 4480
rect 4115 4440 4160 4468
rect 3237 4431 3295 4437
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 5184 4468 5212 4508
rect 5258 4496 5264 4548
rect 5316 4536 5322 4548
rect 5598 4539 5656 4545
rect 5598 4536 5610 4539
rect 5316 4508 5610 4536
rect 5316 4496 5322 4508
rect 5598 4505 5610 4508
rect 5644 4505 5656 4539
rect 6932 4536 6960 4564
rect 5598 4499 5656 4505
rect 5727 4508 6960 4536
rect 7644 4539 7702 4545
rect 5727 4468 5755 4508
rect 7644 4505 7656 4539
rect 7690 4536 7702 4539
rect 8570 4536 8576 4548
rect 7690 4508 8576 4536
rect 7690 4505 7702 4508
rect 7644 4499 7702 4505
rect 8570 4496 8576 4508
rect 8628 4496 8634 4548
rect 5184 4440 5755 4468
rect 5810 4428 5816 4480
rect 5868 4468 5874 4480
rect 6733 4471 6791 4477
rect 6733 4468 6745 4471
rect 5868 4440 6745 4468
rect 5868 4428 5874 4440
rect 6733 4437 6745 4440
rect 6779 4437 6791 4471
rect 6733 4431 6791 4437
rect 6914 4428 6920 4480
rect 6972 4468 6978 4480
rect 8772 4477 8800 4576
rect 9122 4564 9128 4576
rect 9180 4604 9186 4616
rect 9585 4607 9643 4613
rect 9585 4604 9597 4607
rect 9180 4576 9597 4604
rect 9180 4564 9186 4576
rect 9585 4573 9597 4576
rect 9631 4573 9643 4607
rect 9585 4567 9643 4573
rect 9674 4564 9680 4616
rect 9732 4604 9738 4616
rect 9861 4607 9919 4613
rect 9861 4604 9873 4607
rect 9732 4576 9873 4604
rect 9732 4564 9738 4576
rect 9861 4573 9873 4576
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 10137 4607 10195 4613
rect 10137 4573 10149 4607
rect 10183 4604 10195 4607
rect 11146 4604 11152 4616
rect 10183 4576 11152 4604
rect 10183 4573 10195 4576
rect 10137 4567 10195 4573
rect 11146 4564 11152 4576
rect 11204 4564 11210 4616
rect 11532 4604 11560 4771
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 13446 4808 13452 4820
rect 12676 4780 13452 4808
rect 12676 4768 12682 4780
rect 13446 4768 13452 4780
rect 13504 4768 13510 4820
rect 13541 4811 13599 4817
rect 13541 4777 13553 4811
rect 13587 4808 13599 4811
rect 17126 4808 17132 4820
rect 13587 4780 17132 4808
rect 13587 4777 13599 4780
rect 13541 4771 13599 4777
rect 17126 4768 17132 4780
rect 17184 4768 17190 4820
rect 18414 4808 18420 4820
rect 18375 4780 18420 4808
rect 18414 4768 18420 4780
rect 18472 4768 18478 4820
rect 11790 4700 11796 4752
rect 11848 4740 11854 4752
rect 13722 4740 13728 4752
rect 11848 4712 13728 4740
rect 11848 4700 11854 4712
rect 13722 4700 13728 4712
rect 13780 4700 13786 4752
rect 13817 4743 13875 4749
rect 13817 4709 13829 4743
rect 13863 4740 13875 4743
rect 18138 4740 18144 4752
rect 13863 4712 18144 4740
rect 13863 4709 13875 4712
rect 13817 4703 13875 4709
rect 18138 4700 18144 4712
rect 18196 4700 18202 4752
rect 11882 4632 11888 4684
rect 11940 4672 11946 4684
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 11940 4644 12357 4672
rect 11940 4632 11946 4644
rect 12345 4641 12357 4644
rect 12391 4641 12403 4675
rect 12345 4635 12403 4641
rect 12434 4632 12440 4684
rect 12492 4672 12498 4684
rect 14185 4675 14243 4681
rect 14185 4672 14197 4675
rect 12492 4644 14197 4672
rect 12492 4632 12498 4644
rect 14185 4641 14197 4644
rect 14231 4641 14243 4675
rect 14185 4635 14243 4641
rect 15378 4632 15384 4684
rect 15436 4672 15442 4684
rect 16117 4675 16175 4681
rect 16117 4672 16129 4675
rect 15436 4644 16129 4672
rect 15436 4632 15442 4644
rect 16117 4641 16129 4644
rect 16163 4641 16175 4675
rect 16298 4672 16304 4684
rect 16259 4644 16304 4672
rect 16117 4635 16175 4641
rect 16298 4632 16304 4644
rect 16356 4632 16362 4684
rect 16850 4672 16856 4684
rect 16811 4644 16856 4672
rect 16850 4632 16856 4644
rect 16908 4632 16914 4684
rect 18049 4675 18107 4681
rect 18049 4641 18061 4675
rect 18095 4672 18107 4675
rect 18690 4672 18696 4684
rect 18095 4644 18696 4672
rect 18095 4641 18107 4644
rect 18049 4635 18107 4641
rect 18690 4632 18696 4644
rect 18748 4632 18754 4684
rect 11609 4607 11667 4613
rect 11609 4604 11621 4607
rect 11532 4576 11621 4604
rect 11609 4573 11621 4576
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 12250 4564 12256 4616
rect 12308 4604 12314 4616
rect 12529 4607 12587 4613
rect 12529 4604 12541 4607
rect 12308 4576 12541 4604
rect 12308 4564 12314 4576
rect 12529 4573 12541 4576
rect 12575 4573 12587 4607
rect 12529 4567 12587 4573
rect 12710 4564 12716 4616
rect 12768 4604 12774 4616
rect 13081 4607 13139 4613
rect 13081 4604 13093 4607
rect 12768 4576 13093 4604
rect 12768 4564 12774 4576
rect 13081 4573 13093 4576
rect 13127 4573 13139 4607
rect 13081 4567 13139 4573
rect 13170 4564 13176 4616
rect 13228 4604 13234 4616
rect 13357 4607 13415 4613
rect 13357 4604 13369 4607
rect 13228 4576 13369 4604
rect 13228 4564 13234 4576
rect 13357 4573 13369 4576
rect 13403 4573 13415 4607
rect 13630 4604 13636 4616
rect 13591 4576 13636 4604
rect 13357 4567 13415 4573
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 16022 4604 16028 4616
rect 15983 4576 16028 4604
rect 16022 4564 16028 4576
rect 16080 4564 16086 4616
rect 18233 4607 18291 4613
rect 18233 4573 18245 4607
rect 18279 4604 18291 4607
rect 18322 4604 18328 4616
rect 18279 4576 18328 4604
rect 18279 4573 18291 4576
rect 18233 4567 18291 4573
rect 18322 4564 18328 4576
rect 18380 4564 18386 4616
rect 10404 4539 10462 4545
rect 10404 4505 10416 4539
rect 10450 4536 10462 4539
rect 10962 4536 10968 4548
rect 10450 4508 10968 4536
rect 10450 4505 10462 4508
rect 10404 4499 10462 4505
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 14369 4539 14427 4545
rect 13280 4508 14320 4536
rect 7009 4471 7067 4477
rect 7009 4468 7021 4471
rect 6972 4440 7021 4468
rect 6972 4428 6978 4440
rect 7009 4437 7021 4440
rect 7055 4437 7067 4471
rect 7009 4431 7067 4437
rect 8757 4471 8815 4477
rect 8757 4437 8769 4471
rect 8803 4437 8815 4471
rect 8757 4431 8815 4437
rect 10045 4471 10103 4477
rect 10045 4437 10057 4471
rect 10091 4468 10103 4471
rect 10870 4468 10876 4480
rect 10091 4440 10876 4468
rect 10091 4437 10103 4440
rect 10045 4431 10103 4437
rect 10870 4428 10876 4440
rect 10928 4428 10934 4480
rect 11882 4428 11888 4480
rect 11940 4468 11946 4480
rect 12253 4471 12311 4477
rect 12253 4468 12265 4471
rect 11940 4440 12265 4468
rect 11940 4428 11946 4440
rect 12253 4437 12265 4440
rect 12299 4437 12311 4471
rect 12253 4431 12311 4437
rect 12989 4471 13047 4477
rect 12989 4437 13001 4471
rect 13035 4468 13047 4471
rect 13170 4468 13176 4480
rect 13035 4440 13176 4468
rect 13035 4437 13047 4440
rect 12989 4431 13047 4437
rect 13170 4428 13176 4440
rect 13228 4428 13234 4480
rect 13280 4477 13308 4508
rect 13265 4471 13323 4477
rect 13265 4437 13277 4471
rect 13311 4437 13323 4471
rect 14292 4468 14320 4508
rect 14369 4505 14381 4539
rect 14415 4536 14427 4539
rect 15102 4536 15108 4548
rect 14415 4508 15108 4536
rect 14415 4505 14427 4508
rect 14369 4499 14427 4505
rect 15102 4496 15108 4508
rect 15160 4496 15166 4548
rect 15378 4468 15384 4480
rect 14292 4440 15384 4468
rect 13265 4431 13323 4437
rect 15378 4428 15384 4440
rect 15436 4428 15442 4480
rect 1104 4378 18860 4400
rect 1104 4326 5398 4378
rect 5450 4326 5462 4378
rect 5514 4326 5526 4378
rect 5578 4326 5590 4378
rect 5642 4326 5654 4378
rect 5706 4326 9846 4378
rect 9898 4326 9910 4378
rect 9962 4326 9974 4378
rect 10026 4326 10038 4378
rect 10090 4326 10102 4378
rect 10154 4326 14294 4378
rect 14346 4326 14358 4378
rect 14410 4326 14422 4378
rect 14474 4326 14486 4378
rect 14538 4326 14550 4378
rect 14602 4326 18860 4378
rect 1104 4304 18860 4326
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 3513 4267 3571 4273
rect 3513 4264 3525 4267
rect 2832 4236 3525 4264
rect 2832 4224 2838 4236
rect 3513 4233 3525 4236
rect 3559 4233 3571 4267
rect 4249 4267 4307 4273
rect 3513 4227 3571 4233
rect 3620 4236 4200 4264
rect 3620 4196 3648 4236
rect 4172 4196 4200 4236
rect 4249 4233 4261 4267
rect 4295 4264 4307 4267
rect 4522 4264 4528 4276
rect 4295 4236 4528 4264
rect 4295 4233 4307 4236
rect 4249 4227 4307 4233
rect 4522 4224 4528 4236
rect 4580 4224 4586 4276
rect 4985 4267 5043 4273
rect 4985 4233 4997 4267
rect 5031 4264 5043 4267
rect 5166 4264 5172 4276
rect 5031 4236 5172 4264
rect 5031 4233 5043 4236
rect 4985 4227 5043 4233
rect 5166 4224 5172 4236
rect 5224 4224 5230 4276
rect 5445 4267 5503 4273
rect 5445 4233 5457 4267
rect 5491 4264 5503 4267
rect 5994 4264 6000 4276
rect 5491 4236 6000 4264
rect 5491 4233 5503 4236
rect 5445 4227 5503 4233
rect 5552 4208 5580 4236
rect 5994 4224 6000 4236
rect 6052 4224 6058 4276
rect 9398 4264 9404 4276
rect 9311 4236 9404 4264
rect 9398 4224 9404 4236
rect 9456 4264 9462 4276
rect 12066 4264 12072 4276
rect 9456 4236 12072 4264
rect 9456 4224 9462 4236
rect 12066 4224 12072 4236
rect 12124 4264 12130 4276
rect 12250 4264 12256 4276
rect 12124 4236 12256 4264
rect 12124 4224 12130 4236
rect 12250 4224 12256 4236
rect 12308 4224 12314 4276
rect 12437 4267 12495 4273
rect 12437 4233 12449 4267
rect 12483 4264 12495 4267
rect 12894 4264 12900 4276
rect 12483 4236 12900 4264
rect 12483 4233 12495 4236
rect 12437 4227 12495 4233
rect 12894 4224 12900 4236
rect 12952 4224 12958 4276
rect 15562 4224 15568 4276
rect 15620 4264 15626 4276
rect 15930 4264 15936 4276
rect 15620 4236 15936 4264
rect 15620 4224 15626 4236
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 16114 4224 16120 4276
rect 16172 4264 16178 4276
rect 17313 4267 17371 4273
rect 17313 4264 17325 4267
rect 16172 4236 17325 4264
rect 16172 4224 16178 4236
rect 17313 4233 17325 4236
rect 17359 4233 17371 4267
rect 17313 4227 17371 4233
rect 4706 4196 4712 4208
rect 3344 4168 3648 4196
rect 3712 4168 3924 4196
rect 4172 4168 4712 4196
rect 1673 4131 1731 4137
rect 1673 4097 1685 4131
rect 1719 4097 1731 4131
rect 1673 4091 1731 4097
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4128 2099 4131
rect 2130 4128 2136 4140
rect 2087 4100 2136 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 1688 4060 1716 4091
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2222 4088 2228 4140
rect 2280 4128 2286 4140
rect 2317 4131 2375 4137
rect 2317 4128 2329 4131
rect 2280 4100 2329 4128
rect 2280 4088 2286 4100
rect 2317 4097 2329 4100
rect 2363 4097 2375 4131
rect 2317 4091 2375 4097
rect 2593 4131 2651 4137
rect 2593 4097 2605 4131
rect 2639 4128 2651 4131
rect 2774 4128 2780 4140
rect 2639 4100 2780 4128
rect 2639 4097 2651 4100
rect 2593 4091 2651 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 2869 4131 2927 4137
rect 2869 4097 2881 4131
rect 2915 4128 2927 4131
rect 3145 4131 3203 4137
rect 2915 4100 3096 4128
rect 2915 4097 2927 4100
rect 2869 4091 2927 4097
rect 2958 4060 2964 4072
rect 1688 4032 2964 4060
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3068 4060 3096 4100
rect 3145 4097 3157 4131
rect 3191 4128 3203 4131
rect 3344 4128 3372 4168
rect 3191 4100 3372 4128
rect 3421 4131 3479 4137
rect 3191 4097 3203 4100
rect 3145 4091 3203 4097
rect 3421 4097 3433 4131
rect 3467 4128 3479 4131
rect 3602 4128 3608 4140
rect 3467 4100 3608 4128
rect 3467 4097 3479 4100
rect 3421 4091 3479 4097
rect 3602 4088 3608 4100
rect 3660 4088 3666 4140
rect 3712 4137 3740 4168
rect 3896 4140 3924 4168
rect 4706 4156 4712 4168
rect 4764 4156 4770 4208
rect 4908 4168 5120 4196
rect 3697 4131 3755 4137
rect 3697 4097 3709 4131
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 3786 4088 3792 4140
rect 3844 4088 3850 4140
rect 3878 4088 3884 4140
rect 3936 4088 3942 4140
rect 4154 4128 4160 4140
rect 4115 4100 4160 4128
rect 4154 4088 4160 4100
rect 4212 4088 4218 4140
rect 4908 4128 4936 4168
rect 5092 4137 5120 4168
rect 5534 4156 5540 4208
rect 5592 4156 5598 4208
rect 7374 4156 7380 4208
rect 7432 4196 7438 4208
rect 7432 4168 8064 4196
rect 7432 4156 7438 4168
rect 4264 4100 4936 4128
rect 5077 4131 5135 4137
rect 3804 4060 3832 4088
rect 4264 4060 4292 4100
rect 5077 4097 5089 4131
rect 5123 4097 5135 4131
rect 5077 4091 5135 4097
rect 5721 4131 5779 4137
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 5767 4100 6040 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 3068 4032 3372 4060
rect 3804 4032 4292 4060
rect 4433 4063 4491 4069
rect 2038 3952 2044 4004
rect 2096 3992 2102 4004
rect 3237 3995 3295 4001
rect 3237 3992 3249 3995
rect 2096 3964 3249 3992
rect 2096 3952 2102 3964
rect 3237 3961 3249 3964
rect 3283 3961 3295 3995
rect 3237 3955 3295 3961
rect 1486 3924 1492 3936
rect 1447 3896 1492 3924
rect 1486 3884 1492 3896
rect 1544 3884 1550 3936
rect 1578 3884 1584 3936
rect 1636 3924 1642 3936
rect 1857 3927 1915 3933
rect 1857 3924 1869 3927
rect 1636 3896 1869 3924
rect 1636 3884 1642 3896
rect 1857 3893 1869 3896
rect 1903 3893 1915 3927
rect 1857 3887 1915 3893
rect 1946 3884 1952 3936
rect 2004 3924 2010 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 2004 3896 2145 3924
rect 2004 3884 2010 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 2133 3887 2191 3893
rect 2222 3884 2228 3936
rect 2280 3924 2286 3936
rect 2409 3927 2467 3933
rect 2409 3924 2421 3927
rect 2280 3896 2421 3924
rect 2280 3884 2286 3896
rect 2409 3893 2421 3896
rect 2455 3893 2467 3927
rect 2409 3887 2467 3893
rect 2498 3884 2504 3936
rect 2556 3924 2562 3936
rect 2685 3927 2743 3933
rect 2685 3924 2697 3927
rect 2556 3896 2697 3924
rect 2556 3884 2562 3896
rect 2685 3893 2697 3896
rect 2731 3893 2743 3927
rect 2958 3924 2964 3936
rect 2919 3896 2964 3924
rect 2685 3887 2743 3893
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 3344 3924 3372 4032
rect 4433 4029 4445 4063
rect 4479 4060 4491 4063
rect 5261 4063 5319 4069
rect 4479 4032 4936 4060
rect 4479 4029 4491 4032
rect 4433 4023 4491 4029
rect 3786 3992 3792 4004
rect 3747 3964 3792 3992
rect 3786 3952 3792 3964
rect 3844 3952 3850 4004
rect 4614 3992 4620 4004
rect 4575 3964 4620 3992
rect 4614 3952 4620 3964
rect 4672 3952 4678 4004
rect 4908 3992 4936 4032
rect 5261 4029 5273 4063
rect 5307 4060 5319 4063
rect 5350 4060 5356 4072
rect 5307 4032 5356 4060
rect 5307 4029 5319 4032
rect 5261 4023 5319 4029
rect 5350 4020 5356 4032
rect 5408 4020 5414 4072
rect 5810 4020 5816 4072
rect 5868 4020 5874 4072
rect 6012 4060 6040 4100
rect 6086 4088 6092 4140
rect 6144 4128 6150 4140
rect 6457 4131 6515 4137
rect 6457 4128 6469 4131
rect 6144 4100 6469 4128
rect 6144 4088 6150 4100
rect 6457 4097 6469 4100
rect 6503 4097 6515 4131
rect 6457 4091 6515 4097
rect 6546 4088 6552 4140
rect 6604 4088 6610 4140
rect 6730 4137 6736 4140
rect 6724 4091 6736 4137
rect 6788 4128 6794 4140
rect 7929 4131 7987 4137
rect 7929 4128 7941 4131
rect 6788 4100 6824 4128
rect 7852 4100 7941 4128
rect 6730 4088 6736 4091
rect 6788 4088 6794 4100
rect 6564 4060 6592 4088
rect 6012 4032 6592 4060
rect 5828 3992 5856 4020
rect 4908 3964 5856 3992
rect 6181 3995 6239 4001
rect 6181 3961 6193 3995
rect 6227 3992 6239 3995
rect 6270 3992 6276 4004
rect 6227 3964 6276 3992
rect 6227 3961 6239 3964
rect 6181 3955 6239 3961
rect 6270 3952 6276 3964
rect 6328 3952 6334 4004
rect 7852 4001 7880 4100
rect 7929 4097 7941 4100
rect 7975 4097 7987 4131
rect 7929 4091 7987 4097
rect 8036 4060 8064 4168
rect 10060 4168 12112 4196
rect 8570 4128 8576 4140
rect 8531 4100 8576 4128
rect 8570 4088 8576 4100
rect 8628 4088 8634 4140
rect 8665 4131 8723 4137
rect 8665 4097 8677 4131
rect 8711 4128 8723 4131
rect 8941 4131 8999 4137
rect 8941 4128 8953 4131
rect 8711 4100 8953 4128
rect 8711 4097 8723 4100
rect 8665 4091 8723 4097
rect 8941 4097 8953 4100
rect 8987 4097 8999 4131
rect 8941 4091 8999 4097
rect 9585 4131 9643 4137
rect 9585 4097 9597 4131
rect 9631 4097 9643 4131
rect 9585 4091 9643 4097
rect 8680 4060 8708 4091
rect 9600 4060 9628 4091
rect 9674 4088 9680 4140
rect 9732 4128 9738 4140
rect 10060 4128 10088 4168
rect 10226 4128 10232 4140
rect 9732 4100 10088 4128
rect 10187 4100 10232 4128
rect 9732 4088 9738 4100
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 10502 4128 10508 4140
rect 10415 4100 10508 4128
rect 10502 4088 10508 4100
rect 10560 4088 10566 4140
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4128 11207 4131
rect 11238 4128 11244 4140
rect 11195 4100 11244 4128
rect 11195 4097 11207 4100
rect 11149 4091 11207 4097
rect 11238 4088 11244 4100
rect 11296 4088 11302 4140
rect 11701 4131 11759 4137
rect 11701 4097 11713 4131
rect 11747 4097 11759 4131
rect 11974 4128 11980 4140
rect 11935 4100 11980 4128
rect 11701 4091 11759 4097
rect 10520 4060 10548 4088
rect 10870 4060 10876 4072
rect 8036 4032 8708 4060
rect 8864 4032 10876 4060
rect 7837 3995 7895 4001
rect 7837 3961 7849 3995
rect 7883 3992 7895 3995
rect 8018 3992 8024 4004
rect 7883 3964 8024 3992
rect 7883 3961 7895 3964
rect 7837 3955 7895 3961
rect 8018 3952 8024 3964
rect 8076 3952 8082 4004
rect 8864 4001 8892 4032
rect 10870 4020 10876 4032
rect 10928 4020 10934 4072
rect 10965 4063 11023 4069
rect 10965 4029 10977 4063
rect 11011 4060 11023 4063
rect 11054 4060 11060 4072
rect 11011 4032 11060 4060
rect 11011 4029 11023 4032
rect 10965 4023 11023 4029
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 11514 4020 11520 4072
rect 11572 4060 11578 4072
rect 11716 4060 11744 4091
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 12084 4128 12112 4168
rect 13630 4156 13636 4208
rect 13688 4196 13694 4208
rect 15010 4196 15016 4208
rect 13688 4168 15016 4196
rect 13688 4156 13694 4168
rect 15010 4156 15016 4168
rect 15068 4156 15074 4208
rect 15381 4199 15439 4205
rect 15381 4165 15393 4199
rect 15427 4196 15439 4199
rect 15427 4168 15976 4196
rect 15427 4165 15439 4168
rect 15381 4159 15439 4165
rect 12253 4131 12311 4137
rect 12253 4128 12265 4131
rect 12084 4100 12265 4128
rect 12253 4097 12265 4100
rect 12299 4097 12311 4131
rect 12526 4128 12532 4140
rect 12487 4100 12532 4128
rect 12253 4091 12311 4097
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 14642 4128 14648 4140
rect 14603 4100 14648 4128
rect 14642 4088 14648 4100
rect 14700 4088 14706 4140
rect 15102 4088 15108 4140
rect 15160 4128 15166 4140
rect 15519 4131 15577 4137
rect 15519 4128 15531 4131
rect 15160 4100 15531 4128
rect 15160 4088 15166 4100
rect 15519 4097 15531 4100
rect 15565 4097 15577 4131
rect 15519 4091 15577 4097
rect 15622 4131 15680 4137
rect 15622 4097 15634 4131
rect 15668 4128 15680 4131
rect 15841 4131 15899 4137
rect 15668 4097 15700 4128
rect 15622 4091 15700 4097
rect 15841 4097 15853 4131
rect 15887 4097 15899 4131
rect 15841 4091 15899 4097
rect 12618 4060 12624 4072
rect 11572 4032 11744 4060
rect 11900 4032 12624 4060
rect 11572 4020 11578 4032
rect 8849 3995 8907 4001
rect 8849 3961 8861 3995
rect 8895 3961 8907 3995
rect 10318 3992 10324 4004
rect 8849 3955 8907 3961
rect 9876 3964 10324 3992
rect 5534 3924 5540 3936
rect 3344 3896 5540 3924
rect 5534 3884 5540 3896
rect 5592 3884 5598 3936
rect 5902 3924 5908 3936
rect 5815 3896 5908 3924
rect 5902 3884 5908 3896
rect 5960 3924 5966 3936
rect 6822 3924 6828 3936
rect 5960 3896 6828 3924
rect 5960 3884 5966 3896
rect 6822 3884 6828 3896
rect 6880 3884 6886 3936
rect 9122 3924 9128 3936
rect 9083 3896 9128 3924
rect 9122 3884 9128 3896
rect 9180 3884 9186 3936
rect 9876 3933 9904 3964
rect 10318 3952 10324 3964
rect 10376 3952 10382 4004
rect 10413 3995 10471 4001
rect 10413 3961 10425 3995
rect 10459 3992 10471 3995
rect 11238 3992 11244 4004
rect 10459 3964 11244 3992
rect 10459 3961 10471 3964
rect 10413 3955 10471 3961
rect 11238 3952 11244 3964
rect 11296 3952 11302 4004
rect 11900 4001 11928 4032
rect 12618 4020 12624 4032
rect 12676 4020 12682 4072
rect 12802 4060 12808 4072
rect 12763 4032 12808 4060
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 12986 4060 12992 4072
rect 12947 4032 12992 4060
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 13906 4020 13912 4072
rect 13964 4060 13970 4072
rect 14737 4063 14795 4069
rect 14737 4060 14749 4063
rect 13964 4032 14749 4060
rect 13964 4020 13970 4032
rect 14737 4029 14749 4032
rect 14783 4029 14795 4063
rect 14918 4060 14924 4072
rect 14879 4032 14924 4060
rect 14737 4023 14795 4029
rect 14918 4020 14924 4032
rect 14976 4060 14982 4072
rect 15672 4060 15700 4091
rect 14976 4032 15700 4060
rect 14976 4020 14982 4032
rect 11333 3995 11391 4001
rect 11333 3961 11345 3995
rect 11379 3992 11391 3995
rect 11885 3995 11943 4001
rect 11379 3964 11836 3992
rect 11379 3961 11391 3964
rect 11333 3955 11391 3961
rect 9861 3927 9919 3933
rect 9861 3893 9873 3927
rect 9907 3893 9919 3927
rect 9861 3887 9919 3893
rect 10045 3927 10103 3933
rect 10045 3893 10057 3927
rect 10091 3924 10103 3927
rect 10134 3924 10140 3936
rect 10091 3896 10140 3924
rect 10091 3893 10103 3896
rect 10045 3887 10103 3893
rect 10134 3884 10140 3896
rect 10192 3884 10198 3936
rect 10778 3924 10784 3936
rect 10739 3896 10784 3924
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 11609 3927 11667 3933
rect 11609 3893 11621 3927
rect 11655 3924 11667 3927
rect 11698 3924 11704 3936
rect 11655 3896 11704 3924
rect 11655 3893 11667 3896
rect 11609 3887 11667 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 11808 3924 11836 3964
rect 11885 3961 11897 3995
rect 11931 3961 11943 3995
rect 15856 3992 15884 4091
rect 15948 4060 15976 4168
rect 16390 4088 16396 4140
rect 16448 4128 16454 4140
rect 16485 4131 16543 4137
rect 16485 4128 16497 4131
rect 16448 4100 16497 4128
rect 16448 4088 16454 4100
rect 16485 4097 16497 4100
rect 16531 4097 16543 4131
rect 17034 4128 17040 4140
rect 16485 4091 16543 4097
rect 16592 4100 17040 4128
rect 16592 4060 16620 4100
rect 17034 4088 17040 4100
rect 17092 4088 17098 4140
rect 17497 4131 17555 4137
rect 17497 4097 17509 4131
rect 17543 4097 17555 4131
rect 17497 4091 17555 4097
rect 15948 4032 16620 4060
rect 16666 4020 16672 4072
rect 16724 4060 16730 4072
rect 16724 4032 16769 4060
rect 16724 4020 16730 4032
rect 16850 4020 16856 4072
rect 16908 4060 16914 4072
rect 16908 4032 16953 4060
rect 16908 4020 16914 4032
rect 17512 3992 17540 4091
rect 17586 4088 17592 4140
rect 17644 4128 17650 4140
rect 17865 4131 17923 4137
rect 17865 4128 17877 4131
rect 17644 4100 17877 4128
rect 17644 4088 17650 4100
rect 17865 4097 17877 4100
rect 17911 4097 17923 4131
rect 18230 4128 18236 4140
rect 18191 4100 18236 4128
rect 17865 4091 17923 4097
rect 18230 4088 18236 4100
rect 18288 4088 18294 4140
rect 11885 3955 11943 3961
rect 11992 3964 15884 3992
rect 15948 3964 17540 3992
rect 11992 3924 12020 3964
rect 11808 3896 12020 3924
rect 12161 3927 12219 3933
rect 12161 3893 12173 3927
rect 12207 3924 12219 3927
rect 12434 3924 12440 3936
rect 12207 3896 12440 3924
rect 12207 3893 12219 3896
rect 12161 3887 12219 3893
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 12710 3924 12716 3936
rect 12671 3896 12716 3924
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 15948 3924 15976 3964
rect 17862 3952 17868 4004
rect 17920 3992 17926 4004
rect 18049 3995 18107 4001
rect 18049 3992 18061 3995
rect 17920 3964 18061 3992
rect 17920 3952 17926 3964
rect 18049 3961 18061 3964
rect 18095 3961 18107 3995
rect 18049 3955 18107 3961
rect 12952 3896 15976 3924
rect 12952 3884 12958 3896
rect 16022 3884 16028 3936
rect 16080 3924 16086 3936
rect 16298 3924 16304 3936
rect 16080 3896 16125 3924
rect 16259 3896 16304 3924
rect 16080 3884 16086 3896
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 17678 3924 17684 3936
rect 17639 3896 17684 3924
rect 17678 3884 17684 3896
rect 17736 3884 17742 3936
rect 17770 3884 17776 3936
rect 17828 3924 17834 3936
rect 18417 3927 18475 3933
rect 18417 3924 18429 3927
rect 17828 3896 18429 3924
rect 17828 3884 17834 3896
rect 18417 3893 18429 3896
rect 18463 3893 18475 3927
rect 18417 3887 18475 3893
rect 1104 3834 18860 3856
rect 1104 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 3430 3834
rect 3482 3782 7622 3834
rect 7674 3782 7686 3834
rect 7738 3782 7750 3834
rect 7802 3782 7814 3834
rect 7866 3782 7878 3834
rect 7930 3782 12070 3834
rect 12122 3782 12134 3834
rect 12186 3782 12198 3834
rect 12250 3782 12262 3834
rect 12314 3782 12326 3834
rect 12378 3782 16518 3834
rect 16570 3782 16582 3834
rect 16634 3782 16646 3834
rect 16698 3782 16710 3834
rect 16762 3782 16774 3834
rect 16826 3782 18860 3834
rect 1104 3760 18860 3782
rect 2866 3680 2872 3732
rect 2924 3720 2930 3732
rect 3329 3723 3387 3729
rect 3329 3720 3341 3723
rect 2924 3692 3341 3720
rect 2924 3680 2930 3692
rect 3329 3689 3341 3692
rect 3375 3689 3387 3723
rect 3878 3720 3884 3732
rect 3839 3692 3884 3720
rect 3329 3683 3387 3689
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 5350 3720 5356 3732
rect 5311 3692 5356 3720
rect 5350 3680 5356 3692
rect 5408 3680 5414 3732
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 6917 3723 6975 3729
rect 6917 3720 6929 3723
rect 6788 3692 6929 3720
rect 6788 3680 6794 3692
rect 6917 3689 6929 3692
rect 6963 3689 6975 3723
rect 6917 3683 6975 3689
rect 7929 3723 7987 3729
rect 7929 3689 7941 3723
rect 7975 3720 7987 3723
rect 8018 3720 8024 3732
rect 7975 3692 8024 3720
rect 7975 3689 7987 3692
rect 7929 3683 7987 3689
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 9585 3723 9643 3729
rect 9585 3689 9597 3723
rect 9631 3720 9643 3723
rect 10226 3720 10232 3732
rect 9631 3692 10232 3720
rect 9631 3689 9643 3692
rect 9585 3683 9643 3689
rect 10226 3680 10232 3692
rect 10284 3680 10290 3732
rect 12667 3723 12725 3729
rect 12667 3689 12679 3723
rect 12713 3720 12725 3723
rect 12986 3720 12992 3732
rect 12713 3692 12992 3720
rect 12713 3689 12725 3692
rect 12667 3683 12725 3689
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 17218 3720 17224 3732
rect 13648 3692 17224 3720
rect 3053 3655 3111 3661
rect 3053 3652 3065 3655
rect 2746 3624 3065 3652
rect 2222 3584 2228 3596
rect 1688 3556 2228 3584
rect 1688 3525 1716 3556
rect 2222 3544 2228 3556
rect 2280 3544 2286 3596
rect 2746 3584 2774 3624
rect 3053 3621 3065 3624
rect 3099 3621 3111 3655
rect 3053 3615 3111 3621
rect 6825 3655 6883 3661
rect 6825 3621 6837 3655
rect 6871 3621 6883 3655
rect 6825 3615 6883 3621
rect 8113 3655 8171 3661
rect 8113 3621 8125 3655
rect 8159 3652 8171 3655
rect 8159 3624 9628 3652
rect 8159 3621 8171 3624
rect 8113 3615 8171 3621
rect 2424 3556 2774 3584
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 2041 3519 2099 3525
rect 2041 3485 2053 3519
rect 2087 3516 2099 3519
rect 2424 3516 2452 3556
rect 2590 3516 2596 3528
rect 2087 3488 2452 3516
rect 2551 3488 2596 3516
rect 2087 3485 2099 3488
rect 2041 3479 2099 3485
rect 2590 3476 2596 3488
rect 2648 3476 2654 3528
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3516 3019 3519
rect 3142 3516 3148 3528
rect 3007 3488 3148 3516
rect 3007 3485 3019 3488
rect 2961 3479 3019 3485
rect 3142 3476 3148 3488
rect 3200 3476 3206 3528
rect 3237 3519 3295 3525
rect 3237 3485 3249 3519
rect 3283 3516 3295 3519
rect 3418 3516 3424 3528
rect 3283 3488 3424 3516
rect 3283 3485 3295 3488
rect 3237 3479 3295 3485
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 3513 3519 3571 3525
rect 3513 3485 3525 3519
rect 3559 3516 3571 3519
rect 3878 3516 3884 3528
rect 3559 3488 3884 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 3878 3476 3884 3488
rect 3936 3476 3942 3528
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3516 4031 3519
rect 5445 3519 5503 3525
rect 5445 3516 5457 3519
rect 4019 3488 5457 3516
rect 4019 3485 4031 3488
rect 3973 3479 4031 3485
rect 5445 3485 5457 3488
rect 5491 3516 5503 3519
rect 6086 3516 6092 3528
rect 5491 3488 6092 3516
rect 5491 3485 5503 3488
rect 5445 3479 5503 3485
rect 6086 3476 6092 3488
rect 6144 3476 6150 3528
rect 6840 3516 6868 3615
rect 7006 3544 7012 3596
rect 7064 3584 7070 3596
rect 8018 3584 8024 3596
rect 7064 3556 8024 3584
rect 7064 3544 7070 3556
rect 8018 3544 8024 3556
rect 8076 3544 8082 3596
rect 7098 3516 7104 3528
rect 6840 3488 7104 3516
rect 7098 3476 7104 3488
rect 7156 3516 7162 3528
rect 8220 3525 8248 3624
rect 8846 3544 8852 3596
rect 8904 3584 8910 3596
rect 8941 3587 8999 3593
rect 8941 3584 8953 3587
rect 8904 3556 8953 3584
rect 8904 3544 8910 3556
rect 8941 3553 8953 3556
rect 8987 3553 8999 3587
rect 9600 3584 9628 3624
rect 9674 3612 9680 3664
rect 9732 3652 9738 3664
rect 9953 3655 10011 3661
rect 9953 3652 9965 3655
rect 9732 3624 9965 3652
rect 9732 3612 9738 3624
rect 9953 3621 9965 3624
rect 9999 3621 10011 3655
rect 9953 3615 10011 3621
rect 10042 3612 10048 3664
rect 10100 3652 10106 3664
rect 10318 3652 10324 3664
rect 10100 3624 10324 3652
rect 10100 3612 10106 3624
rect 10318 3612 10324 3624
rect 10376 3612 10382 3664
rect 12434 3612 12440 3664
rect 12492 3652 12498 3664
rect 13648 3652 13676 3692
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 18414 3720 18420 3732
rect 18375 3692 18420 3720
rect 18414 3680 18420 3692
rect 18472 3680 18478 3732
rect 12492 3624 13676 3652
rect 12492 3612 12498 3624
rect 13722 3612 13728 3664
rect 13780 3652 13786 3664
rect 14461 3655 14519 3661
rect 14461 3652 14473 3655
rect 13780 3624 14473 3652
rect 13780 3612 13786 3624
rect 14461 3621 14473 3624
rect 14507 3621 14519 3655
rect 14461 3615 14519 3621
rect 16298 3612 16304 3664
rect 16356 3652 16362 3664
rect 18598 3652 18604 3664
rect 16356 3624 18604 3652
rect 16356 3612 16362 3624
rect 18598 3612 18604 3624
rect 18656 3612 18662 3664
rect 11054 3584 11060 3596
rect 9600 3556 11060 3584
rect 8941 3547 8999 3553
rect 11054 3544 11060 3556
rect 11112 3544 11118 3596
rect 13906 3544 13912 3596
rect 13964 3584 13970 3596
rect 14277 3587 14335 3593
rect 14277 3584 14289 3587
rect 13964 3556 14289 3584
rect 13964 3544 13970 3556
rect 14277 3553 14289 3556
rect 14323 3553 14335 3587
rect 15286 3584 15292 3596
rect 15247 3556 15292 3584
rect 14277 3547 14335 3553
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 15470 3584 15476 3596
rect 15431 3556 15476 3584
rect 15470 3544 15476 3556
rect 15528 3544 15534 3596
rect 17586 3584 17592 3596
rect 16684 3556 17592 3584
rect 7561 3519 7619 3525
rect 7561 3516 7573 3519
rect 7156 3488 7573 3516
rect 7156 3476 7162 3488
rect 7561 3485 7573 3488
rect 7607 3485 7619 3519
rect 7561 3479 7619 3485
rect 7653 3519 7711 3525
rect 7653 3485 7665 3519
rect 7699 3485 7711 3519
rect 7653 3479 7711 3485
rect 8205 3519 8263 3525
rect 8205 3485 8217 3519
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 2317 3451 2375 3457
rect 2317 3417 2329 3451
rect 2363 3448 2375 3451
rect 4240 3451 4298 3457
rect 2363 3420 4016 3448
rect 2363 3417 2375 3420
rect 2317 3411 2375 3417
rect 1486 3380 1492 3392
rect 1447 3352 1492 3380
rect 1486 3340 1492 3352
rect 1544 3340 1550 3392
rect 1854 3380 1860 3392
rect 1815 3352 1860 3380
rect 1854 3340 1860 3352
rect 1912 3340 1918 3392
rect 2774 3340 2780 3392
rect 2832 3380 2838 3392
rect 3988 3380 4016 3420
rect 4240 3417 4252 3451
rect 4286 3448 4298 3451
rect 4706 3448 4712 3460
rect 4286 3420 4712 3448
rect 4286 3417 4298 3420
rect 4240 3411 4298 3417
rect 4706 3408 4712 3420
rect 4764 3408 4770 3460
rect 5712 3451 5770 3457
rect 5712 3417 5724 3451
rect 5758 3448 5770 3451
rect 5758 3420 6868 3448
rect 5758 3417 5770 3420
rect 5712 3411 5770 3417
rect 5166 3380 5172 3392
rect 2832 3352 2877 3380
rect 3988 3352 5172 3380
rect 2832 3340 2838 3352
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 6840 3380 6868 3420
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 7668 3448 7696 3479
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 8608 3519 8666 3525
rect 8608 3516 8620 3519
rect 8352 3488 8620 3516
rect 8352 3476 8358 3488
rect 8608 3485 8620 3488
rect 8654 3516 8666 3519
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 8654 3488 9137 3516
rect 8654 3485 8666 3488
rect 8608 3479 8666 3485
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9728 3519 9786 3525
rect 9728 3516 9740 3519
rect 9125 3479 9183 3485
rect 9232 3488 9740 3516
rect 6972 3420 7696 3448
rect 6972 3408 6978 3420
rect 7926 3408 7932 3460
rect 7984 3448 7990 3460
rect 9232 3448 9260 3488
rect 9728 3485 9740 3488
rect 9774 3516 9786 3519
rect 10042 3516 10048 3528
rect 9774 3488 10048 3516
rect 9774 3485 9786 3488
rect 9728 3479 9786 3485
rect 10042 3476 10048 3488
rect 10100 3476 10106 3528
rect 10137 3519 10195 3525
rect 10137 3485 10149 3519
rect 10183 3516 10195 3519
rect 10226 3516 10232 3528
rect 10183 3488 10232 3516
rect 10183 3485 10195 3488
rect 10137 3479 10195 3485
rect 10226 3476 10232 3488
rect 10284 3476 10290 3528
rect 10413 3519 10471 3525
rect 10413 3485 10425 3519
rect 10459 3516 10471 3519
rect 10962 3516 10968 3528
rect 10459 3488 10968 3516
rect 10459 3485 10471 3488
rect 10413 3479 10471 3485
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11146 3476 11152 3528
rect 11204 3516 11210 3528
rect 12161 3519 12219 3525
rect 12161 3516 12173 3519
rect 11204 3488 12173 3516
rect 11204 3476 11210 3488
rect 12161 3485 12173 3488
rect 12207 3485 12219 3519
rect 12161 3479 12219 3485
rect 12250 3476 12256 3528
rect 12308 3525 12314 3528
rect 12308 3519 12346 3525
rect 12334 3485 12346 3519
rect 12308 3479 12346 3485
rect 12564 3519 12622 3525
rect 12564 3485 12576 3519
rect 12610 3485 12622 3519
rect 12564 3479 12622 3485
rect 12308 3476 12314 3479
rect 7984 3420 9260 3448
rect 7984 3408 7990 3420
rect 9490 3408 9496 3460
rect 9548 3448 9554 3460
rect 9815 3451 9873 3457
rect 9548 3420 9720 3448
rect 9548 3408 9554 3420
rect 7190 3380 7196 3392
rect 6840 3352 7196 3380
rect 7190 3340 7196 3352
rect 7248 3340 7254 3392
rect 8386 3380 8392 3392
rect 8347 3352 8392 3380
rect 8386 3340 8392 3352
rect 8444 3340 8450 3392
rect 8711 3383 8769 3389
rect 8711 3349 8723 3383
rect 8757 3380 8769 3383
rect 9582 3380 9588 3392
rect 8757 3352 9588 3380
rect 8757 3349 8769 3352
rect 8711 3343 8769 3349
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 9692 3380 9720 3420
rect 9815 3417 9827 3451
rect 9861 3448 9873 3451
rect 11698 3448 11704 3460
rect 9861 3420 11704 3448
rect 9861 3417 9873 3420
rect 9815 3411 9873 3417
rect 11698 3408 11704 3420
rect 11756 3408 11762 3460
rect 11882 3408 11888 3460
rect 11940 3457 11946 3460
rect 11940 3448 11952 3457
rect 11940 3420 11985 3448
rect 11940 3411 11952 3420
rect 11940 3408 11946 3411
rect 12066 3408 12072 3460
rect 12124 3448 12130 3460
rect 12579 3448 12607 3479
rect 12710 3476 12716 3528
rect 12768 3516 12774 3528
rect 12805 3519 12863 3525
rect 12805 3516 12817 3519
rect 12768 3488 12817 3516
rect 12768 3476 12774 3488
rect 12805 3485 12817 3488
rect 12851 3485 12863 3519
rect 12805 3479 12863 3485
rect 12986 3476 12992 3528
rect 13044 3516 13050 3528
rect 13081 3519 13139 3525
rect 13081 3516 13093 3519
rect 13044 3488 13093 3516
rect 13044 3476 13050 3488
rect 13081 3485 13093 3488
rect 13127 3485 13139 3519
rect 13081 3479 13139 3485
rect 13170 3476 13176 3528
rect 13228 3516 13234 3528
rect 13449 3519 13507 3525
rect 13449 3516 13461 3519
rect 13228 3488 13461 3516
rect 13228 3476 13234 3488
rect 13449 3485 13461 3488
rect 13495 3485 13507 3519
rect 13449 3479 13507 3485
rect 13538 3476 13544 3528
rect 13596 3516 13602 3528
rect 13725 3519 13783 3525
rect 13725 3516 13737 3519
rect 13596 3488 13737 3516
rect 13596 3476 13602 3488
rect 13725 3485 13737 3488
rect 13771 3485 13783 3519
rect 14090 3516 14096 3528
rect 14051 3488 14096 3516
rect 13725 3479 13783 3485
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 15194 3516 15200 3528
rect 15155 3488 15200 3516
rect 15194 3476 15200 3488
rect 15252 3476 15258 3528
rect 14182 3448 14188 3460
rect 12124 3420 12607 3448
rect 13004 3420 14188 3448
rect 12124 3408 12130 3420
rect 10229 3383 10287 3389
rect 10229 3380 10241 3383
rect 9692 3352 10241 3380
rect 10229 3349 10241 3352
rect 10275 3349 10287 3383
rect 10594 3380 10600 3392
rect 10555 3352 10600 3380
rect 10229 3343 10287 3349
rect 10594 3340 10600 3352
rect 10652 3340 10658 3392
rect 10778 3380 10784 3392
rect 10739 3352 10784 3380
rect 10778 3340 10784 3352
rect 10836 3340 10842 3392
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 11514 3380 11520 3392
rect 11204 3352 11520 3380
rect 11204 3340 11210 3352
rect 11514 3340 11520 3352
rect 11572 3340 11578 3392
rect 12391 3383 12449 3389
rect 12391 3349 12403 3383
rect 12437 3380 12449 3383
rect 12894 3380 12900 3392
rect 12437 3352 12900 3380
rect 12437 3349 12449 3352
rect 12391 3343 12449 3349
rect 12894 3340 12900 3352
rect 12952 3340 12958 3392
rect 13004 3389 13032 3420
rect 14182 3408 14188 3420
rect 14240 3408 14246 3460
rect 16684 3448 16712 3556
rect 17586 3544 17592 3556
rect 17644 3544 17650 3596
rect 17221 3519 17279 3525
rect 17221 3485 17233 3519
rect 17267 3516 17279 3519
rect 17310 3516 17316 3528
rect 17267 3488 17316 3516
rect 17267 3485 17279 3488
rect 17221 3479 17279 3485
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 17402 3476 17408 3528
rect 17460 3516 17466 3528
rect 17497 3519 17555 3525
rect 17497 3516 17509 3519
rect 17460 3488 17509 3516
rect 17460 3476 17466 3488
rect 17497 3485 17509 3488
rect 17543 3485 17555 3519
rect 17497 3479 17555 3485
rect 17678 3476 17684 3528
rect 17736 3516 17742 3528
rect 17865 3519 17923 3525
rect 17865 3516 17877 3519
rect 17736 3488 17877 3516
rect 17736 3476 17742 3488
rect 17865 3485 17877 3488
rect 17911 3485 17923 3519
rect 17865 3479 17923 3485
rect 18138 3476 18144 3528
rect 18196 3516 18202 3528
rect 18233 3519 18291 3525
rect 18233 3516 18245 3519
rect 18196 3488 18245 3516
rect 18196 3476 18202 3488
rect 18233 3485 18245 3488
rect 18279 3485 18291 3519
rect 18233 3479 18291 3485
rect 17126 3448 17132 3460
rect 14936 3420 16712 3448
rect 17087 3420 17132 3448
rect 12989 3383 13047 3389
rect 12989 3349 13001 3383
rect 13035 3349 13047 3383
rect 12989 3343 13047 3349
rect 13265 3383 13323 3389
rect 13265 3349 13277 3383
rect 13311 3380 13323 3383
rect 13354 3380 13360 3392
rect 13311 3352 13360 3380
rect 13311 3349 13323 3352
rect 13265 3343 13323 3349
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 13630 3380 13636 3392
rect 13591 3352 13636 3380
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 13909 3383 13967 3389
rect 13909 3349 13921 3383
rect 13955 3380 13967 3383
rect 14936 3380 14964 3420
rect 17126 3408 17132 3420
rect 17184 3408 17190 3460
rect 19610 3448 19616 3460
rect 17328 3420 19616 3448
rect 13955 3352 14964 3380
rect 15013 3383 15071 3389
rect 13955 3349 13967 3352
rect 13909 3343 13967 3349
rect 15013 3349 15025 3383
rect 15059 3380 15071 3383
rect 17328 3380 17356 3420
rect 19610 3408 19616 3420
rect 19668 3408 19674 3460
rect 15059 3352 17356 3380
rect 17405 3383 17463 3389
rect 15059 3349 15071 3352
rect 15013 3343 15071 3349
rect 17405 3349 17417 3383
rect 17451 3380 17463 3383
rect 17494 3380 17500 3392
rect 17451 3352 17500 3380
rect 17451 3349 17463 3352
rect 17405 3343 17463 3349
rect 17494 3340 17500 3352
rect 17552 3340 17558 3392
rect 17586 3340 17592 3392
rect 17644 3380 17650 3392
rect 17681 3383 17739 3389
rect 17681 3380 17693 3383
rect 17644 3352 17693 3380
rect 17644 3340 17650 3352
rect 17681 3349 17693 3352
rect 17727 3349 17739 3383
rect 18046 3380 18052 3392
rect 18007 3352 18052 3380
rect 17681 3343 17739 3349
rect 18046 3340 18052 3352
rect 18104 3340 18110 3392
rect 1104 3290 18860 3312
rect 1104 3238 5398 3290
rect 5450 3238 5462 3290
rect 5514 3238 5526 3290
rect 5578 3238 5590 3290
rect 5642 3238 5654 3290
rect 5706 3238 9846 3290
rect 9898 3238 9910 3290
rect 9962 3238 9974 3290
rect 10026 3238 10038 3290
rect 10090 3238 10102 3290
rect 10154 3238 14294 3290
rect 14346 3238 14358 3290
rect 14410 3238 14422 3290
rect 14474 3238 14486 3290
rect 14538 3238 14550 3290
rect 14602 3238 18860 3290
rect 1104 3216 18860 3238
rect 198 3136 204 3188
rect 256 3176 262 3188
rect 2225 3179 2283 3185
rect 2225 3176 2237 3179
rect 256 3148 2237 3176
rect 256 3136 262 3148
rect 2225 3145 2237 3148
rect 2271 3145 2283 3179
rect 2225 3139 2283 3145
rect 3142 3136 3148 3188
rect 3200 3176 3206 3188
rect 3605 3179 3663 3185
rect 3605 3176 3617 3179
rect 3200 3148 3617 3176
rect 3200 3136 3206 3148
rect 3605 3145 3617 3148
rect 3651 3145 3663 3179
rect 4614 3176 4620 3188
rect 4575 3148 4620 3176
rect 3605 3139 3663 3145
rect 4614 3136 4620 3148
rect 4672 3136 4678 3188
rect 4890 3136 4896 3188
rect 4948 3176 4954 3188
rect 5077 3179 5135 3185
rect 5077 3176 5089 3179
rect 4948 3148 5089 3176
rect 4948 3136 4954 3148
rect 5077 3145 5089 3148
rect 5123 3145 5135 3179
rect 5258 3176 5264 3188
rect 5219 3148 5264 3176
rect 5077 3139 5135 3145
rect 5258 3136 5264 3148
rect 5316 3136 5322 3188
rect 6549 3179 6607 3185
rect 6549 3145 6561 3179
rect 6595 3176 6607 3179
rect 7190 3176 7196 3188
rect 6595 3148 7196 3176
rect 6595 3145 6607 3148
rect 6549 3139 6607 3145
rect 7190 3136 7196 3148
rect 7248 3136 7254 3188
rect 7377 3179 7435 3185
rect 7377 3145 7389 3179
rect 7423 3176 7435 3179
rect 7423 3148 10180 3176
rect 7423 3145 7435 3148
rect 7377 3139 7435 3145
rect 3050 3108 3056 3120
rect 2792 3080 3056 3108
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3040 1731 3043
rect 1946 3040 1952 3052
rect 1719 3012 1952 3040
rect 1719 3009 1731 3012
rect 1673 3003 1731 3009
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 2038 3000 2044 3052
rect 2096 3040 2102 3052
rect 2406 3040 2412 3052
rect 2096 3012 2141 3040
rect 2367 3012 2412 3040
rect 2096 3000 2102 3012
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 2792 3049 2820 3080
rect 3050 3068 3056 3080
rect 3108 3068 3114 3120
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3009 2835 3043
rect 2777 3003 2835 3009
rect 2958 3000 2964 3052
rect 3016 3040 3022 3052
rect 3145 3043 3203 3049
rect 3145 3040 3157 3043
rect 3016 3012 3157 3040
rect 3016 3000 3022 3012
rect 3145 3009 3157 3012
rect 3191 3009 3203 3043
rect 3145 3003 3203 3009
rect 3234 3000 3240 3052
rect 3292 3040 3298 3052
rect 3789 3043 3847 3049
rect 3292 3012 3337 3040
rect 3292 3000 3298 3012
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 4062 3040 4068 3052
rect 3835 3012 4068 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3040 4215 3043
rect 4246 3040 4252 3052
rect 4203 3012 4252 3040
rect 4203 3009 4215 3012
rect 4157 3003 4215 3009
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 4632 3040 4660 3136
rect 7392 3108 7420 3139
rect 9398 3108 9404 3120
rect 6656 3080 7420 3108
rect 8220 3080 9404 3108
rect 6656 3049 6684 3080
rect 4479 3012 4660 3040
rect 5997 3043 6055 3049
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 5997 3009 6009 3043
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3009 6699 3043
rect 6914 3040 6920 3052
rect 6875 3012 6920 3040
rect 6641 3003 6699 3009
rect 658 2932 664 2984
rect 716 2972 722 2984
rect 716 2944 2636 2972
rect 716 2932 722 2944
rect 1118 2864 1124 2916
rect 1176 2904 1182 2916
rect 2608 2913 2636 2944
rect 3418 2932 3424 2984
rect 3476 2972 3482 2984
rect 4893 2975 4951 2981
rect 4893 2972 4905 2975
rect 3476 2944 4905 2972
rect 3476 2932 3482 2944
rect 4893 2941 4905 2944
rect 4939 2941 4951 2975
rect 5902 2972 5908 2984
rect 5863 2944 5908 2972
rect 4893 2935 4951 2941
rect 5902 2932 5908 2944
rect 5960 2932 5966 2984
rect 1857 2907 1915 2913
rect 1857 2904 1869 2907
rect 1176 2876 1869 2904
rect 1176 2864 1182 2876
rect 1857 2873 1869 2876
rect 1903 2873 1915 2907
rect 1857 2867 1915 2873
rect 2593 2907 2651 2913
rect 2593 2873 2605 2907
rect 2639 2873 2651 2907
rect 2593 2867 2651 2873
rect 1486 2836 1492 2848
rect 1447 2808 1492 2836
rect 1486 2796 1492 2808
rect 1544 2796 1550 2848
rect 2958 2836 2964 2848
rect 2919 2808 2964 2836
rect 2958 2796 2964 2808
rect 3016 2796 3022 2848
rect 3050 2796 3056 2848
rect 3108 2836 3114 2848
rect 3421 2839 3479 2845
rect 3421 2836 3433 2839
rect 3108 2808 3433 2836
rect 3108 2796 3114 2808
rect 3421 2805 3433 2808
rect 3467 2805 3479 2839
rect 3970 2836 3976 2848
rect 3931 2808 3976 2836
rect 3421 2799 3479 2805
rect 3970 2796 3976 2808
rect 4028 2796 4034 2848
rect 4246 2836 4252 2848
rect 4207 2808 4252 2836
rect 4246 2796 4252 2808
rect 4304 2796 4310 2848
rect 4614 2796 4620 2848
rect 4672 2836 4678 2848
rect 4709 2839 4767 2845
rect 4709 2836 4721 2839
rect 4672 2808 4721 2836
rect 4672 2796 4678 2808
rect 4709 2805 4721 2808
rect 4755 2805 4767 2839
rect 4709 2799 4767 2805
rect 5629 2839 5687 2845
rect 5629 2805 5641 2839
rect 5675 2836 5687 2839
rect 5718 2836 5724 2848
rect 5675 2808 5724 2836
rect 5675 2805 5687 2808
rect 5629 2799 5687 2805
rect 5718 2796 5724 2808
rect 5776 2796 5782 2848
rect 6012 2836 6040 3003
rect 6380 2972 6408 3003
rect 6914 3000 6920 3012
rect 6972 3040 6978 3052
rect 8220 3049 8248 3080
rect 9398 3068 9404 3080
rect 9456 3068 9462 3120
rect 10152 3108 10180 3148
rect 10226 3136 10232 3188
rect 10284 3176 10290 3188
rect 14918 3176 14924 3188
rect 10284 3148 14924 3176
rect 10284 3136 10290 3148
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 15010 3136 15016 3188
rect 15068 3176 15074 3188
rect 15381 3179 15439 3185
rect 15381 3176 15393 3179
rect 15068 3148 15393 3176
rect 15068 3136 15074 3148
rect 15381 3145 15393 3148
rect 15427 3145 15439 3179
rect 15381 3139 15439 3145
rect 16485 3179 16543 3185
rect 16485 3145 16497 3179
rect 16531 3176 16543 3179
rect 18322 3176 18328 3188
rect 16531 3148 18328 3176
rect 16531 3145 16543 3148
rect 16485 3139 16543 3145
rect 18322 3136 18328 3148
rect 18380 3136 18386 3188
rect 12250 3108 12256 3120
rect 10152 3080 12256 3108
rect 12250 3068 12256 3080
rect 12308 3068 12314 3120
rect 12894 3068 12900 3120
rect 12952 3108 12958 3120
rect 13633 3111 13691 3117
rect 13633 3108 13645 3111
rect 12952 3080 13645 3108
rect 12952 3068 12958 3080
rect 13633 3077 13645 3080
rect 13679 3077 13691 3111
rect 13633 3071 13691 3077
rect 16022 3068 16028 3120
rect 16080 3108 16086 3120
rect 19150 3108 19156 3120
rect 16080 3080 19156 3108
rect 16080 3068 16086 3080
rect 19150 3068 19156 3080
rect 19208 3068 19214 3120
rect 7469 3043 7527 3049
rect 7469 3040 7481 3043
rect 6972 3012 7481 3040
rect 6972 3000 6978 3012
rect 7469 3009 7481 3012
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 8205 3043 8263 3049
rect 8205 3009 8217 3043
rect 8251 3009 8263 3043
rect 8205 3003 8263 3009
rect 8481 3043 8539 3049
rect 8481 3009 8493 3043
rect 8527 3040 8539 3043
rect 9030 3040 9036 3052
rect 8527 3012 9036 3040
rect 8527 3009 8539 3012
rect 8481 3003 8539 3009
rect 9030 3000 9036 3012
rect 9088 3000 9094 3052
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3040 10747 3043
rect 10870 3040 10876 3052
rect 10735 3012 10876 3040
rect 10735 3009 10747 3012
rect 10689 3003 10747 3009
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 11241 3043 11299 3049
rect 11241 3040 11253 3043
rect 11204 3012 11253 3040
rect 11204 3000 11210 3012
rect 11241 3009 11253 3012
rect 11287 3009 11299 3043
rect 11241 3003 11299 3009
rect 11330 3000 11336 3052
rect 11388 3040 11394 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11388 3012 11529 3040
rect 11388 3000 11394 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 13446 3040 13452 3052
rect 13407 3012 13452 3040
rect 11517 3003 11575 3009
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 15562 3040 15568 3052
rect 15523 3012 15568 3040
rect 15562 3000 15568 3012
rect 15620 3000 15626 3052
rect 15654 3000 15660 3052
rect 15712 3040 15718 3052
rect 15749 3043 15807 3049
rect 15749 3040 15761 3043
rect 15712 3012 15761 3040
rect 15712 3000 15718 3012
rect 15749 3009 15761 3012
rect 15795 3009 15807 3043
rect 16298 3040 16304 3052
rect 16259 3012 16304 3040
rect 15749 3003 15807 3009
rect 16298 3000 16304 3012
rect 16356 3000 16362 3052
rect 16761 3043 16819 3049
rect 16761 3009 16773 3043
rect 16807 3040 16819 3043
rect 16942 3040 16948 3052
rect 16807 3012 16948 3040
rect 16807 3009 16819 3012
rect 16761 3003 16819 3009
rect 16942 3000 16948 3012
rect 17000 3000 17006 3052
rect 17126 3040 17132 3052
rect 17087 3012 17132 3040
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 17494 3040 17500 3052
rect 17455 3012 17500 3040
rect 17494 3000 17500 3012
rect 17552 3000 17558 3052
rect 17862 3040 17868 3052
rect 17823 3012 17868 3040
rect 17862 3000 17868 3012
rect 17920 3000 17926 3052
rect 17954 3000 17960 3052
rect 18012 3040 18018 3052
rect 18233 3043 18291 3049
rect 18233 3040 18245 3043
rect 18012 3012 18245 3040
rect 18012 3000 18018 3012
rect 18233 3009 18245 3012
rect 18279 3009 18291 3043
rect 18233 3003 18291 3009
rect 7926 2972 7932 2984
rect 6380 2944 7932 2972
rect 7926 2932 7932 2944
rect 7984 2932 7990 2984
rect 9214 2972 9220 2984
rect 9175 2944 9220 2972
rect 9214 2932 9220 2944
rect 9272 2932 9278 2984
rect 9582 2932 9588 2984
rect 9640 2972 9646 2984
rect 10413 2975 10471 2981
rect 10413 2972 10425 2975
rect 9640 2944 10425 2972
rect 9640 2932 9646 2944
rect 10413 2941 10425 2944
rect 10459 2941 10471 2975
rect 10413 2935 10471 2941
rect 10597 2975 10655 2981
rect 10597 2941 10609 2975
rect 10643 2972 10655 2975
rect 10962 2972 10968 2984
rect 10643 2944 10968 2972
rect 10643 2941 10655 2944
rect 10597 2935 10655 2941
rect 10962 2932 10968 2944
rect 11020 2932 11026 2984
rect 11698 2932 11704 2984
rect 11756 2972 11762 2984
rect 11756 2944 11801 2972
rect 11756 2932 11762 2944
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12492 2944 12537 2972
rect 12492 2932 12498 2944
rect 13262 2932 13268 2984
rect 13320 2972 13326 2984
rect 13906 2972 13912 2984
rect 13320 2944 13912 2972
rect 13320 2932 13326 2944
rect 13906 2932 13912 2944
rect 13964 2932 13970 2984
rect 15102 2972 15108 2984
rect 15063 2944 15108 2972
rect 15102 2932 15108 2944
rect 15160 2932 15166 2984
rect 6181 2907 6239 2913
rect 6181 2873 6193 2907
rect 6227 2904 6239 2907
rect 6730 2904 6736 2916
rect 6227 2876 6736 2904
rect 6227 2873 6239 2876
rect 6181 2867 6239 2873
rect 6730 2864 6736 2876
rect 6788 2864 6794 2916
rect 6825 2907 6883 2913
rect 6825 2873 6837 2907
rect 6871 2904 6883 2907
rect 7282 2904 7288 2916
rect 6871 2876 7288 2904
rect 6871 2873 6883 2876
rect 6825 2867 6883 2873
rect 7282 2864 7288 2876
rect 7340 2864 7346 2916
rect 7374 2864 7380 2916
rect 7432 2904 7438 2916
rect 8021 2907 8079 2913
rect 8021 2904 8033 2907
rect 7432 2876 8033 2904
rect 7432 2864 7438 2876
rect 8021 2873 8033 2876
rect 8067 2873 8079 2907
rect 8021 2867 8079 2873
rect 8202 2864 8208 2916
rect 8260 2904 8266 2916
rect 10778 2904 10784 2916
rect 8260 2876 10784 2904
rect 8260 2864 8266 2876
rect 10778 2864 10784 2876
rect 10836 2904 10842 2916
rect 11146 2904 11152 2916
rect 10836 2876 10916 2904
rect 11107 2876 11152 2904
rect 10836 2864 10842 2876
rect 6914 2836 6920 2848
rect 6012 2808 6920 2836
rect 6914 2796 6920 2808
rect 6972 2796 6978 2848
rect 7098 2836 7104 2848
rect 7059 2808 7104 2836
rect 7098 2796 7104 2808
rect 7156 2796 7162 2848
rect 7466 2796 7472 2848
rect 7524 2836 7530 2848
rect 7561 2839 7619 2845
rect 7561 2836 7573 2839
rect 7524 2808 7573 2836
rect 7524 2796 7530 2808
rect 7561 2805 7573 2808
rect 7607 2805 7619 2839
rect 7561 2799 7619 2805
rect 8389 2839 8447 2845
rect 8389 2805 8401 2839
rect 8435 2836 8447 2839
rect 8478 2836 8484 2848
rect 8435 2808 8484 2836
rect 8435 2805 8447 2808
rect 8389 2799 8447 2805
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 8665 2839 8723 2845
rect 8665 2805 8677 2839
rect 8711 2836 8723 2839
rect 9030 2836 9036 2848
rect 8711 2808 9036 2836
rect 8711 2805 8723 2808
rect 8665 2799 8723 2805
rect 9030 2796 9036 2808
rect 9088 2796 9094 2848
rect 10888 2845 10916 2876
rect 11146 2864 11152 2876
rect 11204 2864 11210 2916
rect 12894 2904 12900 2916
rect 11624 2876 12900 2904
rect 10873 2839 10931 2845
rect 10873 2805 10885 2839
rect 10919 2805 10931 2839
rect 10873 2799 10931 2805
rect 11054 2796 11060 2848
rect 11112 2836 11118 2848
rect 11624 2836 11652 2876
rect 12894 2864 12900 2876
rect 12952 2864 12958 2916
rect 12986 2864 12992 2916
rect 13044 2904 13050 2916
rect 13538 2904 13544 2916
rect 13044 2876 13544 2904
rect 13044 2864 13050 2876
rect 13538 2864 13544 2876
rect 13596 2904 13602 2916
rect 15010 2904 15016 2916
rect 13596 2876 15016 2904
rect 13596 2864 13602 2876
rect 15010 2864 15016 2876
rect 15068 2864 15074 2916
rect 15838 2864 15844 2916
rect 15896 2904 15902 2916
rect 15933 2907 15991 2913
rect 15933 2904 15945 2907
rect 15896 2876 15945 2904
rect 15896 2864 15902 2876
rect 15933 2873 15945 2876
rect 15979 2873 15991 2907
rect 15933 2867 15991 2873
rect 16942 2836 16948 2848
rect 11112 2808 11652 2836
rect 16903 2808 16948 2836
rect 11112 2796 11118 2808
rect 16942 2796 16948 2808
rect 17000 2796 17006 2848
rect 17310 2836 17316 2848
rect 17271 2808 17316 2836
rect 17310 2796 17316 2808
rect 17368 2796 17374 2848
rect 17681 2839 17739 2845
rect 17681 2805 17693 2839
rect 17727 2836 17739 2839
rect 17770 2836 17776 2848
rect 17727 2808 17776 2836
rect 17727 2805 17739 2808
rect 17681 2799 17739 2805
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 17862 2796 17868 2848
rect 17920 2836 17926 2848
rect 18049 2839 18107 2845
rect 18049 2836 18061 2839
rect 17920 2808 18061 2836
rect 17920 2796 17926 2808
rect 18049 2805 18061 2808
rect 18095 2805 18107 2839
rect 18414 2836 18420 2848
rect 18375 2808 18420 2836
rect 18049 2799 18107 2805
rect 18414 2796 18420 2808
rect 18472 2796 18478 2848
rect 1104 2746 18860 2768
rect 1104 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 3430 2746
rect 3482 2694 7622 2746
rect 7674 2694 7686 2746
rect 7738 2694 7750 2746
rect 7802 2694 7814 2746
rect 7866 2694 7878 2746
rect 7930 2694 12070 2746
rect 12122 2694 12134 2746
rect 12186 2694 12198 2746
rect 12250 2694 12262 2746
rect 12314 2694 12326 2746
rect 12378 2694 16518 2746
rect 16570 2694 16582 2746
rect 16634 2694 16646 2746
rect 16698 2694 16710 2746
rect 16762 2694 16774 2746
rect 16826 2694 18860 2746
rect 1104 2672 18860 2694
rect 2314 2592 2320 2644
rect 2372 2632 2378 2644
rect 2593 2635 2651 2641
rect 2593 2632 2605 2635
rect 2372 2604 2605 2632
rect 2372 2592 2378 2604
rect 2593 2601 2605 2604
rect 2639 2601 2651 2635
rect 4706 2632 4712 2644
rect 4667 2604 4712 2632
rect 2593 2595 2651 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 5902 2632 5908 2644
rect 5863 2604 5908 2632
rect 5902 2592 5908 2604
rect 5960 2592 5966 2644
rect 10962 2592 10968 2644
rect 11020 2632 11026 2644
rect 11793 2635 11851 2641
rect 11793 2632 11805 2635
rect 11020 2604 11805 2632
rect 11020 2592 11026 2604
rect 11793 2601 11805 2604
rect 11839 2601 11851 2635
rect 12526 2632 12532 2644
rect 12487 2604 12532 2632
rect 11793 2595 11851 2601
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 12802 2592 12808 2644
rect 12860 2632 12866 2644
rect 13265 2635 13323 2641
rect 13265 2632 13277 2635
rect 12860 2604 13277 2632
rect 12860 2592 12866 2604
rect 13265 2601 13277 2604
rect 13311 2601 13323 2635
rect 13265 2595 13323 2601
rect 15102 2592 15108 2644
rect 15160 2632 15166 2644
rect 16393 2635 16451 2641
rect 16393 2632 16405 2635
rect 15160 2604 16405 2632
rect 15160 2592 15166 2604
rect 16393 2601 16405 2604
rect 16439 2601 16451 2635
rect 18966 2632 18972 2644
rect 16393 2595 16451 2601
rect 16500 2604 18972 2632
rect 2498 2564 2504 2576
rect 1688 2536 2504 2564
rect 1688 2437 1716 2536
rect 2498 2524 2504 2536
rect 2556 2524 2562 2576
rect 3878 2524 3884 2576
rect 3936 2564 3942 2576
rect 4985 2567 5043 2573
rect 4985 2564 4997 2567
rect 3936 2536 4997 2564
rect 3936 2524 3942 2536
rect 4985 2533 4997 2536
rect 5031 2533 5043 2567
rect 4985 2527 5043 2533
rect 10226 2524 10232 2576
rect 10284 2564 10290 2576
rect 11241 2567 11299 2573
rect 11241 2564 11253 2567
rect 10284 2536 11253 2564
rect 10284 2524 10290 2536
rect 11241 2533 11253 2536
rect 11287 2533 11299 2567
rect 11241 2527 11299 2533
rect 11517 2567 11575 2573
rect 11517 2533 11529 2567
rect 11563 2533 11575 2567
rect 15654 2564 15660 2576
rect 11517 2527 11575 2533
rect 11716 2536 15660 2564
rect 3970 2496 3976 2508
rect 2056 2468 3976 2496
rect 2056 2437 2084 2468
rect 3970 2456 3976 2468
rect 4028 2456 4034 2508
rect 4614 2456 4620 2508
rect 4672 2496 4678 2508
rect 8202 2496 8208 2508
rect 4672 2468 4936 2496
rect 4672 2456 4678 2468
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2397 1731 2431
rect 1673 2391 1731 2397
rect 2041 2431 2099 2437
rect 2041 2397 2053 2431
rect 2087 2397 2099 2431
rect 2041 2391 2099 2397
rect 2501 2431 2559 2437
rect 2501 2397 2513 2431
rect 2547 2397 2559 2431
rect 2501 2391 2559 2397
rect 2516 2360 2544 2391
rect 2682 2388 2688 2440
rect 2740 2428 2746 2440
rect 2777 2431 2835 2437
rect 2777 2428 2789 2431
rect 2740 2400 2789 2428
rect 2740 2388 2746 2400
rect 2777 2397 2789 2400
rect 2823 2397 2835 2431
rect 3510 2428 3516 2440
rect 3471 2400 3516 2428
rect 2777 2391 2835 2397
rect 3510 2388 3516 2400
rect 3568 2388 3574 2440
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2428 4123 2431
rect 4246 2428 4252 2440
rect 4111 2400 4252 2428
rect 4111 2397 4123 2400
rect 4065 2391 4123 2397
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2428 4583 2431
rect 4798 2428 4804 2440
rect 4571 2400 4804 2428
rect 4571 2397 4583 2400
rect 4525 2391 4583 2397
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 4908 2437 4936 2468
rect 5552 2468 8208 2496
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 5166 2428 5172 2440
rect 5127 2400 5172 2428
rect 4893 2391 4951 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5552 2437 5580 2468
rect 8202 2456 8208 2468
rect 8260 2456 8266 2508
rect 9766 2496 9772 2508
rect 9727 2468 9772 2496
rect 9766 2456 9772 2468
rect 9824 2456 9830 2508
rect 9953 2499 10011 2505
rect 9953 2465 9965 2499
rect 9999 2496 10011 2499
rect 10318 2496 10324 2508
rect 9999 2468 10324 2496
rect 9999 2465 10011 2468
rect 9953 2459 10011 2465
rect 10318 2456 10324 2468
rect 10376 2456 10382 2508
rect 11532 2496 11560 2527
rect 10888 2468 11560 2496
rect 5537 2431 5595 2437
rect 5537 2397 5549 2431
rect 5583 2397 5595 2431
rect 5718 2428 5724 2440
rect 5679 2400 5724 2428
rect 5537 2391 5595 2397
rect 5718 2388 5724 2400
rect 5776 2388 5782 2440
rect 6638 2428 6644 2440
rect 6599 2400 6644 2428
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 7190 2428 7196 2440
rect 6788 2400 6833 2428
rect 7151 2400 7196 2428
rect 6788 2388 6794 2400
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 7282 2388 7288 2440
rect 7340 2428 7346 2440
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 7340 2400 7757 2428
rect 7340 2388 7346 2400
rect 7745 2397 7757 2400
rect 7791 2397 7803 2431
rect 8386 2428 8392 2440
rect 8347 2400 8392 2428
rect 7745 2391 7803 2397
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 8478 2388 8484 2440
rect 8536 2428 8542 2440
rect 9030 2428 9036 2440
rect 8536 2400 8581 2428
rect 8991 2400 9036 2428
rect 8536 2388 8542 2400
rect 9030 2388 9036 2400
rect 9088 2388 9094 2440
rect 9674 2428 9680 2440
rect 9635 2400 9680 2428
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 10594 2388 10600 2440
rect 10652 2388 10658 2440
rect 10888 2424 10916 2468
rect 10965 2431 11023 2437
rect 10965 2424 10977 2431
rect 10888 2397 10977 2424
rect 11011 2397 11023 2431
rect 10888 2396 11023 2397
rect 10965 2391 11023 2396
rect 11057 2431 11115 2437
rect 11057 2397 11069 2431
rect 11103 2397 11115 2431
rect 11057 2391 11115 2397
rect 2866 2360 2872 2372
rect 2516 2332 2872 2360
rect 2866 2320 2872 2332
rect 2924 2320 2930 2372
rect 10410 2360 10416 2372
rect 10371 2332 10416 2360
rect 10410 2320 10416 2332
rect 10468 2320 10474 2372
rect 10612 2360 10640 2388
rect 11072 2360 11100 2391
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11716 2437 11744 2536
rect 15654 2524 15660 2536
rect 15712 2524 15718 2576
rect 16500 2564 16528 2604
rect 18966 2592 18972 2604
rect 19024 2592 19030 2644
rect 15948 2536 16528 2564
rect 12342 2496 12348 2508
rect 12303 2468 12348 2496
rect 12342 2456 12348 2468
rect 12400 2456 12406 2508
rect 12618 2456 12624 2508
rect 12676 2496 12682 2508
rect 14090 2496 14096 2508
rect 12676 2468 13676 2496
rect 14051 2468 14096 2496
rect 12676 2456 12682 2468
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11204 2400 11713 2428
rect 11204 2388 11210 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 11882 2388 11888 2440
rect 11940 2428 11946 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11940 2400 11989 2428
rect 11940 2388 11946 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12161 2431 12219 2437
rect 12161 2397 12173 2431
rect 12207 2397 12219 2431
rect 12161 2391 12219 2397
rect 10612 2332 11100 2360
rect 1486 2292 1492 2304
rect 1447 2264 1492 2292
rect 1486 2252 1492 2264
rect 1544 2252 1550 2304
rect 1670 2252 1676 2304
rect 1728 2292 1734 2304
rect 1857 2295 1915 2301
rect 1857 2292 1869 2295
rect 1728 2264 1869 2292
rect 1728 2252 1734 2264
rect 1857 2261 1869 2264
rect 1903 2261 1915 2295
rect 1857 2255 1915 2261
rect 2130 2252 2136 2304
rect 2188 2292 2194 2304
rect 2317 2295 2375 2301
rect 2317 2292 2329 2295
rect 2188 2264 2329 2292
rect 2188 2252 2194 2264
rect 2317 2261 2329 2264
rect 2363 2261 2375 2295
rect 2317 2255 2375 2261
rect 2682 2252 2688 2304
rect 2740 2292 2746 2304
rect 2961 2295 3019 2301
rect 2961 2292 2973 2295
rect 2740 2264 2973 2292
rect 2740 2252 2746 2264
rect 2961 2261 2973 2264
rect 3007 2261 3019 2295
rect 2961 2255 3019 2261
rect 3142 2252 3148 2304
rect 3200 2292 3206 2304
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 3200 2264 3341 2292
rect 3200 2252 3206 2264
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3329 2255 3387 2261
rect 3602 2252 3608 2304
rect 3660 2292 3666 2304
rect 3881 2295 3939 2301
rect 3881 2292 3893 2295
rect 3660 2264 3893 2292
rect 3660 2252 3666 2264
rect 3881 2261 3893 2264
rect 3927 2261 3939 2295
rect 3881 2255 3939 2261
rect 4154 2252 4160 2304
rect 4212 2292 4218 2304
rect 4341 2295 4399 2301
rect 4341 2292 4353 2295
rect 4212 2264 4353 2292
rect 4212 2252 4218 2264
rect 4341 2261 4353 2264
rect 4387 2261 4399 2295
rect 4341 2255 4399 2261
rect 5166 2252 5172 2304
rect 5224 2292 5230 2304
rect 5353 2295 5411 2301
rect 5353 2292 5365 2295
rect 5224 2264 5365 2292
rect 5224 2252 5230 2264
rect 5353 2261 5365 2264
rect 5399 2261 5411 2295
rect 6086 2292 6092 2304
rect 6047 2264 6092 2292
rect 5353 2255 5411 2261
rect 6086 2252 6092 2264
rect 6144 2252 6150 2304
rect 6178 2252 6184 2304
rect 6236 2292 6242 2304
rect 6457 2295 6515 2301
rect 6457 2292 6469 2295
rect 6236 2264 6469 2292
rect 6236 2252 6242 2264
rect 6457 2261 6469 2264
rect 6503 2261 6515 2295
rect 6457 2255 6515 2261
rect 6638 2252 6644 2304
rect 6696 2292 6702 2304
rect 6917 2295 6975 2301
rect 6917 2292 6929 2295
rect 6696 2264 6929 2292
rect 6696 2252 6702 2264
rect 6917 2261 6929 2264
rect 6963 2261 6975 2295
rect 6917 2255 6975 2261
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7377 2295 7435 2301
rect 7377 2292 7389 2295
rect 7156 2264 7389 2292
rect 7156 2252 7162 2264
rect 7377 2261 7389 2264
rect 7423 2261 7435 2295
rect 7558 2292 7564 2304
rect 7519 2264 7564 2292
rect 7377 2255 7435 2261
rect 7558 2252 7564 2264
rect 7616 2252 7622 2304
rect 7650 2252 7656 2304
rect 7708 2292 7714 2304
rect 7929 2295 7987 2301
rect 7929 2292 7941 2295
rect 7708 2264 7941 2292
rect 7708 2252 7714 2264
rect 7929 2261 7941 2264
rect 7975 2261 7987 2295
rect 7929 2255 7987 2261
rect 8110 2252 8116 2304
rect 8168 2292 8174 2304
rect 8205 2295 8263 2301
rect 8205 2292 8217 2295
rect 8168 2264 8217 2292
rect 8168 2252 8174 2264
rect 8205 2261 8217 2264
rect 8251 2261 8263 2295
rect 8662 2292 8668 2304
rect 8623 2264 8668 2292
rect 8205 2255 8263 2261
rect 8662 2252 8668 2264
rect 8720 2252 8726 2304
rect 9122 2252 9128 2304
rect 9180 2292 9186 2304
rect 9217 2295 9275 2301
rect 9217 2292 9229 2295
rect 9180 2264 9229 2292
rect 9180 2252 9186 2264
rect 9217 2261 9229 2264
rect 9263 2261 9275 2295
rect 9217 2255 9275 2261
rect 9493 2295 9551 2301
rect 9493 2261 9505 2295
rect 9539 2292 9551 2295
rect 9674 2292 9680 2304
rect 9539 2264 9680 2292
rect 9539 2261 9551 2264
rect 9493 2255 9551 2261
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 10502 2292 10508 2304
rect 10463 2264 10508 2292
rect 10502 2252 10508 2264
rect 10560 2252 10566 2304
rect 10594 2252 10600 2304
rect 10652 2292 10658 2304
rect 10781 2295 10839 2301
rect 10781 2292 10793 2295
rect 10652 2264 10793 2292
rect 10652 2252 10658 2264
rect 10781 2261 10793 2264
rect 10827 2261 10839 2295
rect 10781 2255 10839 2261
rect 10870 2252 10876 2304
rect 10928 2292 10934 2304
rect 12176 2292 12204 2391
rect 12894 2388 12900 2440
rect 12952 2428 12958 2440
rect 13024 2431 13082 2437
rect 13024 2428 13036 2431
rect 12952 2400 13036 2428
rect 12952 2388 12958 2400
rect 13024 2397 13036 2400
rect 13070 2428 13082 2431
rect 13262 2428 13268 2440
rect 13070 2400 13268 2428
rect 13070 2397 13082 2400
rect 13024 2391 13082 2397
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 13446 2428 13452 2440
rect 13407 2400 13452 2428
rect 13446 2388 13452 2400
rect 13504 2388 13510 2440
rect 13648 2437 13676 2468
rect 14090 2456 14096 2468
rect 14148 2456 14154 2508
rect 15948 2505 15976 2536
rect 16666 2524 16672 2576
rect 16724 2564 16730 2576
rect 16853 2567 16911 2573
rect 16853 2564 16865 2567
rect 16724 2536 16865 2564
rect 16724 2524 16730 2536
rect 16853 2533 16865 2536
rect 16899 2533 16911 2567
rect 16853 2527 16911 2533
rect 17126 2524 17132 2576
rect 17184 2564 17190 2576
rect 17589 2567 17647 2573
rect 17589 2564 17601 2567
rect 17184 2536 17601 2564
rect 17184 2524 17190 2536
rect 17589 2533 17601 2536
rect 17635 2533 17647 2567
rect 17589 2527 17647 2533
rect 15933 2499 15991 2505
rect 15933 2465 15945 2499
rect 15979 2465 15991 2499
rect 15933 2459 15991 2465
rect 13633 2431 13691 2437
rect 13633 2397 13645 2431
rect 13679 2397 13691 2431
rect 16022 2428 16028 2440
rect 15983 2400 16028 2428
rect 13633 2391 13691 2397
rect 16022 2388 16028 2400
rect 16080 2388 16086 2440
rect 16666 2388 16672 2440
rect 16724 2428 16730 2440
rect 16724 2400 16769 2428
rect 16724 2388 16730 2400
rect 16850 2388 16856 2440
rect 16908 2428 16914 2440
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 16908 2400 17049 2428
rect 16908 2388 16914 2400
rect 17037 2397 17049 2400
rect 17083 2397 17095 2431
rect 17037 2391 17095 2397
rect 17218 2388 17224 2440
rect 17276 2428 17282 2440
rect 17405 2431 17463 2437
rect 17405 2428 17417 2431
rect 17276 2400 17417 2428
rect 17276 2388 17282 2400
rect 17405 2397 17417 2400
rect 17451 2397 17463 2431
rect 17405 2391 17463 2397
rect 17494 2388 17500 2440
rect 17552 2428 17558 2440
rect 17773 2431 17831 2437
rect 17773 2428 17785 2431
rect 17552 2400 17785 2428
rect 17552 2388 17558 2400
rect 17773 2397 17785 2400
rect 17819 2397 17831 2431
rect 18230 2428 18236 2440
rect 18191 2400 18236 2428
rect 17773 2391 17831 2397
rect 18230 2388 18236 2400
rect 18288 2388 18294 2440
rect 13127 2363 13185 2369
rect 13127 2329 13139 2363
rect 13173 2360 13185 2363
rect 14277 2363 14335 2369
rect 14277 2360 14289 2363
rect 13173 2332 14289 2360
rect 13173 2329 13185 2332
rect 13127 2323 13185 2329
rect 14277 2329 14289 2332
rect 14323 2329 14335 2363
rect 14277 2323 14335 2329
rect 16684 2332 17264 2360
rect 16684 2304 16712 2332
rect 10928 2264 12204 2292
rect 13817 2295 13875 2301
rect 10928 2252 10934 2264
rect 13817 2261 13829 2295
rect 13863 2292 13875 2295
rect 15194 2292 15200 2304
rect 13863 2264 15200 2292
rect 13863 2261 13875 2264
rect 13817 2255 13875 2261
rect 15194 2252 15200 2264
rect 15252 2252 15258 2304
rect 15654 2252 15660 2304
rect 15712 2292 15718 2304
rect 16209 2295 16267 2301
rect 16209 2292 16221 2295
rect 15712 2264 16221 2292
rect 15712 2252 15718 2264
rect 16209 2261 16221 2264
rect 16255 2261 16267 2295
rect 16209 2255 16267 2261
rect 16666 2252 16672 2304
rect 16724 2252 16730 2304
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 17034 2292 17040 2304
rect 16816 2264 17040 2292
rect 16816 2252 16822 2264
rect 17034 2252 17040 2264
rect 17092 2252 17098 2304
rect 17236 2301 17264 2332
rect 17221 2295 17279 2301
rect 17221 2261 17233 2295
rect 17267 2261 17279 2295
rect 17221 2255 17279 2261
rect 17678 2252 17684 2304
rect 17736 2292 17742 2304
rect 17957 2295 18015 2301
rect 17957 2292 17969 2295
rect 17736 2264 17969 2292
rect 17736 2252 17742 2264
rect 17957 2261 17969 2264
rect 18003 2261 18015 2295
rect 17957 2255 18015 2261
rect 18138 2252 18144 2304
rect 18196 2292 18202 2304
rect 18417 2295 18475 2301
rect 18417 2292 18429 2295
rect 18196 2264 18429 2292
rect 18196 2252 18202 2264
rect 18417 2261 18429 2264
rect 18463 2261 18475 2295
rect 18417 2255 18475 2261
rect 1104 2202 18860 2224
rect 1104 2150 5398 2202
rect 5450 2150 5462 2202
rect 5514 2150 5526 2202
rect 5578 2150 5590 2202
rect 5642 2150 5654 2202
rect 5706 2150 9846 2202
rect 9898 2150 9910 2202
rect 9962 2150 9974 2202
rect 10026 2150 10038 2202
rect 10090 2150 10102 2202
rect 10154 2150 14294 2202
rect 14346 2150 14358 2202
rect 14410 2150 14422 2202
rect 14474 2150 14486 2202
rect 14538 2150 14550 2202
rect 14602 2150 18860 2202
rect 1104 2128 18860 2150
rect 10502 2048 10508 2100
rect 10560 2088 10566 2100
rect 12618 2088 12624 2100
rect 10560 2060 12624 2088
rect 10560 2048 10566 2060
rect 12618 2048 12624 2060
rect 12676 2048 12682 2100
rect 15378 2048 15384 2100
rect 15436 2088 15442 2100
rect 18230 2088 18236 2100
rect 15436 2060 18236 2088
rect 15436 2048 15442 2060
rect 18230 2048 18236 2060
rect 18288 2048 18294 2100
rect 6086 1980 6092 2032
rect 6144 2020 6150 2032
rect 13170 2020 13176 2032
rect 6144 1992 13176 2020
rect 6144 1980 6150 1992
rect 13170 1980 13176 1992
rect 13228 2020 13234 2032
rect 13446 2020 13452 2032
rect 13228 1992 13452 2020
rect 13228 1980 13234 1992
rect 13446 1980 13452 1992
rect 13504 1980 13510 2032
rect 13630 1980 13636 2032
rect 13688 2020 13694 2032
rect 17494 2020 17500 2032
rect 13688 1992 17500 2020
rect 13688 1980 13694 1992
rect 17494 1980 17500 1992
rect 17552 1980 17558 2032
rect 7558 1912 7564 1964
rect 7616 1952 7622 1964
rect 11146 1952 11152 1964
rect 7616 1924 11152 1952
rect 7616 1912 7622 1924
rect 11146 1912 11152 1924
rect 11204 1952 11210 1964
rect 11882 1952 11888 1964
rect 11204 1924 11888 1952
rect 11204 1912 11210 1924
rect 11882 1912 11888 1924
rect 11940 1912 11946 1964
rect 13814 1844 13820 1896
rect 13872 1884 13878 1896
rect 16850 1884 16856 1896
rect 13872 1856 16856 1884
rect 13872 1844 13878 1856
rect 16850 1844 16856 1856
rect 16908 1844 16914 1896
rect 10410 1776 10416 1828
rect 10468 1816 10474 1828
rect 12986 1816 12992 1828
rect 10468 1788 12992 1816
rect 10468 1776 10474 1788
rect 12986 1776 12992 1788
rect 13044 1776 13050 1828
rect 11238 1708 11244 1760
rect 11296 1748 11302 1760
rect 16022 1748 16028 1760
rect 11296 1720 16028 1748
rect 11296 1708 11302 1720
rect 16022 1708 16028 1720
rect 16080 1708 16086 1760
<< via1 >>
rect 15936 16056 15988 16108
rect 16396 16056 16448 16108
rect 3792 15172 3844 15224
rect 5540 15172 5592 15224
rect 4436 15036 4488 15088
rect 3608 14968 3660 15020
rect 7288 14968 7340 15020
rect 14188 14968 14240 15020
rect 3884 14900 3936 14952
rect 5080 14900 5132 14952
rect 5172 14900 5224 14952
rect 15200 14900 15252 14952
rect 3700 14832 3752 14884
rect 6644 14832 6696 14884
rect 9128 14832 9180 14884
rect 17040 14832 17092 14884
rect 1216 14764 1268 14816
rect 4068 14764 4120 14816
rect 4160 14764 4212 14816
rect 7472 14764 7524 14816
rect 8116 14764 8168 14816
rect 17960 14764 18012 14816
rect 3174 14662 3226 14714
rect 3238 14662 3290 14714
rect 3302 14662 3354 14714
rect 3366 14662 3418 14714
rect 3430 14662 3482 14714
rect 7622 14662 7674 14714
rect 7686 14662 7738 14714
rect 7750 14662 7802 14714
rect 7814 14662 7866 14714
rect 7878 14662 7930 14714
rect 12070 14662 12122 14714
rect 12134 14662 12186 14714
rect 12198 14662 12250 14714
rect 12262 14662 12314 14714
rect 12326 14662 12378 14714
rect 16518 14662 16570 14714
rect 16582 14662 16634 14714
rect 16646 14662 16698 14714
rect 16710 14662 16762 14714
rect 16774 14662 16826 14714
rect 3516 14560 3568 14612
rect 5448 14560 5500 14612
rect 5816 14560 5868 14612
rect 4068 14492 4120 14544
rect 6920 14560 6972 14612
rect 7380 14603 7432 14612
rect 7380 14569 7389 14603
rect 7389 14569 7423 14603
rect 7423 14569 7432 14603
rect 7380 14560 7432 14569
rect 7472 14560 7524 14612
rect 8668 14603 8720 14612
rect 8668 14569 8677 14603
rect 8677 14569 8711 14603
rect 8711 14569 8720 14603
rect 8668 14560 8720 14569
rect 9312 14603 9364 14612
rect 9312 14569 9321 14603
rect 9321 14569 9355 14603
rect 9355 14569 9364 14603
rect 9312 14560 9364 14569
rect 9956 14603 10008 14612
rect 9956 14569 9965 14603
rect 9965 14569 9999 14603
rect 9999 14569 10008 14603
rect 9956 14560 10008 14569
rect 10600 14603 10652 14612
rect 10600 14569 10609 14603
rect 10609 14569 10643 14603
rect 10643 14569 10652 14603
rect 10600 14560 10652 14569
rect 11888 14560 11940 14612
rect 8208 14535 8260 14544
rect 8208 14501 8217 14535
rect 8217 14501 8251 14535
rect 8251 14501 8260 14535
rect 8208 14492 8260 14501
rect 11980 14492 12032 14544
rect 2688 14424 2740 14476
rect 2964 14424 3016 14476
rect 3700 14424 3752 14476
rect 4160 14424 4212 14476
rect 5724 14424 5776 14476
rect 2228 14399 2280 14408
rect 2228 14365 2237 14399
rect 2237 14365 2271 14399
rect 2271 14365 2280 14399
rect 2228 14356 2280 14365
rect 3424 14288 3476 14340
rect 4528 14356 4580 14408
rect 5540 14399 5592 14408
rect 5540 14365 5549 14399
rect 5549 14365 5583 14399
rect 5583 14365 5592 14399
rect 5540 14356 5592 14365
rect 6000 14399 6052 14408
rect 6000 14365 6009 14399
rect 6009 14365 6043 14399
rect 6043 14365 6052 14399
rect 6000 14356 6052 14365
rect 6184 14356 6236 14408
rect 6552 14356 6604 14408
rect 7380 14356 7432 14408
rect 8668 14356 8720 14408
rect 9312 14356 9364 14408
rect 9956 14356 10008 14408
rect 10600 14356 10652 14408
rect 11520 14399 11572 14408
rect 11520 14365 11529 14399
rect 11529 14365 11563 14399
rect 11563 14365 11572 14399
rect 12532 14603 12584 14612
rect 12532 14569 12541 14603
rect 12541 14569 12575 14603
rect 12575 14569 12584 14603
rect 12532 14560 12584 14569
rect 13176 14603 13228 14612
rect 13176 14569 13185 14603
rect 13185 14569 13219 14603
rect 13219 14569 13228 14603
rect 13176 14560 13228 14569
rect 13268 14560 13320 14612
rect 12348 14492 12400 14544
rect 15844 14492 15896 14544
rect 16488 14492 16540 14544
rect 17408 14424 17460 14476
rect 17960 14467 18012 14476
rect 17960 14433 17969 14467
rect 17969 14433 18003 14467
rect 18003 14433 18012 14467
rect 17960 14424 18012 14433
rect 11520 14356 11572 14365
rect 12532 14356 12584 14408
rect 13176 14356 13228 14408
rect 13820 14356 13872 14408
rect 14832 14356 14884 14408
rect 15568 14399 15620 14408
rect 15568 14365 15577 14399
rect 15577 14365 15611 14399
rect 15611 14365 15620 14399
rect 15568 14356 15620 14365
rect 16028 14356 16080 14408
rect 15660 14288 15712 14340
rect 16120 14288 16172 14340
rect 17684 14399 17736 14408
rect 17684 14365 17693 14399
rect 17693 14365 17727 14399
rect 17727 14365 17736 14399
rect 17684 14356 17736 14365
rect 5724 14220 5776 14272
rect 6460 14220 6512 14272
rect 7196 14220 7248 14272
rect 8852 14220 8904 14272
rect 9772 14220 9824 14272
rect 10692 14220 10744 14272
rect 10876 14263 10928 14272
rect 10876 14229 10885 14263
rect 10885 14229 10919 14263
rect 10919 14229 10928 14263
rect 10876 14220 10928 14229
rect 11888 14220 11940 14272
rect 12808 14263 12860 14272
rect 12808 14229 12817 14263
rect 12817 14229 12851 14263
rect 12851 14229 12860 14263
rect 12808 14220 12860 14229
rect 13452 14263 13504 14272
rect 13452 14229 13461 14263
rect 13461 14229 13495 14263
rect 13495 14229 13504 14263
rect 13452 14220 13504 14229
rect 15108 14220 15160 14272
rect 15752 14220 15804 14272
rect 16488 14220 16540 14272
rect 5398 14118 5450 14170
rect 5462 14118 5514 14170
rect 5526 14118 5578 14170
rect 5590 14118 5642 14170
rect 5654 14118 5706 14170
rect 9846 14118 9898 14170
rect 9910 14118 9962 14170
rect 9974 14118 10026 14170
rect 10038 14118 10090 14170
rect 10102 14118 10154 14170
rect 14294 14118 14346 14170
rect 14358 14118 14410 14170
rect 14422 14118 14474 14170
rect 14486 14118 14538 14170
rect 14550 14118 14602 14170
rect 4160 14016 4212 14068
rect 4344 14059 4396 14068
rect 4344 14025 4353 14059
rect 4353 14025 4387 14059
rect 4387 14025 4396 14059
rect 4344 14016 4396 14025
rect 4804 14016 4856 14068
rect 4068 13948 4120 14000
rect 3608 13880 3660 13932
rect 3976 13880 4028 13932
rect 4436 13880 4488 13932
rect 4804 13923 4856 13932
rect 4804 13889 4813 13923
rect 4813 13889 4847 13923
rect 4847 13889 4856 13923
rect 4804 13880 4856 13889
rect 5172 13923 5224 13932
rect 5172 13889 5181 13923
rect 5181 13889 5215 13923
rect 5215 13889 5224 13923
rect 5172 13880 5224 13889
rect 5540 13923 5592 13932
rect 5540 13889 5549 13923
rect 5549 13889 5583 13923
rect 5583 13889 5592 13923
rect 5540 13880 5592 13889
rect 6552 14059 6604 14068
rect 6552 14025 6561 14059
rect 6561 14025 6595 14059
rect 6595 14025 6604 14059
rect 6552 14016 6604 14025
rect 6644 14016 6696 14068
rect 9312 14016 9364 14068
rect 13268 14016 13320 14068
rect 5724 13948 5776 14000
rect 14188 14016 14240 14068
rect 15568 14016 15620 14068
rect 6184 13923 6236 13932
rect 6184 13889 6193 13923
rect 6193 13889 6227 13923
rect 6227 13889 6236 13923
rect 6184 13880 6236 13889
rect 6276 13880 6328 13932
rect 6460 13880 6512 13932
rect 7012 13923 7064 13932
rect 7012 13889 7021 13923
rect 7021 13889 7055 13923
rect 7055 13889 7064 13923
rect 7380 13923 7432 13932
rect 7012 13880 7064 13889
rect 2044 13812 2096 13864
rect 2780 13812 2832 13864
rect 3700 13812 3752 13864
rect 3884 13812 3936 13864
rect 1584 13744 1636 13796
rect 3976 13744 4028 13796
rect 6000 13812 6052 13864
rect 7380 13889 7389 13923
rect 7389 13889 7423 13923
rect 7423 13889 7432 13923
rect 7380 13880 7432 13889
rect 8208 13880 8260 13932
rect 14832 13948 14884 14000
rect 9128 13812 9180 13864
rect 11612 13812 11664 13864
rect 12348 13812 12400 13864
rect 14924 13880 14976 13932
rect 14740 13812 14792 13864
rect 15016 13812 15068 13864
rect 296 13676 348 13728
rect 6736 13744 6788 13796
rect 8116 13744 8168 13796
rect 4436 13676 4488 13728
rect 5080 13676 5132 13728
rect 6552 13676 6604 13728
rect 6644 13719 6696 13728
rect 6644 13685 6653 13719
rect 6653 13685 6687 13719
rect 6687 13685 6696 13719
rect 15384 13880 15436 13932
rect 15844 13880 15896 13932
rect 16304 13880 16356 13932
rect 16856 13880 16908 13932
rect 15200 13812 15252 13864
rect 16304 13744 16356 13796
rect 17040 13855 17092 13864
rect 17040 13821 17049 13855
rect 17049 13821 17083 13855
rect 17083 13821 17092 13855
rect 17040 13812 17092 13821
rect 17684 13855 17736 13864
rect 17684 13821 17693 13855
rect 17693 13821 17727 13855
rect 17727 13821 17736 13855
rect 17684 13812 17736 13821
rect 18052 13812 18104 13864
rect 6644 13676 6696 13685
rect 16028 13676 16080 13728
rect 3174 13574 3226 13626
rect 3238 13574 3290 13626
rect 3302 13574 3354 13626
rect 3366 13574 3418 13626
rect 3430 13574 3482 13626
rect 7622 13574 7674 13626
rect 7686 13574 7738 13626
rect 7750 13574 7802 13626
rect 7814 13574 7866 13626
rect 7878 13574 7930 13626
rect 12070 13574 12122 13626
rect 12134 13574 12186 13626
rect 12198 13574 12250 13626
rect 12262 13574 12314 13626
rect 12326 13574 12378 13626
rect 16518 13574 16570 13626
rect 16582 13574 16634 13626
rect 16646 13574 16698 13626
rect 16710 13574 16762 13626
rect 16774 13574 16826 13626
rect 2872 13472 2924 13524
rect 5540 13472 5592 13524
rect 15660 13472 15712 13524
rect 16120 13472 16172 13524
rect 16856 13472 16908 13524
rect 2504 13336 2556 13388
rect 1952 13311 2004 13320
rect 1952 13277 1961 13311
rect 1961 13277 1995 13311
rect 1995 13277 2004 13311
rect 1952 13268 2004 13277
rect 2228 13311 2280 13320
rect 2228 13277 2237 13311
rect 2237 13277 2271 13311
rect 2271 13277 2280 13311
rect 2228 13268 2280 13277
rect 2964 13268 3016 13320
rect 3240 13268 3292 13320
rect 2228 13132 2280 13184
rect 3608 13336 3660 13388
rect 4160 13336 4212 13388
rect 6552 13404 6604 13456
rect 16304 13447 16356 13456
rect 16304 13413 16313 13447
rect 16313 13413 16347 13447
rect 16347 13413 16356 13447
rect 16304 13404 16356 13413
rect 4436 13268 4488 13320
rect 16396 13336 16448 13388
rect 15936 13311 15988 13320
rect 3792 13200 3844 13252
rect 4344 13200 4396 13252
rect 5080 13200 5132 13252
rect 3516 13132 3568 13184
rect 3884 13132 3936 13184
rect 4252 13132 4304 13184
rect 5172 13132 5224 13184
rect 5264 13175 5316 13184
rect 5264 13141 5273 13175
rect 5273 13141 5307 13175
rect 5307 13141 5316 13175
rect 15936 13277 15945 13311
rect 15945 13277 15979 13311
rect 15979 13277 15988 13311
rect 15936 13268 15988 13277
rect 17224 13268 17276 13320
rect 17684 13311 17736 13320
rect 17684 13277 17693 13311
rect 17693 13277 17727 13311
rect 17727 13277 17736 13311
rect 17684 13268 17736 13277
rect 6368 13243 6420 13252
rect 6368 13209 6377 13243
rect 6377 13209 6411 13243
rect 6411 13209 6420 13243
rect 6368 13200 6420 13209
rect 15200 13200 15252 13252
rect 5264 13132 5316 13141
rect 17408 13132 17460 13184
rect 5398 13030 5450 13082
rect 5462 13030 5514 13082
rect 5526 13030 5578 13082
rect 5590 13030 5642 13082
rect 5654 13030 5706 13082
rect 9846 13030 9898 13082
rect 9910 13030 9962 13082
rect 9974 13030 10026 13082
rect 10038 13030 10090 13082
rect 10102 13030 10154 13082
rect 14294 13030 14346 13082
rect 14358 13030 14410 13082
rect 14422 13030 14474 13082
rect 14486 13030 14538 13082
rect 14550 13030 14602 13082
rect 2136 12724 2188 12776
rect 2228 12767 2280 12776
rect 2228 12733 2237 12767
rect 2237 12733 2271 12767
rect 2271 12733 2280 12767
rect 3148 12835 3200 12844
rect 3148 12801 3157 12835
rect 3157 12801 3191 12835
rect 3191 12801 3200 12835
rect 3148 12792 3200 12801
rect 3424 12860 3476 12912
rect 3608 12903 3660 12912
rect 3608 12869 3642 12903
rect 3642 12869 3660 12903
rect 4068 12928 4120 12980
rect 4988 12928 5040 12980
rect 5172 12971 5224 12980
rect 5172 12937 5181 12971
rect 5181 12937 5215 12971
rect 5215 12937 5224 12971
rect 5172 12928 5224 12937
rect 5908 12971 5960 12980
rect 5908 12937 5917 12971
rect 5917 12937 5951 12971
rect 5951 12937 5960 12971
rect 5908 12928 5960 12937
rect 16396 12928 16448 12980
rect 3608 12860 3660 12869
rect 17500 12903 17552 12912
rect 17500 12869 17509 12903
rect 17509 12869 17543 12903
rect 17543 12869 17552 12903
rect 17500 12860 17552 12869
rect 2228 12724 2280 12733
rect 2964 12724 3016 12776
rect 4896 12792 4948 12844
rect 4988 12792 5040 12844
rect 4528 12724 4580 12776
rect 5724 12767 5776 12776
rect 4712 12699 4764 12708
rect 4712 12665 4721 12699
rect 4721 12665 4755 12699
rect 4755 12665 4764 12699
rect 5724 12733 5733 12767
rect 5733 12733 5767 12767
rect 5767 12733 5776 12767
rect 14556 12792 14608 12844
rect 19616 12792 19668 12844
rect 5724 12724 5776 12733
rect 17684 12767 17736 12776
rect 17684 12733 17693 12767
rect 17693 12733 17727 12767
rect 17727 12733 17736 12767
rect 17684 12724 17736 12733
rect 17960 12767 18012 12776
rect 17960 12733 17969 12767
rect 17969 12733 18003 12767
rect 18003 12733 18012 12767
rect 17960 12724 18012 12733
rect 4712 12656 4764 12665
rect 10968 12656 11020 12708
rect 4804 12631 4856 12640
rect 4804 12597 4813 12631
rect 4813 12597 4847 12631
rect 4847 12597 4856 12631
rect 4804 12588 4856 12597
rect 5080 12588 5132 12640
rect 11060 12588 11112 12640
rect 15200 12588 15252 12640
rect 18328 12588 18380 12640
rect 3174 12486 3226 12538
rect 3238 12486 3290 12538
rect 3302 12486 3354 12538
rect 3366 12486 3418 12538
rect 3430 12486 3482 12538
rect 7622 12486 7674 12538
rect 7686 12486 7738 12538
rect 7750 12486 7802 12538
rect 7814 12486 7866 12538
rect 7878 12486 7930 12538
rect 12070 12486 12122 12538
rect 12134 12486 12186 12538
rect 12198 12486 12250 12538
rect 12262 12486 12314 12538
rect 12326 12486 12378 12538
rect 16518 12486 16570 12538
rect 16582 12486 16634 12538
rect 16646 12486 16698 12538
rect 16710 12486 16762 12538
rect 16774 12486 16826 12538
rect 2780 12384 2832 12436
rect 4068 12384 4120 12436
rect 4528 12427 4580 12436
rect 4528 12393 4537 12427
rect 4537 12393 4571 12427
rect 4571 12393 4580 12427
rect 4528 12384 4580 12393
rect 4896 12427 4948 12436
rect 4896 12393 4905 12427
rect 4905 12393 4939 12427
rect 4939 12393 4948 12427
rect 4896 12384 4948 12393
rect 17592 12384 17644 12436
rect 4712 12316 4764 12368
rect 3608 12248 3660 12300
rect 15844 12248 15896 12300
rect 18144 12248 18196 12300
rect 2596 12180 2648 12232
rect 3240 12223 3292 12232
rect 3240 12189 3249 12223
rect 3249 12189 3283 12223
rect 3283 12189 3292 12223
rect 3240 12180 3292 12189
rect 3516 12180 3568 12232
rect 3976 12180 4028 12232
rect 5356 12223 5408 12232
rect 5356 12189 5390 12223
rect 5390 12189 5408 12223
rect 5356 12180 5408 12189
rect 6920 12180 6972 12232
rect 17316 12180 17368 12232
rect 17684 12223 17736 12232
rect 17684 12189 17693 12223
rect 17693 12189 17727 12223
rect 17727 12189 17736 12223
rect 17684 12180 17736 12189
rect 2504 12112 2556 12164
rect 3700 12112 3752 12164
rect 2320 12087 2372 12096
rect 2320 12053 2329 12087
rect 2329 12053 2363 12087
rect 2363 12053 2372 12087
rect 2320 12044 2372 12053
rect 2412 12044 2464 12096
rect 3976 12044 4028 12096
rect 4344 12044 4396 12096
rect 6460 12087 6512 12096
rect 6460 12053 6469 12087
rect 6469 12053 6503 12087
rect 6503 12053 6512 12087
rect 6460 12044 6512 12053
rect 8576 12155 8628 12164
rect 8576 12121 8585 12155
rect 8585 12121 8619 12155
rect 8619 12121 8628 12155
rect 8576 12112 8628 12121
rect 14924 12112 14976 12164
rect 17960 12112 18012 12164
rect 10232 12044 10284 12096
rect 13820 12044 13872 12096
rect 17408 12087 17460 12096
rect 17408 12053 17417 12087
rect 17417 12053 17451 12087
rect 17451 12053 17460 12087
rect 17408 12044 17460 12053
rect 17868 12044 17920 12096
rect 5398 11942 5450 11994
rect 5462 11942 5514 11994
rect 5526 11942 5578 11994
rect 5590 11942 5642 11994
rect 5654 11942 5706 11994
rect 9846 11942 9898 11994
rect 9910 11942 9962 11994
rect 9974 11942 10026 11994
rect 10038 11942 10090 11994
rect 10102 11942 10154 11994
rect 14294 11942 14346 11994
rect 14358 11942 14410 11994
rect 14422 11942 14474 11994
rect 14486 11942 14538 11994
rect 14550 11942 14602 11994
rect 2412 11883 2464 11892
rect 2412 11849 2421 11883
rect 2421 11849 2455 11883
rect 2455 11849 2464 11883
rect 2412 11840 2464 11849
rect 2964 11840 3016 11892
rect 3792 11840 3844 11892
rect 3976 11840 4028 11892
rect 8300 11840 8352 11892
rect 13636 11840 13688 11892
rect 17132 11840 17184 11892
rect 18052 11840 18104 11892
rect 2872 11772 2924 11824
rect 3700 11704 3752 11756
rect 3884 11772 3936 11824
rect 3976 11704 4028 11756
rect 4712 11704 4764 11756
rect 6460 11772 6512 11824
rect 7012 11772 7064 11824
rect 6368 11747 6420 11756
rect 6368 11713 6377 11747
rect 6377 11713 6411 11747
rect 6411 11713 6420 11747
rect 6368 11704 6420 11713
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 12808 11772 12860 11824
rect 14004 11772 14056 11824
rect 15844 11704 15896 11756
rect 17500 11747 17552 11756
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 17776 11704 17828 11756
rect 2228 11679 2280 11688
rect 2228 11645 2237 11679
rect 2237 11645 2271 11679
rect 2271 11645 2280 11679
rect 2228 11636 2280 11645
rect 2872 11679 2924 11688
rect 2872 11645 2881 11679
rect 2881 11645 2915 11679
rect 2915 11645 2924 11679
rect 2872 11636 2924 11645
rect 3056 11679 3108 11688
rect 3056 11645 3065 11679
rect 3065 11645 3099 11679
rect 3099 11645 3108 11679
rect 3056 11636 3108 11645
rect 3608 11636 3660 11688
rect 15752 11636 15804 11688
rect 17316 11636 17368 11688
rect 17960 11679 18012 11688
rect 17960 11645 17969 11679
rect 17969 11645 18003 11679
rect 18003 11645 18012 11679
rect 17960 11636 18012 11645
rect 2964 11500 3016 11552
rect 3608 11500 3660 11552
rect 4160 11500 4212 11552
rect 15108 11568 15160 11620
rect 17776 11568 17828 11620
rect 6092 11500 6144 11552
rect 7472 11500 7524 11552
rect 8116 11500 8168 11552
rect 10232 11500 10284 11552
rect 15660 11500 15712 11552
rect 17408 11543 17460 11552
rect 17408 11509 17417 11543
rect 17417 11509 17451 11543
rect 17451 11509 17460 11543
rect 17408 11500 17460 11509
rect 3174 11398 3226 11450
rect 3238 11398 3290 11450
rect 3302 11398 3354 11450
rect 3366 11398 3418 11450
rect 3430 11398 3482 11450
rect 7622 11398 7674 11450
rect 7686 11398 7738 11450
rect 7750 11398 7802 11450
rect 7814 11398 7866 11450
rect 7878 11398 7930 11450
rect 12070 11398 12122 11450
rect 12134 11398 12186 11450
rect 12198 11398 12250 11450
rect 12262 11398 12314 11450
rect 12326 11398 12378 11450
rect 16518 11398 16570 11450
rect 16582 11398 16634 11450
rect 16646 11398 16698 11450
rect 16710 11398 16762 11450
rect 16774 11398 16826 11450
rect 2504 11339 2556 11348
rect 2504 11305 2513 11339
rect 2513 11305 2547 11339
rect 2547 11305 2556 11339
rect 2504 11296 2556 11305
rect 3516 11296 3568 11348
rect 3700 11296 3752 11348
rect 4068 11296 4120 11348
rect 3976 11228 4028 11280
rect 4252 11228 4304 11280
rect 2964 11203 3016 11212
rect 2964 11169 2973 11203
rect 2973 11169 3007 11203
rect 3007 11169 3016 11203
rect 2964 11160 3016 11169
rect 3056 11203 3108 11212
rect 3056 11169 3065 11203
rect 3065 11169 3099 11203
rect 3099 11169 3108 11203
rect 3056 11160 3108 11169
rect 3424 11160 3476 11212
rect 8392 11296 8444 11348
rect 11152 11296 11204 11348
rect 12716 11296 12768 11348
rect 17592 11296 17644 11348
rect 1952 11135 2004 11144
rect 1952 11101 1961 11135
rect 1961 11101 1995 11135
rect 1995 11101 2004 11135
rect 1952 11092 2004 11101
rect 2228 11135 2280 11144
rect 2228 11101 2237 11135
rect 2237 11101 2271 11135
rect 2271 11101 2280 11135
rect 2228 11092 2280 11101
rect 4896 11135 4948 11144
rect 4896 11101 4905 11135
rect 4905 11101 4939 11135
rect 4939 11101 4948 11135
rect 4896 11092 4948 11101
rect 5816 11135 5868 11144
rect 5816 11101 5825 11135
rect 5825 11101 5859 11135
rect 5859 11101 5868 11135
rect 5816 11092 5868 11101
rect 3056 11024 3108 11076
rect 5724 11024 5776 11076
rect 6736 11228 6788 11280
rect 15752 11271 15804 11280
rect 15752 11237 15761 11271
rect 15761 11237 15795 11271
rect 15795 11237 15804 11271
rect 15752 11228 15804 11237
rect 15844 11228 15896 11280
rect 14648 11160 14700 11212
rect 6368 11092 6420 11144
rect 14188 11092 14240 11144
rect 15476 11135 15528 11144
rect 15476 11101 15485 11135
rect 15485 11101 15519 11135
rect 15519 11101 15528 11135
rect 15476 11092 15528 11101
rect 16396 11092 16448 11144
rect 17224 11092 17276 11144
rect 17408 11092 17460 11144
rect 17592 11135 17644 11144
rect 17592 11101 17601 11135
rect 17601 11101 17635 11135
rect 17635 11101 17644 11135
rect 17592 11092 17644 11101
rect 17684 11135 17736 11144
rect 17684 11101 17693 11135
rect 17693 11101 17727 11135
rect 17727 11101 17736 11135
rect 17684 11092 17736 11101
rect 6828 11024 6880 11076
rect 7472 11024 7524 11076
rect 2412 10999 2464 11008
rect 2412 10965 2421 10999
rect 2421 10965 2455 10999
rect 2455 10965 2464 10999
rect 2412 10956 2464 10965
rect 4988 10999 5040 11008
rect 4988 10965 4997 10999
rect 4997 10965 5031 10999
rect 5031 10965 5040 10999
rect 4988 10956 5040 10965
rect 5080 10956 5132 11008
rect 6276 10999 6328 11008
rect 6276 10965 6285 10999
rect 6285 10965 6319 10999
rect 6319 10965 6328 10999
rect 6276 10956 6328 10965
rect 7288 10956 7340 11008
rect 9036 10956 9088 11008
rect 10692 10956 10744 11008
rect 13452 11024 13504 11076
rect 15292 11024 15344 11076
rect 12900 10956 12952 11008
rect 15844 11024 15896 11076
rect 16672 10999 16724 11008
rect 16672 10965 16681 10999
rect 16681 10965 16715 10999
rect 16715 10965 16724 10999
rect 16672 10956 16724 10965
rect 17132 10999 17184 11008
rect 17132 10965 17141 10999
rect 17141 10965 17175 10999
rect 17175 10965 17184 10999
rect 17132 10956 17184 10965
rect 17224 10956 17276 11008
rect 5398 10854 5450 10906
rect 5462 10854 5514 10906
rect 5526 10854 5578 10906
rect 5590 10854 5642 10906
rect 5654 10854 5706 10906
rect 9846 10854 9898 10906
rect 9910 10854 9962 10906
rect 9974 10854 10026 10906
rect 10038 10854 10090 10906
rect 10102 10854 10154 10906
rect 14294 10854 14346 10906
rect 14358 10854 14410 10906
rect 14422 10854 14474 10906
rect 14486 10854 14538 10906
rect 14550 10854 14602 10906
rect 2320 10752 2372 10804
rect 3148 10752 3200 10804
rect 4160 10752 4212 10804
rect 4896 10752 4948 10804
rect 5080 10795 5132 10804
rect 5080 10761 5089 10795
rect 5089 10761 5123 10795
rect 5123 10761 5132 10795
rect 5080 10752 5132 10761
rect 1584 10659 1636 10668
rect 1584 10625 1593 10659
rect 1593 10625 1627 10659
rect 1627 10625 1636 10659
rect 1584 10616 1636 10625
rect 3516 10684 3568 10736
rect 6276 10752 6328 10804
rect 8392 10795 8444 10804
rect 8392 10761 8401 10795
rect 8401 10761 8435 10795
rect 8435 10761 8444 10795
rect 8392 10752 8444 10761
rect 12716 10795 12768 10804
rect 12716 10761 12725 10795
rect 12725 10761 12759 10795
rect 12759 10761 12768 10795
rect 12716 10752 12768 10761
rect 13544 10795 13596 10804
rect 13544 10761 13553 10795
rect 13553 10761 13587 10795
rect 13587 10761 13596 10795
rect 13544 10752 13596 10761
rect 17960 10752 18012 10804
rect 7288 10727 7340 10736
rect 4804 10616 4856 10668
rect 3884 10591 3936 10600
rect 3884 10557 3893 10591
rect 3893 10557 3927 10591
rect 3927 10557 3936 10591
rect 3884 10548 3936 10557
rect 5448 10548 5500 10600
rect 7288 10693 7322 10727
rect 7322 10693 7340 10727
rect 7288 10684 7340 10693
rect 14096 10684 14148 10736
rect 17132 10727 17184 10736
rect 5908 10659 5960 10668
rect 5908 10625 5917 10659
rect 5917 10625 5951 10659
rect 5951 10625 5960 10659
rect 5908 10616 5960 10625
rect 6368 10616 6420 10668
rect 6828 10616 6880 10668
rect 6736 10548 6788 10600
rect 8484 10616 8536 10668
rect 9036 10659 9088 10668
rect 9036 10625 9045 10659
rect 9045 10625 9079 10659
rect 9079 10625 9088 10659
rect 9036 10616 9088 10625
rect 11336 10616 11388 10668
rect 13636 10659 13688 10668
rect 13636 10625 13645 10659
rect 13645 10625 13679 10659
rect 13679 10625 13688 10659
rect 13636 10616 13688 10625
rect 15568 10659 15620 10668
rect 15568 10625 15577 10659
rect 15577 10625 15611 10659
rect 15611 10625 15620 10659
rect 15568 10616 15620 10625
rect 16856 10616 16908 10668
rect 17132 10693 17141 10727
rect 17141 10693 17175 10727
rect 17175 10693 17184 10727
rect 17132 10684 17184 10693
rect 18604 10616 18656 10668
rect 10508 10591 10560 10600
rect 10508 10557 10517 10591
rect 10517 10557 10551 10591
rect 10551 10557 10560 10591
rect 10508 10548 10560 10557
rect 10692 10591 10744 10600
rect 10692 10557 10701 10591
rect 10701 10557 10735 10591
rect 10735 10557 10744 10591
rect 10692 10548 10744 10557
rect 11704 10548 11756 10600
rect 11980 10591 12032 10600
rect 11980 10557 11989 10591
rect 11989 10557 12023 10591
rect 12023 10557 12032 10591
rect 11980 10548 12032 10557
rect 12900 10591 12952 10600
rect 1400 10455 1452 10464
rect 1400 10421 1409 10455
rect 1409 10421 1443 10455
rect 1443 10421 1452 10455
rect 1400 10412 1452 10421
rect 2688 10412 2740 10464
rect 3700 10412 3752 10464
rect 10324 10480 10376 10532
rect 12900 10557 12909 10591
rect 12909 10557 12943 10591
rect 12943 10557 12952 10591
rect 12900 10548 12952 10557
rect 13452 10548 13504 10600
rect 15752 10591 15804 10600
rect 15752 10557 15761 10591
rect 15761 10557 15795 10591
rect 15795 10557 15804 10591
rect 15752 10548 15804 10557
rect 16120 10548 16172 10600
rect 17684 10591 17736 10600
rect 17684 10557 17693 10591
rect 17693 10557 17727 10591
rect 17727 10557 17736 10591
rect 17684 10548 17736 10557
rect 17960 10591 18012 10600
rect 17960 10557 17969 10591
rect 17969 10557 18003 10591
rect 18003 10557 18012 10591
rect 17960 10548 18012 10557
rect 14096 10480 14148 10532
rect 15200 10523 15252 10532
rect 15200 10489 15209 10523
rect 15209 10489 15243 10523
rect 15243 10489 15252 10523
rect 15200 10480 15252 10489
rect 16212 10480 16264 10532
rect 4528 10412 4580 10464
rect 5816 10412 5868 10464
rect 5908 10412 5960 10464
rect 8208 10412 8260 10464
rect 9956 10412 10008 10464
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 13084 10412 13136 10464
rect 16304 10455 16356 10464
rect 16304 10421 16313 10455
rect 16313 10421 16347 10455
rect 16347 10421 16356 10455
rect 16304 10412 16356 10421
rect 17500 10412 17552 10464
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 3430 10310 3482 10362
rect 7622 10310 7674 10362
rect 7686 10310 7738 10362
rect 7750 10310 7802 10362
rect 7814 10310 7866 10362
rect 7878 10310 7930 10362
rect 12070 10310 12122 10362
rect 12134 10310 12186 10362
rect 12198 10310 12250 10362
rect 12262 10310 12314 10362
rect 12326 10310 12378 10362
rect 16518 10310 16570 10362
rect 16582 10310 16634 10362
rect 16646 10310 16698 10362
rect 16710 10310 16762 10362
rect 16774 10310 16826 10362
rect 2044 10208 2096 10260
rect 2872 10208 2924 10260
rect 4528 10208 4580 10260
rect 4988 10208 5040 10260
rect 3976 10140 4028 10192
rect 8576 10208 8628 10260
rect 10508 10251 10560 10260
rect 10508 10217 10517 10251
rect 10517 10217 10551 10251
rect 10551 10217 10560 10251
rect 10508 10208 10560 10217
rect 11336 10251 11388 10260
rect 11336 10217 11345 10251
rect 11345 10217 11379 10251
rect 11379 10217 11388 10251
rect 11336 10208 11388 10217
rect 11980 10208 12032 10260
rect 15568 10208 15620 10260
rect 2504 10072 2556 10124
rect 3516 10072 3568 10124
rect 5448 10115 5500 10124
rect 5448 10081 5457 10115
rect 5457 10081 5491 10115
rect 5491 10081 5500 10115
rect 5448 10072 5500 10081
rect 6736 10140 6788 10192
rect 1492 10047 1544 10056
rect 1492 10013 1501 10047
rect 1501 10013 1535 10047
rect 1535 10013 1544 10047
rect 1492 10004 1544 10013
rect 1860 10047 1912 10056
rect 1860 10013 1869 10047
rect 1869 10013 1903 10047
rect 1903 10013 1912 10047
rect 1860 10004 1912 10013
rect 2320 10047 2372 10056
rect 2320 10013 2329 10047
rect 2329 10013 2363 10047
rect 2363 10013 2372 10047
rect 2320 10004 2372 10013
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 3700 10004 3752 10056
rect 2228 9936 2280 9988
rect 2044 9868 2096 9920
rect 3792 9936 3844 9988
rect 4528 9936 4580 9988
rect 5816 10004 5868 10056
rect 6000 10047 6052 10056
rect 6000 10013 6009 10047
rect 6009 10013 6043 10047
rect 6043 10013 6052 10047
rect 6000 10004 6052 10013
rect 6276 10072 6328 10124
rect 8484 10140 8536 10192
rect 10692 10140 10744 10192
rect 13544 10140 13596 10192
rect 16948 10140 17000 10192
rect 9036 10072 9088 10124
rect 10416 10072 10468 10124
rect 10968 10115 11020 10124
rect 10968 10081 10977 10115
rect 10977 10081 11011 10115
rect 11011 10081 11020 10115
rect 10968 10072 11020 10081
rect 12900 10072 12952 10124
rect 13636 10072 13688 10124
rect 17500 10115 17552 10124
rect 17500 10081 17509 10115
rect 17509 10081 17543 10115
rect 17543 10081 17552 10115
rect 17500 10072 17552 10081
rect 6736 10004 6788 10056
rect 6828 10004 6880 10056
rect 8116 10004 8168 10056
rect 9956 10047 10008 10056
rect 9956 10013 9965 10047
rect 9965 10013 9999 10047
rect 9999 10013 10008 10047
rect 9956 10004 10008 10013
rect 11520 10004 11572 10056
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 12808 10004 12860 10056
rect 3700 9868 3752 9920
rect 9680 9936 9732 9988
rect 10232 9936 10284 9988
rect 11612 9936 11664 9988
rect 14188 10004 14240 10056
rect 16120 10004 16172 10056
rect 16304 10004 16356 10056
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 6092 9911 6144 9920
rect 6092 9877 6101 9911
rect 6101 9877 6135 9911
rect 6135 9877 6144 9911
rect 6092 9868 6144 9877
rect 7196 9868 7248 9920
rect 8668 9868 8720 9920
rect 10416 9868 10468 9920
rect 18236 9979 18288 9988
rect 12624 9911 12676 9920
rect 12624 9877 12633 9911
rect 12633 9877 12667 9911
rect 12667 9877 12676 9911
rect 12624 9868 12676 9877
rect 13452 9868 13504 9920
rect 18236 9945 18245 9979
rect 18245 9945 18279 9979
rect 18279 9945 18288 9979
rect 18236 9936 18288 9945
rect 16304 9868 16356 9920
rect 16948 9911 17000 9920
rect 16948 9877 16957 9911
rect 16957 9877 16991 9911
rect 16991 9877 17000 9911
rect 16948 9868 17000 9877
rect 17408 9911 17460 9920
rect 17408 9877 17417 9911
rect 17417 9877 17451 9911
rect 17451 9877 17460 9911
rect 17408 9868 17460 9877
rect 17684 9868 17736 9920
rect 5398 9766 5450 9818
rect 5462 9766 5514 9818
rect 5526 9766 5578 9818
rect 5590 9766 5642 9818
rect 5654 9766 5706 9818
rect 9846 9766 9898 9818
rect 9910 9766 9962 9818
rect 9974 9766 10026 9818
rect 10038 9766 10090 9818
rect 10102 9766 10154 9818
rect 14294 9766 14346 9818
rect 14358 9766 14410 9818
rect 14422 9766 14474 9818
rect 14486 9766 14538 9818
rect 14550 9766 14602 9818
rect 3884 9664 3936 9716
rect 5816 9707 5868 9716
rect 5816 9673 5825 9707
rect 5825 9673 5859 9707
rect 5859 9673 5868 9707
rect 5816 9664 5868 9673
rect 6092 9664 6144 9716
rect 1308 9392 1360 9444
rect 4620 9596 4672 9648
rect 5448 9596 5500 9648
rect 6552 9596 6604 9648
rect 12716 9664 12768 9716
rect 12808 9664 12860 9716
rect 7012 9596 7064 9648
rect 8668 9639 8720 9648
rect 8668 9605 8686 9639
rect 8686 9605 8720 9639
rect 8668 9596 8720 9605
rect 9588 9596 9640 9648
rect 10232 9596 10284 9648
rect 2320 9528 2372 9580
rect 2872 9528 2924 9580
rect 3608 9571 3660 9580
rect 3608 9537 3617 9571
rect 3617 9537 3651 9571
rect 3651 9537 3660 9571
rect 3608 9528 3660 9537
rect 4528 9571 4580 9580
rect 4528 9537 4537 9571
rect 4537 9537 4571 9571
rect 4571 9537 4580 9571
rect 4528 9528 4580 9537
rect 4988 9528 5040 9580
rect 1768 9503 1820 9512
rect 1768 9469 1777 9503
rect 1777 9469 1811 9503
rect 1811 9469 1820 9503
rect 1768 9460 1820 9469
rect 2964 9460 3016 9512
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 3056 9392 3108 9444
rect 3792 9460 3844 9512
rect 5172 9528 5224 9580
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 5356 9460 5408 9512
rect 2964 9324 3016 9376
rect 3516 9324 3568 9376
rect 4804 9324 4856 9376
rect 5816 9460 5868 9512
rect 6736 9460 6788 9512
rect 6000 9392 6052 9444
rect 6276 9392 6328 9444
rect 6460 9324 6512 9376
rect 6736 9324 6788 9376
rect 11980 9528 12032 9580
rect 12716 9528 12768 9580
rect 13636 9528 13688 9580
rect 14188 9571 14240 9580
rect 14188 9537 14197 9571
rect 14197 9537 14231 9571
rect 14231 9537 14240 9571
rect 14188 9528 14240 9537
rect 15752 9664 15804 9716
rect 16304 9707 16356 9716
rect 16304 9673 16313 9707
rect 16313 9673 16347 9707
rect 16347 9673 16356 9707
rect 16304 9664 16356 9673
rect 16856 9664 16908 9716
rect 8944 9503 8996 9512
rect 8944 9469 8953 9503
rect 8953 9469 8987 9503
rect 8987 9469 8996 9503
rect 8944 9460 8996 9469
rect 10968 9460 11020 9512
rect 12992 9503 13044 9512
rect 9680 9392 9732 9444
rect 11152 9392 11204 9444
rect 12716 9392 12768 9444
rect 12992 9469 13001 9503
rect 13001 9469 13035 9503
rect 13035 9469 13044 9503
rect 12992 9460 13044 9469
rect 13268 9503 13320 9512
rect 13268 9469 13277 9503
rect 13277 9469 13311 9503
rect 13311 9469 13320 9503
rect 13268 9460 13320 9469
rect 16856 9528 16908 9580
rect 17040 9571 17092 9580
rect 17040 9537 17049 9571
rect 17049 9537 17083 9571
rect 17083 9537 17092 9571
rect 17040 9528 17092 9537
rect 16948 9460 17000 9512
rect 17132 9503 17184 9512
rect 17132 9469 17141 9503
rect 17141 9469 17175 9503
rect 17175 9469 17184 9503
rect 17132 9460 17184 9469
rect 12900 9392 12952 9444
rect 13452 9392 13504 9444
rect 13636 9392 13688 9444
rect 17776 9460 17828 9512
rect 8668 9324 8720 9376
rect 8760 9324 8812 9376
rect 10232 9324 10284 9376
rect 10784 9324 10836 9376
rect 12440 9324 12492 9376
rect 12808 9324 12860 9376
rect 13912 9367 13964 9376
rect 13912 9333 13921 9367
rect 13921 9333 13955 9367
rect 13955 9333 13964 9367
rect 13912 9324 13964 9333
rect 15568 9324 15620 9376
rect 15936 9324 15988 9376
rect 18328 9392 18380 9444
rect 17592 9367 17644 9376
rect 17592 9333 17601 9367
rect 17601 9333 17635 9367
rect 17635 9333 17644 9367
rect 17592 9324 17644 9333
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 3430 9222 3482 9274
rect 7622 9222 7674 9274
rect 7686 9222 7738 9274
rect 7750 9222 7802 9274
rect 7814 9222 7866 9274
rect 7878 9222 7930 9274
rect 12070 9222 12122 9274
rect 12134 9222 12186 9274
rect 12198 9222 12250 9274
rect 12262 9222 12314 9274
rect 12326 9222 12378 9274
rect 16518 9222 16570 9274
rect 16582 9222 16634 9274
rect 16646 9222 16698 9274
rect 16710 9222 16762 9274
rect 16774 9222 16826 9274
rect 1860 9120 1912 9172
rect 2688 9120 2740 9172
rect 3608 9120 3660 9172
rect 4528 9120 4580 9172
rect 5356 9120 5408 9172
rect 8484 9120 8536 9172
rect 8576 9120 8628 9172
rect 9496 9120 9548 9172
rect 12532 9120 12584 9172
rect 12624 9120 12676 9172
rect 13728 9120 13780 9172
rect 15292 9120 15344 9172
rect 6000 9052 6052 9104
rect 1584 8916 1636 8968
rect 1768 8916 1820 8968
rect 3056 8959 3108 8968
rect 3056 8925 3065 8959
rect 3065 8925 3099 8959
rect 3099 8925 3108 8959
rect 3056 8916 3108 8925
rect 5448 8984 5500 9036
rect 8576 9027 8628 9036
rect 8024 8916 8076 8968
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 2688 8891 2740 8900
rect 2688 8857 2706 8891
rect 2706 8857 2740 8891
rect 3424 8891 3476 8900
rect 2688 8848 2740 8857
rect 3424 8857 3433 8891
rect 3433 8857 3467 8891
rect 3467 8857 3476 8891
rect 3424 8848 3476 8857
rect 3884 8780 3936 8832
rect 4528 8780 4580 8832
rect 4896 8891 4948 8900
rect 4896 8857 4914 8891
rect 4914 8857 4948 8891
rect 4896 8848 4948 8857
rect 7104 8848 7156 8900
rect 7564 8848 7616 8900
rect 6000 8780 6052 8832
rect 7472 8780 7524 8832
rect 8576 8993 8585 9027
rect 8585 8993 8619 9027
rect 8619 8993 8628 9027
rect 8576 8984 8628 8993
rect 11520 9052 11572 9104
rect 12808 9052 12860 9104
rect 13912 9052 13964 9104
rect 16120 9120 16172 9172
rect 16856 9120 16908 9172
rect 17040 9120 17092 9172
rect 17408 9120 17460 9172
rect 17500 9120 17552 9172
rect 9588 8984 9640 9036
rect 8760 8916 8812 8968
rect 13268 8984 13320 9036
rect 13452 9027 13504 9036
rect 13452 8993 13461 9027
rect 13461 8993 13495 9027
rect 13495 8993 13504 9027
rect 13452 8984 13504 8993
rect 13544 8984 13596 9036
rect 13820 9027 13872 9036
rect 13820 8993 13829 9027
rect 13829 8993 13863 9027
rect 13863 8993 13872 9027
rect 13820 8984 13872 8993
rect 16120 8984 16172 9036
rect 16488 8984 16540 9036
rect 8760 8780 8812 8832
rect 9496 8848 9548 8900
rect 9312 8780 9364 8832
rect 14188 8916 14240 8968
rect 12716 8848 12768 8900
rect 12992 8848 13044 8900
rect 14832 8891 14884 8900
rect 14832 8857 14866 8891
rect 14866 8857 14884 8891
rect 14832 8848 14884 8857
rect 17592 8984 17644 9036
rect 17684 8959 17736 8968
rect 17684 8925 17693 8959
rect 17693 8925 17727 8959
rect 17727 8925 17736 8959
rect 17684 8916 17736 8925
rect 18788 8984 18840 9036
rect 17500 8848 17552 8900
rect 10232 8780 10284 8832
rect 10416 8823 10468 8832
rect 10416 8789 10425 8823
rect 10425 8789 10459 8823
rect 10459 8789 10468 8823
rect 10416 8780 10468 8789
rect 11152 8780 11204 8832
rect 13176 8780 13228 8832
rect 13544 8780 13596 8832
rect 13820 8780 13872 8832
rect 15752 8780 15804 8832
rect 16120 8780 16172 8832
rect 16672 8780 16724 8832
rect 16948 8780 17000 8832
rect 18420 8823 18472 8832
rect 18420 8789 18429 8823
rect 18429 8789 18463 8823
rect 18463 8789 18472 8823
rect 18420 8780 18472 8789
rect 5398 8678 5450 8730
rect 5462 8678 5514 8730
rect 5526 8678 5578 8730
rect 5590 8678 5642 8730
rect 5654 8678 5706 8730
rect 9846 8678 9898 8730
rect 9910 8678 9962 8730
rect 9974 8678 10026 8730
rect 10038 8678 10090 8730
rect 10102 8678 10154 8730
rect 14294 8678 14346 8730
rect 14358 8678 14410 8730
rect 14422 8678 14474 8730
rect 14486 8678 14538 8730
rect 14550 8678 14602 8730
rect 2596 8619 2648 8628
rect 2596 8585 2605 8619
rect 2605 8585 2639 8619
rect 2639 8585 2648 8619
rect 2596 8576 2648 8585
rect 2964 8576 3016 8628
rect 3700 8576 3752 8628
rect 4068 8576 4120 8628
rect 5264 8576 5316 8628
rect 2688 8508 2740 8560
rect 1584 8415 1636 8424
rect 1584 8381 1593 8415
rect 1593 8381 1627 8415
rect 1627 8381 1636 8415
rect 1584 8372 1636 8381
rect 2688 8415 2740 8424
rect 2688 8381 2697 8415
rect 2697 8381 2731 8415
rect 2731 8381 2740 8415
rect 2688 8372 2740 8381
rect 3884 8508 3936 8560
rect 5540 8508 5592 8560
rect 6000 8576 6052 8628
rect 6736 8619 6788 8628
rect 6736 8585 6745 8619
rect 6745 8585 6779 8619
rect 6779 8585 6788 8619
rect 6736 8576 6788 8585
rect 5908 8508 5960 8560
rect 6828 8508 6880 8560
rect 7012 8576 7064 8628
rect 7564 8576 7616 8628
rect 7656 8508 7708 8560
rect 8116 8576 8168 8628
rect 10784 8576 10836 8628
rect 8300 8551 8352 8560
rect 8300 8517 8309 8551
rect 8309 8517 8343 8551
rect 8343 8517 8352 8551
rect 8300 8508 8352 8517
rect 8484 8508 8536 8560
rect 4344 8483 4396 8492
rect 4344 8449 4353 8483
rect 4353 8449 4387 8483
rect 4387 8449 4396 8483
rect 4344 8440 4396 8449
rect 5172 8440 5224 8492
rect 8024 8440 8076 8492
rect 8116 8440 8168 8492
rect 14648 8576 14700 8628
rect 14832 8576 14884 8628
rect 13728 8551 13780 8560
rect 13728 8517 13737 8551
rect 13737 8517 13771 8551
rect 13771 8517 13780 8551
rect 13728 8508 13780 8517
rect 13820 8551 13872 8560
rect 13820 8517 13829 8551
rect 13829 8517 13863 8551
rect 13863 8517 13872 8551
rect 13820 8508 13872 8517
rect 14188 8508 14240 8560
rect 16948 8576 17000 8628
rect 17132 8576 17184 8628
rect 17500 8619 17552 8628
rect 17500 8585 17509 8619
rect 17509 8585 17543 8619
rect 17543 8585 17552 8619
rect 17500 8576 17552 8585
rect 17868 8576 17920 8628
rect 9772 8440 9824 8492
rect 11980 8483 12032 8492
rect 11980 8449 11989 8483
rect 11989 8449 12023 8483
rect 12023 8449 12032 8483
rect 11980 8440 12032 8449
rect 13636 8440 13688 8492
rect 14832 8440 14884 8492
rect 15844 8483 15896 8492
rect 17316 8508 17368 8560
rect 15844 8449 15862 8483
rect 15862 8449 15896 8483
rect 15844 8440 15896 8449
rect 16304 8483 16356 8492
rect 16304 8449 16313 8483
rect 16313 8449 16347 8483
rect 16347 8449 16356 8483
rect 16304 8440 16356 8449
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 17960 8440 18012 8492
rect 3056 8372 3108 8424
rect 3884 8372 3936 8424
rect 4436 8415 4488 8424
rect 4436 8381 4445 8415
rect 4445 8381 4479 8415
rect 4479 8381 4488 8415
rect 4436 8372 4488 8381
rect 4528 8415 4580 8424
rect 4528 8381 4537 8415
rect 4537 8381 4571 8415
rect 4571 8381 4580 8415
rect 4528 8372 4580 8381
rect 6460 8415 6512 8424
rect 5080 8304 5132 8356
rect 2964 8236 3016 8288
rect 4068 8236 4120 8288
rect 4160 8236 4212 8288
rect 5264 8304 5316 8356
rect 6460 8381 6469 8415
rect 6469 8381 6503 8415
rect 6503 8381 6512 8415
rect 6460 8372 6512 8381
rect 7104 8372 7156 8424
rect 8392 8415 8444 8424
rect 6828 8304 6880 8356
rect 7196 8304 7248 8356
rect 8392 8381 8401 8415
rect 8401 8381 8435 8415
rect 8435 8381 8444 8415
rect 8392 8372 8444 8381
rect 8484 8415 8536 8424
rect 8484 8381 8493 8415
rect 8493 8381 8527 8415
rect 8527 8381 8536 8415
rect 8484 8372 8536 8381
rect 13176 8415 13228 8424
rect 13176 8381 13185 8415
rect 13185 8381 13219 8415
rect 13219 8381 13228 8415
rect 13176 8372 13228 8381
rect 13452 8372 13504 8424
rect 10416 8304 10468 8356
rect 11520 8347 11572 8356
rect 11520 8313 11529 8347
rect 11529 8313 11563 8347
rect 11563 8313 11572 8347
rect 11520 8304 11572 8313
rect 12532 8347 12584 8356
rect 12532 8313 12541 8347
rect 12541 8313 12575 8347
rect 12575 8313 12584 8347
rect 12532 8304 12584 8313
rect 12716 8304 12768 8356
rect 14280 8372 14332 8424
rect 16488 8372 16540 8424
rect 16948 8415 17000 8424
rect 16948 8381 16957 8415
rect 16957 8381 16991 8415
rect 16991 8381 17000 8415
rect 16948 8372 17000 8381
rect 14556 8304 14608 8356
rect 16396 8304 16448 8356
rect 18328 8347 18380 8356
rect 18328 8313 18337 8347
rect 18337 8313 18371 8347
rect 18371 8313 18380 8347
rect 18328 8304 18380 8313
rect 6092 8236 6144 8288
rect 6460 8236 6512 8288
rect 8116 8236 8168 8288
rect 8208 8236 8260 8288
rect 10232 8236 10284 8288
rect 11336 8279 11388 8288
rect 11336 8245 11345 8279
rect 11345 8245 11379 8279
rect 11379 8245 11388 8279
rect 11336 8236 11388 8245
rect 12440 8279 12492 8288
rect 12440 8245 12449 8279
rect 12449 8245 12483 8279
rect 12483 8245 12492 8279
rect 12440 8236 12492 8245
rect 13912 8236 13964 8288
rect 15936 8236 15988 8288
rect 18052 8236 18104 8288
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 3430 8134 3482 8186
rect 7622 8134 7674 8186
rect 7686 8134 7738 8186
rect 7750 8134 7802 8186
rect 7814 8134 7866 8186
rect 7878 8134 7930 8186
rect 12070 8134 12122 8186
rect 12134 8134 12186 8186
rect 12198 8134 12250 8186
rect 12262 8134 12314 8186
rect 12326 8134 12378 8186
rect 16518 8134 16570 8186
rect 16582 8134 16634 8186
rect 16646 8134 16698 8186
rect 16710 8134 16762 8186
rect 16774 8134 16826 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 2320 8075 2372 8084
rect 2320 8041 2329 8075
rect 2329 8041 2363 8075
rect 2363 8041 2372 8075
rect 2320 8032 2372 8041
rect 2688 8075 2740 8084
rect 2688 8041 2697 8075
rect 2697 8041 2731 8075
rect 2731 8041 2740 8075
rect 2688 8032 2740 8041
rect 2504 7964 2556 8016
rect 5908 8032 5960 8084
rect 6000 8032 6052 8084
rect 8760 8032 8812 8084
rect 8944 8032 8996 8084
rect 13820 8032 13872 8084
rect 14188 8032 14240 8084
rect 15844 8075 15896 8084
rect 15844 8041 15853 8075
rect 15853 8041 15887 8075
rect 15887 8041 15896 8075
rect 15844 8032 15896 8041
rect 3976 7964 4028 8016
rect 8392 7964 8444 8016
rect 3332 7939 3384 7948
rect 3332 7905 3341 7939
rect 3341 7905 3375 7939
rect 3375 7905 3384 7939
rect 3332 7896 3384 7905
rect 5264 7896 5316 7948
rect 7288 7939 7340 7948
rect 7288 7905 7297 7939
rect 7297 7905 7331 7939
rect 7331 7905 7340 7939
rect 7288 7896 7340 7905
rect 7472 7939 7524 7948
rect 7472 7905 7481 7939
rect 7481 7905 7515 7939
rect 7515 7905 7524 7939
rect 7472 7896 7524 7905
rect 9772 7964 9824 8016
rect 9588 7939 9640 7948
rect 9588 7905 9597 7939
rect 9597 7905 9631 7939
rect 9631 7905 9640 7939
rect 9588 7896 9640 7905
rect 10048 7964 10100 8016
rect 10232 8007 10284 8016
rect 10232 7973 10241 8007
rect 10241 7973 10275 8007
rect 10275 7973 10284 8007
rect 10232 7964 10284 7973
rect 12256 7964 12308 8016
rect 13636 7964 13688 8016
rect 1584 7828 1636 7880
rect 2688 7828 2740 7880
rect 2780 7828 2832 7880
rect 3148 7871 3200 7880
rect 3148 7837 3157 7871
rect 3157 7837 3191 7871
rect 3191 7837 3200 7871
rect 3148 7828 3200 7837
rect 2320 7760 2372 7812
rect 5816 7828 5868 7880
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 8024 7828 8076 7880
rect 8208 7828 8260 7880
rect 1768 7692 1820 7744
rect 5540 7760 5592 7812
rect 6276 7760 6328 7812
rect 5080 7692 5132 7744
rect 5724 7735 5776 7744
rect 5724 7701 5733 7735
rect 5733 7701 5767 7735
rect 5767 7701 5776 7735
rect 5724 7692 5776 7701
rect 8760 7828 8812 7880
rect 9680 7828 9732 7880
rect 10416 7871 10468 7880
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 11152 7828 11204 7880
rect 13636 7828 13688 7880
rect 11336 7760 11388 7812
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 14280 7760 14332 7812
rect 16948 8032 17000 8084
rect 17040 8032 17092 8084
rect 15660 7896 15712 7948
rect 17500 7964 17552 8016
rect 14924 7871 14976 7880
rect 14924 7837 14933 7871
rect 14933 7837 14967 7871
rect 14967 7837 14976 7871
rect 14924 7828 14976 7837
rect 15108 7828 15160 7880
rect 15936 7871 15988 7880
rect 15936 7837 15945 7871
rect 15945 7837 15979 7871
rect 15979 7837 15988 7871
rect 15936 7828 15988 7837
rect 16948 7896 17000 7948
rect 17316 7939 17368 7948
rect 17316 7905 17325 7939
rect 17325 7905 17359 7939
rect 17359 7905 17368 7939
rect 17316 7896 17368 7905
rect 16212 7828 16264 7880
rect 13912 7735 13964 7744
rect 13912 7701 13921 7735
rect 13921 7701 13955 7735
rect 13955 7701 13964 7735
rect 13912 7692 13964 7701
rect 14188 7692 14240 7744
rect 15844 7760 15896 7812
rect 17132 7828 17184 7880
rect 17960 7871 18012 7880
rect 17960 7837 17969 7871
rect 17969 7837 18003 7871
rect 18003 7837 18012 7871
rect 17960 7828 18012 7837
rect 18236 7828 18288 7880
rect 15200 7692 15252 7744
rect 16396 7692 16448 7744
rect 16856 7692 16908 7744
rect 17224 7735 17276 7744
rect 17224 7701 17233 7735
rect 17233 7701 17267 7735
rect 17267 7701 17276 7735
rect 18052 7735 18104 7744
rect 17224 7692 17276 7701
rect 18052 7701 18061 7735
rect 18061 7701 18095 7735
rect 18095 7701 18104 7735
rect 18052 7692 18104 7701
rect 18696 7692 18748 7744
rect 5398 7590 5450 7642
rect 5462 7590 5514 7642
rect 5526 7590 5578 7642
rect 5590 7590 5642 7642
rect 5654 7590 5706 7642
rect 9846 7590 9898 7642
rect 9910 7590 9962 7642
rect 9974 7590 10026 7642
rect 10038 7590 10090 7642
rect 10102 7590 10154 7642
rect 14294 7590 14346 7642
rect 14358 7590 14410 7642
rect 14422 7590 14474 7642
rect 14486 7590 14538 7642
rect 14550 7590 14602 7642
rect 1676 7488 1728 7540
rect 1860 7531 1912 7540
rect 1860 7497 1869 7531
rect 1869 7497 1903 7531
rect 1903 7497 1912 7531
rect 1860 7488 1912 7497
rect 2596 7488 2648 7540
rect 3056 7531 3108 7540
rect 3056 7497 3065 7531
rect 3065 7497 3099 7531
rect 3099 7497 3108 7531
rect 3056 7488 3108 7497
rect 4160 7488 4212 7540
rect 4436 7488 4488 7540
rect 5080 7531 5132 7540
rect 5080 7497 5089 7531
rect 5089 7497 5123 7531
rect 5123 7497 5132 7531
rect 5080 7488 5132 7497
rect 5908 7531 5960 7540
rect 3884 7420 3936 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 2044 7395 2096 7404
rect 2044 7361 2053 7395
rect 2053 7361 2087 7395
rect 2087 7361 2096 7395
rect 2044 7352 2096 7361
rect 2228 7259 2280 7268
rect 2228 7225 2237 7259
rect 2237 7225 2271 7259
rect 2271 7225 2280 7259
rect 2228 7216 2280 7225
rect 2596 7395 2648 7404
rect 2596 7361 2605 7395
rect 2605 7361 2639 7395
rect 2639 7361 2648 7395
rect 3148 7395 3200 7404
rect 2596 7352 2648 7361
rect 3148 7361 3157 7395
rect 3157 7361 3191 7395
rect 3191 7361 3200 7395
rect 3148 7352 3200 7361
rect 4068 7352 4120 7404
rect 5908 7497 5917 7531
rect 5917 7497 5951 7531
rect 5951 7497 5960 7531
rect 5908 7488 5960 7497
rect 7288 7488 7340 7540
rect 7012 7420 7064 7472
rect 8484 7420 8536 7472
rect 5908 7352 5960 7404
rect 3332 7327 3384 7336
rect 3332 7293 3341 7327
rect 3341 7293 3375 7327
rect 3375 7293 3384 7327
rect 3332 7284 3384 7293
rect 4896 7284 4948 7336
rect 8116 7395 8168 7404
rect 8116 7361 8125 7395
rect 8125 7361 8159 7395
rect 8159 7361 8168 7395
rect 8116 7352 8168 7361
rect 9772 7488 9824 7540
rect 11060 7531 11112 7540
rect 11060 7497 11069 7531
rect 11069 7497 11103 7531
rect 11103 7497 11112 7531
rect 11060 7488 11112 7497
rect 11796 7488 11848 7540
rect 10508 7420 10560 7472
rect 12440 7420 12492 7472
rect 9680 7352 9732 7404
rect 12532 7352 12584 7404
rect 4344 7216 4396 7268
rect 5264 7216 5316 7268
rect 11152 7284 11204 7336
rect 11980 7284 12032 7336
rect 13544 7352 13596 7404
rect 13820 7395 13872 7404
rect 13820 7361 13829 7395
rect 13829 7361 13863 7395
rect 13863 7361 13872 7395
rect 13820 7352 13872 7361
rect 14188 7488 14240 7540
rect 14924 7488 14976 7540
rect 16764 7488 16816 7540
rect 17960 7531 18012 7540
rect 17960 7497 17969 7531
rect 17969 7497 18003 7531
rect 18003 7497 18012 7531
rect 17960 7488 18012 7497
rect 18420 7531 18472 7540
rect 18420 7497 18429 7531
rect 18429 7497 18463 7531
rect 18463 7497 18472 7531
rect 18420 7488 18472 7497
rect 17868 7420 17920 7472
rect 15292 7395 15344 7404
rect 13452 7327 13504 7336
rect 11704 7216 11756 7268
rect 13452 7293 13461 7327
rect 13461 7293 13495 7327
rect 13495 7293 13504 7327
rect 13452 7284 13504 7293
rect 13636 7284 13688 7336
rect 15292 7361 15301 7395
rect 15301 7361 15335 7395
rect 15335 7361 15344 7395
rect 15292 7352 15344 7361
rect 15476 7352 15528 7404
rect 15660 7352 15712 7404
rect 16120 7395 16172 7404
rect 6828 7148 6880 7200
rect 12256 7216 12308 7268
rect 15752 7284 15804 7336
rect 16120 7361 16129 7395
rect 16129 7361 16163 7395
rect 16163 7361 16172 7395
rect 16120 7352 16172 7361
rect 16856 7352 16908 7404
rect 17408 7395 17460 7404
rect 17408 7361 17417 7395
rect 17417 7361 17451 7395
rect 17451 7361 17460 7395
rect 17408 7352 17460 7361
rect 18144 7395 18196 7404
rect 18144 7361 18153 7395
rect 18153 7361 18187 7395
rect 18187 7361 18196 7395
rect 18144 7352 18196 7361
rect 18236 7395 18288 7404
rect 18236 7361 18245 7395
rect 18245 7361 18279 7395
rect 18279 7361 18288 7395
rect 18236 7352 18288 7361
rect 16764 7284 16816 7336
rect 15936 7216 15988 7268
rect 12716 7191 12768 7200
rect 12716 7157 12725 7191
rect 12725 7157 12759 7191
rect 12759 7157 12768 7191
rect 12716 7148 12768 7157
rect 13728 7191 13780 7200
rect 13728 7157 13737 7191
rect 13737 7157 13771 7191
rect 13771 7157 13780 7191
rect 13728 7148 13780 7157
rect 15108 7148 15160 7200
rect 15568 7148 15620 7200
rect 15752 7191 15804 7200
rect 15752 7157 15761 7191
rect 15761 7157 15795 7191
rect 15795 7157 15804 7191
rect 15752 7148 15804 7157
rect 18052 7284 18104 7336
rect 17776 7216 17828 7268
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 3430 7046 3482 7098
rect 7622 7046 7674 7098
rect 7686 7046 7738 7098
rect 7750 7046 7802 7098
rect 7814 7046 7866 7098
rect 7878 7046 7930 7098
rect 12070 7046 12122 7098
rect 12134 7046 12186 7098
rect 12198 7046 12250 7098
rect 12262 7046 12314 7098
rect 12326 7046 12378 7098
rect 16518 7046 16570 7098
rect 16582 7046 16634 7098
rect 16646 7046 16698 7098
rect 16710 7046 16762 7098
rect 16774 7046 16826 7098
rect 1492 6987 1544 6996
rect 1492 6953 1501 6987
rect 1501 6953 1535 6987
rect 1535 6953 1544 6987
rect 1492 6944 1544 6953
rect 2596 6987 2648 6996
rect 2596 6953 2605 6987
rect 2605 6953 2639 6987
rect 2639 6953 2648 6987
rect 2596 6944 2648 6953
rect 5264 6944 5316 6996
rect 8300 6944 8352 6996
rect 8392 6944 8444 6996
rect 10508 6944 10560 6996
rect 11980 6987 12032 6996
rect 11980 6953 11989 6987
rect 11989 6953 12023 6987
rect 12023 6953 12032 6987
rect 11980 6944 12032 6953
rect 12440 6944 12492 6996
rect 2320 6919 2372 6928
rect 2320 6885 2329 6919
rect 2329 6885 2363 6919
rect 2363 6885 2372 6919
rect 2320 6876 2372 6885
rect 5908 6876 5960 6928
rect 6736 6876 6788 6928
rect 1768 6740 1820 6792
rect 2136 6783 2188 6792
rect 2136 6749 2145 6783
rect 2145 6749 2179 6783
rect 2179 6749 2188 6783
rect 2136 6740 2188 6749
rect 2596 6740 2648 6792
rect 3240 6672 3292 6724
rect 1860 6647 1912 6656
rect 1860 6613 1869 6647
rect 1869 6613 1903 6647
rect 1903 6613 1912 6647
rect 1860 6604 1912 6613
rect 3516 6604 3568 6656
rect 6920 6808 6972 6860
rect 7288 6876 7340 6928
rect 8944 6919 8996 6928
rect 7196 6808 7248 6860
rect 7656 6808 7708 6860
rect 8944 6885 8953 6919
rect 8953 6885 8987 6919
rect 8987 6885 8996 6919
rect 8944 6876 8996 6885
rect 11796 6876 11848 6928
rect 8484 6808 8536 6860
rect 11980 6808 12032 6860
rect 3884 6740 3936 6792
rect 4344 6740 4396 6792
rect 5724 6740 5776 6792
rect 7380 6740 7432 6792
rect 4160 6672 4212 6724
rect 6920 6672 6972 6724
rect 8944 6672 8996 6724
rect 9404 6715 9456 6724
rect 7932 6604 7984 6656
rect 8024 6604 8076 6656
rect 8760 6647 8812 6656
rect 8760 6613 8769 6647
rect 8769 6613 8803 6647
rect 8803 6613 8812 6647
rect 9404 6681 9413 6715
rect 9413 6681 9447 6715
rect 9447 6681 9456 6715
rect 9404 6672 9456 6681
rect 9312 6647 9364 6656
rect 8760 6604 8812 6613
rect 9312 6613 9321 6647
rect 9321 6613 9355 6647
rect 9355 6613 9364 6647
rect 9312 6604 9364 6613
rect 9680 6740 9732 6792
rect 11152 6740 11204 6792
rect 12440 6808 12492 6860
rect 13268 6808 13320 6860
rect 15476 6944 15528 6996
rect 13820 6876 13872 6928
rect 14740 6876 14792 6928
rect 16488 6876 16540 6928
rect 13636 6808 13688 6860
rect 13912 6808 13964 6860
rect 12900 6740 12952 6792
rect 14832 6783 14884 6792
rect 14832 6749 14841 6783
rect 14841 6749 14875 6783
rect 14875 6749 14884 6783
rect 14832 6740 14884 6749
rect 16672 6808 16724 6860
rect 16856 6851 16908 6860
rect 16856 6817 16865 6851
rect 16865 6817 16899 6851
rect 16899 6817 16908 6851
rect 16856 6808 16908 6817
rect 13268 6715 13320 6724
rect 11428 6604 11480 6656
rect 12440 6647 12492 6656
rect 12440 6613 12449 6647
rect 12449 6613 12483 6647
rect 12483 6613 12492 6647
rect 12440 6604 12492 6613
rect 12624 6604 12676 6656
rect 13268 6681 13277 6715
rect 13277 6681 13311 6715
rect 13311 6681 13320 6715
rect 13268 6672 13320 6681
rect 13820 6672 13872 6724
rect 15660 6672 15712 6724
rect 13452 6604 13504 6656
rect 14740 6647 14792 6656
rect 14740 6613 14749 6647
rect 14749 6613 14783 6647
rect 14783 6613 14792 6647
rect 14740 6604 14792 6613
rect 16120 6604 16172 6656
rect 16856 6672 16908 6724
rect 17224 6944 17276 6996
rect 18420 6987 18472 6996
rect 18420 6953 18429 6987
rect 18429 6953 18463 6987
rect 18463 6953 18472 6987
rect 18420 6944 18472 6953
rect 17408 6876 17460 6928
rect 17224 6808 17276 6860
rect 16304 6647 16356 6656
rect 16304 6613 16313 6647
rect 16313 6613 16347 6647
rect 16347 6613 16356 6647
rect 16672 6647 16724 6656
rect 16304 6604 16356 6613
rect 16672 6613 16681 6647
rect 16681 6613 16715 6647
rect 16715 6613 16724 6647
rect 16672 6604 16724 6613
rect 17408 6604 17460 6656
rect 17684 6604 17736 6656
rect 17960 6647 18012 6656
rect 17960 6613 17969 6647
rect 17969 6613 18003 6647
rect 18003 6613 18012 6647
rect 17960 6604 18012 6613
rect 5398 6502 5450 6554
rect 5462 6502 5514 6554
rect 5526 6502 5578 6554
rect 5590 6502 5642 6554
rect 5654 6502 5706 6554
rect 9846 6502 9898 6554
rect 9910 6502 9962 6554
rect 9974 6502 10026 6554
rect 10038 6502 10090 6554
rect 10102 6502 10154 6554
rect 14294 6502 14346 6554
rect 14358 6502 14410 6554
rect 14422 6502 14474 6554
rect 14486 6502 14538 6554
rect 14550 6502 14602 6554
rect 2136 6400 2188 6452
rect 2688 6400 2740 6452
rect 3240 6400 3292 6452
rect 7012 6400 7064 6452
rect 3884 6332 3936 6384
rect 1676 6307 1728 6316
rect 1676 6273 1685 6307
rect 1685 6273 1719 6307
rect 1719 6273 1728 6307
rect 1676 6264 1728 6273
rect 1860 6307 1912 6316
rect 1860 6273 1869 6307
rect 1869 6273 1903 6307
rect 1903 6273 1912 6307
rect 1860 6264 1912 6273
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 2504 6264 2556 6316
rect 5540 6332 5592 6384
rect 6920 6332 6972 6384
rect 7472 6400 7524 6452
rect 7656 6443 7708 6452
rect 7656 6409 7665 6443
rect 7665 6409 7699 6443
rect 7699 6409 7708 6443
rect 7656 6400 7708 6409
rect 8024 6443 8076 6452
rect 8024 6409 8033 6443
rect 8033 6409 8067 6443
rect 8067 6409 8076 6443
rect 8024 6400 8076 6409
rect 9312 6400 9364 6452
rect 4160 6264 4212 6316
rect 4528 6307 4580 6316
rect 4528 6273 4537 6307
rect 4537 6273 4571 6307
rect 4571 6273 4580 6307
rect 4528 6264 4580 6273
rect 5816 6307 5868 6316
rect 5816 6273 5834 6307
rect 5834 6273 5868 6307
rect 5816 6264 5868 6273
rect 6092 6239 6144 6248
rect 1492 6103 1544 6112
rect 1492 6069 1501 6103
rect 1501 6069 1535 6103
rect 1535 6069 1544 6103
rect 1492 6060 1544 6069
rect 2136 6103 2188 6112
rect 2136 6069 2145 6103
rect 2145 6069 2179 6103
rect 2179 6069 2188 6103
rect 2136 6060 2188 6069
rect 2596 6103 2648 6112
rect 2596 6069 2605 6103
rect 2605 6069 2639 6103
rect 2639 6069 2648 6103
rect 2596 6060 2648 6069
rect 4068 6103 4120 6112
rect 4068 6069 4077 6103
rect 4077 6069 4111 6103
rect 4111 6069 4120 6103
rect 4068 6060 4120 6069
rect 6092 6205 6101 6239
rect 6101 6205 6135 6239
rect 6135 6205 6144 6239
rect 6092 6196 6144 6205
rect 8484 6332 8536 6384
rect 8944 6332 8996 6384
rect 10692 6400 10744 6452
rect 12900 6443 12952 6452
rect 12900 6409 12909 6443
rect 12909 6409 12943 6443
rect 12943 6409 12952 6443
rect 12900 6400 12952 6409
rect 13820 6400 13872 6452
rect 16304 6400 16356 6452
rect 16672 6443 16724 6452
rect 16672 6409 16681 6443
rect 16681 6409 16715 6443
rect 16715 6409 16724 6443
rect 16672 6400 16724 6409
rect 17960 6400 18012 6452
rect 18144 6400 18196 6452
rect 9772 6332 9824 6384
rect 10232 6332 10284 6384
rect 10324 6375 10376 6384
rect 10324 6341 10342 6375
rect 10342 6341 10376 6375
rect 10324 6332 10376 6341
rect 8300 6264 8352 6316
rect 10692 6307 10744 6316
rect 5724 6060 5776 6112
rect 5816 6060 5868 6112
rect 6368 6103 6420 6112
rect 6368 6069 6377 6103
rect 6377 6069 6411 6103
rect 6411 6069 6420 6103
rect 6368 6060 6420 6069
rect 6920 6060 6972 6112
rect 8944 6196 8996 6248
rect 7748 6128 7800 6180
rect 8760 6128 8812 6180
rect 10692 6273 10701 6307
rect 10701 6273 10735 6307
rect 10735 6273 10744 6307
rect 10692 6264 10744 6273
rect 11152 6196 11204 6248
rect 12072 6264 12124 6316
rect 14280 6332 14332 6384
rect 14832 6332 14884 6384
rect 16488 6332 16540 6384
rect 14740 6264 14792 6316
rect 15108 6196 15160 6248
rect 8392 6060 8444 6112
rect 10232 6060 10284 6112
rect 11428 6060 11480 6112
rect 14464 6103 14516 6112
rect 14464 6069 14473 6103
rect 14473 6069 14507 6103
rect 14507 6069 14516 6103
rect 14464 6060 14516 6069
rect 16856 6264 16908 6316
rect 17040 6264 17092 6316
rect 16120 6239 16172 6248
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16488 6239 16540 6248
rect 16120 6196 16172 6205
rect 16488 6205 16497 6239
rect 16497 6205 16531 6239
rect 16531 6205 16540 6239
rect 16488 6196 16540 6205
rect 16764 6196 16816 6248
rect 17316 6264 17368 6316
rect 17224 6239 17276 6248
rect 17224 6205 17233 6239
rect 17233 6205 17267 6239
rect 17267 6205 17276 6239
rect 18328 6264 18380 6316
rect 18604 6264 18656 6316
rect 17224 6196 17276 6205
rect 17040 6128 17092 6180
rect 17316 6128 17368 6180
rect 16212 6060 16264 6112
rect 17684 6060 17736 6112
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 3430 5958 3482 6010
rect 7622 5958 7674 6010
rect 7686 5958 7738 6010
rect 7750 5958 7802 6010
rect 7814 5958 7866 6010
rect 7878 5958 7930 6010
rect 12070 5958 12122 6010
rect 12134 5958 12186 6010
rect 12198 5958 12250 6010
rect 12262 5958 12314 6010
rect 12326 5958 12378 6010
rect 16518 5958 16570 6010
rect 16582 5958 16634 6010
rect 16646 5958 16698 6010
rect 16710 5958 16762 6010
rect 16774 5958 16826 6010
rect 3884 5856 3936 5908
rect 4068 5788 4120 5840
rect 4712 5788 4764 5840
rect 5540 5788 5592 5840
rect 6092 5788 6144 5840
rect 6828 5788 6880 5840
rect 12440 5856 12492 5908
rect 15660 5899 15712 5908
rect 15660 5865 15669 5899
rect 15669 5865 15703 5899
rect 15703 5865 15712 5899
rect 15660 5856 15712 5865
rect 16212 5899 16264 5908
rect 16212 5865 16221 5899
rect 16221 5865 16255 5899
rect 16255 5865 16264 5899
rect 16212 5856 16264 5865
rect 17040 5899 17092 5908
rect 17040 5865 17049 5899
rect 17049 5865 17083 5899
rect 17083 5865 17092 5899
rect 17040 5856 17092 5865
rect 18052 5899 18104 5908
rect 18052 5865 18061 5899
rect 18061 5865 18095 5899
rect 18095 5865 18104 5899
rect 18052 5856 18104 5865
rect 18420 5899 18472 5908
rect 18420 5865 18429 5899
rect 18429 5865 18463 5899
rect 18463 5865 18472 5899
rect 18420 5856 18472 5865
rect 2504 5720 2556 5772
rect 2596 5720 2648 5772
rect 3700 5720 3752 5772
rect 4160 5720 4212 5772
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 1768 5652 1820 5661
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 1952 5559 2004 5568
rect 1952 5525 1961 5559
rect 1961 5525 1995 5559
rect 1995 5525 2004 5559
rect 1952 5516 2004 5525
rect 2504 5516 2556 5568
rect 2872 5559 2924 5568
rect 2872 5525 2881 5559
rect 2881 5525 2915 5559
rect 2915 5525 2924 5559
rect 3240 5559 3292 5568
rect 2872 5516 2924 5525
rect 3240 5525 3249 5559
rect 3249 5525 3283 5559
rect 3283 5525 3292 5559
rect 3240 5516 3292 5525
rect 4528 5584 4580 5636
rect 5816 5720 5868 5772
rect 8944 5720 8996 5772
rect 7104 5652 7156 5704
rect 7472 5652 7524 5704
rect 6828 5584 6880 5636
rect 4620 5516 4672 5568
rect 4896 5559 4948 5568
rect 4896 5525 4905 5559
rect 4905 5525 4939 5559
rect 4939 5525 4948 5559
rect 4896 5516 4948 5525
rect 6092 5516 6144 5568
rect 6552 5516 6604 5568
rect 6736 5516 6788 5568
rect 7104 5559 7156 5568
rect 7104 5525 7113 5559
rect 7113 5525 7147 5559
rect 7147 5525 7156 5559
rect 7104 5516 7156 5525
rect 7656 5584 7708 5636
rect 13820 5788 13872 5840
rect 11152 5720 11204 5772
rect 12716 5763 12768 5772
rect 12716 5729 12725 5763
rect 12725 5729 12759 5763
rect 12759 5729 12768 5763
rect 12716 5720 12768 5729
rect 12900 5763 12952 5772
rect 12900 5729 12909 5763
rect 12909 5729 12943 5763
rect 12943 5729 12952 5763
rect 12900 5720 12952 5729
rect 13636 5763 13688 5772
rect 13636 5729 13645 5763
rect 13645 5729 13679 5763
rect 13679 5729 13688 5763
rect 13636 5720 13688 5729
rect 15936 5788 15988 5840
rect 17224 5720 17276 5772
rect 10232 5652 10284 5704
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 14280 5695 14332 5704
rect 14280 5661 14289 5695
rect 14289 5661 14323 5695
rect 14323 5661 14332 5695
rect 14280 5652 14332 5661
rect 11520 5584 11572 5636
rect 12624 5627 12676 5636
rect 12624 5593 12633 5627
rect 12633 5593 12667 5627
rect 12667 5593 12676 5627
rect 12624 5584 12676 5593
rect 13452 5627 13504 5636
rect 13452 5593 13461 5627
rect 13461 5593 13495 5627
rect 13495 5593 13504 5627
rect 13452 5584 13504 5593
rect 13728 5584 13780 5636
rect 8208 5516 8260 5568
rect 10324 5516 10376 5568
rect 11060 5516 11112 5568
rect 14004 5516 14056 5568
rect 14464 5584 14516 5636
rect 16856 5652 16908 5704
rect 17776 5720 17828 5772
rect 17316 5584 17368 5636
rect 17684 5584 17736 5636
rect 15292 5516 15344 5568
rect 15936 5559 15988 5568
rect 15936 5525 15945 5559
rect 15945 5525 15979 5559
rect 15979 5525 15988 5559
rect 15936 5516 15988 5525
rect 16580 5559 16632 5568
rect 16580 5525 16589 5559
rect 16589 5525 16623 5559
rect 16623 5525 16632 5559
rect 16580 5516 16632 5525
rect 16672 5559 16724 5568
rect 16672 5525 16681 5559
rect 16681 5525 16715 5559
rect 16715 5525 16724 5559
rect 16672 5516 16724 5525
rect 17500 5559 17552 5568
rect 17500 5525 17509 5559
rect 17509 5525 17543 5559
rect 17543 5525 17552 5559
rect 17500 5516 17552 5525
rect 5398 5414 5450 5466
rect 5462 5414 5514 5466
rect 5526 5414 5578 5466
rect 5590 5414 5642 5466
rect 5654 5414 5706 5466
rect 9846 5414 9898 5466
rect 9910 5414 9962 5466
rect 9974 5414 10026 5466
rect 10038 5414 10090 5466
rect 10102 5414 10154 5466
rect 14294 5414 14346 5466
rect 14358 5414 14410 5466
rect 14422 5414 14474 5466
rect 14486 5414 14538 5466
rect 14550 5414 14602 5466
rect 1676 5312 1728 5364
rect 2320 5312 2372 5364
rect 3240 5312 3292 5364
rect 6368 5312 6420 5364
rect 6552 5312 6604 5364
rect 8208 5312 8260 5364
rect 9588 5312 9640 5364
rect 4344 5287 4396 5296
rect 4344 5253 4353 5287
rect 4353 5253 4387 5287
rect 4387 5253 4396 5287
rect 4344 5244 4396 5253
rect 4436 5244 4488 5296
rect 1768 5176 1820 5228
rect 2044 5219 2096 5228
rect 2044 5185 2053 5219
rect 2053 5185 2087 5219
rect 2087 5185 2096 5219
rect 2044 5176 2096 5185
rect 2320 5219 2372 5228
rect 2320 5185 2329 5219
rect 2329 5185 2363 5219
rect 2363 5185 2372 5219
rect 2320 5176 2372 5185
rect 6000 5244 6052 5296
rect 6092 5244 6144 5296
rect 5724 5176 5776 5228
rect 8484 5244 8536 5296
rect 11060 5244 11112 5296
rect 11428 5312 11480 5364
rect 14096 5312 14148 5364
rect 14832 5312 14884 5364
rect 1860 5108 1912 5160
rect 2412 5108 2464 5160
rect 2596 5151 2648 5160
rect 2596 5117 2605 5151
rect 2605 5117 2639 5151
rect 2639 5117 2648 5151
rect 2596 5108 2648 5117
rect 5264 5151 5316 5160
rect 5264 5117 5273 5151
rect 5273 5117 5307 5151
rect 5307 5117 5316 5151
rect 5264 5108 5316 5117
rect 8116 5176 8168 5228
rect 8392 5176 8444 5228
rect 8944 5176 8996 5228
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 11428 5176 11480 5228
rect 11704 5176 11756 5228
rect 1492 5083 1544 5092
rect 1492 5049 1501 5083
rect 1501 5049 1535 5083
rect 1535 5049 1544 5083
rect 1492 5040 1544 5049
rect 2780 5040 2832 5092
rect 4160 5040 4212 5092
rect 5172 5040 5224 5092
rect 1860 5015 1912 5024
rect 1860 4981 1869 5015
rect 1869 4981 1903 5015
rect 1903 4981 1912 5015
rect 1860 4972 1912 4981
rect 3056 4972 3108 5024
rect 4068 4972 4120 5024
rect 4528 4972 4580 5024
rect 10508 5108 10560 5160
rect 11612 5108 11664 5160
rect 15016 5244 15068 5296
rect 7564 5040 7616 5092
rect 7104 4972 7156 5024
rect 7472 4972 7524 5024
rect 9036 4972 9088 5024
rect 9588 4972 9640 5024
rect 12624 5040 12676 5092
rect 10692 4972 10744 5024
rect 10968 5015 11020 5024
rect 10968 4981 10977 5015
rect 10977 4981 11011 5015
rect 11011 4981 11020 5015
rect 10968 4972 11020 4981
rect 11336 5015 11388 5024
rect 11336 4981 11345 5015
rect 11345 4981 11379 5015
rect 11379 4981 11388 5015
rect 11336 4972 11388 4981
rect 12440 4972 12492 5024
rect 12716 5015 12768 5024
rect 12716 4981 12725 5015
rect 12725 4981 12759 5015
rect 12759 4981 12768 5015
rect 12716 4972 12768 4981
rect 13268 5151 13320 5160
rect 13268 5117 13277 5151
rect 13277 5117 13311 5151
rect 13311 5117 13320 5151
rect 13268 5108 13320 5117
rect 13820 5108 13872 5160
rect 14740 5176 14792 5228
rect 15660 5219 15712 5228
rect 15660 5185 15668 5219
rect 15668 5185 15712 5219
rect 15660 5176 15712 5185
rect 16304 5312 16356 5364
rect 16672 5312 16724 5364
rect 17132 5355 17184 5364
rect 17132 5321 17141 5355
rect 17141 5321 17175 5355
rect 17175 5321 17184 5355
rect 17132 5312 17184 5321
rect 17500 5312 17552 5364
rect 18512 5312 18564 5364
rect 16212 5176 16264 5228
rect 17316 5244 17368 5296
rect 17868 5176 17920 5228
rect 14924 5108 14976 5160
rect 15292 5040 15344 5092
rect 14004 4972 14056 5024
rect 15384 5015 15436 5024
rect 15384 4981 15393 5015
rect 15393 4981 15427 5015
rect 15427 4981 15436 5015
rect 15384 4972 15436 4981
rect 15476 4972 15528 5024
rect 17316 5151 17368 5160
rect 17316 5117 17325 5151
rect 17325 5117 17359 5151
rect 17359 5117 17368 5151
rect 18052 5151 18104 5160
rect 17316 5108 17368 5117
rect 18052 5117 18061 5151
rect 18061 5117 18095 5151
rect 18095 5117 18104 5151
rect 18052 5108 18104 5117
rect 18788 5176 18840 5228
rect 18236 5040 18288 5092
rect 16304 4972 16356 5024
rect 18144 4972 18196 5024
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 3430 4870 3482 4922
rect 7622 4870 7674 4922
rect 7686 4870 7738 4922
rect 7750 4870 7802 4922
rect 7814 4870 7866 4922
rect 7878 4870 7930 4922
rect 12070 4870 12122 4922
rect 12134 4870 12186 4922
rect 12198 4870 12250 4922
rect 12262 4870 12314 4922
rect 12326 4870 12378 4922
rect 16518 4870 16570 4922
rect 16582 4870 16634 4922
rect 16646 4870 16698 4922
rect 16710 4870 16762 4922
rect 16774 4870 16826 4922
rect 1768 4811 1820 4820
rect 1768 4777 1777 4811
rect 1777 4777 1811 4811
rect 1811 4777 1820 4811
rect 1768 4768 1820 4777
rect 2044 4811 2096 4820
rect 2044 4777 2053 4811
rect 2053 4777 2087 4811
rect 2087 4777 2096 4811
rect 2044 4768 2096 4777
rect 3700 4768 3752 4820
rect 4068 4811 4120 4820
rect 4068 4777 4077 4811
rect 4077 4777 4111 4811
rect 4111 4777 4120 4811
rect 4068 4768 4120 4777
rect 4436 4811 4488 4820
rect 4436 4777 4445 4811
rect 4445 4777 4479 4811
rect 4479 4777 4488 4811
rect 4436 4768 4488 4777
rect 4896 4768 4948 4820
rect 8484 4768 8536 4820
rect 8944 4811 8996 4820
rect 8944 4777 8953 4811
rect 8953 4777 8987 4811
rect 8987 4777 8996 4811
rect 8944 4768 8996 4777
rect 9680 4811 9732 4820
rect 9680 4777 9689 4811
rect 9689 4777 9723 4811
rect 9723 4777 9732 4811
rect 9680 4768 9732 4777
rect 10784 4768 10836 4820
rect 2044 4564 2096 4616
rect 2228 4607 2280 4616
rect 2228 4573 2237 4607
rect 2237 4573 2271 4607
rect 2271 4573 2280 4607
rect 2228 4564 2280 4573
rect 2780 4564 2832 4616
rect 7288 4700 7340 4752
rect 2964 4632 3016 4684
rect 4988 4675 5040 4684
rect 4988 4641 4997 4675
rect 4997 4641 5031 4675
rect 5031 4641 5040 4675
rect 4988 4632 5040 4641
rect 5264 4632 5316 4684
rect 4712 4564 4764 4616
rect 6092 4564 6144 4616
rect 6920 4564 6972 4616
rect 7288 4564 7340 4616
rect 8116 4564 8168 4616
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 2412 4428 2464 4480
rect 2688 4471 2740 4480
rect 2688 4437 2697 4471
rect 2697 4437 2731 4471
rect 2731 4437 2740 4471
rect 2688 4428 2740 4437
rect 2780 4428 2832 4480
rect 2964 4471 3016 4480
rect 2964 4437 2973 4471
rect 2973 4437 3007 4471
rect 3007 4437 3016 4471
rect 2964 4428 3016 4437
rect 3056 4428 3108 4480
rect 4160 4471 4212 4480
rect 4160 4437 4169 4471
rect 4169 4437 4203 4471
rect 4203 4437 4212 4471
rect 4160 4428 4212 4437
rect 5264 4496 5316 4548
rect 8576 4496 8628 4548
rect 5816 4428 5868 4480
rect 6920 4428 6972 4480
rect 9128 4564 9180 4616
rect 9680 4564 9732 4616
rect 11152 4564 11204 4616
rect 12624 4768 12676 4820
rect 13452 4768 13504 4820
rect 17132 4768 17184 4820
rect 18420 4811 18472 4820
rect 18420 4777 18429 4811
rect 18429 4777 18463 4811
rect 18463 4777 18472 4811
rect 18420 4768 18472 4777
rect 11796 4700 11848 4752
rect 13728 4700 13780 4752
rect 18144 4700 18196 4752
rect 11888 4632 11940 4684
rect 12440 4632 12492 4684
rect 15384 4632 15436 4684
rect 16304 4675 16356 4684
rect 16304 4641 16313 4675
rect 16313 4641 16347 4675
rect 16347 4641 16356 4675
rect 16304 4632 16356 4641
rect 16856 4675 16908 4684
rect 16856 4641 16865 4675
rect 16865 4641 16899 4675
rect 16899 4641 16908 4675
rect 16856 4632 16908 4641
rect 18696 4632 18748 4684
rect 12256 4564 12308 4616
rect 12716 4564 12768 4616
rect 13176 4564 13228 4616
rect 13636 4607 13688 4616
rect 13636 4573 13645 4607
rect 13645 4573 13679 4607
rect 13679 4573 13688 4607
rect 13636 4564 13688 4573
rect 16028 4607 16080 4616
rect 16028 4573 16037 4607
rect 16037 4573 16071 4607
rect 16071 4573 16080 4607
rect 16028 4564 16080 4573
rect 18328 4564 18380 4616
rect 10968 4496 11020 4548
rect 10876 4428 10928 4480
rect 11888 4428 11940 4480
rect 13176 4428 13228 4480
rect 15108 4496 15160 4548
rect 15384 4428 15436 4480
rect 5398 4326 5450 4378
rect 5462 4326 5514 4378
rect 5526 4326 5578 4378
rect 5590 4326 5642 4378
rect 5654 4326 5706 4378
rect 9846 4326 9898 4378
rect 9910 4326 9962 4378
rect 9974 4326 10026 4378
rect 10038 4326 10090 4378
rect 10102 4326 10154 4378
rect 14294 4326 14346 4378
rect 14358 4326 14410 4378
rect 14422 4326 14474 4378
rect 14486 4326 14538 4378
rect 14550 4326 14602 4378
rect 2780 4224 2832 4276
rect 4528 4224 4580 4276
rect 5172 4224 5224 4276
rect 6000 4224 6052 4276
rect 9404 4267 9456 4276
rect 9404 4233 9413 4267
rect 9413 4233 9447 4267
rect 9447 4233 9456 4267
rect 9404 4224 9456 4233
rect 12072 4224 12124 4276
rect 12256 4224 12308 4276
rect 12900 4224 12952 4276
rect 15568 4224 15620 4276
rect 15936 4224 15988 4276
rect 16120 4224 16172 4276
rect 2136 4088 2188 4140
rect 2228 4088 2280 4140
rect 2780 4088 2832 4140
rect 2964 4020 3016 4072
rect 3608 4088 3660 4140
rect 4712 4156 4764 4208
rect 3792 4088 3844 4140
rect 3884 4088 3936 4140
rect 4160 4131 4212 4140
rect 4160 4097 4169 4131
rect 4169 4097 4203 4131
rect 4203 4097 4212 4131
rect 4160 4088 4212 4097
rect 5540 4156 5592 4208
rect 7380 4156 7432 4208
rect 2044 3952 2096 4004
rect 1492 3927 1544 3936
rect 1492 3893 1501 3927
rect 1501 3893 1535 3927
rect 1535 3893 1544 3927
rect 1492 3884 1544 3893
rect 1584 3884 1636 3936
rect 1952 3884 2004 3936
rect 2228 3884 2280 3936
rect 2504 3884 2556 3936
rect 2964 3927 3016 3936
rect 2964 3893 2973 3927
rect 2973 3893 3007 3927
rect 3007 3893 3016 3927
rect 2964 3884 3016 3893
rect 3792 3995 3844 4004
rect 3792 3961 3801 3995
rect 3801 3961 3835 3995
rect 3835 3961 3844 3995
rect 3792 3952 3844 3961
rect 4620 3995 4672 4004
rect 4620 3961 4629 3995
rect 4629 3961 4663 3995
rect 4663 3961 4672 3995
rect 4620 3952 4672 3961
rect 5356 4020 5408 4072
rect 5816 4020 5868 4072
rect 6092 4088 6144 4140
rect 6552 4088 6604 4140
rect 6736 4131 6788 4140
rect 6736 4097 6770 4131
rect 6770 4097 6788 4131
rect 6736 4088 6788 4097
rect 6276 3952 6328 4004
rect 8576 4131 8628 4140
rect 8576 4097 8585 4131
rect 8585 4097 8619 4131
rect 8619 4097 8628 4131
rect 8576 4088 8628 4097
rect 9680 4088 9732 4140
rect 10232 4131 10284 4140
rect 10232 4097 10241 4131
rect 10241 4097 10275 4131
rect 10275 4097 10284 4131
rect 10232 4088 10284 4097
rect 10508 4131 10560 4140
rect 10508 4097 10517 4131
rect 10517 4097 10551 4131
rect 10551 4097 10560 4131
rect 10508 4088 10560 4097
rect 11244 4088 11296 4140
rect 11980 4131 12032 4140
rect 8024 3952 8076 4004
rect 10876 4020 10928 4072
rect 11060 4020 11112 4072
rect 11520 4020 11572 4072
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 13636 4156 13688 4208
rect 15016 4156 15068 4208
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 14648 4131 14700 4140
rect 14648 4097 14657 4131
rect 14657 4097 14691 4131
rect 14691 4097 14700 4131
rect 14648 4088 14700 4097
rect 15108 4088 15160 4140
rect 5540 3884 5592 3936
rect 5908 3927 5960 3936
rect 5908 3893 5917 3927
rect 5917 3893 5951 3927
rect 5951 3893 5960 3927
rect 5908 3884 5960 3893
rect 6828 3884 6880 3936
rect 9128 3927 9180 3936
rect 9128 3893 9137 3927
rect 9137 3893 9171 3927
rect 9171 3893 9180 3927
rect 9128 3884 9180 3893
rect 10324 3952 10376 4004
rect 11244 3952 11296 4004
rect 12624 4020 12676 4072
rect 12808 4063 12860 4072
rect 12808 4029 12817 4063
rect 12817 4029 12851 4063
rect 12851 4029 12860 4063
rect 12808 4020 12860 4029
rect 12992 4063 13044 4072
rect 12992 4029 13001 4063
rect 13001 4029 13035 4063
rect 13035 4029 13044 4063
rect 12992 4020 13044 4029
rect 13912 4020 13964 4072
rect 14924 4063 14976 4072
rect 14924 4029 14933 4063
rect 14933 4029 14967 4063
rect 14967 4029 14976 4063
rect 14924 4020 14976 4029
rect 10140 3884 10192 3936
rect 10784 3927 10836 3936
rect 10784 3893 10793 3927
rect 10793 3893 10827 3927
rect 10827 3893 10836 3927
rect 10784 3884 10836 3893
rect 11704 3884 11756 3936
rect 16396 4088 16448 4140
rect 17040 4088 17092 4140
rect 16672 4063 16724 4072
rect 16672 4029 16681 4063
rect 16681 4029 16715 4063
rect 16715 4029 16724 4063
rect 16672 4020 16724 4029
rect 16856 4063 16908 4072
rect 16856 4029 16865 4063
rect 16865 4029 16899 4063
rect 16899 4029 16908 4063
rect 16856 4020 16908 4029
rect 17592 4088 17644 4140
rect 18236 4131 18288 4140
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 12440 3884 12492 3936
rect 12716 3927 12768 3936
rect 12716 3893 12725 3927
rect 12725 3893 12759 3927
rect 12759 3893 12768 3927
rect 12716 3884 12768 3893
rect 12900 3884 12952 3936
rect 17868 3952 17920 4004
rect 16028 3927 16080 3936
rect 16028 3893 16037 3927
rect 16037 3893 16071 3927
rect 16071 3893 16080 3927
rect 16304 3927 16356 3936
rect 16028 3884 16080 3893
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 17684 3927 17736 3936
rect 17684 3893 17693 3927
rect 17693 3893 17727 3927
rect 17727 3893 17736 3927
rect 17684 3884 17736 3893
rect 17776 3884 17828 3936
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 3430 3782 3482 3834
rect 7622 3782 7674 3834
rect 7686 3782 7738 3834
rect 7750 3782 7802 3834
rect 7814 3782 7866 3834
rect 7878 3782 7930 3834
rect 12070 3782 12122 3834
rect 12134 3782 12186 3834
rect 12198 3782 12250 3834
rect 12262 3782 12314 3834
rect 12326 3782 12378 3834
rect 16518 3782 16570 3834
rect 16582 3782 16634 3834
rect 16646 3782 16698 3834
rect 16710 3782 16762 3834
rect 16774 3782 16826 3834
rect 2872 3680 2924 3732
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 5356 3723 5408 3732
rect 5356 3689 5365 3723
rect 5365 3689 5399 3723
rect 5399 3689 5408 3723
rect 5356 3680 5408 3689
rect 6736 3680 6788 3732
rect 8024 3680 8076 3732
rect 10232 3680 10284 3732
rect 12992 3680 13044 3732
rect 2228 3544 2280 3596
rect 2596 3519 2648 3528
rect 2596 3485 2605 3519
rect 2605 3485 2639 3519
rect 2639 3485 2648 3519
rect 2596 3476 2648 3485
rect 3148 3476 3200 3528
rect 3424 3476 3476 3528
rect 3884 3476 3936 3528
rect 6092 3476 6144 3528
rect 7012 3544 7064 3596
rect 8024 3544 8076 3596
rect 7104 3476 7156 3528
rect 8852 3544 8904 3596
rect 9680 3612 9732 3664
rect 10048 3612 10100 3664
rect 10324 3612 10376 3664
rect 12440 3612 12492 3664
rect 17224 3680 17276 3732
rect 18420 3723 18472 3732
rect 18420 3689 18429 3723
rect 18429 3689 18463 3723
rect 18463 3689 18472 3723
rect 18420 3680 18472 3689
rect 13728 3612 13780 3664
rect 16304 3612 16356 3664
rect 18604 3612 18656 3664
rect 11060 3544 11112 3596
rect 13912 3544 13964 3596
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 15476 3587 15528 3596
rect 15476 3553 15485 3587
rect 15485 3553 15519 3587
rect 15519 3553 15528 3587
rect 15476 3544 15528 3553
rect 1492 3383 1544 3392
rect 1492 3349 1501 3383
rect 1501 3349 1535 3383
rect 1535 3349 1544 3383
rect 1492 3340 1544 3349
rect 1860 3383 1912 3392
rect 1860 3349 1869 3383
rect 1869 3349 1903 3383
rect 1903 3349 1912 3383
rect 1860 3340 1912 3349
rect 2780 3383 2832 3392
rect 2780 3349 2789 3383
rect 2789 3349 2823 3383
rect 2823 3349 2832 3383
rect 4712 3408 4764 3460
rect 2780 3340 2832 3349
rect 5172 3340 5224 3392
rect 6920 3408 6972 3460
rect 8300 3476 8352 3528
rect 7932 3408 7984 3460
rect 10048 3476 10100 3528
rect 10232 3476 10284 3528
rect 10968 3476 11020 3528
rect 11152 3476 11204 3528
rect 12256 3519 12308 3528
rect 12256 3485 12300 3519
rect 12300 3485 12308 3519
rect 12256 3476 12308 3485
rect 9496 3408 9548 3460
rect 7196 3340 7248 3392
rect 8392 3383 8444 3392
rect 8392 3349 8401 3383
rect 8401 3349 8435 3383
rect 8435 3349 8444 3383
rect 8392 3340 8444 3349
rect 9588 3340 9640 3392
rect 11704 3408 11756 3460
rect 11888 3451 11940 3460
rect 11888 3417 11906 3451
rect 11906 3417 11940 3451
rect 11888 3408 11940 3417
rect 12072 3408 12124 3460
rect 12716 3476 12768 3528
rect 12992 3476 13044 3528
rect 13176 3476 13228 3528
rect 13544 3476 13596 3528
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 15200 3519 15252 3528
rect 15200 3485 15209 3519
rect 15209 3485 15243 3519
rect 15243 3485 15252 3519
rect 15200 3476 15252 3485
rect 10600 3383 10652 3392
rect 10600 3349 10609 3383
rect 10609 3349 10643 3383
rect 10643 3349 10652 3383
rect 10600 3340 10652 3349
rect 10784 3383 10836 3392
rect 10784 3349 10793 3383
rect 10793 3349 10827 3383
rect 10827 3349 10836 3383
rect 10784 3340 10836 3349
rect 11152 3340 11204 3392
rect 11520 3340 11572 3392
rect 12900 3340 12952 3392
rect 14188 3408 14240 3460
rect 17592 3544 17644 3596
rect 17316 3476 17368 3528
rect 17408 3476 17460 3528
rect 17684 3476 17736 3528
rect 18144 3476 18196 3528
rect 17132 3451 17184 3460
rect 13360 3340 13412 3392
rect 13636 3383 13688 3392
rect 13636 3349 13645 3383
rect 13645 3349 13679 3383
rect 13679 3349 13688 3383
rect 13636 3340 13688 3349
rect 17132 3417 17141 3451
rect 17141 3417 17175 3451
rect 17175 3417 17184 3451
rect 17132 3408 17184 3417
rect 19616 3408 19668 3460
rect 17500 3340 17552 3392
rect 17592 3340 17644 3392
rect 18052 3383 18104 3392
rect 18052 3349 18061 3383
rect 18061 3349 18095 3383
rect 18095 3349 18104 3383
rect 18052 3340 18104 3349
rect 5398 3238 5450 3290
rect 5462 3238 5514 3290
rect 5526 3238 5578 3290
rect 5590 3238 5642 3290
rect 5654 3238 5706 3290
rect 9846 3238 9898 3290
rect 9910 3238 9962 3290
rect 9974 3238 10026 3290
rect 10038 3238 10090 3290
rect 10102 3238 10154 3290
rect 14294 3238 14346 3290
rect 14358 3238 14410 3290
rect 14422 3238 14474 3290
rect 14486 3238 14538 3290
rect 14550 3238 14602 3290
rect 204 3136 256 3188
rect 3148 3136 3200 3188
rect 4620 3179 4672 3188
rect 4620 3145 4629 3179
rect 4629 3145 4663 3179
rect 4663 3145 4672 3179
rect 4620 3136 4672 3145
rect 4896 3136 4948 3188
rect 5264 3179 5316 3188
rect 5264 3145 5273 3179
rect 5273 3145 5307 3179
rect 5307 3145 5316 3179
rect 5264 3136 5316 3145
rect 7196 3136 7248 3188
rect 1952 3000 2004 3052
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2412 3043 2464 3052
rect 2044 3000 2096 3009
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 3056 3068 3108 3120
rect 2964 3000 3016 3052
rect 3240 3043 3292 3052
rect 3240 3009 3249 3043
rect 3249 3009 3283 3043
rect 3283 3009 3292 3043
rect 3240 3000 3292 3009
rect 4068 3000 4120 3052
rect 4252 3000 4304 3052
rect 6920 3043 6972 3052
rect 664 2932 716 2984
rect 1124 2864 1176 2916
rect 3424 2932 3476 2984
rect 5908 2975 5960 2984
rect 5908 2941 5917 2975
rect 5917 2941 5951 2975
rect 5951 2941 5960 2975
rect 5908 2932 5960 2941
rect 1492 2839 1544 2848
rect 1492 2805 1501 2839
rect 1501 2805 1535 2839
rect 1535 2805 1544 2839
rect 1492 2796 1544 2805
rect 2964 2839 3016 2848
rect 2964 2805 2973 2839
rect 2973 2805 3007 2839
rect 3007 2805 3016 2839
rect 2964 2796 3016 2805
rect 3056 2796 3108 2848
rect 3976 2839 4028 2848
rect 3976 2805 3985 2839
rect 3985 2805 4019 2839
rect 4019 2805 4028 2839
rect 3976 2796 4028 2805
rect 4252 2839 4304 2848
rect 4252 2805 4261 2839
rect 4261 2805 4295 2839
rect 4295 2805 4304 2839
rect 4252 2796 4304 2805
rect 4620 2796 4672 2848
rect 5724 2796 5776 2848
rect 6920 3009 6929 3043
rect 6929 3009 6963 3043
rect 6963 3009 6972 3043
rect 9404 3068 9456 3120
rect 10232 3136 10284 3188
rect 14924 3136 14976 3188
rect 15016 3136 15068 3188
rect 18328 3136 18380 3188
rect 12256 3068 12308 3120
rect 12900 3068 12952 3120
rect 16028 3068 16080 3120
rect 19156 3068 19208 3120
rect 6920 3000 6972 3009
rect 9036 3000 9088 3052
rect 10876 3000 10928 3052
rect 11152 3000 11204 3052
rect 11336 3000 11388 3052
rect 13452 3043 13504 3052
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 15568 3043 15620 3052
rect 15568 3009 15577 3043
rect 15577 3009 15611 3043
rect 15611 3009 15620 3043
rect 15568 3000 15620 3009
rect 15660 3000 15712 3052
rect 16304 3043 16356 3052
rect 16304 3009 16313 3043
rect 16313 3009 16347 3043
rect 16347 3009 16356 3043
rect 16304 3000 16356 3009
rect 16948 3000 17000 3052
rect 17132 3043 17184 3052
rect 17132 3009 17141 3043
rect 17141 3009 17175 3043
rect 17175 3009 17184 3043
rect 17132 3000 17184 3009
rect 17500 3043 17552 3052
rect 17500 3009 17509 3043
rect 17509 3009 17543 3043
rect 17543 3009 17552 3043
rect 17500 3000 17552 3009
rect 17868 3043 17920 3052
rect 17868 3009 17877 3043
rect 17877 3009 17911 3043
rect 17911 3009 17920 3043
rect 17868 3000 17920 3009
rect 17960 3000 18012 3052
rect 7932 2975 7984 2984
rect 7932 2941 7941 2975
rect 7941 2941 7975 2975
rect 7975 2941 7984 2975
rect 7932 2932 7984 2941
rect 9220 2975 9272 2984
rect 9220 2941 9229 2975
rect 9229 2941 9263 2975
rect 9263 2941 9272 2975
rect 9220 2932 9272 2941
rect 9588 2932 9640 2984
rect 10968 2932 11020 2984
rect 11704 2975 11756 2984
rect 11704 2941 11713 2975
rect 11713 2941 11747 2975
rect 11747 2941 11756 2975
rect 11704 2932 11756 2941
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 13268 2932 13320 2984
rect 13912 2932 13964 2984
rect 15108 2975 15160 2984
rect 15108 2941 15117 2975
rect 15117 2941 15151 2975
rect 15151 2941 15160 2975
rect 15108 2932 15160 2941
rect 6736 2864 6788 2916
rect 7288 2864 7340 2916
rect 7380 2864 7432 2916
rect 8208 2864 8260 2916
rect 10784 2864 10836 2916
rect 11152 2907 11204 2916
rect 6920 2796 6972 2848
rect 7104 2839 7156 2848
rect 7104 2805 7113 2839
rect 7113 2805 7147 2839
rect 7147 2805 7156 2839
rect 7104 2796 7156 2805
rect 7472 2796 7524 2848
rect 8484 2796 8536 2848
rect 9036 2796 9088 2848
rect 11152 2873 11161 2907
rect 11161 2873 11195 2907
rect 11195 2873 11204 2907
rect 11152 2864 11204 2873
rect 11060 2796 11112 2848
rect 12900 2864 12952 2916
rect 12992 2864 13044 2916
rect 13544 2864 13596 2916
rect 15016 2864 15068 2916
rect 15844 2864 15896 2916
rect 16948 2839 17000 2848
rect 16948 2805 16957 2839
rect 16957 2805 16991 2839
rect 16991 2805 17000 2839
rect 16948 2796 17000 2805
rect 17316 2839 17368 2848
rect 17316 2805 17325 2839
rect 17325 2805 17359 2839
rect 17359 2805 17368 2839
rect 17316 2796 17368 2805
rect 17776 2796 17828 2848
rect 17868 2796 17920 2848
rect 18420 2839 18472 2848
rect 18420 2805 18429 2839
rect 18429 2805 18463 2839
rect 18463 2805 18472 2839
rect 18420 2796 18472 2805
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 3430 2694 3482 2746
rect 7622 2694 7674 2746
rect 7686 2694 7738 2746
rect 7750 2694 7802 2746
rect 7814 2694 7866 2746
rect 7878 2694 7930 2746
rect 12070 2694 12122 2746
rect 12134 2694 12186 2746
rect 12198 2694 12250 2746
rect 12262 2694 12314 2746
rect 12326 2694 12378 2746
rect 16518 2694 16570 2746
rect 16582 2694 16634 2746
rect 16646 2694 16698 2746
rect 16710 2694 16762 2746
rect 16774 2694 16826 2746
rect 2320 2592 2372 2644
rect 4712 2635 4764 2644
rect 4712 2601 4721 2635
rect 4721 2601 4755 2635
rect 4755 2601 4764 2635
rect 4712 2592 4764 2601
rect 5908 2635 5960 2644
rect 5908 2601 5917 2635
rect 5917 2601 5951 2635
rect 5951 2601 5960 2635
rect 5908 2592 5960 2601
rect 10968 2592 11020 2644
rect 12532 2635 12584 2644
rect 12532 2601 12541 2635
rect 12541 2601 12575 2635
rect 12575 2601 12584 2635
rect 12532 2592 12584 2601
rect 12808 2592 12860 2644
rect 15108 2592 15160 2644
rect 2504 2524 2556 2576
rect 3884 2524 3936 2576
rect 10232 2524 10284 2576
rect 3976 2456 4028 2508
rect 4620 2456 4672 2508
rect 2688 2388 2740 2440
rect 3516 2431 3568 2440
rect 3516 2397 3525 2431
rect 3525 2397 3559 2431
rect 3559 2397 3568 2431
rect 3516 2388 3568 2397
rect 4252 2388 4304 2440
rect 4804 2388 4856 2440
rect 5172 2431 5224 2440
rect 5172 2397 5181 2431
rect 5181 2397 5215 2431
rect 5215 2397 5224 2431
rect 5172 2388 5224 2397
rect 8208 2456 8260 2508
rect 9772 2499 9824 2508
rect 9772 2465 9781 2499
rect 9781 2465 9815 2499
rect 9815 2465 9824 2499
rect 9772 2456 9824 2465
rect 10324 2456 10376 2508
rect 5724 2431 5776 2440
rect 5724 2397 5733 2431
rect 5733 2397 5767 2431
rect 5767 2397 5776 2431
rect 5724 2388 5776 2397
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 7196 2431 7248 2440
rect 6736 2388 6788 2397
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 7288 2388 7340 2440
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 9036 2431 9088 2440
rect 8484 2388 8536 2397
rect 9036 2397 9045 2431
rect 9045 2397 9079 2431
rect 9079 2397 9088 2431
rect 9036 2388 9088 2397
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 10600 2388 10652 2440
rect 2872 2320 2924 2372
rect 10416 2363 10468 2372
rect 10416 2329 10425 2363
rect 10425 2329 10459 2363
rect 10459 2329 10468 2363
rect 10416 2320 10468 2329
rect 11152 2388 11204 2440
rect 15660 2524 15712 2576
rect 18972 2592 19024 2644
rect 12348 2499 12400 2508
rect 12348 2465 12357 2499
rect 12357 2465 12391 2499
rect 12391 2465 12400 2499
rect 12348 2456 12400 2465
rect 12624 2456 12676 2508
rect 14096 2499 14148 2508
rect 11888 2388 11940 2440
rect 1492 2295 1544 2304
rect 1492 2261 1501 2295
rect 1501 2261 1535 2295
rect 1535 2261 1544 2295
rect 1492 2252 1544 2261
rect 1676 2252 1728 2304
rect 2136 2252 2188 2304
rect 2688 2252 2740 2304
rect 3148 2252 3200 2304
rect 3608 2252 3660 2304
rect 4160 2252 4212 2304
rect 5172 2252 5224 2304
rect 6092 2295 6144 2304
rect 6092 2261 6101 2295
rect 6101 2261 6135 2295
rect 6135 2261 6144 2295
rect 6092 2252 6144 2261
rect 6184 2252 6236 2304
rect 6644 2252 6696 2304
rect 7104 2252 7156 2304
rect 7564 2295 7616 2304
rect 7564 2261 7573 2295
rect 7573 2261 7607 2295
rect 7607 2261 7616 2295
rect 7564 2252 7616 2261
rect 7656 2252 7708 2304
rect 8116 2252 8168 2304
rect 8668 2295 8720 2304
rect 8668 2261 8677 2295
rect 8677 2261 8711 2295
rect 8711 2261 8720 2295
rect 8668 2252 8720 2261
rect 9128 2252 9180 2304
rect 9680 2252 9732 2304
rect 10508 2295 10560 2304
rect 10508 2261 10517 2295
rect 10517 2261 10551 2295
rect 10551 2261 10560 2295
rect 10508 2252 10560 2261
rect 10600 2252 10652 2304
rect 10876 2252 10928 2304
rect 12900 2388 12952 2440
rect 13268 2388 13320 2440
rect 13452 2431 13504 2440
rect 13452 2397 13461 2431
rect 13461 2397 13495 2431
rect 13495 2397 13504 2431
rect 13452 2388 13504 2397
rect 14096 2465 14105 2499
rect 14105 2465 14139 2499
rect 14139 2465 14148 2499
rect 14096 2456 14148 2465
rect 16672 2524 16724 2576
rect 17132 2524 17184 2576
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 16672 2431 16724 2440
rect 16672 2397 16681 2431
rect 16681 2397 16715 2431
rect 16715 2397 16724 2431
rect 16672 2388 16724 2397
rect 16856 2388 16908 2440
rect 17224 2388 17276 2440
rect 17500 2388 17552 2440
rect 18236 2431 18288 2440
rect 18236 2397 18245 2431
rect 18245 2397 18279 2431
rect 18279 2397 18288 2431
rect 18236 2388 18288 2397
rect 15200 2252 15252 2304
rect 15660 2252 15712 2304
rect 16672 2252 16724 2304
rect 16764 2252 16816 2304
rect 17040 2252 17092 2304
rect 17684 2252 17736 2304
rect 18144 2252 18196 2304
rect 5398 2150 5450 2202
rect 5462 2150 5514 2202
rect 5526 2150 5578 2202
rect 5590 2150 5642 2202
rect 5654 2150 5706 2202
rect 9846 2150 9898 2202
rect 9910 2150 9962 2202
rect 9974 2150 10026 2202
rect 10038 2150 10090 2202
rect 10102 2150 10154 2202
rect 14294 2150 14346 2202
rect 14358 2150 14410 2202
rect 14422 2150 14474 2202
rect 14486 2150 14538 2202
rect 14550 2150 14602 2202
rect 10508 2048 10560 2100
rect 12624 2048 12676 2100
rect 15384 2048 15436 2100
rect 18236 2048 18288 2100
rect 6092 1980 6144 2032
rect 13176 1980 13228 2032
rect 13452 1980 13504 2032
rect 13636 1980 13688 2032
rect 17500 1980 17552 2032
rect 7564 1912 7616 1964
rect 11152 1912 11204 1964
rect 11888 1912 11940 1964
rect 13820 1844 13872 1896
rect 16856 1844 16908 1896
rect 10416 1776 10468 1828
rect 12992 1776 13044 1828
rect 11244 1708 11296 1760
rect 16028 1708 16080 1760
<< metal2 >>
rect 294 16400 350 17200
rect 938 16538 994 17200
rect 938 16510 1256 16538
rect 938 16400 994 16510
rect 308 13734 336 16400
rect 1228 14822 1256 16510
rect 1582 16400 1638 17200
rect 2226 16538 2282 17200
rect 2226 16510 2544 16538
rect 2226 16400 2282 16510
rect 1216 14816 1268 14822
rect 1216 14758 1268 14764
rect 1596 13802 1624 16400
rect 2226 14512 2282 14521
rect 2226 14447 2282 14456
rect 2240 14414 2268 14447
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2240 13977 2268 14350
rect 2226 13968 2282 13977
rect 2226 13903 2282 13912
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1584 13796 1636 13802
rect 1584 13738 1636 13744
rect 296 13728 348 13734
rect 296 13670 348 13676
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 1964 12889 1992 13262
rect 1950 12880 2006 12889
rect 1950 12815 2006 12824
rect 1952 11144 2004 11150
rect 1950 11112 1952 11121
rect 2004 11112 2006 11121
rect 1950 11047 2006 11056
rect 1582 10704 1638 10713
rect 1582 10639 1584 10648
rect 1636 10639 1638 10648
rect 1584 10610 1636 10616
rect 1490 10568 1546 10577
rect 1490 10503 1546 10512
rect 1400 10464 1452 10470
rect 1400 10406 1452 10412
rect 1308 9444 1360 9450
rect 1308 9386 1360 9392
rect 1320 9353 1348 9386
rect 1306 9344 1362 9353
rect 1306 9279 1362 9288
rect 1412 7410 1440 10406
rect 1504 10062 1532 10503
rect 2056 10266 2084 13806
rect 2516 13394 2544 16510
rect 2870 16400 2926 17200
rect 3514 16400 3570 17200
rect 3790 16824 3846 16833
rect 3790 16759 3846 16768
rect 2688 14476 2740 14482
rect 2688 14418 2740 14424
rect 2700 13410 2728 14418
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13569 2820 13806
rect 2778 13560 2834 13569
rect 2884 13530 2912 16400
rect 3054 16008 3110 16017
rect 3054 15943 3110 15952
rect 2962 14784 3018 14793
rect 2962 14719 3018 14728
rect 2976 14482 3004 14719
rect 2964 14476 3016 14482
rect 3068 14464 3096 15943
rect 3174 14716 3482 14736
rect 3174 14714 3180 14716
rect 3236 14714 3260 14716
rect 3316 14714 3340 14716
rect 3396 14714 3420 14716
rect 3476 14714 3482 14716
rect 3236 14662 3238 14714
rect 3418 14662 3420 14714
rect 3174 14660 3180 14662
rect 3236 14660 3260 14662
rect 3316 14660 3340 14662
rect 3396 14660 3420 14662
rect 3476 14660 3482 14662
rect 3174 14640 3482 14660
rect 3528 14618 3556 16400
rect 3804 15230 3832 16759
rect 4158 16538 4214 17200
rect 4158 16510 4384 16538
rect 3882 16416 3938 16425
rect 4158 16400 4214 16510
rect 3882 16351 3938 16360
rect 3792 15224 3844 15230
rect 3606 15192 3662 15201
rect 3792 15166 3844 15172
rect 3606 15127 3662 15136
rect 3620 15026 3648 15127
rect 3608 15020 3660 15026
rect 3608 14962 3660 14968
rect 3516 14612 3568 14618
rect 3516 14554 3568 14560
rect 3068 14436 3556 14464
rect 2964 14418 3016 14424
rect 3054 14376 3110 14385
rect 3054 14311 3110 14320
rect 3422 14376 3478 14385
rect 3422 14311 3424 14320
rect 2778 13495 2834 13504
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 3068 13444 3096 14311
rect 3476 14311 3478 14320
rect 3424 14282 3476 14288
rect 3174 13628 3482 13648
rect 3174 13626 3180 13628
rect 3236 13626 3260 13628
rect 3316 13626 3340 13628
rect 3396 13626 3420 13628
rect 3476 13626 3482 13628
rect 3236 13574 3238 13626
rect 3418 13574 3420 13626
rect 3174 13572 3180 13574
rect 3236 13572 3260 13574
rect 3316 13572 3340 13574
rect 3396 13572 3420 13574
rect 3476 13572 3482 13574
rect 3174 13552 3482 13572
rect 2962 13424 3018 13433
rect 2504 13388 2556 13394
rect 2700 13382 2912 13410
rect 2504 13330 2556 13336
rect 2228 13320 2280 13326
rect 2228 13262 2280 13268
rect 2778 13288 2834 13297
rect 2240 13190 2268 13262
rect 2778 13223 2834 13232
rect 2228 13184 2280 13190
rect 2226 13152 2228 13161
rect 2280 13152 2282 13161
rect 2226 13087 2282 13096
rect 2240 13061 2268 13087
rect 2136 12776 2188 12782
rect 2228 12776 2280 12782
rect 2136 12718 2188 12724
rect 2226 12744 2228 12753
rect 2280 12744 2282 12753
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 1858 10160 1914 10169
rect 1858 10095 1914 10104
rect 1872 10062 1900 10095
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1860 10056 1912 10062
rect 1860 9998 1912 10004
rect 1504 8090 1532 9998
rect 1768 9512 1820 9518
rect 1768 9454 1820 9460
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 8974 1624 9318
rect 1780 8974 1808 9454
rect 1872 9178 1900 9998
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 1860 9172 1912 9178
rect 1860 9114 1912 9120
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1596 8430 1624 8774
rect 1674 8528 1730 8537
rect 1674 8463 1730 8472
rect 1584 8424 1636 8430
rect 1584 8366 1636 8372
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1596 7886 1624 8366
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1490 7712 1546 7721
rect 1490 7647 1546 7656
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1504 7002 1532 7647
rect 1688 7546 1716 8463
rect 1858 8120 1914 8129
rect 1858 8055 1914 8064
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1492 6996 1544 7002
rect 1492 6938 1544 6944
rect 1780 6798 1808 7686
rect 1872 7546 1900 8055
rect 1950 7848 2006 7857
rect 1950 7783 2006 7792
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 1872 6497 1900 6598
rect 1858 6488 1914 6497
rect 1858 6423 1914 6432
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1860 6316 1912 6322
rect 1860 6258 1912 6264
rect 1492 6112 1544 6118
rect 1490 6080 1492 6089
rect 1544 6080 1546 6089
rect 1490 6015 1546 6024
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 1544 5536 1546 5545
rect 1490 5471 1546 5480
rect 1688 5370 1716 6258
rect 1872 6225 1900 6258
rect 1858 6216 1914 6225
rect 1858 6151 1914 6160
rect 1768 5704 1820 5710
rect 1766 5672 1768 5681
rect 1820 5672 1822 5681
rect 1964 5658 1992 7783
rect 2056 7410 2084 9862
rect 2148 8537 2176 12718
rect 2226 12679 2282 12688
rect 2792 12594 2820 13223
rect 2700 12566 2820 12594
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2228 11688 2280 11694
rect 2228 11630 2280 11636
rect 2240 11393 2268 11630
rect 2226 11384 2282 11393
rect 2226 11319 2282 11328
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2240 10985 2268 11086
rect 2226 10976 2282 10985
rect 2226 10911 2282 10920
rect 2332 10810 2360 12038
rect 2424 11898 2452 12038
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2516 11354 2544 12106
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2320 10804 2372 10810
rect 2320 10746 2372 10752
rect 2424 10062 2452 10950
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2320 10056 2372 10062
rect 2318 10024 2320 10033
rect 2412 10056 2464 10062
rect 2372 10024 2374 10033
rect 2228 9988 2280 9994
rect 2412 9998 2464 10004
rect 2318 9959 2374 9968
rect 2228 9930 2280 9936
rect 2134 8528 2190 8537
rect 2134 8463 2190 8472
rect 2240 7993 2268 9930
rect 2424 9761 2452 9998
rect 2410 9752 2466 9761
rect 2410 9687 2466 9696
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2332 8090 2360 9522
rect 2410 9072 2466 9081
rect 2410 9007 2466 9016
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2226 7984 2282 7993
rect 2226 7919 2282 7928
rect 2320 7812 2372 7818
rect 2320 7754 2372 7760
rect 2044 7404 2096 7410
rect 2044 7346 2096 7352
rect 2226 7304 2282 7313
rect 2226 7239 2228 7248
rect 2280 7239 2282 7248
rect 2228 7210 2280 7216
rect 2332 7154 2360 7754
rect 2240 7126 2360 7154
rect 2136 6792 2188 6798
rect 2136 6734 2188 6740
rect 2148 6458 2176 6734
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2240 6338 2268 7126
rect 2320 6928 2372 6934
rect 2318 6896 2320 6905
rect 2372 6896 2374 6905
rect 2318 6831 2374 6840
rect 2240 6322 2360 6338
rect 2240 6316 2372 6322
rect 2240 6310 2320 6316
rect 2320 6258 2372 6264
rect 2136 6112 2188 6118
rect 2136 6054 2188 6060
rect 1766 5607 1822 5616
rect 1872 5630 1992 5658
rect 1676 5364 1728 5370
rect 1676 5306 1728 5312
rect 1768 5228 1820 5234
rect 1768 5170 1820 5176
rect 1490 5128 1546 5137
rect 1490 5063 1492 5072
rect 1544 5063 1546 5072
rect 1492 5034 1544 5040
rect 1780 4826 1808 5170
rect 1872 5166 1900 5630
rect 1952 5568 2004 5574
rect 1952 5510 2004 5516
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1860 5024 1912 5030
rect 1860 4966 1912 4972
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 1872 4729 1900 4966
rect 1858 4720 1914 4729
rect 1858 4655 1914 4664
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1504 4321 1532 4422
rect 1490 4312 1546 4321
rect 1490 4247 1546 4256
rect 1964 4026 1992 5510
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 2056 4826 2084 5170
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 2044 4616 2096 4622
rect 2042 4584 2044 4593
rect 2096 4584 2098 4593
rect 2042 4519 2098 4528
rect 2148 4146 2176 6054
rect 2332 5370 2360 6258
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2424 5250 2452 9007
rect 2516 8022 2544 10066
rect 2608 9625 2636 12174
rect 2700 11778 2728 12566
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2792 11937 2820 12378
rect 2778 11928 2834 11937
rect 2778 11863 2834 11872
rect 2884 11830 2912 13382
rect 3068 13416 3188 13444
rect 2962 13359 3018 13368
rect 2976 13326 3004 13359
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 3160 12850 3188 13416
rect 3528 13410 3556 14436
rect 3620 13938 3648 14962
rect 3896 14958 3924 16351
rect 4158 15600 4214 15609
rect 4158 15535 4214 15544
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 3700 14884 3752 14890
rect 3700 14826 3752 14832
rect 3712 14482 3740 14826
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 3608 13932 3660 13938
rect 3608 13874 3660 13880
rect 3896 13870 3924 14894
rect 4172 14822 4200 15535
rect 4068 14816 4120 14822
rect 4068 14758 4120 14764
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4080 14550 4108 14758
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 4172 14482 4200 14758
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 4356 14074 4384 16510
rect 4802 16400 4858 17200
rect 5446 16400 5502 17200
rect 6090 16538 6146 17200
rect 6012 16510 6146 16538
rect 4436 15088 4488 15094
rect 4436 15030 4488 15036
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4344 14068 4396 14074
rect 4344 14010 4396 14016
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 3976 13932 4028 13938
rect 3976 13874 4028 13880
rect 3700 13864 3752 13870
rect 3700 13806 3752 13812
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 3252 13382 3556 13410
rect 3252 13326 3280 13382
rect 3240 13320 3292 13326
rect 3528 13297 3556 13382
rect 3608 13388 3660 13394
rect 3608 13330 3660 13336
rect 3240 13262 3292 13268
rect 3514 13288 3570 13297
rect 3514 13223 3570 13232
rect 3516 13184 3568 13190
rect 3436 13132 3516 13138
rect 3436 13126 3568 13132
rect 3436 13110 3556 13126
rect 3436 12918 3464 13110
rect 3620 12918 3648 13330
rect 3424 12912 3476 12918
rect 3424 12854 3476 12860
rect 3608 12912 3660 12918
rect 3608 12854 3660 12860
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2976 12073 3004 12718
rect 3174 12540 3482 12560
rect 3174 12538 3180 12540
rect 3236 12538 3260 12540
rect 3316 12538 3340 12540
rect 3396 12538 3420 12540
rect 3476 12538 3482 12540
rect 3236 12486 3238 12538
rect 3418 12486 3420 12538
rect 3174 12484 3180 12486
rect 3236 12484 3260 12486
rect 3316 12484 3340 12486
rect 3396 12484 3420 12486
rect 3476 12484 3482 12486
rect 3174 12464 3482 12484
rect 3238 12336 3294 12345
rect 3620 12306 3648 12854
rect 3238 12271 3294 12280
rect 3608 12300 3660 12306
rect 3252 12238 3280 12271
rect 3608 12242 3660 12248
rect 3240 12232 3292 12238
rect 3240 12174 3292 12180
rect 3516 12232 3568 12238
rect 3516 12174 3568 12180
rect 2962 12064 3018 12073
rect 2962 11999 3018 12008
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2872 11824 2924 11830
rect 2700 11750 2820 11778
rect 2872 11766 2924 11772
rect 2688 10464 2740 10470
rect 2688 10406 2740 10412
rect 2594 9616 2650 9625
rect 2594 9551 2650 9560
rect 2700 9178 2728 10406
rect 2688 9172 2740 9178
rect 2688 9114 2740 9120
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2504 8016 2556 8022
rect 2504 7958 2556 7964
rect 2608 7546 2636 8570
rect 2700 8566 2728 8842
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2688 8424 2740 8430
rect 2688 8366 2740 8372
rect 2700 8090 2728 8366
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2792 7886 2820 11750
rect 2872 11688 2924 11694
rect 2872 11630 2924 11636
rect 2884 10266 2912 11630
rect 2976 11558 3004 11834
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 3068 11234 3096 11630
rect 3174 11452 3482 11472
rect 3174 11450 3180 11452
rect 3236 11450 3260 11452
rect 3316 11450 3340 11452
rect 3396 11450 3420 11452
rect 3476 11450 3482 11452
rect 3236 11398 3238 11450
rect 3418 11398 3420 11450
rect 3174 11396 3180 11398
rect 3236 11396 3260 11398
rect 3316 11396 3340 11398
rect 3396 11396 3420 11398
rect 3476 11396 3482 11398
rect 3174 11376 3482 11396
rect 3528 11354 3556 12174
rect 3620 11694 3648 12242
rect 3712 12170 3740 13806
rect 3988 13802 4016 13874
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3792 13252 3844 13258
rect 3792 13194 3844 13200
rect 3700 12164 3752 12170
rect 3700 12106 3752 12112
rect 3804 11898 3832 13194
rect 3884 13184 3936 13190
rect 3884 13126 3936 13132
rect 3896 12220 3924 13126
rect 4080 12986 4108 13942
rect 4172 13818 4200 14010
rect 4448 13938 4476 15030
rect 4528 14408 4580 14414
rect 4580 14368 4660 14396
rect 4528 14350 4580 14356
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4172 13790 4384 13818
rect 4160 13388 4212 13394
rect 4160 13330 4212 13336
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 3976 12232 4028 12238
rect 3896 12192 3976 12220
rect 3792 11892 3844 11898
rect 3792 11834 3844 11840
rect 3896 11830 3924 12192
rect 3976 12174 4028 12180
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3988 11898 4016 12038
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3884 11824 3936 11830
rect 3698 11792 3754 11801
rect 3884 11766 3936 11772
rect 3698 11727 3700 11736
rect 3752 11727 3754 11736
rect 3700 11698 3752 11704
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3608 11552 3660 11558
rect 3608 11494 3660 11500
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 3422 11248 3478 11257
rect 3068 11218 3188 11234
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 3056 11212 3188 11218
rect 3108 11206 3188 11212
rect 3056 11154 3108 11160
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2596 7540 2648 7546
rect 2596 7482 2648 7488
rect 2700 7426 2728 7822
rect 2608 7410 2728 7426
rect 2596 7404 2728 7410
rect 2648 7398 2728 7404
rect 2596 7346 2648 7352
rect 2608 7002 2636 7346
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2792 6914 2820 7822
rect 2700 6886 2820 6914
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2504 6316 2556 6322
rect 2504 6258 2556 6264
rect 2516 5778 2544 6258
rect 2608 6118 2636 6734
rect 2700 6458 2728 6886
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2596 6112 2648 6118
rect 2596 6054 2648 6060
rect 2608 5778 2636 6054
rect 2504 5772 2556 5778
rect 2504 5714 2556 5720
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2884 5658 2912 9522
rect 2976 9518 3004 11154
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 2964 9512 3016 9518
rect 2964 9454 3016 9460
rect 3068 9450 3096 11018
rect 3160 10810 3188 11206
rect 3422 11183 3424 11192
rect 3476 11183 3478 11192
rect 3424 11154 3476 11160
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3516 10736 3568 10742
rect 3516 10678 3568 10684
rect 3174 10364 3482 10384
rect 3174 10362 3180 10364
rect 3236 10362 3260 10364
rect 3316 10362 3340 10364
rect 3396 10362 3420 10364
rect 3476 10362 3482 10364
rect 3236 10310 3238 10362
rect 3418 10310 3420 10362
rect 3174 10308 3180 10310
rect 3236 10308 3260 10310
rect 3316 10308 3340 10310
rect 3396 10308 3420 10310
rect 3476 10308 3482 10310
rect 3174 10288 3482 10308
rect 3528 10130 3556 10678
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 3528 9382 3556 10066
rect 3620 9908 3648 11494
rect 3712 11354 3740 11698
rect 3700 11348 3752 11354
rect 3700 11290 3752 11296
rect 3896 10606 3924 11766
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3988 11665 4016 11698
rect 3974 11656 4030 11665
rect 3974 11591 4030 11600
rect 3988 11286 4016 11591
rect 4080 11354 4108 12378
rect 4172 11558 4200 13330
rect 4356 13258 4384 13790
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4448 13326 4476 13670
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4344 13252 4396 13258
rect 4344 13194 4396 13200
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4264 12220 4292 13126
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4540 12442 4568 12718
rect 4528 12436 4580 12442
rect 4528 12378 4580 12384
rect 4264 12192 4476 12220
rect 4344 12096 4396 12102
rect 4344 12038 4396 12044
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3976 11280 4028 11286
rect 3976 11222 4028 11228
rect 4066 11248 4122 11257
rect 4066 11183 4122 11192
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3700 10464 3752 10470
rect 3700 10406 3752 10412
rect 3712 10169 3740 10406
rect 3698 10160 3754 10169
rect 3698 10095 3754 10104
rect 3712 10062 3740 10095
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3792 9988 3844 9994
rect 3792 9930 3844 9936
rect 3700 9920 3752 9926
rect 3620 9880 3700 9908
rect 3700 9862 3752 9868
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3620 9489 3648 9522
rect 3606 9480 3662 9489
rect 3606 9415 3662 9424
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 3516 9376 3568 9382
rect 3516 9318 3568 9324
rect 2976 8634 3004 9318
rect 3174 9276 3482 9296
rect 3174 9274 3180 9276
rect 3236 9274 3260 9276
rect 3316 9274 3340 9276
rect 3396 9274 3420 9276
rect 3476 9274 3482 9276
rect 3236 9222 3238 9274
rect 3418 9222 3420 9274
rect 3174 9220 3180 9222
rect 3236 9220 3260 9222
rect 3316 9220 3340 9222
rect 3396 9220 3420 9222
rect 3476 9220 3482 9222
rect 3174 9200 3482 9220
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3056 8968 3108 8974
rect 3054 8936 3056 8945
rect 3108 8936 3110 8945
rect 3054 8871 3110 8880
rect 3422 8936 3478 8945
rect 3422 8871 3424 8880
rect 3476 8871 3478 8880
rect 3424 8842 3476 8848
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2792 5630 2912 5658
rect 2504 5568 2556 5574
rect 2504 5510 2556 5516
rect 2332 5234 2452 5250
rect 2320 5228 2452 5234
rect 2372 5222 2452 5228
rect 2320 5170 2372 5176
rect 2226 5128 2282 5137
rect 2226 5063 2282 5072
rect 2240 4622 2268 5063
rect 2228 4616 2280 4622
rect 2228 4558 2280 4564
rect 2136 4140 2188 4146
rect 2136 4082 2188 4088
rect 2228 4140 2280 4146
rect 2228 4082 2280 4088
rect 2240 4026 2268 4082
rect 1872 3998 1992 4026
rect 2044 4004 2096 4010
rect 1492 3936 1544 3942
rect 1490 3904 1492 3913
rect 1584 3936 1636 3942
rect 1544 3904 1546 3913
rect 1584 3878 1636 3884
rect 1490 3839 1546 3848
rect 1490 3496 1546 3505
rect 1490 3431 1546 3440
rect 1504 3398 1532 3431
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 204 3188 256 3194
rect 204 3130 256 3136
rect 216 800 244 3130
rect 664 2984 716 2990
rect 664 2926 716 2932
rect 676 800 704 2926
rect 1124 2916 1176 2922
rect 1124 2858 1176 2864
rect 1136 800 1164 2858
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 1504 2689 1532 2790
rect 1490 2680 1546 2689
rect 1490 2615 1546 2624
rect 1492 2304 1544 2310
rect 1490 2272 1492 2281
rect 1544 2272 1546 2281
rect 1490 2207 1546 2216
rect 1596 1057 1624 3878
rect 1872 3505 1900 3998
rect 2044 3946 2096 3952
rect 2148 3998 2268 4026
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1858 3496 1914 3505
rect 1858 3431 1914 3440
rect 1860 3392 1912 3398
rect 1860 3334 1912 3340
rect 1872 3097 1900 3334
rect 1858 3088 1914 3097
rect 1964 3058 1992 3878
rect 2056 3058 2084 3946
rect 2148 3369 2176 3998
rect 2228 3936 2280 3942
rect 2228 3878 2280 3884
rect 2240 3602 2268 3878
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2134 3360 2190 3369
rect 2134 3295 2190 3304
rect 1858 3023 1914 3032
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 2332 2650 2360 5170
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2424 4593 2452 5102
rect 2410 4584 2466 4593
rect 2410 4519 2466 4528
rect 2412 4480 2464 4486
rect 2412 4422 2464 4428
rect 2424 3058 2452 4422
rect 2516 4321 2544 5510
rect 2596 5160 2648 5166
rect 2596 5102 2648 5108
rect 2502 4312 2558 4321
rect 2502 4247 2558 4256
rect 2504 3936 2556 3942
rect 2504 3878 2556 3884
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2516 2582 2544 3878
rect 2608 3534 2636 5102
rect 2792 5098 2820 5630
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 2780 4616 2832 4622
rect 2884 4604 2912 5510
rect 2976 4690 3004 8230
rect 3068 7546 3096 8366
rect 3174 8188 3482 8208
rect 3174 8186 3180 8188
rect 3236 8186 3260 8188
rect 3316 8186 3340 8188
rect 3396 8186 3420 8188
rect 3476 8186 3482 8188
rect 3236 8134 3238 8186
rect 3418 8134 3420 8186
rect 3174 8132 3180 8134
rect 3236 8132 3260 8134
rect 3316 8132 3340 8134
rect 3396 8132 3420 8134
rect 3476 8132 3482 8134
rect 3174 8112 3482 8132
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3148 7880 3200 7886
rect 3146 7848 3148 7857
rect 3200 7848 3202 7857
rect 3146 7783 3202 7792
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 3146 7440 3202 7449
rect 3146 7375 3148 7384
rect 3200 7375 3202 7384
rect 3148 7346 3200 7352
rect 3344 7342 3372 7890
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3174 7100 3482 7120
rect 3174 7098 3180 7100
rect 3236 7098 3260 7100
rect 3316 7098 3340 7100
rect 3396 7098 3420 7100
rect 3476 7098 3482 7100
rect 3236 7046 3238 7098
rect 3418 7046 3420 7098
rect 3174 7044 3180 7046
rect 3236 7044 3260 7046
rect 3316 7044 3340 7046
rect 3396 7044 3420 7046
rect 3476 7044 3482 7046
rect 3174 7024 3482 7044
rect 3240 6724 3292 6730
rect 3240 6666 3292 6672
rect 3252 6458 3280 6666
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3174 6012 3482 6032
rect 3174 6010 3180 6012
rect 3236 6010 3260 6012
rect 3316 6010 3340 6012
rect 3396 6010 3420 6012
rect 3476 6010 3482 6012
rect 3236 5958 3238 6010
rect 3418 5958 3420 6010
rect 3174 5956 3180 5958
rect 3236 5956 3260 5958
rect 3316 5956 3340 5958
rect 3396 5956 3420 5958
rect 3476 5956 3482 5958
rect 3174 5936 3482 5956
rect 3054 5672 3110 5681
rect 3054 5607 3110 5616
rect 3068 5030 3096 5607
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3252 5370 3280 5510
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 3174 4924 3482 4944
rect 3174 4922 3180 4924
rect 3236 4922 3260 4924
rect 3316 4922 3340 4924
rect 3396 4922 3420 4924
rect 3476 4922 3482 4924
rect 3236 4870 3238 4922
rect 3418 4870 3420 4922
rect 3174 4868 3180 4870
rect 3236 4868 3260 4870
rect 3316 4868 3340 4870
rect 3396 4868 3420 4870
rect 3476 4868 3482 4870
rect 3174 4848 3482 4868
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2832 4576 2912 4604
rect 2780 4558 2832 4564
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 2596 3528 2648 3534
rect 2596 3470 2648 3476
rect 2504 2576 2556 2582
rect 2504 2518 2556 2524
rect 2700 2446 2728 4422
rect 2792 4282 2820 4422
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2792 3641 2820 4082
rect 2976 4078 3004 4422
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2778 3632 2834 3641
rect 2778 3567 2834 3576
rect 2780 3392 2832 3398
rect 2780 3334 2832 3340
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 1676 2304 1728 2310
rect 1676 2246 1728 2252
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2688 2304 2740 2310
rect 2688 2246 2740 2252
rect 1582 1048 1638 1057
rect 1582 983 1638 992
rect 1688 800 1716 2246
rect 2148 800 2176 2246
rect 2700 800 2728 2246
rect 2792 1465 2820 3334
rect 2884 2378 2912 3674
rect 2976 3058 3004 3878
rect 3068 3126 3096 4422
rect 3174 3836 3482 3856
rect 3174 3834 3180 3836
rect 3236 3834 3260 3836
rect 3316 3834 3340 3836
rect 3396 3834 3420 3836
rect 3476 3834 3482 3836
rect 3236 3782 3238 3834
rect 3418 3782 3420 3834
rect 3174 3780 3180 3782
rect 3236 3780 3260 3782
rect 3316 3780 3340 3782
rect 3396 3780 3420 3782
rect 3476 3780 3482 3782
rect 3174 3760 3482 3780
rect 3148 3528 3200 3534
rect 3424 3528 3476 3534
rect 3148 3470 3200 3476
rect 3238 3496 3294 3505
rect 3160 3194 3188 3470
rect 3238 3431 3294 3440
rect 3422 3496 3424 3505
rect 3476 3496 3478 3505
rect 3422 3431 3478 3440
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 3252 3058 3280 3431
rect 2964 3052 3016 3058
rect 2964 2994 3016 3000
rect 3240 3052 3292 3058
rect 3240 2994 3292 3000
rect 3436 2990 3464 3431
rect 3424 2984 3476 2990
rect 3424 2926 3476 2932
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 2976 921 3004 2790
rect 3068 1873 3096 2790
rect 3174 2748 3482 2768
rect 3174 2746 3180 2748
rect 3236 2746 3260 2748
rect 3316 2746 3340 2748
rect 3396 2746 3420 2748
rect 3476 2746 3482 2748
rect 3236 2694 3238 2746
rect 3418 2694 3420 2746
rect 3174 2692 3180 2694
rect 3236 2692 3260 2694
rect 3316 2692 3340 2694
rect 3396 2692 3420 2694
rect 3476 2692 3482 2694
rect 3174 2672 3482 2692
rect 3528 2446 3556 6598
rect 3620 4146 3648 9114
rect 3712 8945 3740 9862
rect 3804 9518 3832 9930
rect 3896 9722 3924 10542
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 3884 9716 3936 9722
rect 3884 9658 3936 9664
rect 3792 9512 3844 9518
rect 3792 9454 3844 9460
rect 3698 8936 3754 8945
rect 3698 8871 3754 8880
rect 3700 8628 3752 8634
rect 3700 8570 3752 8576
rect 3712 5778 3740 8570
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3698 5536 3754 5545
rect 3698 5471 3754 5480
rect 3712 4826 3740 5471
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 3804 4146 3832 9454
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3896 8566 3924 8774
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 3884 8424 3936 8430
rect 3882 8392 3884 8401
rect 3988 8412 4016 10134
rect 4080 8634 4108 11183
rect 4172 10810 4200 11494
rect 4252 11280 4304 11286
rect 4356 11257 4384 12038
rect 4252 11222 4304 11228
rect 4342 11248 4398 11257
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 3936 8392 4016 8412
rect 3938 8384 4016 8392
rect 3882 8327 3938 8336
rect 3896 7478 3924 8327
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 4160 8288 4212 8294
rect 4160 8230 4212 8236
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3896 6390 3924 6734
rect 3884 6384 3936 6390
rect 3884 6326 3936 6332
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3896 4146 3924 5850
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3792 4140 3844 4146
rect 3792 4082 3844 4088
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3790 4040 3846 4049
rect 3790 3975 3792 3984
rect 3844 3975 3846 3984
rect 3792 3946 3844 3952
rect 3896 3738 3924 4082
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3884 3528 3936 3534
rect 3988 3516 4016 7958
rect 4080 7410 4108 8230
rect 4172 7546 4200 8230
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4080 6746 4108 7346
rect 4080 6730 4200 6746
rect 4080 6724 4212 6730
rect 4080 6718 4160 6724
rect 4160 6666 4212 6672
rect 4160 6316 4212 6322
rect 4160 6258 4212 6264
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4080 5846 4108 6054
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 4172 5778 4200 6258
rect 4160 5772 4212 5778
rect 4160 5714 4212 5720
rect 4066 5672 4122 5681
rect 4066 5607 4122 5616
rect 4080 5030 4108 5607
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4080 4826 4108 4966
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4172 4706 4200 5034
rect 3936 3488 4016 3516
rect 4080 4678 4200 4706
rect 3884 3470 3936 3476
rect 4080 3058 4108 4678
rect 4160 4480 4212 4486
rect 4158 4448 4160 4457
rect 4212 4448 4214 4457
rect 4158 4383 4214 4392
rect 4172 4185 4200 4383
rect 4158 4176 4214 4185
rect 4158 4111 4160 4120
rect 4212 4111 4214 4120
rect 4160 4082 4212 4088
rect 4172 4051 4200 4082
rect 4264 3058 4292 11222
rect 4342 11183 4398 11192
rect 4448 10033 4476 12192
rect 4526 12064 4582 12073
rect 4526 11999 4582 12008
rect 4540 10470 4568 11999
rect 4528 10464 4580 10470
rect 4528 10406 4580 10412
rect 4540 10266 4568 10406
rect 4528 10260 4580 10266
rect 4528 10202 4580 10208
rect 4434 10024 4490 10033
rect 4434 9959 4490 9968
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4540 9586 4568 9930
rect 4632 9738 4660 14368
rect 4816 14074 4844 16400
rect 5080 14952 5132 14958
rect 5080 14894 5132 14900
rect 5172 14952 5224 14958
rect 5172 14894 5224 14900
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4804 13932 4856 13938
rect 4804 13874 4856 13880
rect 4816 13841 4844 13874
rect 4802 13832 4858 13841
rect 4802 13767 4858 13776
rect 5092 13734 5120 14894
rect 5184 13938 5212 14894
rect 5460 14618 5488 16400
rect 5540 15224 5592 15230
rect 5540 15166 5592 15172
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5552 14600 5580 15166
rect 5816 14612 5868 14618
rect 5552 14572 5816 14600
rect 5552 14414 5580 14572
rect 5816 14554 5868 14560
rect 5724 14476 5776 14482
rect 5776 14436 5856 14464
rect 5724 14418 5776 14424
rect 5540 14408 5592 14414
rect 5540 14350 5592 14356
rect 5724 14272 5776 14278
rect 5724 14214 5776 14220
rect 5398 14172 5706 14192
rect 5398 14170 5404 14172
rect 5460 14170 5484 14172
rect 5540 14170 5564 14172
rect 5620 14170 5644 14172
rect 5700 14170 5706 14172
rect 5460 14118 5462 14170
rect 5642 14118 5644 14170
rect 5398 14116 5404 14118
rect 5460 14116 5484 14118
rect 5540 14116 5564 14118
rect 5620 14116 5644 14118
rect 5700 14116 5706 14118
rect 5398 14096 5706 14116
rect 5736 14006 5764 14214
rect 5724 14000 5776 14006
rect 5724 13942 5776 13948
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5080 13728 5132 13734
rect 5080 13670 5132 13676
rect 5552 13530 5580 13874
rect 5722 13832 5778 13841
rect 5722 13767 5778 13776
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 4988 12980 5040 12986
rect 4988 12922 5040 12928
rect 5000 12850 5028 12922
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 4712 12708 4764 12714
rect 4712 12650 4764 12656
rect 4724 12374 4752 12650
rect 4804 12640 4856 12646
rect 4804 12582 4856 12588
rect 4712 12368 4764 12374
rect 4712 12310 4764 12316
rect 4724 11762 4752 12310
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4816 10674 4844 12582
rect 4908 12442 4936 12786
rect 5092 12646 5120 13194
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 5184 12986 5212 13126
rect 5172 12980 5224 12986
rect 5172 12922 5224 12928
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 4896 12436 4948 12442
rect 4896 12378 4948 12384
rect 5276 12220 5304 13126
rect 5398 13084 5706 13104
rect 5398 13082 5404 13084
rect 5460 13082 5484 13084
rect 5540 13082 5564 13084
rect 5620 13082 5644 13084
rect 5700 13082 5706 13084
rect 5460 13030 5462 13082
rect 5642 13030 5644 13082
rect 5398 13028 5404 13030
rect 5460 13028 5484 13030
rect 5540 13028 5564 13030
rect 5620 13028 5644 13030
rect 5700 13028 5706 13030
rect 5398 13008 5706 13028
rect 5736 12782 5764 13767
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5356 12232 5408 12238
rect 5276 12192 5356 12220
rect 5356 12174 5408 12180
rect 5398 11996 5706 12016
rect 5398 11994 5404 11996
rect 5460 11994 5484 11996
rect 5540 11994 5564 11996
rect 5620 11994 5644 11996
rect 5700 11994 5706 11996
rect 5460 11942 5462 11994
rect 5642 11942 5644 11994
rect 5398 11940 5404 11942
rect 5460 11940 5484 11942
rect 5540 11940 5564 11942
rect 5620 11940 5644 11942
rect 5700 11940 5706 11942
rect 5398 11920 5706 11940
rect 5828 11257 5856 14436
rect 6012 14414 6040 16510
rect 6090 16400 6146 16510
rect 6734 16538 6790 17200
rect 6734 16510 6868 16538
rect 6734 16400 6790 16510
rect 6644 14884 6696 14890
rect 6644 14826 6696 14832
rect 6000 14408 6052 14414
rect 6184 14408 6236 14414
rect 6000 14350 6052 14356
rect 6104 14368 6184 14396
rect 6012 13870 6040 14350
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 5906 13288 5962 13297
rect 5906 13223 5962 13232
rect 5920 12986 5948 13223
rect 5908 12980 5960 12986
rect 5908 12922 5960 12928
rect 6104 11558 6132 14368
rect 6184 14350 6236 14356
rect 6552 14408 6604 14414
rect 6552 14350 6604 14356
rect 6460 14272 6512 14278
rect 6460 14214 6512 14220
rect 6182 13968 6238 13977
rect 6472 13938 6500 14214
rect 6564 14074 6592 14350
rect 6656 14074 6684 14826
rect 6840 14600 6868 16510
rect 7378 16400 7434 17200
rect 8022 16400 8078 17200
rect 8666 16400 8722 17200
rect 9310 16400 9366 17200
rect 9954 16400 10010 17200
rect 10598 16400 10654 17200
rect 11242 16538 11298 17200
rect 11242 16510 11560 16538
rect 11242 16400 11298 16510
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 6920 14612 6972 14618
rect 6840 14572 6920 14600
rect 6920 14554 6972 14560
rect 7102 14376 7158 14385
rect 7102 14311 7158 14320
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 7010 13968 7066 13977
rect 6182 13903 6184 13912
rect 6236 13903 6238 13912
rect 6276 13932 6328 13938
rect 6184 13874 6236 13880
rect 6276 13874 6328 13880
rect 6460 13932 6512 13938
rect 7010 13903 7012 13912
rect 6460 13874 6512 13880
rect 7064 13903 7066 13912
rect 7012 13874 7064 13880
rect 6288 12434 6316 13874
rect 6736 13796 6788 13802
rect 6736 13738 6788 13744
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 6564 13462 6592 13670
rect 6552 13456 6604 13462
rect 6552 13398 6604 13404
rect 6366 13288 6422 13297
rect 6366 13223 6368 13232
rect 6420 13223 6422 13232
rect 6368 13194 6420 13200
rect 6196 12406 6316 12434
rect 6092 11552 6144 11558
rect 6092 11494 6144 11500
rect 5814 11248 5870 11257
rect 5814 11183 5870 11192
rect 5828 11150 5856 11183
rect 4896 11144 4948 11150
rect 5816 11144 5868 11150
rect 4896 11086 4948 11092
rect 5262 11112 5318 11121
rect 4908 10810 4936 11086
rect 5816 11086 5868 11092
rect 5262 11047 5318 11056
rect 5724 11076 5776 11082
rect 4988 11008 5040 11014
rect 4988 10950 5040 10956
rect 5080 11008 5132 11014
rect 5080 10950 5132 10956
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 5000 10266 5028 10950
rect 5092 10810 5120 10950
rect 5080 10804 5132 10810
rect 5080 10746 5132 10752
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4632 9710 4752 9738
rect 4620 9648 4672 9654
rect 4620 9590 4672 9596
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4540 9178 4568 9522
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4356 7274 4384 8434
rect 4540 8430 4568 8774
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4448 7546 4476 8366
rect 4526 7984 4582 7993
rect 4526 7919 4582 7928
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4344 7268 4396 7274
rect 4344 7210 4396 7216
rect 4344 6792 4396 6798
rect 4540 6780 4568 7919
rect 4344 6734 4396 6740
rect 4448 6752 4568 6780
rect 4356 5302 4384 6734
rect 4448 5302 4476 6752
rect 4526 6352 4582 6361
rect 4526 6287 4528 6296
rect 4580 6287 4582 6296
rect 4528 6258 4580 6264
rect 4540 5642 4568 6258
rect 4632 5658 4660 9590
rect 4724 5846 4752 9710
rect 5170 9616 5226 9625
rect 4988 9580 5040 9586
rect 5170 9551 5172 9560
rect 4988 9522 5040 9528
rect 5224 9551 5226 9560
rect 5172 9522 5224 9528
rect 4804 9376 4856 9382
rect 4804 9318 4856 9324
rect 4712 5840 4764 5846
rect 4712 5782 4764 5788
rect 4528 5636 4580 5642
rect 4632 5630 4752 5658
rect 4528 5578 4580 5584
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 4436 5296 4488 5302
rect 4436 5238 4488 5244
rect 4448 4826 4476 5238
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4540 4282 4568 4966
rect 4528 4276 4580 4282
rect 4528 4218 4580 4224
rect 4632 4010 4660 5510
rect 4724 4622 4752 5630
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4724 4214 4752 4558
rect 4712 4208 4764 4214
rect 4712 4150 4764 4156
rect 4620 4004 4672 4010
rect 4620 3946 4672 3952
rect 4618 3496 4674 3505
rect 4618 3431 4674 3440
rect 4712 3460 4764 3466
rect 4632 3194 4660 3431
rect 4712 3402 4764 3408
rect 4620 3188 4672 3194
rect 4620 3130 4672 3136
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 3976 2848 4028 2854
rect 3976 2790 4028 2796
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 3884 2576 3936 2582
rect 3884 2518 3936 2524
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 3054 1864 3110 1873
rect 3054 1799 3110 1808
rect 2962 912 3018 921
rect 2962 847 3018 856
rect 3160 800 3188 2246
rect 3620 800 3648 2246
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1674 0 1730 800
rect 2134 0 2190 800
rect 2686 0 2742 800
rect 3146 0 3202 800
rect 3606 0 3662 800
rect 3896 241 3924 2518
rect 3988 2514 4016 2790
rect 3976 2508 4028 2514
rect 3976 2450 4028 2456
rect 4264 2446 4292 2790
rect 4632 2514 4660 2790
rect 4724 2650 4752 3402
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4620 2508 4672 2514
rect 4620 2450 4672 2456
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4172 800 4200 2246
rect 4632 800 4660 2450
rect 4816 2446 4844 9318
rect 4896 8900 4948 8906
rect 4896 8842 4948 8848
rect 4908 7342 4936 8842
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4908 4826 4936 5510
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 5000 4690 5028 9522
rect 5276 8634 5304 11047
rect 5724 11018 5776 11024
rect 5398 10908 5706 10928
rect 5398 10906 5404 10908
rect 5460 10906 5484 10908
rect 5540 10906 5564 10908
rect 5620 10906 5644 10908
rect 5700 10906 5706 10908
rect 5460 10854 5462 10906
rect 5642 10854 5644 10906
rect 5398 10852 5404 10854
rect 5460 10852 5484 10854
rect 5540 10852 5564 10854
rect 5620 10852 5644 10854
rect 5700 10852 5706 10854
rect 5398 10832 5706 10852
rect 5448 10600 5500 10606
rect 5448 10542 5500 10548
rect 5460 10130 5488 10542
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5398 9820 5706 9840
rect 5398 9818 5404 9820
rect 5460 9818 5484 9820
rect 5540 9818 5564 9820
rect 5620 9818 5644 9820
rect 5700 9818 5706 9820
rect 5460 9766 5462 9818
rect 5642 9766 5644 9818
rect 5398 9764 5404 9766
rect 5460 9764 5484 9766
rect 5540 9764 5564 9766
rect 5620 9764 5644 9766
rect 5700 9764 5706 9766
rect 5398 9744 5706 9764
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5368 9178 5396 9454
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5460 9042 5488 9590
rect 5736 9081 5764 11018
rect 5906 10704 5962 10713
rect 5906 10639 5908 10648
rect 5960 10639 5962 10648
rect 5908 10610 5960 10616
rect 5920 10470 5948 10610
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5828 10062 5856 10406
rect 5816 10056 5868 10062
rect 5816 9998 5868 10004
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5828 9518 5856 9658
rect 6012 9568 6040 9998
rect 6092 9920 6144 9926
rect 6092 9862 6144 9868
rect 6104 9722 6132 9862
rect 6092 9716 6144 9722
rect 6092 9658 6144 9664
rect 6012 9540 6132 9568
rect 5816 9512 5868 9518
rect 5816 9454 5868 9460
rect 5722 9072 5778 9081
rect 5448 9036 5500 9042
rect 5722 9007 5778 9016
rect 5448 8978 5500 8984
rect 5398 8732 5706 8752
rect 5398 8730 5404 8732
rect 5460 8730 5484 8732
rect 5540 8730 5564 8732
rect 5620 8730 5644 8732
rect 5700 8730 5706 8732
rect 5460 8678 5462 8730
rect 5642 8678 5644 8730
rect 5398 8676 5404 8678
rect 5460 8676 5484 8678
rect 5540 8676 5564 8678
rect 5620 8676 5644 8678
rect 5700 8676 5706 8678
rect 5398 8656 5706 8676
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5276 8537 5304 8570
rect 5540 8560 5592 8566
rect 5078 8528 5134 8537
rect 5262 8528 5318 8537
rect 5078 8463 5134 8472
rect 5172 8492 5224 8498
rect 5092 8362 5120 8463
rect 5540 8502 5592 8508
rect 5262 8463 5318 8472
rect 5172 8434 5224 8440
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 5092 7546 5120 7686
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5184 7426 5212 8434
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5276 7954 5304 8298
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5092 7398 5212 7426
rect 4988 4684 5040 4690
rect 4988 4626 5040 4632
rect 4894 4584 4950 4593
rect 4894 4519 4950 4528
rect 4908 3194 4936 4519
rect 5092 3369 5120 7398
rect 5276 7274 5304 7890
rect 5552 7818 5580 8502
rect 5828 7886 5856 9454
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 6012 9110 6040 9386
rect 6000 9104 6052 9110
rect 6000 9046 6052 9052
rect 6012 8838 6040 9046
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 6012 8634 6040 8774
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5908 8560 5960 8566
rect 5908 8502 5960 8508
rect 5920 8090 5948 8502
rect 6104 8294 6132 9540
rect 6092 8288 6144 8294
rect 6092 8230 6144 8236
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5398 7644 5706 7664
rect 5398 7642 5404 7644
rect 5460 7642 5484 7644
rect 5540 7642 5564 7644
rect 5620 7642 5644 7644
rect 5700 7642 5706 7644
rect 5460 7590 5462 7642
rect 5642 7590 5644 7642
rect 5398 7588 5404 7590
rect 5460 7588 5484 7590
rect 5540 7588 5564 7590
rect 5620 7588 5644 7590
rect 5700 7588 5706 7590
rect 5398 7568 5706 7588
rect 5264 7268 5316 7274
rect 5264 7210 5316 7216
rect 5276 7002 5304 7210
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5736 6798 5764 7686
rect 5920 7546 5948 8026
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5920 6934 5948 7346
rect 5908 6928 5960 6934
rect 5908 6870 5960 6876
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5398 6556 5706 6576
rect 5398 6554 5404 6556
rect 5460 6554 5484 6556
rect 5540 6554 5564 6556
rect 5620 6554 5644 6556
rect 5700 6554 5706 6556
rect 5460 6502 5462 6554
rect 5642 6502 5644 6554
rect 5398 6500 5404 6502
rect 5460 6500 5484 6502
rect 5540 6500 5564 6502
rect 5620 6500 5644 6502
rect 5700 6500 5706 6502
rect 5398 6480 5706 6500
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5552 5846 5580 6326
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5828 6118 5856 6258
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5816 6112 5868 6118
rect 5816 6054 5868 6060
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5398 5468 5706 5488
rect 5398 5466 5404 5468
rect 5460 5466 5484 5468
rect 5540 5466 5564 5468
rect 5620 5466 5644 5468
rect 5700 5466 5706 5468
rect 5460 5414 5462 5466
rect 5642 5414 5644 5466
rect 5398 5412 5404 5414
rect 5460 5412 5484 5414
rect 5540 5412 5564 5414
rect 5620 5412 5644 5414
rect 5700 5412 5706 5414
rect 5398 5392 5706 5412
rect 5736 5234 5764 6054
rect 5828 5778 5856 6054
rect 5816 5772 5868 5778
rect 5816 5714 5868 5720
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 5264 5160 5316 5166
rect 5264 5102 5316 5108
rect 5172 5092 5224 5098
rect 5172 5034 5224 5040
rect 5184 4282 5212 5034
rect 5276 4690 5304 5102
rect 5264 4684 5316 4690
rect 5264 4626 5316 4632
rect 5276 4554 5304 4626
rect 5264 4548 5316 4554
rect 5264 4490 5316 4496
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5276 4060 5304 4490
rect 5828 4486 5856 5714
rect 5920 5681 5948 6870
rect 5906 5672 5962 5681
rect 5906 5607 5962 5616
rect 6012 5302 6040 8026
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6104 5846 6132 6190
rect 6092 5840 6144 5846
rect 6092 5782 6144 5788
rect 6104 5574 6132 5782
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6104 5302 6132 5510
rect 6000 5296 6052 5302
rect 6000 5238 6052 5244
rect 6092 5296 6144 5302
rect 6092 5238 6144 5244
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5398 4380 5706 4400
rect 5398 4378 5404 4380
rect 5460 4378 5484 4380
rect 5540 4378 5564 4380
rect 5620 4378 5644 4380
rect 5700 4378 5706 4380
rect 5460 4326 5462 4378
rect 5642 4326 5644 4378
rect 5398 4324 5404 4326
rect 5460 4324 5484 4326
rect 5540 4324 5564 4326
rect 5620 4324 5644 4326
rect 5700 4324 5706 4326
rect 5398 4304 5706 4324
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5356 4072 5408 4078
rect 5276 4032 5356 4060
rect 5356 4014 5408 4020
rect 5368 3738 5396 4014
rect 5552 3942 5580 4150
rect 5828 4078 5856 4422
rect 6012 4282 6040 5238
rect 6104 4622 6132 5238
rect 6092 4616 6144 4622
rect 6092 4558 6144 4564
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 6104 4146 6132 4558
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5908 3936 5960 3942
rect 5908 3878 5960 3884
rect 5356 3732 5408 3738
rect 5356 3674 5408 3680
rect 5920 3641 5948 3878
rect 5906 3632 5962 3641
rect 5906 3567 5962 3576
rect 6104 3534 6132 4082
rect 6092 3528 6144 3534
rect 6092 3470 6144 3476
rect 5172 3392 5224 3398
rect 5078 3360 5134 3369
rect 5172 3334 5224 3340
rect 5262 3360 5318 3369
rect 5078 3295 5134 3304
rect 4896 3188 4948 3194
rect 4896 3130 4948 3136
rect 5184 2446 5212 3334
rect 5262 3295 5318 3304
rect 5276 3194 5304 3295
rect 5398 3292 5706 3312
rect 5398 3290 5404 3292
rect 5460 3290 5484 3292
rect 5540 3290 5564 3292
rect 5620 3290 5644 3292
rect 5700 3290 5706 3292
rect 5460 3238 5462 3290
rect 5642 3238 5644 3290
rect 5398 3236 5404 3238
rect 5460 3236 5484 3238
rect 5540 3236 5564 3238
rect 5620 3236 5644 3238
rect 5700 3236 5706 3238
rect 5398 3216 5706 3236
rect 5264 3188 5316 3194
rect 5264 3130 5316 3136
rect 5908 2984 5960 2990
rect 5906 2952 5908 2961
rect 5960 2952 5962 2961
rect 5906 2887 5962 2896
rect 5724 2848 5776 2854
rect 5724 2790 5776 2796
rect 5736 2446 5764 2790
rect 6196 2774 6224 12406
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6472 11830 6500 12038
rect 6460 11824 6512 11830
rect 6460 11766 6512 11772
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6380 11150 6408 11698
rect 6368 11144 6420 11150
rect 6368 11086 6420 11092
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6288 10810 6316 10950
rect 6276 10804 6328 10810
rect 6276 10746 6328 10752
rect 6380 10674 6408 11086
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 6288 9450 6316 10066
rect 6276 9444 6328 9450
rect 6276 9386 6328 9392
rect 6472 9382 6500 11766
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6460 9376 6512 9382
rect 6460 9318 6512 9324
rect 6472 8430 6500 9318
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 6288 4010 6316 7754
rect 6368 6112 6420 6118
rect 6368 6054 6420 6060
rect 6380 5370 6408 6054
rect 6368 5364 6420 5370
rect 6368 5306 6420 5312
rect 6276 4004 6328 4010
rect 6276 3946 6328 3952
rect 6472 2961 6500 8230
rect 6564 5574 6592 9590
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6564 5137 6592 5306
rect 6550 5128 6606 5137
rect 6550 5063 6606 5072
rect 6564 4146 6592 5063
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6458 2952 6514 2961
rect 6458 2887 6514 2896
rect 5920 2746 6224 2774
rect 5920 2650 5948 2746
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 6656 2446 6684 13670
rect 6748 11286 6776 13738
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 6828 11076 6880 11082
rect 6828 11018 6880 11024
rect 6840 10792 6868 11018
rect 6748 10764 6868 10792
rect 6748 10606 6776 10764
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6736 10600 6788 10606
rect 6736 10542 6788 10548
rect 6748 10198 6776 10542
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6748 10062 6776 10134
rect 6840 10062 6868 10610
rect 6736 10056 6788 10062
rect 6736 9998 6788 10004
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6748 9382 6776 9454
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6840 9081 6868 9522
rect 6826 9072 6882 9081
rect 6826 9007 6882 9016
rect 6734 8800 6790 8809
rect 6734 8735 6790 8744
rect 6748 8634 6776 8735
rect 6826 8664 6882 8673
rect 6736 8628 6788 8634
rect 6826 8599 6882 8608
rect 6736 8570 6788 8576
rect 6748 6934 6776 8570
rect 6840 8566 6868 8599
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6840 7206 6868 8298
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6932 6866 6960 12174
rect 7012 11824 7064 11830
rect 7012 11766 7064 11772
rect 7024 9654 7052 11766
rect 7116 10588 7144 14311
rect 7196 14272 7248 14278
rect 7196 14214 7248 14220
rect 7208 12434 7236 14214
rect 7300 13954 7328 14962
rect 7392 14618 7420 16400
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7484 14618 7512 14758
rect 7622 14716 7930 14736
rect 7622 14714 7628 14716
rect 7684 14714 7708 14716
rect 7764 14714 7788 14716
rect 7844 14714 7868 14716
rect 7924 14714 7930 14716
rect 7684 14662 7686 14714
rect 7866 14662 7868 14714
rect 7622 14660 7628 14662
rect 7684 14660 7708 14662
rect 7764 14660 7788 14662
rect 7844 14660 7868 14662
rect 7924 14660 7930 14662
rect 7622 14640 7930 14660
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7392 14414 7420 14554
rect 7380 14408 7432 14414
rect 7380 14350 7432 14356
rect 7300 13938 7420 13954
rect 7300 13932 7432 13938
rect 7300 13926 7380 13932
rect 7380 13874 7432 13880
rect 7622 13628 7930 13648
rect 7622 13626 7628 13628
rect 7684 13626 7708 13628
rect 7764 13626 7788 13628
rect 7844 13626 7868 13628
rect 7924 13626 7930 13628
rect 7684 13574 7686 13626
rect 7866 13574 7868 13626
rect 7622 13572 7628 13574
rect 7684 13572 7708 13574
rect 7764 13572 7788 13574
rect 7844 13572 7868 13574
rect 7924 13572 7930 13574
rect 7622 13552 7930 13572
rect 7622 12540 7930 12560
rect 7622 12538 7628 12540
rect 7684 12538 7708 12540
rect 7764 12538 7788 12540
rect 7844 12538 7868 12540
rect 7924 12538 7930 12540
rect 7684 12486 7686 12538
rect 7866 12486 7868 12538
rect 7622 12484 7628 12486
rect 7684 12484 7708 12486
rect 7764 12484 7788 12486
rect 7844 12484 7868 12486
rect 7924 12484 7930 12486
rect 7622 12464 7930 12484
rect 7208 12406 7420 12434
rect 7288 11008 7340 11014
rect 7288 10950 7340 10956
rect 7300 10742 7328 10950
rect 7288 10736 7340 10742
rect 7288 10678 7340 10684
rect 7116 10560 7328 10588
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7012 9648 7064 9654
rect 7012 9590 7064 9596
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7024 7886 7052 8570
rect 7116 8430 7144 8842
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 7012 7880 7064 7886
rect 7012 7822 7064 7828
rect 7012 7472 7064 7478
rect 7012 7414 7064 7420
rect 6920 6860 6972 6866
rect 6920 6802 6972 6808
rect 6920 6724 6972 6730
rect 6920 6666 6972 6672
rect 6932 6390 6960 6666
rect 7024 6458 7052 7414
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6920 6384 6972 6390
rect 6920 6326 6972 6332
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 6840 5642 6868 5782
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6748 4298 6776 5510
rect 6932 4622 6960 6054
rect 7116 5710 7144 8366
rect 7208 8362 7236 9862
rect 7196 8356 7248 8362
rect 7196 8298 7248 8304
rect 7300 8072 7328 10560
rect 7208 8044 7328 8072
rect 7208 6866 7236 8044
rect 7288 7948 7340 7954
rect 7288 7890 7340 7896
rect 7300 7546 7328 7890
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7300 6934 7328 7482
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 7196 6860 7248 6866
rect 7196 6802 7248 6808
rect 7208 5760 7236 6802
rect 7392 6798 7420 12406
rect 7472 11552 7524 11558
rect 7472 11494 7524 11500
rect 7484 11082 7512 11494
rect 7622 11452 7930 11472
rect 7622 11450 7628 11452
rect 7684 11450 7708 11452
rect 7764 11450 7788 11452
rect 7844 11450 7868 11452
rect 7924 11450 7930 11452
rect 7684 11398 7686 11450
rect 7866 11398 7868 11450
rect 7622 11396 7628 11398
rect 7684 11396 7708 11398
rect 7764 11396 7788 11398
rect 7844 11396 7868 11398
rect 7924 11396 7930 11398
rect 7622 11376 7930 11396
rect 7472 11076 7524 11082
rect 7472 11018 7524 11024
rect 7622 10364 7930 10384
rect 7622 10362 7628 10364
rect 7684 10362 7708 10364
rect 7764 10362 7788 10364
rect 7844 10362 7868 10364
rect 7924 10362 7930 10364
rect 7684 10310 7686 10362
rect 7866 10310 7868 10362
rect 7622 10308 7628 10310
rect 7684 10308 7708 10310
rect 7764 10308 7788 10310
rect 7844 10308 7868 10310
rect 7924 10308 7930 10310
rect 7622 10288 7930 10308
rect 7622 9276 7930 9296
rect 7622 9274 7628 9276
rect 7684 9274 7708 9276
rect 7764 9274 7788 9276
rect 7844 9274 7868 9276
rect 7924 9274 7930 9276
rect 7684 9222 7686 9274
rect 7866 9222 7868 9274
rect 7622 9220 7628 9222
rect 7684 9220 7708 9222
rect 7764 9220 7788 9222
rect 7844 9220 7868 9222
rect 7924 9220 7930 9222
rect 7622 9200 7930 9220
rect 8036 8974 8064 16400
rect 8116 14816 8168 14822
rect 8116 14758 8168 14764
rect 8128 13802 8156 14758
rect 8680 14618 8708 16400
rect 9128 14884 9180 14890
rect 9128 14826 9180 14832
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8208 14544 8260 14550
rect 8206 14512 8208 14521
rect 8260 14512 8262 14521
rect 8206 14447 8262 14456
rect 8680 14414 8708 14554
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8208 13932 8260 13938
rect 8208 13874 8260 13880
rect 8116 13796 8168 13802
rect 8116 13738 8168 13744
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 8128 10062 8156 11494
rect 8220 10470 8248 13874
rect 8576 12164 8628 12170
rect 8576 12106 8628 12112
rect 8300 11892 8352 11898
rect 8300 11834 8352 11840
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8024 8968 8076 8974
rect 8024 8910 8076 8916
rect 7564 8900 7616 8906
rect 7564 8842 7616 8848
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 7954 7512 8774
rect 7576 8634 7604 8842
rect 8206 8800 8262 8809
rect 8206 8735 8262 8744
rect 8114 8664 8170 8673
rect 7564 8628 7616 8634
rect 8114 8599 8116 8608
rect 7564 8570 7616 8576
rect 8168 8599 8170 8608
rect 8116 8570 8168 8576
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7668 8294 7696 8502
rect 8024 8492 8076 8498
rect 8116 8492 8168 8498
rect 8076 8452 8116 8480
rect 8024 8434 8076 8440
rect 8116 8434 8168 8440
rect 8220 8294 8248 8735
rect 8312 8673 8340 11834
rect 8392 11756 8444 11762
rect 8392 11698 8444 11704
rect 8404 11354 8432 11698
rect 8482 11520 8538 11529
rect 8482 11455 8538 11464
rect 8392 11348 8444 11354
rect 8392 11290 8444 11296
rect 8404 10810 8432 11290
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8496 10674 8524 11455
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8588 10418 8616 12106
rect 8404 10390 8616 10418
rect 8298 8664 8354 8673
rect 8298 8599 8354 8608
rect 8312 8566 8340 8599
rect 8300 8560 8352 8566
rect 8404 8548 8432 10390
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8484 10192 8536 10198
rect 8484 10134 8536 10140
rect 8496 9178 8524 10134
rect 8588 9178 8616 10202
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8680 9654 8708 9862
rect 8668 9648 8720 9654
rect 8668 9590 8720 9596
rect 8668 9376 8720 9382
rect 8668 9318 8720 9324
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8680 9058 8708 9318
rect 8588 9042 8708 9058
rect 8576 9036 8708 9042
rect 8628 9030 8708 9036
rect 8576 8978 8628 8984
rect 8484 8560 8536 8566
rect 8404 8520 8484 8548
rect 8300 8502 8352 8508
rect 8484 8502 8536 8508
rect 7668 8276 7972 8294
rect 8116 8288 8168 8294
rect 7668 8266 8064 8276
rect 7944 8248 8064 8266
rect 7622 8188 7930 8208
rect 7622 8186 7628 8188
rect 7684 8186 7708 8188
rect 7764 8186 7788 8188
rect 7844 8186 7868 8188
rect 7924 8186 7930 8188
rect 7684 8134 7686 8186
rect 7866 8134 7868 8186
rect 7622 8132 7628 8134
rect 7684 8132 7708 8134
rect 7764 8132 7788 8134
rect 7844 8132 7868 8134
rect 7924 8132 7930 8134
rect 7622 8112 7930 8132
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 8036 7886 8064 8248
rect 8116 8230 8168 8236
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8128 8106 8156 8230
rect 8312 8106 8340 8502
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8484 8424 8536 8430
rect 8588 8412 8616 8978
rect 8772 8974 8800 9318
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8760 8832 8812 8838
rect 8758 8800 8760 8809
rect 8812 8800 8814 8809
rect 8758 8735 8814 8744
rect 8536 8384 8616 8412
rect 8484 8366 8536 8372
rect 8128 8078 8340 8106
rect 8404 8022 8432 8366
rect 8392 8016 8444 8022
rect 8206 7984 8262 7993
rect 8392 7958 8444 7964
rect 8206 7919 8262 7928
rect 8220 7886 8248 7919
rect 8024 7880 8076 7886
rect 8024 7822 8076 7828
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 7622 7100 7930 7120
rect 7622 7098 7628 7100
rect 7684 7098 7708 7100
rect 7764 7098 7788 7100
rect 7844 7098 7868 7100
rect 7924 7098 7930 7100
rect 7684 7046 7686 7098
rect 7866 7046 7868 7098
rect 7622 7044 7628 7046
rect 7684 7044 7708 7046
rect 7764 7044 7788 7046
rect 7844 7044 7868 7046
rect 7924 7044 7930 7046
rect 7622 7024 7930 7044
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7380 6792 7432 6798
rect 7668 6769 7696 6802
rect 7380 6734 7432 6740
rect 7654 6760 7710 6769
rect 7208 5732 7328 5760
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7116 5030 7144 5510
rect 7194 5264 7250 5273
rect 7194 5199 7250 5208
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 6920 4616 6972 4622
rect 6920 4558 6972 4564
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 6748 4270 6868 4298
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6748 3738 6776 4082
rect 6840 3942 6868 4270
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6932 3466 6960 4422
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6932 3058 6960 3402
rect 6920 3052 6972 3058
rect 6920 2994 6972 3000
rect 6736 2916 6788 2922
rect 6736 2858 6788 2864
rect 6748 2446 6776 2858
rect 6920 2848 6972 2854
rect 7024 2836 7052 3538
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7116 2854 7144 3470
rect 7208 3398 7236 5199
rect 7300 4758 7328 5732
rect 7288 4752 7340 4758
rect 7288 4694 7340 4700
rect 7288 4616 7340 4622
rect 7392 4604 7420 6734
rect 7654 6695 7710 6704
rect 7668 6458 7696 6695
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 8024 6656 8076 6662
rect 8024 6598 8076 6604
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7484 6225 7512 6394
rect 7746 6352 7802 6361
rect 7746 6287 7802 6296
rect 7470 6216 7526 6225
rect 7760 6186 7788 6287
rect 7470 6151 7526 6160
rect 7748 6180 7800 6186
rect 7484 5794 7512 6151
rect 7748 6122 7800 6128
rect 7944 6100 7972 6598
rect 8036 6458 8064 6598
rect 8024 6452 8076 6458
rect 8024 6394 8076 6400
rect 7944 6072 8064 6100
rect 7622 6012 7930 6032
rect 7622 6010 7628 6012
rect 7684 6010 7708 6012
rect 7764 6010 7788 6012
rect 7844 6010 7868 6012
rect 7924 6010 7930 6012
rect 7684 5958 7686 6010
rect 7866 5958 7868 6010
rect 7622 5956 7628 5958
rect 7684 5956 7708 5958
rect 7764 5956 7788 5958
rect 7844 5956 7868 5958
rect 7924 5956 7930 5958
rect 7622 5936 7930 5956
rect 7484 5766 7604 5794
rect 7472 5704 7524 5710
rect 7472 5646 7524 5652
rect 7484 5030 7512 5646
rect 7576 5098 7604 5766
rect 7656 5636 7708 5642
rect 7656 5578 7708 5584
rect 7668 5273 7696 5578
rect 7654 5264 7710 5273
rect 7654 5199 7710 5208
rect 7564 5092 7616 5098
rect 7564 5034 7616 5040
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7340 4576 7420 4604
rect 7288 4558 7340 4564
rect 7392 4214 7420 4576
rect 7380 4208 7432 4214
rect 7286 4176 7342 4185
rect 7380 4150 7432 4156
rect 7286 4111 7342 4120
rect 7300 3505 7328 4111
rect 7286 3496 7342 3505
rect 7286 3431 7342 3440
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 6972 2808 7052 2836
rect 7104 2848 7156 2854
rect 6920 2790 6972 2796
rect 7104 2790 7156 2796
rect 7208 2446 7236 3130
rect 7300 3040 7328 3431
rect 7300 3012 7420 3040
rect 7392 2922 7420 3012
rect 7288 2916 7340 2922
rect 7288 2858 7340 2864
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7300 2446 7328 2858
rect 7484 2854 7512 4966
rect 7622 4924 7930 4944
rect 7622 4922 7628 4924
rect 7684 4922 7708 4924
rect 7764 4922 7788 4924
rect 7844 4922 7868 4924
rect 7924 4922 7930 4924
rect 7684 4870 7686 4922
rect 7866 4870 7868 4922
rect 7622 4868 7628 4870
rect 7684 4868 7708 4870
rect 7764 4868 7788 4870
rect 7844 4868 7868 4870
rect 7924 4868 7930 4870
rect 7622 4848 7930 4868
rect 8036 4128 8064 6072
rect 8128 5234 8156 7346
rect 8404 7002 8432 7686
rect 8496 7478 8524 8366
rect 8760 8084 8812 8090
rect 8760 8026 8812 8032
rect 8772 7886 8800 8026
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8484 7472 8536 7478
rect 8484 7414 8536 7420
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8206 6352 8262 6361
rect 8312 6322 8340 6938
rect 8496 6866 8524 7414
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8496 6390 8524 6802
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8206 6287 8262 6296
rect 8300 6316 8352 6322
rect 8220 5574 8248 6287
rect 8300 6258 8352 6264
rect 8772 6186 8800 6598
rect 8760 6180 8812 6186
rect 8760 6122 8812 6128
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 8220 5370 8248 5510
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 8404 5234 8432 6054
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8116 5228 8168 5234
rect 8116 5170 8168 5176
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8128 4622 8156 5170
rect 8496 4826 8524 5238
rect 8484 4820 8536 4826
rect 8484 4762 8536 4768
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8588 4146 8616 4490
rect 8576 4140 8628 4146
rect 8036 4100 8248 4128
rect 8024 4004 8076 4010
rect 8024 3946 8076 3952
rect 7622 3836 7930 3856
rect 7622 3834 7628 3836
rect 7684 3834 7708 3836
rect 7764 3834 7788 3836
rect 7844 3834 7868 3836
rect 7924 3834 7930 3836
rect 7684 3782 7686 3834
rect 7866 3782 7868 3834
rect 7622 3780 7628 3782
rect 7684 3780 7708 3782
rect 7764 3780 7788 3782
rect 7844 3780 7868 3782
rect 7924 3780 7930 3782
rect 7622 3760 7930 3780
rect 8036 3738 8064 3946
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 8024 3596 8076 3602
rect 8220 3584 8248 4100
rect 8576 4082 8628 4088
rect 8864 3602 8892 14214
rect 9140 13870 9168 14826
rect 9324 14618 9352 16400
rect 9968 14618 9996 16400
rect 10612 14618 10640 16400
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 9324 14414 9352 14554
rect 9968 14414 9996 14554
rect 10612 14414 10640 14554
rect 11532 14414 11560 16510
rect 11886 16400 11942 17200
rect 12530 16400 12586 17200
rect 13174 16400 13230 17200
rect 13818 16400 13874 17200
rect 14462 16538 14518 17200
rect 14462 16510 14780 16538
rect 14462 16400 14518 16510
rect 11900 14618 11928 16400
rect 12070 14716 12378 14736
rect 12070 14714 12076 14716
rect 12132 14714 12156 14716
rect 12212 14714 12236 14716
rect 12292 14714 12316 14716
rect 12372 14714 12378 14716
rect 12132 14662 12134 14714
rect 12314 14662 12316 14714
rect 12070 14660 12076 14662
rect 12132 14660 12156 14662
rect 12212 14660 12236 14662
rect 12292 14660 12316 14662
rect 12372 14660 12378 14662
rect 12070 14640 12378 14660
rect 12544 14618 12572 16400
rect 13188 14618 13216 16400
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 12532 14612 12584 14618
rect 12532 14554 12584 14560
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 12348 14544 12400 14550
rect 12348 14486 12400 14492
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9956 14408 10008 14414
rect 9956 14350 10008 14356
rect 10600 14408 10652 14414
rect 10600 14350 10652 14356
rect 11520 14408 11572 14414
rect 11520 14350 11572 14356
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10876 14272 10928 14278
rect 11888 14272 11940 14278
rect 10876 14214 10928 14220
rect 11808 14232 11888 14260
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9140 12434 9168 13806
rect 9324 12434 9352 14010
rect 9140 12406 9260 12434
rect 9324 12406 9444 12434
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9048 10674 9076 10950
rect 9036 10668 9088 10674
rect 9036 10610 9088 10616
rect 9048 10130 9076 10610
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 8944 9512 8996 9518
rect 8944 9454 8996 9460
rect 8956 8090 8984 9454
rect 9126 9072 9182 9081
rect 9126 9007 9182 9016
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 8956 6730 8984 6870
rect 8944 6724 8996 6730
rect 8944 6666 8996 6672
rect 8944 6384 8996 6390
rect 8944 6326 8996 6332
rect 8956 6254 8984 6326
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8956 5778 8984 6190
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 9140 5545 9168 9007
rect 9126 5536 9182 5545
rect 9126 5471 9182 5480
rect 8944 5228 8996 5234
rect 8944 5170 8996 5176
rect 8956 4826 8984 5170
rect 9036 5024 9088 5030
rect 9036 4966 9088 4972
rect 8944 4820 8996 4826
rect 8944 4762 8996 4768
rect 8076 3556 8248 3584
rect 8024 3538 8076 3544
rect 8220 3516 8248 3556
rect 8852 3596 8904 3602
rect 8852 3538 8904 3544
rect 8300 3528 8352 3534
rect 8220 3488 8300 3516
rect 8300 3470 8352 3476
rect 7932 3460 7984 3466
rect 7932 3402 7984 3408
rect 7944 2990 7972 3402
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 7932 2984 7984 2990
rect 7932 2926 7984 2932
rect 8208 2916 8260 2922
rect 8208 2858 8260 2864
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 7622 2748 7930 2768
rect 7622 2746 7628 2748
rect 7684 2746 7708 2748
rect 7764 2746 7788 2748
rect 7844 2746 7868 2748
rect 7924 2746 7930 2748
rect 7684 2694 7686 2746
rect 7866 2694 7868 2746
rect 7622 2692 7628 2694
rect 7684 2692 7708 2694
rect 7764 2692 7788 2694
rect 7844 2692 7868 2694
rect 7924 2692 7930 2694
rect 7622 2672 7930 2692
rect 8220 2514 8248 2858
rect 8208 2508 8260 2514
rect 8208 2450 8260 2456
rect 8404 2446 8432 3334
rect 9048 3058 9076 4966
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9140 3942 9168 4558
rect 9128 3936 9180 3942
rect 9128 3878 9180 3884
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 9232 2990 9260 12406
rect 9312 8832 9364 8838
rect 9310 8800 9312 8809
rect 9364 8800 9366 8809
rect 9310 8735 9366 8744
rect 9416 6730 9444 12406
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9508 8906 9536 9114
rect 9600 9042 9628 9590
rect 9692 9450 9720 9930
rect 9680 9444 9732 9450
rect 9680 9386 9732 9392
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9496 8900 9548 8906
rect 9496 8842 9548 8848
rect 9494 8664 9550 8673
rect 9494 8599 9550 8608
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 6458 9352 6598
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9404 4276 9456 4282
rect 9404 4218 9456 4224
rect 9416 3126 9444 4218
rect 9508 4128 9536 8599
rect 9600 7954 9628 8978
rect 9784 8616 9812 14214
rect 9846 14172 10154 14192
rect 9846 14170 9852 14172
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 10148 14170 10154 14172
rect 9908 14118 9910 14170
rect 10090 14118 10092 14170
rect 9846 14116 9852 14118
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 10148 14116 10154 14118
rect 9846 14096 10154 14116
rect 9846 13084 10154 13104
rect 9846 13082 9852 13084
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 10148 13082 10154 13084
rect 9908 13030 9910 13082
rect 10090 13030 10092 13082
rect 9846 13028 9852 13030
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 10148 13028 10154 13030
rect 9846 13008 10154 13028
rect 10704 12434 10732 14214
rect 10612 12406 10732 12434
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 9846 11996 10154 12016
rect 9846 11994 9852 11996
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 10148 11994 10154 11996
rect 9908 11942 9910 11994
rect 10090 11942 10092 11994
rect 9846 11940 9852 11942
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 10148 11940 10154 11942
rect 9846 11920 10154 11940
rect 10244 11558 10272 12038
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 9846 10908 10154 10928
rect 9846 10906 9852 10908
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 10148 10906 10154 10908
rect 9908 10854 9910 10906
rect 10090 10854 10092 10906
rect 9846 10852 9852 10854
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 10148 10852 10154 10854
rect 9846 10832 10154 10852
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 10062 9996 10406
rect 9956 10056 10008 10062
rect 9956 9998 10008 10004
rect 10244 9994 10272 11494
rect 10414 11112 10470 11121
rect 10414 11047 10470 11056
rect 10324 10532 10376 10538
rect 10324 10474 10376 10480
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 9846 9820 10154 9840
rect 9846 9818 9852 9820
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 10148 9818 10154 9820
rect 9908 9766 9910 9818
rect 10090 9766 10092 9818
rect 9846 9764 9852 9766
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 10148 9764 10154 9766
rect 9846 9744 10154 9764
rect 10244 9654 10272 9930
rect 10232 9648 10284 9654
rect 10232 9590 10284 9596
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10244 8838 10272 9318
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 9846 8732 10154 8752
rect 9846 8730 9852 8732
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 10148 8730 10154 8732
rect 9908 8678 9910 8730
rect 10090 8678 10092 8730
rect 9846 8676 9852 8678
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 10148 8676 10154 8678
rect 9846 8656 10154 8676
rect 9784 8588 9996 8616
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 9784 8022 9812 8434
rect 9772 8016 9824 8022
rect 9678 7984 9734 7993
rect 9588 7948 9640 7954
rect 9772 7958 9824 7964
rect 9678 7919 9734 7928
rect 9588 7890 9640 7896
rect 9692 7886 9720 7919
rect 9680 7880 9732 7886
rect 9680 7822 9732 7828
rect 9784 7546 9812 7958
rect 9968 7868 9996 8588
rect 10232 8288 10284 8294
rect 10232 8230 10284 8236
rect 10244 8022 10272 8230
rect 10048 8016 10100 8022
rect 10046 7984 10048 7993
rect 10232 8016 10284 8022
rect 10100 7984 10102 7993
rect 10232 7958 10284 7964
rect 10046 7919 10102 7928
rect 9968 7840 10272 7868
rect 9846 7644 10154 7664
rect 9846 7642 9852 7644
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 10148 7642 10154 7644
rect 9908 7590 9910 7642
rect 10090 7590 10092 7642
rect 9846 7588 9852 7590
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 10148 7588 10154 7590
rect 9846 7568 10154 7588
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9680 7404 9732 7410
rect 9680 7346 9732 7352
rect 9692 6798 9720 7346
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9846 6556 10154 6576
rect 9846 6554 9852 6556
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 10148 6554 10154 6556
rect 9908 6502 9910 6554
rect 10090 6502 10092 6554
rect 9846 6500 9852 6502
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 10148 6500 10154 6502
rect 9846 6480 10154 6500
rect 10244 6390 10272 7840
rect 10336 6390 10364 10474
rect 10428 10130 10456 11047
rect 10508 10600 10560 10606
rect 10508 10542 10560 10548
rect 10520 10266 10548 10542
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10416 9920 10468 9926
rect 10416 9862 10468 9868
rect 10428 9489 10456 9862
rect 10414 9480 10470 9489
rect 10414 9415 10470 9424
rect 10428 8838 10456 9415
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10428 7886 10456 8298
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10324 6384 10376 6390
rect 10324 6326 10376 6332
rect 9678 5536 9734 5545
rect 9678 5471 9734 5480
rect 9588 5364 9640 5370
rect 9588 5306 9640 5312
rect 9600 5030 9628 5306
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9692 4826 9720 5471
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9692 4622 9720 4762
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9680 4140 9732 4146
rect 9508 4100 9680 4128
rect 9508 3466 9536 4100
rect 9680 4082 9732 4088
rect 9680 3664 9732 3670
rect 9680 3606 9732 3612
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9600 2990 9628 3334
rect 9220 2984 9272 2990
rect 9220 2926 9272 2932
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 8496 2446 8524 2790
rect 9048 2446 9076 2790
rect 9692 2446 9720 3606
rect 9784 2514 9812 6326
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 5710 10272 6054
rect 10428 5710 10456 7822
rect 10508 7472 10560 7478
rect 10508 7414 10560 7420
rect 10520 7002 10548 7414
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10324 5568 10376 5574
rect 10324 5510 10376 5516
rect 9846 5468 10154 5488
rect 9846 5466 9852 5468
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 10148 5466 10154 5468
rect 9908 5414 9910 5466
rect 10090 5414 10092 5466
rect 9846 5412 9852 5414
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 10148 5412 10154 5414
rect 9846 5392 10154 5412
rect 10336 5234 10364 5510
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 9846 4380 10154 4400
rect 9846 4378 9852 4380
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 10148 4378 10154 4380
rect 9908 4326 9910 4378
rect 10090 4326 10092 4378
rect 9846 4324 9852 4326
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 10148 4324 10154 4326
rect 9846 4304 10154 4324
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 10152 3618 10180 3878
rect 10244 3738 10272 4082
rect 10336 4010 10364 5170
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10520 4146 10548 5102
rect 10612 4842 10640 12406
rect 10888 11121 10916 14214
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 10968 12708 11020 12714
rect 10968 12650 11020 12656
rect 10874 11112 10930 11121
rect 10874 11047 10930 11056
rect 10692 11008 10744 11014
rect 10692 10950 10744 10956
rect 10704 10606 10732 10950
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10692 10192 10744 10198
rect 10692 10134 10744 10140
rect 10704 6458 10732 10134
rect 10980 10130 11008 12650
rect 11060 12640 11112 12646
rect 11060 12582 11112 12588
rect 10968 10124 11020 10130
rect 10968 10066 11020 10072
rect 10980 9518 11008 10066
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10796 8634 10824 9318
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 11072 7546 11100 12582
rect 11150 11656 11206 11665
rect 11150 11591 11206 11600
rect 11164 11354 11192 11591
rect 11152 11348 11204 11354
rect 11152 11290 11204 11296
rect 11242 10704 11298 10713
rect 11242 10639 11298 10648
rect 11336 10668 11388 10674
rect 11150 9480 11206 9489
rect 11150 9415 11152 9424
rect 11204 9415 11206 9424
rect 11152 9386 11204 9392
rect 11164 8838 11192 9386
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11152 7880 11204 7886
rect 11256 7857 11284 10639
rect 11336 10610 11388 10616
rect 11348 10266 11376 10610
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11532 10062 11560 10406
rect 11520 10056 11572 10062
rect 11624 10033 11652 13806
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11716 10062 11744 10542
rect 11704 10056 11756 10062
rect 11520 9998 11572 10004
rect 11610 10024 11666 10033
rect 11704 9998 11756 10004
rect 11610 9959 11612 9968
rect 11664 9959 11666 9968
rect 11612 9930 11664 9936
rect 11624 9899 11652 9930
rect 11520 9104 11572 9110
rect 11520 9046 11572 9052
rect 11532 8673 11560 9046
rect 11808 8786 11836 14232
rect 11888 14214 11940 14220
rect 11992 12434 12020 14486
rect 12360 13870 12388 14486
rect 12544 14414 12572 14554
rect 13188 14414 13216 14554
rect 12532 14408 12584 14414
rect 12532 14350 12584 14356
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12070 13628 12378 13648
rect 12070 13626 12076 13628
rect 12132 13626 12156 13628
rect 12212 13626 12236 13628
rect 12292 13626 12316 13628
rect 12372 13626 12378 13628
rect 12132 13574 12134 13626
rect 12314 13574 12316 13626
rect 12070 13572 12076 13574
rect 12132 13572 12156 13574
rect 12212 13572 12236 13574
rect 12292 13572 12316 13574
rect 12372 13572 12378 13574
rect 12070 13552 12378 13572
rect 12070 12540 12378 12560
rect 12070 12538 12076 12540
rect 12132 12538 12156 12540
rect 12212 12538 12236 12540
rect 12292 12538 12316 12540
rect 12372 12538 12378 12540
rect 12132 12486 12134 12538
rect 12314 12486 12316 12538
rect 12070 12484 12076 12486
rect 12132 12484 12156 12486
rect 12212 12484 12236 12486
rect 12292 12484 12316 12486
rect 12372 12484 12378 12486
rect 12070 12464 12378 12484
rect 11624 8758 11836 8786
rect 11900 12406 12020 12434
rect 11518 8664 11574 8673
rect 11518 8599 11574 8608
rect 11520 8356 11572 8362
rect 11520 8298 11572 8304
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11152 7822 11204 7828
rect 11242 7848 11298 7857
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11164 7342 11192 7822
rect 11348 7818 11376 8230
rect 11242 7783 11298 7792
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11152 7336 11204 7342
rect 11152 7278 11204 7284
rect 11164 6798 11192 7278
rect 11532 6905 11560 8298
rect 11518 6896 11574 6905
rect 11518 6831 11574 6840
rect 11152 6792 11204 6798
rect 11152 6734 11204 6740
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10704 5030 10732 6258
rect 11164 6254 11192 6734
rect 11428 6656 11480 6662
rect 11428 6598 11480 6604
rect 11152 6248 11204 6254
rect 11152 6190 11204 6196
rect 11164 5778 11192 6190
rect 11440 6118 11468 6598
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11152 5772 11204 5778
rect 11152 5714 11204 5720
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11072 5302 11100 5510
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 10692 5024 10744 5030
rect 10692 4966 10744 4972
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10612 4814 10732 4842
rect 10508 4140 10560 4146
rect 10508 4082 10560 4088
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 10232 3732 10284 3738
rect 10232 3674 10284 3680
rect 10324 3664 10376 3670
rect 10060 3534 10088 3606
rect 10152 3590 10272 3618
rect 10324 3606 10376 3612
rect 10244 3534 10272 3590
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 9846 3292 10154 3312
rect 9846 3290 9852 3292
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 10148 3290 10154 3292
rect 9908 3238 9910 3290
rect 10090 3238 10092 3290
rect 9846 3236 9852 3238
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 10148 3236 10154 3238
rect 9846 3216 10154 3236
rect 10244 3194 10272 3470
rect 10232 3188 10284 3194
rect 10232 3130 10284 3136
rect 10232 2576 10284 2582
rect 10232 2518 10284 2524
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 5172 2304 5224 2310
rect 5172 2246 5224 2252
rect 5184 800 5212 2246
rect 5398 2204 5706 2224
rect 5398 2202 5404 2204
rect 5460 2202 5484 2204
rect 5540 2202 5564 2204
rect 5620 2202 5644 2204
rect 5700 2202 5706 2204
rect 5460 2150 5462 2202
rect 5642 2150 5644 2202
rect 5398 2148 5404 2150
rect 5460 2148 5484 2150
rect 5540 2148 5564 2150
rect 5620 2148 5644 2150
rect 5700 2148 5706 2150
rect 5398 2128 5706 2148
rect 5736 1714 5764 2382
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 7564 2304 7616 2310
rect 7564 2246 7616 2252
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 6104 2038 6132 2246
rect 6092 2032 6144 2038
rect 6092 1974 6144 1980
rect 5644 1686 5764 1714
rect 5644 800 5672 1686
rect 6196 800 6224 2246
rect 6656 800 6684 2246
rect 7116 800 7144 2246
rect 7576 1970 7604 2246
rect 7564 1964 7616 1970
rect 7564 1906 7616 1912
rect 7668 800 7696 2246
rect 8128 800 8156 2246
rect 8680 800 8708 2246
rect 9140 800 9168 2246
rect 9692 800 9720 2246
rect 9846 2204 10154 2224
rect 9846 2202 9852 2204
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 10148 2202 10154 2204
rect 9908 2150 9910 2202
rect 10090 2150 10092 2202
rect 9846 2148 9852 2150
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 10148 2148 10154 2150
rect 9846 2128 10154 2148
rect 10244 1170 10272 2518
rect 10336 2514 10364 3606
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10324 2508 10376 2514
rect 10324 2450 10376 2456
rect 10612 2446 10640 3334
rect 10704 2774 10732 4814
rect 10784 4820 10836 4826
rect 10784 4762 10836 4768
rect 10796 3942 10824 4762
rect 10980 4554 11008 4966
rect 11058 4720 11114 4729
rect 11058 4655 11114 4664
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10888 4185 10916 4422
rect 10874 4176 10930 4185
rect 10874 4111 10930 4120
rect 11072 4078 11100 4655
rect 11164 4622 11192 5714
rect 11532 5642 11560 6831
rect 11520 5636 11572 5642
rect 11520 5578 11572 5584
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11440 5234 11468 5306
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11242 4584 11298 4593
rect 10876 4072 10928 4078
rect 11060 4072 11112 4078
rect 10876 4014 10928 4020
rect 10980 4032 11060 4060
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10796 2922 10824 3334
rect 10888 3058 10916 4014
rect 10980 3534 11008 4032
rect 11060 4014 11112 4020
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10784 2916 10836 2922
rect 10784 2858 10836 2864
rect 10704 2746 10916 2774
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10416 2372 10468 2378
rect 10416 2314 10468 2320
rect 10428 1834 10456 2314
rect 10888 2310 10916 2746
rect 10980 2650 11008 2926
rect 11072 2854 11100 3538
rect 11164 3534 11192 4558
rect 11242 4519 11298 4528
rect 11256 4146 11284 4519
rect 11244 4140 11296 4146
rect 11244 4082 11296 4088
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 11164 3058 11192 3334
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11152 2916 11204 2922
rect 11152 2858 11204 2864
rect 11060 2848 11112 2854
rect 11060 2790 11112 2796
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 11164 2446 11192 2858
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 10508 2304 10560 2310
rect 10508 2246 10560 2252
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10876 2304 10928 2310
rect 10876 2246 10928 2252
rect 10520 2106 10548 2246
rect 10508 2100 10560 2106
rect 10508 2042 10560 2048
rect 10416 1828 10468 1834
rect 10416 1770 10468 1776
rect 10152 1142 10272 1170
rect 10152 800 10180 1142
rect 10612 800 10640 2246
rect 11152 1964 11204 1970
rect 11152 1906 11204 1912
rect 11164 800 11192 1906
rect 11256 1766 11284 3946
rect 11348 3058 11376 4966
rect 11336 3052 11388 3058
rect 11336 2994 11388 3000
rect 11440 2774 11468 5170
rect 11624 5166 11652 8758
rect 11796 7540 11848 7546
rect 11796 7482 11848 7488
rect 11704 7268 11756 7274
rect 11704 7210 11756 7216
rect 11716 5352 11744 7210
rect 11808 6934 11836 7482
rect 11796 6928 11848 6934
rect 11796 6870 11848 6876
rect 11716 5324 11836 5352
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11612 5160 11664 5166
rect 11612 5102 11664 5108
rect 11520 4072 11572 4078
rect 11518 4040 11520 4049
rect 11572 4040 11574 4049
rect 11518 3975 11574 3984
rect 11532 3398 11560 3975
rect 11716 3942 11744 5170
rect 11808 4758 11836 5324
rect 11796 4752 11848 4758
rect 11796 4694 11848 4700
rect 11900 4690 11928 12406
rect 12820 11830 12848 14214
rect 13280 14074 13308 14554
rect 13832 14414 13860 16400
rect 14188 15020 14240 15026
rect 14188 14962 14240 14968
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13464 12434 13492 14214
rect 14200 14074 14228 14962
rect 14294 14172 14602 14192
rect 14294 14170 14300 14172
rect 14356 14170 14380 14172
rect 14436 14170 14460 14172
rect 14516 14170 14540 14172
rect 14596 14170 14602 14172
rect 14356 14118 14358 14170
rect 14538 14118 14540 14170
rect 14294 14116 14300 14118
rect 14356 14116 14380 14118
rect 14436 14116 14460 14118
rect 14516 14116 14540 14118
rect 14596 14116 14602 14118
rect 14294 14096 14602 14116
rect 14188 14068 14240 14074
rect 14188 14010 14240 14016
rect 14752 13870 14780 16510
rect 15106 16400 15162 17200
rect 15750 16538 15806 17200
rect 16118 16824 16174 16833
rect 15396 16510 15806 16538
rect 14832 14408 14884 14414
rect 15120 14362 15148 16400
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 14832 14350 14884 14356
rect 14844 14006 14872 14350
rect 14936 14334 15148 14362
rect 14832 14000 14884 14006
rect 14832 13942 14884 13948
rect 14936 13938 14964 14334
rect 15108 14272 15160 14278
rect 15108 14214 15160 14220
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14094 13424 14150 13433
rect 14094 13359 14150 13368
rect 13188 12406 13492 12434
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12070 11452 12378 11472
rect 12070 11450 12076 11452
rect 12132 11450 12156 11452
rect 12212 11450 12236 11452
rect 12292 11450 12316 11452
rect 12372 11450 12378 11452
rect 12132 11398 12134 11450
rect 12314 11398 12316 11450
rect 12070 11396 12076 11398
rect 12132 11396 12156 11398
rect 12212 11396 12236 11398
rect 12292 11396 12316 11398
rect 12372 11396 12378 11398
rect 12070 11376 12378 11396
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12728 10810 12756 11290
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12912 10606 12940 10950
rect 11980 10600 12032 10606
rect 11980 10542 12032 10548
rect 12900 10600 12952 10606
rect 12900 10542 12952 10548
rect 11992 10266 12020 10542
rect 12070 10364 12378 10384
rect 12070 10362 12076 10364
rect 12132 10362 12156 10364
rect 12212 10362 12236 10364
rect 12292 10362 12316 10364
rect 12372 10362 12378 10364
rect 12132 10310 12134 10362
rect 12314 10310 12316 10362
rect 12070 10308 12076 10310
rect 12132 10308 12156 10310
rect 12212 10308 12236 10310
rect 12292 10308 12316 10310
rect 12372 10308 12378 10310
rect 12070 10288 12378 10308
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 12912 10130 12940 10542
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11992 8809 12020 9522
rect 12440 9376 12492 9382
rect 12440 9318 12492 9324
rect 12070 9276 12378 9296
rect 12070 9274 12076 9276
rect 12132 9274 12156 9276
rect 12212 9274 12236 9276
rect 12292 9274 12316 9276
rect 12372 9274 12378 9276
rect 12132 9222 12134 9274
rect 12314 9222 12316 9274
rect 12070 9220 12076 9222
rect 12132 9220 12156 9222
rect 12212 9220 12236 9222
rect 12292 9220 12316 9222
rect 12372 9220 12378 9222
rect 12070 9200 12378 9220
rect 12452 9058 12480 9318
rect 12530 9208 12586 9217
rect 12636 9178 12664 9862
rect 12820 9722 12848 9998
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12808 9716 12860 9722
rect 12808 9658 12860 9664
rect 12728 9586 12756 9658
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12992 9512 13044 9518
rect 12728 9450 12940 9466
rect 12992 9454 13044 9460
rect 12716 9444 12952 9450
rect 12768 9438 12900 9444
rect 12716 9386 12768 9392
rect 12900 9386 12952 9392
rect 12808 9376 12860 9382
rect 12806 9344 12808 9353
rect 12860 9344 12862 9353
rect 12806 9279 12862 9288
rect 12898 9208 12954 9217
rect 12530 9143 12532 9152
rect 12584 9143 12586 9152
rect 12624 9172 12676 9178
rect 12532 9114 12584 9120
rect 12898 9143 12954 9152
rect 12624 9114 12676 9120
rect 12808 9104 12860 9110
rect 12452 9052 12808 9058
rect 12452 9046 12860 9052
rect 12452 9030 12848 9046
rect 12716 8900 12768 8906
rect 12716 8842 12768 8848
rect 11978 8800 12034 8809
rect 11978 8735 12034 8744
rect 11978 8528 12034 8537
rect 11978 8463 11980 8472
rect 12032 8463 12034 8472
rect 11980 8434 12032 8440
rect 11992 7857 12020 8434
rect 12728 8362 12756 8842
rect 12912 8786 12940 9143
rect 13004 8906 13032 9454
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 12912 8758 13032 8786
rect 12532 8356 12584 8362
rect 12532 8298 12584 8304
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 12070 8188 12378 8208
rect 12070 8186 12076 8188
rect 12132 8186 12156 8188
rect 12212 8186 12236 8188
rect 12292 8186 12316 8188
rect 12372 8186 12378 8188
rect 12132 8134 12134 8186
rect 12314 8134 12316 8186
rect 12070 8132 12076 8134
rect 12132 8132 12156 8134
rect 12212 8132 12236 8134
rect 12292 8132 12316 8134
rect 12372 8132 12378 8134
rect 12070 8112 12378 8132
rect 12256 8016 12308 8022
rect 12256 7958 12308 7964
rect 11978 7848 12034 7857
rect 11978 7783 12034 7792
rect 11980 7336 12032 7342
rect 11980 7278 12032 7284
rect 11992 7002 12020 7278
rect 12268 7274 12296 7958
rect 12452 7478 12480 8230
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 12544 7410 12572 8298
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 12256 7268 12308 7274
rect 12256 7210 12308 7216
rect 12716 7200 12768 7206
rect 12716 7142 12768 7148
rect 12070 7100 12378 7120
rect 12070 7098 12076 7100
rect 12132 7098 12156 7100
rect 12212 7098 12236 7100
rect 12292 7098 12316 7100
rect 12372 7098 12378 7100
rect 12132 7046 12134 7098
rect 12314 7046 12316 7098
rect 12070 7044 12076 7046
rect 12132 7044 12156 7046
rect 12212 7044 12236 7046
rect 12292 7044 12316 7046
rect 12372 7044 12378 7046
rect 12070 7024 12378 7044
rect 11980 6996 12032 7002
rect 11980 6938 12032 6944
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 11992 6866 12020 6938
rect 12452 6866 12480 6938
rect 11980 6860 12032 6866
rect 11980 6802 12032 6808
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 11992 6304 12020 6802
rect 12440 6656 12492 6662
rect 12440 6598 12492 6604
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12072 6316 12124 6322
rect 11992 6276 12072 6304
rect 12072 6258 12124 6264
rect 12070 6012 12378 6032
rect 12070 6010 12076 6012
rect 12132 6010 12156 6012
rect 12212 6010 12236 6012
rect 12292 6010 12316 6012
rect 12372 6010 12378 6012
rect 12132 5958 12134 6010
rect 12314 5958 12316 6010
rect 12070 5956 12076 5958
rect 12132 5956 12156 5958
rect 12212 5956 12236 5958
rect 12292 5956 12316 5958
rect 12372 5956 12378 5958
rect 12070 5936 12378 5956
rect 12452 5914 12480 6598
rect 12440 5908 12492 5914
rect 12440 5850 12492 5856
rect 12636 5642 12664 6598
rect 12728 5778 12756 7142
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 12912 6458 12940 6734
rect 12900 6452 12952 6458
rect 12900 6394 12952 6400
rect 12912 5778 12940 6394
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12624 5636 12676 5642
rect 12624 5578 12676 5584
rect 13004 5137 13032 8758
rect 13096 5681 13124 10406
rect 13188 8922 13216 12406
rect 13820 12096 13872 12102
rect 13820 12038 13872 12044
rect 13636 11892 13688 11898
rect 13636 11834 13688 11840
rect 13452 11076 13504 11082
rect 13452 11018 13504 11024
rect 13464 10606 13492 11018
rect 13544 10804 13596 10810
rect 13544 10746 13596 10752
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 13358 10024 13414 10033
rect 13358 9959 13414 9968
rect 13268 9512 13320 9518
rect 13268 9454 13320 9460
rect 13280 9042 13308 9454
rect 13268 9036 13320 9042
rect 13268 8978 13320 8984
rect 13188 8894 13308 8922
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13188 8430 13216 8774
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 13280 7698 13308 8894
rect 13372 7993 13400 9959
rect 13464 9926 13492 10542
rect 13556 10198 13584 10746
rect 13648 10674 13676 11834
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13544 10192 13596 10198
rect 13544 10134 13596 10140
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13464 9450 13492 9862
rect 13648 9586 13676 10066
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13648 9450 13676 9522
rect 13452 9444 13504 9450
rect 13452 9386 13504 9392
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13464 9042 13492 9386
rect 13542 9208 13598 9217
rect 13542 9143 13598 9152
rect 13728 9172 13780 9178
rect 13556 9042 13584 9143
rect 13728 9114 13780 9120
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 13556 8838 13584 8978
rect 13544 8832 13596 8838
rect 13740 8809 13768 9114
rect 13832 9042 13860 12038
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13924 9110 13952 9318
rect 13912 9104 13964 9110
rect 13912 9046 13964 9052
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13820 8832 13872 8838
rect 13544 8774 13596 8780
rect 13726 8800 13782 8809
rect 13820 8774 13872 8780
rect 13726 8735 13782 8744
rect 13740 8566 13768 8735
rect 13832 8673 13860 8774
rect 13818 8664 13874 8673
rect 13818 8599 13874 8608
rect 13832 8566 13860 8599
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13452 8424 13504 8430
rect 13452 8366 13504 8372
rect 13358 7984 13414 7993
rect 13358 7919 13414 7928
rect 13280 7670 13400 7698
rect 13266 7304 13322 7313
rect 13266 7239 13322 7248
rect 13280 6866 13308 7239
rect 13268 6860 13320 6866
rect 13268 6802 13320 6808
rect 13280 6730 13308 6802
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13082 5672 13138 5681
rect 13082 5607 13138 5616
rect 13268 5160 13320 5166
rect 12990 5128 13046 5137
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12820 5086 12990 5114
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12070 4924 12378 4944
rect 12070 4922 12076 4924
rect 12132 4922 12156 4924
rect 12212 4922 12236 4924
rect 12292 4922 12316 4924
rect 12372 4922 12378 4924
rect 12132 4870 12134 4922
rect 12314 4870 12316 4922
rect 12070 4868 12076 4870
rect 12132 4868 12156 4870
rect 12212 4868 12236 4870
rect 12292 4868 12316 4870
rect 12372 4868 12378 4870
rect 12070 4848 12378 4868
rect 12452 4690 12480 4966
rect 12636 4826 12664 5034
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12728 4622 12756 4966
rect 12256 4616 12308 4622
rect 12256 4558 12308 4564
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11704 3936 11756 3942
rect 11756 3896 11836 3924
rect 11704 3878 11756 3884
rect 11704 3460 11756 3466
rect 11704 3402 11756 3408
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11716 2990 11744 3402
rect 11808 3346 11836 3896
rect 11900 3466 11928 4422
rect 11978 4312 12034 4321
rect 12268 4282 12296 4558
rect 11978 4247 12034 4256
rect 12072 4276 12124 4282
rect 11992 4146 12020 4247
rect 12072 4218 12124 4224
rect 12256 4276 12308 4282
rect 12256 4218 12308 4224
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 12084 3924 12112 4218
rect 12820 4162 12848 5086
rect 13268 5102 13320 5108
rect 12990 5063 13046 5072
rect 13176 4616 13228 4622
rect 13096 4564 13176 4570
rect 13096 4558 13228 4564
rect 13096 4542 13216 4558
rect 12900 4276 12952 4282
rect 12900 4218 12952 4224
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12728 4134 12848 4162
rect 11992 3896 12112 3924
rect 12440 3936 12492 3942
rect 11888 3460 11940 3466
rect 11992 3448 12020 3896
rect 12440 3878 12492 3884
rect 12070 3836 12378 3856
rect 12070 3834 12076 3836
rect 12132 3834 12156 3836
rect 12212 3834 12236 3836
rect 12292 3834 12316 3836
rect 12372 3834 12378 3836
rect 12132 3782 12134 3834
rect 12314 3782 12316 3834
rect 12070 3780 12076 3782
rect 12132 3780 12156 3782
rect 12212 3780 12236 3782
rect 12292 3780 12316 3782
rect 12372 3780 12378 3782
rect 12070 3760 12378 3780
rect 12452 3670 12480 3878
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12256 3528 12308 3534
rect 12256 3470 12308 3476
rect 12072 3460 12124 3466
rect 11992 3420 12072 3448
rect 11888 3402 11940 3408
rect 12072 3402 12124 3408
rect 11808 3318 12020 3346
rect 11704 2984 11756 2990
rect 11704 2926 11756 2932
rect 11440 2746 11652 2774
rect 11244 1760 11296 1766
rect 11244 1702 11296 1708
rect 11624 800 11652 2746
rect 11992 2632 12020 3318
rect 12268 3126 12296 3470
rect 12438 3360 12494 3369
rect 12438 3295 12494 3304
rect 12256 3120 12308 3126
rect 12256 3062 12308 3068
rect 12268 2836 12296 3062
rect 12452 2990 12480 3295
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12268 2808 12480 2836
rect 12070 2748 12378 2768
rect 12070 2746 12076 2748
rect 12132 2746 12156 2748
rect 12212 2746 12236 2748
rect 12292 2746 12316 2748
rect 12372 2746 12378 2748
rect 12132 2694 12134 2746
rect 12314 2694 12316 2746
rect 12070 2692 12076 2694
rect 12132 2692 12156 2694
rect 12212 2692 12236 2694
rect 12292 2692 12316 2694
rect 12372 2692 12378 2694
rect 12070 2672 12378 2692
rect 11992 2604 12204 2632
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 11900 1970 11928 2382
rect 11888 1964 11940 1970
rect 11888 1906 11940 1912
rect 12176 800 12204 2604
rect 12452 2530 12480 2808
rect 12544 2650 12572 4082
rect 12624 4072 12676 4078
rect 12728 4049 12756 4134
rect 12808 4072 12860 4078
rect 12624 4014 12676 4020
rect 12714 4040 12770 4049
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12360 2514 12480 2530
rect 12636 2514 12664 4014
rect 12808 4014 12860 4020
rect 12714 3975 12770 3984
rect 12716 3936 12768 3942
rect 12714 3904 12716 3913
rect 12768 3904 12770 3913
rect 12714 3839 12770 3848
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12348 2508 12480 2514
rect 12400 2502 12480 2508
rect 12624 2508 12676 2514
rect 12348 2450 12400 2456
rect 12624 2450 12676 2456
rect 12728 2122 12756 3470
rect 12820 2650 12848 4014
rect 12912 3942 12940 4218
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 13004 3738 13032 4014
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12992 3528 13044 3534
rect 12992 3470 13044 3476
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12912 3126 12940 3334
rect 12900 3120 12952 3126
rect 12900 3062 12952 3068
rect 13004 2922 13032 3470
rect 12900 2916 12952 2922
rect 12900 2858 12952 2864
rect 12992 2916 13044 2922
rect 12992 2858 13044 2864
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 12912 2446 12940 2858
rect 13096 2774 13124 4542
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13188 3534 13216 4422
rect 13280 3754 13308 5102
rect 13372 4049 13400 7670
rect 13464 7342 13492 8366
rect 13648 8022 13676 8434
rect 13924 8294 13952 9046
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13648 7562 13676 7822
rect 13648 7534 13768 7562
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 13452 6656 13504 6662
rect 13452 6598 13504 6604
rect 13464 5642 13492 6598
rect 13452 5636 13504 5642
rect 13452 5578 13504 5584
rect 13450 5536 13506 5545
rect 13556 5522 13584 7346
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13648 6866 13676 7278
rect 13740 7206 13768 7534
rect 13832 7410 13860 8026
rect 13912 7744 13964 7750
rect 13912 7686 13964 7692
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13728 7200 13780 7206
rect 13728 7142 13780 7148
rect 13740 6905 13768 7142
rect 13820 6928 13872 6934
rect 13726 6896 13782 6905
rect 13636 6860 13688 6866
rect 13820 6870 13872 6876
rect 13726 6831 13782 6840
rect 13636 6802 13688 6808
rect 13648 5778 13676 6802
rect 13832 6730 13860 6870
rect 13924 6866 13952 7686
rect 13912 6860 13964 6866
rect 13912 6802 13964 6808
rect 14016 6746 14044 11766
rect 14108 10742 14136 13359
rect 14294 13084 14602 13104
rect 14294 13082 14300 13084
rect 14356 13082 14380 13084
rect 14436 13082 14460 13084
rect 14516 13082 14540 13084
rect 14596 13082 14602 13084
rect 14356 13030 14358 13082
rect 14538 13030 14540 13082
rect 14294 13028 14300 13030
rect 14356 13028 14380 13030
rect 14436 13028 14460 13030
rect 14516 13028 14540 13030
rect 14596 13028 14602 13030
rect 14294 13008 14602 13028
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14568 12356 14596 12786
rect 14568 12328 14780 12356
rect 14294 11996 14602 12016
rect 14294 11994 14300 11996
rect 14356 11994 14380 11996
rect 14436 11994 14460 11996
rect 14516 11994 14540 11996
rect 14596 11994 14602 11996
rect 14356 11942 14358 11994
rect 14538 11942 14540 11994
rect 14294 11940 14300 11942
rect 14356 11940 14380 11942
rect 14436 11940 14460 11942
rect 14516 11940 14540 11942
rect 14596 11940 14602 11942
rect 14294 11920 14602 11940
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14096 10532 14148 10538
rect 14096 10474 14148 10480
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13924 6718 14044 6746
rect 13832 6458 13860 6666
rect 13820 6452 13872 6458
rect 13820 6394 13872 6400
rect 13832 5846 13860 6394
rect 13820 5840 13872 5846
rect 13726 5808 13782 5817
rect 13636 5772 13688 5778
rect 13820 5782 13872 5788
rect 13726 5743 13782 5752
rect 13636 5714 13688 5720
rect 13740 5642 13768 5743
rect 13728 5636 13780 5642
rect 13728 5578 13780 5584
rect 13556 5494 13676 5522
rect 13450 5471 13506 5480
rect 13464 5250 13492 5471
rect 13464 5222 13584 5250
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13358 4040 13414 4049
rect 13358 3975 13414 3984
rect 13280 3726 13400 3754
rect 13176 3528 13228 3534
rect 13176 3470 13228 3476
rect 13372 3398 13400 3726
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13464 3058 13492 4762
rect 13556 3534 13584 5222
rect 13648 4622 13676 5494
rect 13820 5160 13872 5166
rect 13820 5102 13872 5108
rect 13832 4842 13860 5102
rect 13740 4814 13860 4842
rect 13740 4758 13768 4814
rect 13728 4752 13780 4758
rect 13728 4694 13780 4700
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13648 4214 13676 4558
rect 13726 4312 13782 4321
rect 13726 4247 13782 4256
rect 13636 4208 13688 4214
rect 13636 4150 13688 4156
rect 13634 4040 13690 4049
rect 13634 3975 13690 3984
rect 13648 3777 13676 3975
rect 13634 3768 13690 3777
rect 13634 3703 13690 3712
rect 13740 3670 13768 4247
rect 13924 4078 13952 6718
rect 14004 5568 14056 5574
rect 14004 5510 14056 5516
rect 14016 5030 14044 5510
rect 14108 5370 14136 10474
rect 14200 10062 14228 11086
rect 14294 10908 14602 10928
rect 14294 10906 14300 10908
rect 14356 10906 14380 10908
rect 14436 10906 14460 10908
rect 14516 10906 14540 10908
rect 14596 10906 14602 10908
rect 14356 10854 14358 10906
rect 14538 10854 14540 10906
rect 14294 10852 14300 10854
rect 14356 10852 14380 10854
rect 14436 10852 14460 10854
rect 14516 10852 14540 10854
rect 14596 10852 14602 10854
rect 14294 10832 14602 10852
rect 14188 10056 14240 10062
rect 14188 9998 14240 10004
rect 14200 9586 14228 9998
rect 14294 9820 14602 9840
rect 14294 9818 14300 9820
rect 14356 9818 14380 9820
rect 14436 9818 14460 9820
rect 14516 9818 14540 9820
rect 14596 9818 14602 9820
rect 14356 9766 14358 9818
rect 14538 9766 14540 9818
rect 14294 9764 14300 9766
rect 14356 9764 14380 9766
rect 14436 9764 14460 9766
rect 14516 9764 14540 9766
rect 14596 9764 14602 9766
rect 14294 9744 14602 9764
rect 14188 9580 14240 9586
rect 14188 9522 14240 9528
rect 14200 8974 14228 9522
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14200 8566 14228 8910
rect 14294 8732 14602 8752
rect 14294 8730 14300 8732
rect 14356 8730 14380 8732
rect 14436 8730 14460 8732
rect 14516 8730 14540 8732
rect 14596 8730 14602 8732
rect 14356 8678 14358 8730
rect 14538 8678 14540 8730
rect 14294 8676 14300 8678
rect 14356 8676 14380 8678
rect 14436 8676 14460 8678
rect 14516 8676 14540 8678
rect 14596 8676 14602 8678
rect 14294 8656 14602 8676
rect 14660 8634 14688 11154
rect 14648 8628 14700 8634
rect 14648 8570 14700 8576
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14200 8090 14228 8502
rect 14280 8424 14332 8430
rect 14280 8366 14332 8372
rect 14188 8084 14240 8090
rect 14188 8026 14240 8032
rect 14292 7818 14320 8366
rect 14556 8356 14608 8362
rect 14556 8298 14608 8304
rect 14568 7993 14596 8298
rect 14752 8242 14780 12328
rect 14924 12164 14976 12170
rect 14924 12106 14976 12112
rect 14832 8900 14884 8906
rect 14832 8842 14884 8848
rect 14844 8634 14872 8842
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 14832 8492 14884 8498
rect 14832 8434 14884 8440
rect 14844 8265 14872 8434
rect 14660 8214 14780 8242
rect 14830 8256 14886 8265
rect 14554 7984 14610 7993
rect 14554 7919 14610 7928
rect 14280 7812 14332 7818
rect 14280 7754 14332 7760
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14200 7546 14228 7686
rect 14294 7644 14602 7664
rect 14294 7642 14300 7644
rect 14356 7642 14380 7644
rect 14436 7642 14460 7644
rect 14516 7642 14540 7644
rect 14596 7642 14602 7644
rect 14356 7590 14358 7642
rect 14538 7590 14540 7642
rect 14294 7588 14300 7590
rect 14356 7588 14380 7590
rect 14436 7588 14460 7590
rect 14516 7588 14540 7590
rect 14596 7588 14602 7590
rect 14294 7568 14602 7588
rect 14188 7540 14240 7546
rect 14188 7482 14240 7488
rect 14294 6556 14602 6576
rect 14294 6554 14300 6556
rect 14356 6554 14380 6556
rect 14436 6554 14460 6556
rect 14516 6554 14540 6556
rect 14596 6554 14602 6556
rect 14356 6502 14358 6554
rect 14538 6502 14540 6554
rect 14294 6500 14300 6502
rect 14356 6500 14380 6502
rect 14436 6500 14460 6502
rect 14516 6500 14540 6502
rect 14596 6500 14602 6502
rect 14294 6480 14602 6500
rect 14280 6384 14332 6390
rect 14280 6326 14332 6332
rect 14292 5710 14320 6326
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14476 5642 14504 6054
rect 14464 5636 14516 5642
rect 14464 5578 14516 5584
rect 14294 5468 14602 5488
rect 14294 5466 14300 5468
rect 14356 5466 14380 5468
rect 14436 5466 14460 5468
rect 14516 5466 14540 5468
rect 14596 5466 14602 5468
rect 14356 5414 14358 5466
rect 14538 5414 14540 5466
rect 14294 5412 14300 5414
rect 14356 5412 14380 5414
rect 14436 5412 14460 5414
rect 14516 5412 14540 5414
rect 14596 5412 14602 5414
rect 14294 5392 14602 5412
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 14004 5024 14056 5030
rect 14004 4966 14056 4972
rect 13912 4072 13964 4078
rect 13912 4014 13964 4020
rect 13818 3904 13874 3913
rect 13818 3839 13874 3848
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13544 3528 13596 3534
rect 13542 3496 13544 3505
rect 13596 3496 13598 3505
rect 13542 3431 13598 3440
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13004 2746 13124 2774
rect 12900 2440 12952 2446
rect 12900 2382 12952 2388
rect 12636 2106 12756 2122
rect 12624 2100 12756 2106
rect 12676 2094 12756 2100
rect 12624 2042 12676 2048
rect 12636 800 12664 2042
rect 13004 1834 13032 2746
rect 13280 2446 13308 2926
rect 13544 2916 13596 2922
rect 13544 2858 13596 2864
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 13464 2038 13492 2382
rect 13176 2032 13228 2038
rect 13176 1974 13228 1980
rect 13452 2032 13504 2038
rect 13452 1974 13504 1980
rect 12992 1828 13044 1834
rect 12992 1770 13044 1776
rect 13188 800 13216 1974
rect 13556 1442 13584 2858
rect 13648 2038 13676 3334
rect 13636 2032 13688 2038
rect 13636 1974 13688 1980
rect 13832 1902 13860 3839
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13924 2990 13952 3538
rect 13912 2984 13964 2990
rect 13912 2926 13964 2932
rect 13820 1896 13872 1902
rect 13820 1838 13872 1844
rect 14016 1442 14044 4966
rect 14294 4380 14602 4400
rect 14294 4378 14300 4380
rect 14356 4378 14380 4380
rect 14436 4378 14460 4380
rect 14516 4378 14540 4380
rect 14596 4378 14602 4380
rect 14356 4326 14358 4378
rect 14538 4326 14540 4378
rect 14294 4324 14300 4326
rect 14356 4324 14380 4326
rect 14436 4324 14460 4326
rect 14516 4324 14540 4326
rect 14596 4324 14602 4326
rect 14294 4304 14602 4324
rect 14660 4146 14688 8214
rect 14830 8191 14886 8200
rect 14936 8072 14964 12106
rect 14752 8044 14964 8072
rect 14752 6934 14780 8044
rect 14830 7984 14886 7993
rect 14830 7919 14886 7928
rect 14740 6928 14792 6934
rect 14740 6870 14792 6876
rect 14844 6882 14872 7919
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 14936 7546 14964 7822
rect 14924 7540 14976 7546
rect 14924 7482 14976 7488
rect 14844 6854 14964 6882
rect 14832 6792 14884 6798
rect 14832 6734 14884 6740
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14752 6322 14780 6598
rect 14844 6390 14872 6734
rect 14832 6384 14884 6390
rect 14832 6326 14884 6332
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14832 5364 14884 5370
rect 14832 5306 14884 5312
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14648 4140 14700 4146
rect 14648 4082 14700 4088
rect 14094 4040 14150 4049
rect 14094 3975 14150 3984
rect 14108 3534 14136 3975
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14188 3460 14240 3466
rect 14188 3402 14240 3408
rect 14200 2774 14228 3402
rect 14294 3292 14602 3312
rect 14294 3290 14300 3292
rect 14356 3290 14380 3292
rect 14436 3290 14460 3292
rect 14516 3290 14540 3292
rect 14596 3290 14602 3292
rect 14356 3238 14358 3290
rect 14538 3238 14540 3290
rect 14294 3236 14300 3238
rect 14356 3236 14380 3238
rect 14436 3236 14460 3238
rect 14516 3236 14540 3238
rect 14596 3236 14602 3238
rect 14294 3216 14602 3236
rect 14752 2774 14780 5170
rect 14108 2746 14228 2774
rect 14660 2746 14780 2774
rect 14108 2514 14136 2746
rect 14096 2508 14148 2514
rect 14096 2450 14148 2456
rect 14294 2204 14602 2224
rect 14294 2202 14300 2204
rect 14356 2202 14380 2204
rect 14436 2202 14460 2204
rect 14516 2202 14540 2204
rect 14596 2202 14602 2204
rect 14356 2150 14358 2202
rect 14538 2150 14540 2202
rect 14294 2148 14300 2150
rect 14356 2148 14380 2150
rect 14436 2148 14460 2150
rect 14516 2148 14540 2150
rect 14596 2148 14602 2150
rect 14294 2128 14602 2148
rect 13556 1414 13676 1442
rect 14016 1414 14136 1442
rect 13648 800 13676 1414
rect 14108 800 14136 1414
rect 14660 800 14688 2746
rect 3882 232 3938 241
rect 3882 167 3938 176
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 5170 0 5226 800
rect 5630 0 5686 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7102 0 7158 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8666 0 8722 800
rect 9126 0 9182 800
rect 9678 0 9734 800
rect 10138 0 10194 800
rect 10598 0 10654 800
rect 11150 0 11206 800
rect 11610 0 11666 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13174 0 13230 800
rect 13634 0 13690 800
rect 14094 0 14150 800
rect 14646 0 14702 800
rect 14844 762 14872 5306
rect 14936 5166 14964 6854
rect 15028 5302 15056 13806
rect 15120 12481 15148 14214
rect 15212 13870 15240 14894
rect 15396 13938 15424 16510
rect 15750 16400 15806 16510
rect 16040 16782 16118 16810
rect 15936 16108 15988 16114
rect 15936 16050 15988 16056
rect 15844 14544 15896 14550
rect 15844 14486 15896 14492
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15580 14074 15608 14350
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15568 14068 15620 14074
rect 15568 14010 15620 14016
rect 15384 13932 15436 13938
rect 15384 13874 15436 13880
rect 15200 13864 15252 13870
rect 15200 13806 15252 13812
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15212 12646 15240 13194
rect 15200 12640 15252 12646
rect 15200 12582 15252 12588
rect 15106 12472 15162 12481
rect 15106 12407 15162 12416
rect 15108 11620 15160 11626
rect 15108 11562 15160 11568
rect 15120 10418 15148 11562
rect 15212 10713 15240 12582
rect 15292 11076 15344 11082
rect 15292 11018 15344 11024
rect 15198 10704 15254 10713
rect 15198 10639 15254 10648
rect 15198 10568 15254 10577
rect 15198 10503 15200 10512
rect 15252 10503 15254 10512
rect 15200 10474 15252 10480
rect 15120 10390 15240 10418
rect 15212 8945 15240 10390
rect 15304 9178 15332 11018
rect 15292 9172 15344 9178
rect 15292 9114 15344 9120
rect 15198 8936 15254 8945
rect 15198 8871 15254 8880
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15290 7848 15346 7857
rect 15120 7206 15148 7822
rect 15290 7783 15346 7792
rect 15200 7744 15252 7750
rect 15200 7686 15252 7692
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15120 6254 15148 7142
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15016 5296 15068 5302
rect 15016 5238 15068 5244
rect 14924 5160 14976 5166
rect 14924 5102 14976 5108
rect 15108 4548 15160 4554
rect 15108 4490 15160 4496
rect 15016 4208 15068 4214
rect 15016 4150 15068 4156
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 14936 3194 14964 4014
rect 15028 3194 15056 4150
rect 15120 4146 15148 4490
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 15106 4040 15162 4049
rect 15106 3975 15162 3984
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 15016 3188 15068 3194
rect 15016 3130 15068 3136
rect 15120 2990 15148 3975
rect 15212 3534 15240 7686
rect 15304 7410 15332 7783
rect 15292 7404 15344 7410
rect 15292 7346 15344 7352
rect 15290 6216 15346 6225
rect 15290 6151 15346 6160
rect 15304 5574 15332 6151
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15396 5409 15424 13874
rect 15672 13530 15700 14282
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15764 11694 15792 14214
rect 15856 13938 15884 14486
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 15948 13326 15976 16050
rect 16040 14414 16068 16782
rect 16118 16759 16174 16768
rect 16302 16416 16358 16425
rect 16394 16400 16450 17200
rect 17038 16400 17094 17200
rect 17682 16538 17738 17200
rect 17328 16510 17738 16538
rect 16302 16351 16358 16360
rect 16118 15600 16174 15609
rect 16118 15535 16174 15544
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 16132 14346 16160 15535
rect 16210 15192 16266 15201
rect 16210 15127 16266 15136
rect 16120 14340 16172 14346
rect 16120 14282 16172 14288
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15844 12300 15896 12306
rect 15844 12242 15896 12248
rect 15856 11762 15884 12242
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15476 11144 15528 11150
rect 15476 11086 15528 11092
rect 15488 9738 15516 11086
rect 15568 10668 15620 10674
rect 15568 10610 15620 10616
rect 15580 10266 15608 10610
rect 15568 10260 15620 10266
rect 15568 10202 15620 10208
rect 15488 9710 15608 9738
rect 15580 9382 15608 9710
rect 15568 9376 15620 9382
rect 15474 9344 15530 9353
rect 15568 9318 15620 9324
rect 15474 9279 15530 9288
rect 15488 7410 15516 9279
rect 15566 8936 15622 8945
rect 15566 8871 15622 8880
rect 15580 7426 15608 8871
rect 15672 7954 15700 11494
rect 15764 11286 15792 11630
rect 15856 11286 15884 11698
rect 15752 11280 15804 11286
rect 15752 11222 15804 11228
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15948 11121 15976 13262
rect 15934 11112 15990 11121
rect 15844 11076 15896 11082
rect 15934 11047 15990 11056
rect 15844 11018 15896 11024
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15764 9722 15792 10542
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15856 9081 15884 11018
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15842 9072 15898 9081
rect 15842 9007 15898 9016
rect 15752 8832 15804 8838
rect 15948 8809 15976 9318
rect 15752 8774 15804 8780
rect 15934 8800 15990 8809
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15764 7857 15792 8774
rect 15934 8735 15990 8744
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15856 8090 15884 8434
rect 15936 8288 15988 8294
rect 15936 8230 15988 8236
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15948 7886 15976 8230
rect 15936 7880 15988 7886
rect 15750 7848 15806 7857
rect 15936 7822 15988 7828
rect 15750 7783 15806 7792
rect 15844 7812 15896 7818
rect 15580 7410 15700 7426
rect 15476 7404 15528 7410
rect 15580 7404 15712 7410
rect 15580 7398 15660 7404
rect 15476 7346 15528 7352
rect 15660 7346 15712 7352
rect 15488 7002 15516 7346
rect 15764 7342 15792 7783
rect 15844 7754 15896 7760
rect 15752 7336 15804 7342
rect 15752 7278 15804 7284
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15752 7200 15804 7206
rect 15752 7142 15804 7148
rect 15476 6996 15528 7002
rect 15476 6938 15528 6944
rect 15382 5400 15438 5409
rect 15382 5335 15438 5344
rect 15292 5092 15344 5098
rect 15292 5034 15344 5040
rect 15304 3602 15332 5034
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15476 5024 15528 5030
rect 15476 4966 15528 4972
rect 15396 4690 15424 4966
rect 15384 4684 15436 4690
rect 15384 4626 15436 4632
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15108 2984 15160 2990
rect 15108 2926 15160 2932
rect 15016 2916 15068 2922
rect 15016 2858 15068 2864
rect 15028 2774 15056 2858
rect 15028 2746 15148 2774
rect 15120 2650 15148 2746
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15028 870 15148 898
rect 15028 762 15056 870
rect 15120 800 15148 870
rect 14844 734 15056 762
rect 15106 0 15162 800
rect 15212 241 15240 2246
rect 15396 2106 15424 4422
rect 15488 3602 15516 4966
rect 15580 4282 15608 7142
rect 15660 6724 15712 6730
rect 15660 6666 15712 6672
rect 15672 5914 15700 6666
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15660 5228 15712 5234
rect 15660 5170 15712 5176
rect 15568 4276 15620 4282
rect 15568 4218 15620 4224
rect 15566 4040 15622 4049
rect 15566 3975 15622 3984
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15580 3058 15608 3975
rect 15672 3058 15700 5170
rect 15764 3097 15792 7142
rect 15750 3088 15806 3097
rect 15568 3052 15620 3058
rect 15568 2994 15620 3000
rect 15660 3052 15712 3058
rect 15750 3023 15806 3032
rect 15660 2994 15712 3000
rect 15672 2582 15700 2994
rect 15856 2922 15884 7754
rect 15936 7268 15988 7274
rect 15936 7210 15988 7216
rect 15948 5846 15976 7210
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 15936 5568 15988 5574
rect 15936 5510 15988 5516
rect 15948 5273 15976 5510
rect 15934 5264 15990 5273
rect 15934 5199 15990 5208
rect 16040 4622 16068 13670
rect 16132 13530 16160 14282
rect 16224 13818 16252 15127
rect 16316 13938 16344 16351
rect 16408 16114 16436 16400
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16394 16008 16450 16017
rect 16394 15943 16450 15952
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16224 13802 16344 13818
rect 16224 13796 16356 13802
rect 16224 13790 16304 13796
rect 16304 13738 16356 13744
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16316 13462 16344 13738
rect 16304 13456 16356 13462
rect 16304 13398 16356 13404
rect 16408 13394 16436 15943
rect 17052 14890 17080 16400
rect 17040 14884 17092 14890
rect 17040 14826 17092 14832
rect 16518 14716 16826 14736
rect 16518 14714 16524 14716
rect 16580 14714 16604 14716
rect 16660 14714 16684 14716
rect 16740 14714 16764 14716
rect 16820 14714 16826 14716
rect 16580 14662 16582 14714
rect 16762 14662 16764 14714
rect 16518 14660 16524 14662
rect 16580 14660 16604 14662
rect 16660 14660 16684 14662
rect 16740 14660 16764 14662
rect 16820 14660 16826 14662
rect 16518 14640 16826 14660
rect 16488 14544 16540 14550
rect 16488 14486 16540 14492
rect 16500 14278 16528 14486
rect 16488 14272 16540 14278
rect 16488 14214 16540 14220
rect 16856 13932 16908 13938
rect 16856 13874 16908 13880
rect 16518 13628 16826 13648
rect 16518 13626 16524 13628
rect 16580 13626 16604 13628
rect 16660 13626 16684 13628
rect 16740 13626 16764 13628
rect 16820 13626 16826 13628
rect 16580 13574 16582 13626
rect 16762 13574 16764 13626
rect 16518 13572 16524 13574
rect 16580 13572 16604 13574
rect 16660 13572 16684 13574
rect 16740 13572 16764 13574
rect 16820 13572 16826 13574
rect 16518 13552 16826 13572
rect 16868 13530 16896 13874
rect 17040 13864 17092 13870
rect 17038 13832 17040 13841
rect 17092 13832 17094 13841
rect 17038 13767 17094 13776
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16408 12986 16436 13330
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16518 12540 16826 12560
rect 16518 12538 16524 12540
rect 16580 12538 16604 12540
rect 16660 12538 16684 12540
rect 16740 12538 16764 12540
rect 16820 12538 16826 12540
rect 16580 12486 16582 12538
rect 16762 12486 16764 12538
rect 16518 12484 16524 12486
rect 16580 12484 16604 12486
rect 16660 12484 16684 12486
rect 16740 12484 16764 12486
rect 16820 12484 16826 12486
rect 16518 12464 16826 12484
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 16518 11452 16826 11472
rect 16518 11450 16524 11452
rect 16580 11450 16604 11452
rect 16660 11450 16684 11452
rect 16740 11450 16764 11452
rect 16820 11450 16826 11452
rect 16580 11398 16582 11450
rect 16762 11398 16764 11450
rect 16518 11396 16524 11398
rect 16580 11396 16604 11398
rect 16660 11396 16684 11398
rect 16740 11396 16764 11398
rect 16820 11396 16826 11398
rect 16518 11376 16826 11396
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 16132 10062 16160 10542
rect 16212 10532 16264 10538
rect 16212 10474 16264 10480
rect 16120 10056 16172 10062
rect 16120 9998 16172 10004
rect 16132 9178 16160 9998
rect 16120 9172 16172 9178
rect 16120 9114 16172 9120
rect 16132 9042 16160 9114
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16132 8673 16160 8774
rect 16118 8664 16174 8673
rect 16118 8599 16174 8608
rect 16224 8242 16252 10474
rect 16304 10464 16356 10470
rect 16304 10406 16356 10412
rect 16316 10062 16344 10406
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16316 9722 16344 9862
rect 16304 9716 16356 9722
rect 16304 9658 16356 9664
rect 16408 9625 16436 11086
rect 17144 11014 17172 11834
rect 17236 11150 17264 13262
rect 17328 12753 17356 16510
rect 17682 16400 17738 16510
rect 18326 16400 18382 17200
rect 18970 16538 19026 17200
rect 18800 16510 19026 16538
rect 17960 14816 18012 14822
rect 17406 14784 17462 14793
rect 17960 14758 18012 14764
rect 17406 14719 17462 14728
rect 17420 14482 17448 14719
rect 17972 14482 18000 14758
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17696 14249 17724 14350
rect 17682 14240 17738 14249
rect 17604 14198 17682 14226
rect 17498 13832 17554 13841
rect 17498 13767 17554 13776
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17314 12744 17370 12753
rect 17314 12679 17370 12688
rect 17316 12232 17368 12238
rect 17316 12174 17368 12180
rect 17328 11914 17356 12174
rect 17420 12102 17448 13126
rect 17512 12918 17540 13767
rect 17500 12912 17552 12918
rect 17500 12854 17552 12860
rect 17604 12442 17632 14198
rect 17682 14175 17738 14184
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 17696 13433 17724 13806
rect 17682 13424 17738 13433
rect 17682 13359 17738 13368
rect 17684 13320 17736 13326
rect 17684 13262 17736 13268
rect 17696 13025 17724 13262
rect 17682 13016 17738 13025
rect 17682 12951 17738 12960
rect 17684 12776 17736 12782
rect 17684 12718 17736 12724
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 17696 12617 17724 12718
rect 17682 12608 17738 12617
rect 17682 12543 17738 12552
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17684 12232 17736 12238
rect 17684 12174 17736 12180
rect 17774 12200 17830 12209
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17328 11886 17448 11914
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 16672 11008 16724 11014
rect 16670 10976 16672 10985
rect 17132 11008 17184 11014
rect 16724 10976 16726 10985
rect 17132 10950 17184 10956
rect 17224 11008 17276 11014
rect 17224 10950 17276 10956
rect 16670 10911 16726 10920
rect 17144 10849 17172 10950
rect 17130 10840 17186 10849
rect 17130 10775 17186 10784
rect 17144 10742 17172 10775
rect 17132 10736 17184 10742
rect 17132 10678 17184 10684
rect 16856 10668 16908 10674
rect 16856 10610 16908 10616
rect 16518 10364 16826 10384
rect 16518 10362 16524 10364
rect 16580 10362 16604 10364
rect 16660 10362 16684 10364
rect 16740 10362 16764 10364
rect 16820 10362 16826 10364
rect 16580 10310 16582 10362
rect 16762 10310 16764 10362
rect 16518 10308 16524 10310
rect 16580 10308 16604 10310
rect 16660 10308 16684 10310
rect 16740 10308 16764 10310
rect 16820 10308 16826 10310
rect 16518 10288 16826 10308
rect 16868 9722 16896 10610
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16960 9926 16988 10134
rect 16948 9920 17000 9926
rect 16948 9862 17000 9868
rect 16856 9716 16908 9722
rect 16856 9658 16908 9664
rect 16394 9616 16450 9625
rect 16394 9551 16450 9560
rect 16856 9580 16908 9586
rect 16302 9480 16358 9489
rect 16302 9415 16358 9424
rect 16316 8498 16344 9415
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16408 8362 16436 9551
rect 16856 9522 16908 9528
rect 16518 9276 16826 9296
rect 16518 9274 16524 9276
rect 16580 9274 16604 9276
rect 16660 9274 16684 9276
rect 16740 9274 16764 9276
rect 16820 9274 16826 9276
rect 16580 9222 16582 9274
rect 16762 9222 16764 9274
rect 16518 9220 16524 9222
rect 16580 9220 16604 9222
rect 16660 9220 16684 9222
rect 16740 9220 16764 9222
rect 16820 9220 16826 9222
rect 16518 9200 16826 9220
rect 16868 9178 16896 9522
rect 16960 9518 16988 9862
rect 17040 9580 17092 9586
rect 17040 9522 17092 9528
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 17052 9178 17080 9522
rect 17132 9512 17184 9518
rect 17132 9454 17184 9460
rect 16856 9172 16908 9178
rect 16856 9114 16908 9120
rect 17040 9172 17092 9178
rect 17040 9114 17092 9120
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16500 8430 16528 8978
rect 16672 8832 16724 8838
rect 16670 8800 16672 8809
rect 16724 8800 16726 8809
rect 16670 8735 16726 8744
rect 16488 8424 16540 8430
rect 16488 8366 16540 8372
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16132 8214 16252 8242
rect 16132 7410 16160 8214
rect 16518 8188 16826 8208
rect 16518 8186 16524 8188
rect 16580 8186 16604 8188
rect 16660 8186 16684 8188
rect 16740 8186 16764 8188
rect 16820 8186 16826 8188
rect 16580 8134 16582 8186
rect 16762 8134 16764 8186
rect 16518 8132 16524 8134
rect 16580 8132 16604 8134
rect 16660 8132 16684 8134
rect 16740 8132 16764 8134
rect 16820 8132 16826 8134
rect 16518 8112 16826 8132
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16132 6769 16160 7346
rect 16118 6760 16174 6769
rect 16118 6695 16174 6704
rect 16120 6656 16172 6662
rect 16120 6598 16172 6604
rect 16132 6254 16160 6598
rect 16224 6338 16252 7822
rect 16868 7750 16896 9114
rect 16948 8832 17000 8838
rect 16948 8774 17000 8780
rect 16960 8634 16988 8774
rect 17144 8634 17172 9454
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16960 8090 16988 8366
rect 17052 8090 17080 8434
rect 16948 8084 17000 8090
rect 16948 8026 17000 8032
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17236 7970 17264 10950
rect 17328 9058 17356 11630
rect 17420 11558 17448 11886
rect 17696 11801 17724 12174
rect 17972 12170 18000 12718
rect 17774 12135 17830 12144
rect 17960 12164 18012 12170
rect 17682 11792 17738 11801
rect 17500 11756 17552 11762
rect 17788 11762 17816 12135
rect 17960 12106 18012 12112
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17682 11727 17738 11736
rect 17776 11756 17828 11762
rect 17500 11698 17552 11704
rect 17776 11698 17828 11704
rect 17408 11552 17460 11558
rect 17406 11520 17408 11529
rect 17460 11520 17462 11529
rect 17406 11455 17462 11464
rect 17512 11257 17540 11698
rect 17776 11620 17828 11626
rect 17776 11562 17828 11568
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17498 11248 17554 11257
rect 17498 11183 17554 11192
rect 17604 11150 17632 11290
rect 17408 11144 17460 11150
rect 17408 11086 17460 11092
rect 17592 11144 17644 11150
rect 17592 11086 17644 11092
rect 17684 11144 17736 11150
rect 17684 11086 17736 11092
rect 17420 10010 17448 11086
rect 17696 10849 17724 11086
rect 17682 10840 17738 10849
rect 17682 10775 17738 10784
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17500 10464 17552 10470
rect 17696 10441 17724 10542
rect 17500 10406 17552 10412
rect 17682 10432 17738 10441
rect 17512 10130 17540 10406
rect 17682 10367 17738 10376
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17420 9982 17540 10010
rect 17408 9920 17460 9926
rect 17408 9862 17460 9868
rect 17420 9178 17448 9862
rect 17512 9178 17540 9982
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17592 9376 17644 9382
rect 17592 9318 17644 9324
rect 17408 9172 17460 9178
rect 17408 9114 17460 9120
rect 17500 9172 17552 9178
rect 17500 9114 17552 9120
rect 17328 9030 17448 9058
rect 17604 9042 17632 9318
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 16948 7948 17000 7954
rect 16948 7890 17000 7896
rect 17052 7942 17264 7970
rect 17328 7954 17356 8502
rect 17316 7948 17368 7954
rect 16396 7744 16448 7750
rect 16396 7686 16448 7692
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16316 6458 16344 6598
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16224 6310 16344 6338
rect 16120 6248 16172 6254
rect 16120 6190 16172 6196
rect 16212 6112 16264 6118
rect 16212 6054 16264 6060
rect 16224 5914 16252 6054
rect 16212 5908 16264 5914
rect 16212 5850 16264 5856
rect 16210 5536 16266 5545
rect 16210 5471 16266 5480
rect 16224 5234 16252 5471
rect 16316 5370 16344 6310
rect 16304 5364 16356 5370
rect 16304 5306 16356 5312
rect 16212 5228 16264 5234
rect 16212 5170 16264 5176
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16316 4690 16344 4966
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16028 4616 16080 4622
rect 16028 4558 16080 4564
rect 16118 4584 16174 4593
rect 16118 4519 16174 4528
rect 16132 4282 16160 4519
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 15948 3233 15976 4218
rect 16408 4146 16436 7686
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 16776 7342 16804 7482
rect 16856 7404 16908 7410
rect 16856 7346 16908 7352
rect 16764 7336 16816 7342
rect 16764 7278 16816 7284
rect 16518 7100 16826 7120
rect 16518 7098 16524 7100
rect 16580 7098 16604 7100
rect 16660 7098 16684 7100
rect 16740 7098 16764 7100
rect 16820 7098 16826 7100
rect 16580 7046 16582 7098
rect 16762 7046 16764 7098
rect 16518 7044 16524 7046
rect 16580 7044 16604 7046
rect 16660 7044 16684 7046
rect 16740 7044 16764 7046
rect 16820 7044 16826 7046
rect 16518 7024 16826 7044
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16670 6896 16726 6905
rect 16500 6390 16528 6870
rect 16868 6866 16896 7346
rect 16670 6831 16672 6840
rect 16724 6831 16726 6840
rect 16856 6860 16908 6866
rect 16672 6802 16724 6808
rect 16856 6802 16908 6808
rect 16868 6730 16896 6802
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16672 6656 16724 6662
rect 16672 6598 16724 6604
rect 16684 6458 16712 6598
rect 16672 6452 16724 6458
rect 16672 6394 16724 6400
rect 16488 6384 16540 6390
rect 16488 6326 16540 6332
rect 16762 6352 16818 6361
rect 16762 6287 16818 6296
rect 16856 6316 16908 6322
rect 16776 6254 16804 6287
rect 16856 6258 16908 6264
rect 16488 6248 16540 6254
rect 16486 6216 16488 6225
rect 16764 6248 16816 6254
rect 16540 6216 16542 6225
rect 16764 6190 16816 6196
rect 16486 6151 16542 6160
rect 16518 6012 16826 6032
rect 16518 6010 16524 6012
rect 16580 6010 16604 6012
rect 16660 6010 16684 6012
rect 16740 6010 16764 6012
rect 16820 6010 16826 6012
rect 16580 5958 16582 6010
rect 16762 5958 16764 6010
rect 16518 5956 16524 5958
rect 16580 5956 16604 5958
rect 16660 5956 16684 5958
rect 16740 5956 16764 5958
rect 16820 5956 16826 5958
rect 16518 5936 16826 5956
rect 16868 5710 16896 6258
rect 16856 5704 16908 5710
rect 16578 5672 16634 5681
rect 16856 5646 16908 5652
rect 16578 5607 16634 5616
rect 16592 5574 16620 5607
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16672 5568 16724 5574
rect 16672 5510 16724 5516
rect 16684 5370 16712 5510
rect 16854 5400 16910 5409
rect 16672 5364 16724 5370
rect 16854 5335 16910 5344
rect 16672 5306 16724 5312
rect 16518 4924 16826 4944
rect 16518 4922 16524 4924
rect 16580 4922 16604 4924
rect 16660 4922 16684 4924
rect 16740 4922 16764 4924
rect 16820 4922 16826 4924
rect 16580 4870 16582 4922
rect 16762 4870 16764 4922
rect 16518 4868 16524 4870
rect 16580 4868 16604 4870
rect 16660 4868 16684 4870
rect 16740 4868 16764 4870
rect 16820 4868 16826 4870
rect 16518 4848 16826 4868
rect 16868 4690 16896 5335
rect 16856 4684 16908 4690
rect 16856 4626 16908 4632
rect 16854 4312 16910 4321
rect 16854 4247 16910 4256
rect 16396 4140 16448 4146
rect 16396 4082 16448 4088
rect 16868 4078 16896 4247
rect 16672 4072 16724 4078
rect 16670 4040 16672 4049
rect 16856 4072 16908 4078
rect 16724 4040 16726 4049
rect 16856 4014 16908 4020
rect 16670 3975 16726 3984
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 15934 3224 15990 3233
rect 15934 3159 15990 3168
rect 16040 3126 16068 3878
rect 16316 3670 16344 3878
rect 16518 3836 16826 3856
rect 16518 3834 16524 3836
rect 16580 3834 16604 3836
rect 16660 3834 16684 3836
rect 16740 3834 16764 3836
rect 16820 3834 16826 3836
rect 16580 3782 16582 3834
rect 16762 3782 16764 3834
rect 16518 3780 16524 3782
rect 16580 3780 16604 3782
rect 16660 3780 16684 3782
rect 16740 3780 16764 3782
rect 16820 3780 16826 3782
rect 16518 3760 16826 3780
rect 16304 3664 16356 3670
rect 16304 3606 16356 3612
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 16960 3058 16988 7890
rect 17052 6322 17080 7942
rect 17316 7890 17368 7896
rect 17132 7880 17184 7886
rect 17420 7834 17448 9030
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17500 8900 17552 8906
rect 17500 8842 17552 8848
rect 17512 8634 17540 8842
rect 17604 8809 17632 8978
rect 17696 8974 17724 9862
rect 17788 9518 17816 11562
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17788 9353 17816 9454
rect 17774 9344 17830 9353
rect 17774 9279 17830 9288
rect 17880 9194 17908 12038
rect 18064 11898 18092 13806
rect 18340 12646 18368 16400
rect 18800 13297 18828 16510
rect 18970 16400 19026 16510
rect 19614 16400 19670 17200
rect 18786 13288 18842 13297
rect 18786 13223 18842 13232
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18800 12434 18828 13223
rect 19628 12850 19656 16400
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 18800 12406 19012 12434
rect 18144 12300 18196 12306
rect 18144 12242 18196 12248
rect 18052 11892 18104 11898
rect 18052 11834 18104 11840
rect 17960 11688 18012 11694
rect 17960 11630 18012 11636
rect 17972 10810 18000 11630
rect 17960 10804 18012 10810
rect 17960 10746 18012 10752
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17972 10033 18000 10542
rect 17958 10024 18014 10033
rect 17958 9959 18014 9968
rect 18156 9674 18184 12242
rect 18604 10668 18656 10674
rect 18604 10610 18656 10616
rect 18420 10056 18472 10062
rect 18418 10024 18420 10033
rect 18472 10024 18474 10033
rect 18236 9988 18288 9994
rect 18418 9959 18474 9968
rect 18236 9930 18288 9936
rect 17788 9166 17908 9194
rect 18064 9646 18184 9674
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17590 8800 17646 8809
rect 17788 8786 17816 9166
rect 17866 9072 17922 9081
rect 17866 9007 17922 9016
rect 17590 8735 17646 8744
rect 17696 8758 17816 8786
rect 17500 8628 17552 8634
rect 17500 8570 17552 8576
rect 17500 8016 17552 8022
rect 17500 7958 17552 7964
rect 17132 7822 17184 7828
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17040 6180 17092 6186
rect 17040 6122 17092 6128
rect 17052 5914 17080 6122
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17144 5794 17172 7822
rect 17328 7806 17448 7834
rect 17224 7744 17276 7750
rect 17222 7712 17224 7721
rect 17276 7712 17278 7721
rect 17222 7647 17278 7656
rect 17236 7002 17264 7647
rect 17224 6996 17276 7002
rect 17224 6938 17276 6944
rect 17224 6860 17276 6866
rect 17224 6802 17276 6808
rect 17236 6254 17264 6802
rect 17328 6322 17356 7806
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17420 7313 17448 7346
rect 17406 7304 17462 7313
rect 17406 7239 17462 7248
rect 17512 6984 17540 7958
rect 17512 6956 17632 6984
rect 17408 6928 17460 6934
rect 17460 6888 17540 6916
rect 17408 6870 17460 6876
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17420 6497 17448 6598
rect 17406 6488 17462 6497
rect 17406 6423 17462 6432
rect 17512 6372 17540 6888
rect 17420 6344 17540 6372
rect 17316 6316 17368 6322
rect 17316 6258 17368 6264
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 17052 5766 17172 5794
rect 17236 5778 17264 6190
rect 17316 6180 17368 6186
rect 17316 6122 17368 6128
rect 17224 5772 17276 5778
rect 17052 4146 17080 5766
rect 17224 5714 17276 5720
rect 17328 5642 17356 6122
rect 17316 5636 17368 5642
rect 17316 5578 17368 5584
rect 17130 5536 17186 5545
rect 17130 5471 17186 5480
rect 17144 5370 17172 5471
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 17328 5302 17356 5578
rect 17316 5296 17368 5302
rect 17316 5238 17368 5244
rect 17328 5166 17356 5238
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17420 5012 17448 6344
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 17512 5370 17540 5510
rect 17500 5364 17552 5370
rect 17500 5306 17552 5312
rect 17328 4984 17448 5012
rect 17132 4820 17184 4826
rect 17132 4762 17184 4768
rect 17040 4140 17092 4146
rect 17040 4082 17092 4088
rect 17144 3618 17172 4762
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17052 3590 17172 3618
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 16316 2961 16344 2994
rect 16302 2952 16358 2961
rect 15844 2916 15896 2922
rect 16302 2887 16358 2896
rect 15844 2858 15896 2864
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16518 2748 16826 2768
rect 16518 2746 16524 2748
rect 16580 2746 16604 2748
rect 16660 2746 16684 2748
rect 16740 2746 16764 2748
rect 16820 2746 16826 2748
rect 16580 2694 16582 2746
rect 16762 2694 16764 2746
rect 16518 2692 16524 2694
rect 16580 2692 16604 2694
rect 16660 2692 16684 2694
rect 16740 2692 16764 2694
rect 16820 2692 16826 2694
rect 16518 2672 16826 2692
rect 15660 2576 15712 2582
rect 16672 2576 16724 2582
rect 15660 2518 15712 2524
rect 16500 2524 16672 2530
rect 16500 2518 16724 2524
rect 16500 2502 16712 2518
rect 16028 2440 16080 2446
rect 16028 2382 16080 2388
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 15384 2100 15436 2106
rect 15384 2042 15436 2048
rect 15672 800 15700 2246
rect 16040 1766 16068 2382
rect 16028 1760 16080 1766
rect 16028 1702 16080 1708
rect 16132 870 16252 898
rect 16132 800 16160 870
rect 15198 232 15254 241
rect 15198 167 15254 176
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16224 762 16252 870
rect 16500 762 16528 2502
rect 16672 2440 16724 2446
rect 16856 2440 16908 2446
rect 16724 2388 16804 2394
rect 16672 2382 16804 2388
rect 16856 2382 16908 2388
rect 16684 2366 16804 2382
rect 16776 2310 16804 2366
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16684 800 16712 2246
rect 16868 1902 16896 2382
rect 16856 1896 16908 1902
rect 16856 1838 16908 1844
rect 16960 1465 16988 2790
rect 17052 2310 17080 3590
rect 17130 3496 17186 3505
rect 17130 3431 17132 3440
rect 17184 3431 17186 3440
rect 17132 3402 17184 3408
rect 17130 3088 17186 3097
rect 17130 3023 17132 3032
rect 17184 3023 17186 3032
rect 17132 2994 17184 3000
rect 17132 2576 17184 2582
rect 17132 2518 17184 2524
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 16946 1456 17002 1465
rect 16946 1391 17002 1400
rect 17144 800 17172 2518
rect 17236 2446 17264 3674
rect 17328 3534 17356 4984
rect 17604 4264 17632 6956
rect 17696 6662 17724 8758
rect 17880 8634 17908 9007
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17960 8492 18012 8498
rect 18064 8480 18092 9646
rect 18012 8452 18092 8480
rect 17960 8434 18012 8440
rect 18052 8288 18104 8294
rect 18052 8230 18104 8236
rect 17960 7880 18012 7886
rect 17958 7848 17960 7857
rect 18012 7848 18014 7857
rect 17958 7783 18014 7792
rect 18064 7750 18092 8230
rect 18248 7886 18276 9930
rect 18328 9444 18380 9450
rect 18328 9386 18380 9392
rect 18340 8362 18368 9386
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18328 8356 18380 8362
rect 18328 8298 18380 8304
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17868 7472 17920 7478
rect 17972 7449 18000 7482
rect 17868 7414 17920 7420
rect 17958 7440 18014 7449
rect 17776 7268 17828 7274
rect 17776 7210 17828 7216
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17696 5642 17724 6054
rect 17788 5778 17816 7210
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17880 5234 17908 7414
rect 17958 7375 18014 7384
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 17960 6656 18012 6662
rect 17960 6598 18012 6604
rect 17972 6458 18000 6598
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 18064 6304 18092 7278
rect 18156 6458 18184 7346
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 17972 6276 18092 6304
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 17774 4856 17830 4865
rect 17774 4791 17830 4800
rect 17420 4236 17632 4264
rect 17420 3534 17448 4236
rect 17498 4176 17554 4185
rect 17498 4111 17554 4120
rect 17592 4140 17644 4146
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17512 3482 17540 4111
rect 17592 4082 17644 4088
rect 17604 3602 17632 4082
rect 17788 3942 17816 4791
rect 17866 4448 17922 4457
rect 17866 4383 17922 4392
rect 17880 4010 17908 4383
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17696 3641 17724 3878
rect 17682 3632 17738 3641
rect 17592 3596 17644 3602
rect 17682 3567 17738 3576
rect 17592 3538 17644 3544
rect 17684 3528 17736 3534
rect 17512 3476 17684 3482
rect 17512 3470 17736 3476
rect 17512 3454 17724 3470
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17512 3058 17540 3334
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17328 1057 17356 2790
rect 17500 2440 17552 2446
rect 17500 2382 17552 2388
rect 17512 2038 17540 2382
rect 17500 2032 17552 2038
rect 17500 1974 17552 1980
rect 17604 1873 17632 3334
rect 17866 3224 17922 3233
rect 17866 3159 17922 3168
rect 17880 3058 17908 3159
rect 17972 3058 18000 6276
rect 18050 6216 18106 6225
rect 18050 6151 18106 6160
rect 18064 5914 18092 6151
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 18248 5250 18276 7346
rect 18340 6322 18368 8298
rect 18432 8265 18460 8774
rect 18510 8664 18566 8673
rect 18510 8599 18566 8608
rect 18418 8256 18474 8265
rect 18418 8191 18474 8200
rect 18418 7848 18474 7857
rect 18418 7783 18474 7792
rect 18432 7546 18460 7783
rect 18420 7540 18472 7546
rect 18420 7482 18472 7488
rect 18418 7032 18474 7041
rect 18418 6967 18420 6976
rect 18472 6967 18474 6976
rect 18420 6938 18472 6944
rect 18418 6624 18474 6633
rect 18418 6559 18474 6568
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 18432 5914 18460 6559
rect 18420 5908 18472 5914
rect 18420 5850 18472 5856
rect 18418 5672 18474 5681
rect 18418 5607 18474 5616
rect 18156 5222 18276 5250
rect 18052 5160 18104 5166
rect 18050 5128 18052 5137
rect 18104 5128 18106 5137
rect 18050 5063 18106 5072
rect 18156 5030 18184 5222
rect 18236 5092 18288 5098
rect 18236 5034 18288 5040
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18144 4752 18196 4758
rect 18144 4694 18196 4700
rect 18156 3534 18184 4694
rect 18248 4146 18276 5034
rect 18432 4826 18460 5607
rect 18524 5370 18552 8599
rect 18616 6322 18644 10610
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18604 6316 18656 6322
rect 18604 6258 18656 6264
rect 18512 5364 18564 5370
rect 18512 5306 18564 5312
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18708 4690 18736 7686
rect 18800 7585 18828 8978
rect 18786 7576 18842 7585
rect 18786 7511 18842 7520
rect 18800 5234 18828 7511
rect 18788 5228 18840 5234
rect 18788 5170 18840 5176
rect 18696 4684 18748 4690
rect 18696 4626 18748 4632
rect 18328 4616 18380 4622
rect 18328 4558 18380 4564
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18064 3233 18092 3334
rect 18050 3224 18106 3233
rect 18340 3194 18368 4558
rect 18418 4040 18474 4049
rect 18418 3975 18474 3984
rect 18432 3738 18460 3975
rect 18420 3732 18472 3738
rect 18420 3674 18472 3680
rect 18604 3664 18656 3670
rect 18604 3606 18656 3612
rect 18050 3159 18106 3168
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17868 2848 17920 2854
rect 17868 2790 17920 2796
rect 18420 2848 18472 2854
rect 18420 2790 18472 2796
rect 17684 2304 17736 2310
rect 17684 2246 17736 2252
rect 17590 1864 17646 1873
rect 17590 1799 17646 1808
rect 17696 1170 17724 2246
rect 17604 1142 17724 1170
rect 17314 1048 17370 1057
rect 17314 983 17370 992
rect 17604 800 17632 1142
rect 17788 921 17816 2790
rect 17880 2281 17908 2790
rect 18432 2689 18460 2790
rect 18418 2680 18474 2689
rect 18418 2615 18474 2624
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 18144 2304 18196 2310
rect 17866 2272 17922 2281
rect 18144 2246 18196 2252
rect 17866 2207 17922 2216
rect 17774 912 17830 921
rect 17774 847 17830 856
rect 18156 800 18184 2246
rect 18248 2106 18276 2382
rect 18236 2100 18288 2106
rect 18236 2042 18288 2048
rect 18616 800 18644 3606
rect 18984 2650 19012 12406
rect 19616 3460 19668 3466
rect 19616 3402 19668 3408
rect 19156 3120 19208 3126
rect 19156 3062 19208 3068
rect 18972 2644 19024 2650
rect 18972 2586 19024 2592
rect 19168 800 19196 3062
rect 19628 800 19656 3402
rect 16224 734 16528 762
rect 16670 0 16726 800
rect 17130 0 17186 800
rect 17590 0 17646 800
rect 18142 0 18198 800
rect 18602 0 18658 800
rect 19154 0 19210 800
rect 19614 0 19670 800
<< via2 >>
rect 2226 14456 2282 14512
rect 2226 13912 2282 13968
rect 1950 12824 2006 12880
rect 1950 11092 1952 11112
rect 1952 11092 2004 11112
rect 2004 11092 2006 11112
rect 1950 11056 2006 11092
rect 1582 10668 1638 10704
rect 1582 10648 1584 10668
rect 1584 10648 1636 10668
rect 1636 10648 1638 10668
rect 1490 10512 1546 10568
rect 1306 9288 1362 9344
rect 3790 16768 3846 16824
rect 2778 13504 2834 13560
rect 3054 15952 3110 16008
rect 2962 14728 3018 14784
rect 3180 14714 3236 14716
rect 3260 14714 3316 14716
rect 3340 14714 3396 14716
rect 3420 14714 3476 14716
rect 3180 14662 3226 14714
rect 3226 14662 3236 14714
rect 3260 14662 3290 14714
rect 3290 14662 3302 14714
rect 3302 14662 3316 14714
rect 3340 14662 3354 14714
rect 3354 14662 3366 14714
rect 3366 14662 3396 14714
rect 3420 14662 3430 14714
rect 3430 14662 3476 14714
rect 3180 14660 3236 14662
rect 3260 14660 3316 14662
rect 3340 14660 3396 14662
rect 3420 14660 3476 14662
rect 3882 16360 3938 16416
rect 3606 15136 3662 15192
rect 3054 14320 3110 14376
rect 3422 14340 3478 14376
rect 3422 14320 3424 14340
rect 3424 14320 3476 14340
rect 3476 14320 3478 14340
rect 3180 13626 3236 13628
rect 3260 13626 3316 13628
rect 3340 13626 3396 13628
rect 3420 13626 3476 13628
rect 3180 13574 3226 13626
rect 3226 13574 3236 13626
rect 3260 13574 3290 13626
rect 3290 13574 3302 13626
rect 3302 13574 3316 13626
rect 3340 13574 3354 13626
rect 3354 13574 3366 13626
rect 3366 13574 3396 13626
rect 3420 13574 3430 13626
rect 3430 13574 3476 13626
rect 3180 13572 3236 13574
rect 3260 13572 3316 13574
rect 3340 13572 3396 13574
rect 3420 13572 3476 13574
rect 2778 13232 2834 13288
rect 2226 13132 2228 13152
rect 2228 13132 2280 13152
rect 2280 13132 2282 13152
rect 2226 13096 2282 13132
rect 2226 12724 2228 12744
rect 2228 12724 2280 12744
rect 2280 12724 2282 12744
rect 1858 10104 1914 10160
rect 1674 8472 1730 8528
rect 1490 7656 1546 7712
rect 1858 8064 1914 8120
rect 1950 7792 2006 7848
rect 1858 6432 1914 6488
rect 1490 6060 1492 6080
rect 1492 6060 1544 6080
rect 1544 6060 1546 6080
rect 1490 6024 1546 6060
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 1858 6160 1914 6216
rect 1766 5652 1768 5672
rect 1768 5652 1820 5672
rect 1820 5652 1822 5672
rect 2226 12688 2282 12724
rect 2226 11328 2282 11384
rect 2226 10920 2282 10976
rect 2318 10004 2320 10024
rect 2320 10004 2372 10024
rect 2372 10004 2374 10024
rect 2318 9968 2374 10004
rect 2134 8472 2190 8528
rect 2410 9696 2466 9752
rect 2410 9016 2466 9072
rect 2226 7928 2282 7984
rect 2226 7268 2282 7304
rect 2226 7248 2228 7268
rect 2228 7248 2280 7268
rect 2280 7248 2282 7268
rect 2318 6876 2320 6896
rect 2320 6876 2372 6896
rect 2372 6876 2374 6896
rect 2318 6840 2374 6876
rect 1766 5616 1822 5652
rect 1490 5092 1546 5128
rect 1490 5072 1492 5092
rect 1492 5072 1544 5092
rect 1544 5072 1546 5092
rect 1858 4664 1914 4720
rect 1490 4256 1546 4312
rect 2042 4564 2044 4584
rect 2044 4564 2096 4584
rect 2096 4564 2098 4584
rect 2042 4528 2098 4564
rect 2778 11872 2834 11928
rect 2962 13368 3018 13424
rect 4158 15544 4214 15600
rect 3514 13232 3570 13288
rect 3180 12538 3236 12540
rect 3260 12538 3316 12540
rect 3340 12538 3396 12540
rect 3420 12538 3476 12540
rect 3180 12486 3226 12538
rect 3226 12486 3236 12538
rect 3260 12486 3290 12538
rect 3290 12486 3302 12538
rect 3302 12486 3316 12538
rect 3340 12486 3354 12538
rect 3354 12486 3366 12538
rect 3366 12486 3396 12538
rect 3420 12486 3430 12538
rect 3430 12486 3476 12538
rect 3180 12484 3236 12486
rect 3260 12484 3316 12486
rect 3340 12484 3396 12486
rect 3420 12484 3476 12486
rect 3238 12280 3294 12336
rect 2962 12008 3018 12064
rect 2594 9560 2650 9616
rect 3180 11450 3236 11452
rect 3260 11450 3316 11452
rect 3340 11450 3396 11452
rect 3420 11450 3476 11452
rect 3180 11398 3226 11450
rect 3226 11398 3236 11450
rect 3260 11398 3290 11450
rect 3290 11398 3302 11450
rect 3302 11398 3316 11450
rect 3340 11398 3354 11450
rect 3354 11398 3366 11450
rect 3366 11398 3396 11450
rect 3420 11398 3430 11450
rect 3430 11398 3476 11450
rect 3180 11396 3236 11398
rect 3260 11396 3316 11398
rect 3340 11396 3396 11398
rect 3420 11396 3476 11398
rect 3698 11756 3754 11792
rect 3698 11736 3700 11756
rect 3700 11736 3752 11756
rect 3752 11736 3754 11756
rect 3422 11212 3478 11248
rect 3422 11192 3424 11212
rect 3424 11192 3476 11212
rect 3476 11192 3478 11212
rect 3180 10362 3236 10364
rect 3260 10362 3316 10364
rect 3340 10362 3396 10364
rect 3420 10362 3476 10364
rect 3180 10310 3226 10362
rect 3226 10310 3236 10362
rect 3260 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3316 10362
rect 3340 10310 3354 10362
rect 3354 10310 3366 10362
rect 3366 10310 3396 10362
rect 3420 10310 3430 10362
rect 3430 10310 3476 10362
rect 3180 10308 3236 10310
rect 3260 10308 3316 10310
rect 3340 10308 3396 10310
rect 3420 10308 3476 10310
rect 3974 11600 4030 11656
rect 4066 11192 4122 11248
rect 3698 10104 3754 10160
rect 3606 9424 3662 9480
rect 3180 9274 3236 9276
rect 3260 9274 3316 9276
rect 3340 9274 3396 9276
rect 3420 9274 3476 9276
rect 3180 9222 3226 9274
rect 3226 9222 3236 9274
rect 3260 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3316 9274
rect 3340 9222 3354 9274
rect 3354 9222 3366 9274
rect 3366 9222 3396 9274
rect 3420 9222 3430 9274
rect 3430 9222 3476 9274
rect 3180 9220 3236 9222
rect 3260 9220 3316 9222
rect 3340 9220 3396 9222
rect 3420 9220 3476 9222
rect 3054 8916 3056 8936
rect 3056 8916 3108 8936
rect 3108 8916 3110 8936
rect 3054 8880 3110 8916
rect 3422 8900 3478 8936
rect 3422 8880 3424 8900
rect 3424 8880 3476 8900
rect 3476 8880 3478 8900
rect 2226 5072 2282 5128
rect 1490 3884 1492 3904
rect 1492 3884 1544 3904
rect 1544 3884 1546 3904
rect 1490 3848 1546 3884
rect 1490 3440 1546 3496
rect 1490 2624 1546 2680
rect 1490 2252 1492 2272
rect 1492 2252 1544 2272
rect 1544 2252 1546 2272
rect 1490 2216 1546 2252
rect 1858 3440 1914 3496
rect 1858 3032 1914 3088
rect 2134 3304 2190 3360
rect 2410 4528 2466 4584
rect 2502 4256 2558 4312
rect 3180 8186 3236 8188
rect 3260 8186 3316 8188
rect 3340 8186 3396 8188
rect 3420 8186 3476 8188
rect 3180 8134 3226 8186
rect 3226 8134 3236 8186
rect 3260 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3316 8186
rect 3340 8134 3354 8186
rect 3354 8134 3366 8186
rect 3366 8134 3396 8186
rect 3420 8134 3430 8186
rect 3430 8134 3476 8186
rect 3180 8132 3236 8134
rect 3260 8132 3316 8134
rect 3340 8132 3396 8134
rect 3420 8132 3476 8134
rect 3146 7828 3148 7848
rect 3148 7828 3200 7848
rect 3200 7828 3202 7848
rect 3146 7792 3202 7828
rect 3146 7404 3202 7440
rect 3146 7384 3148 7404
rect 3148 7384 3200 7404
rect 3200 7384 3202 7404
rect 3180 7098 3236 7100
rect 3260 7098 3316 7100
rect 3340 7098 3396 7100
rect 3420 7098 3476 7100
rect 3180 7046 3226 7098
rect 3226 7046 3236 7098
rect 3260 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3316 7098
rect 3340 7046 3354 7098
rect 3354 7046 3366 7098
rect 3366 7046 3396 7098
rect 3420 7046 3430 7098
rect 3430 7046 3476 7098
rect 3180 7044 3236 7046
rect 3260 7044 3316 7046
rect 3340 7044 3396 7046
rect 3420 7044 3476 7046
rect 3180 6010 3236 6012
rect 3260 6010 3316 6012
rect 3340 6010 3396 6012
rect 3420 6010 3476 6012
rect 3180 5958 3226 6010
rect 3226 5958 3236 6010
rect 3260 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3316 6010
rect 3340 5958 3354 6010
rect 3354 5958 3366 6010
rect 3366 5958 3396 6010
rect 3420 5958 3430 6010
rect 3430 5958 3476 6010
rect 3180 5956 3236 5958
rect 3260 5956 3316 5958
rect 3340 5956 3396 5958
rect 3420 5956 3476 5958
rect 3054 5616 3110 5672
rect 3180 4922 3236 4924
rect 3260 4922 3316 4924
rect 3340 4922 3396 4924
rect 3420 4922 3476 4924
rect 3180 4870 3226 4922
rect 3226 4870 3236 4922
rect 3260 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3316 4922
rect 3340 4870 3354 4922
rect 3354 4870 3366 4922
rect 3366 4870 3396 4922
rect 3420 4870 3430 4922
rect 3430 4870 3476 4922
rect 3180 4868 3236 4870
rect 3260 4868 3316 4870
rect 3340 4868 3396 4870
rect 3420 4868 3476 4870
rect 2778 3576 2834 3632
rect 1582 992 1638 1048
rect 3180 3834 3236 3836
rect 3260 3834 3316 3836
rect 3340 3834 3396 3836
rect 3420 3834 3476 3836
rect 3180 3782 3226 3834
rect 3226 3782 3236 3834
rect 3260 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3316 3834
rect 3340 3782 3354 3834
rect 3354 3782 3366 3834
rect 3366 3782 3396 3834
rect 3420 3782 3430 3834
rect 3430 3782 3476 3834
rect 3180 3780 3236 3782
rect 3260 3780 3316 3782
rect 3340 3780 3396 3782
rect 3420 3780 3476 3782
rect 3238 3440 3294 3496
rect 3422 3476 3424 3496
rect 3424 3476 3476 3496
rect 3476 3476 3478 3496
rect 3422 3440 3478 3476
rect 2778 1400 2834 1456
rect 3180 2746 3236 2748
rect 3260 2746 3316 2748
rect 3340 2746 3396 2748
rect 3420 2746 3476 2748
rect 3180 2694 3226 2746
rect 3226 2694 3236 2746
rect 3260 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3316 2746
rect 3340 2694 3354 2746
rect 3354 2694 3366 2746
rect 3366 2694 3396 2746
rect 3420 2694 3430 2746
rect 3430 2694 3476 2746
rect 3180 2692 3236 2694
rect 3260 2692 3316 2694
rect 3340 2692 3396 2694
rect 3420 2692 3476 2694
rect 3698 8880 3754 8936
rect 3698 5480 3754 5536
rect 3882 8372 3884 8392
rect 3884 8372 3936 8392
rect 3936 8372 3938 8392
rect 3882 8336 3938 8372
rect 3790 4004 3846 4040
rect 3790 3984 3792 4004
rect 3792 3984 3844 4004
rect 3844 3984 3846 4004
rect 4066 5616 4122 5672
rect 4158 4428 4160 4448
rect 4160 4428 4212 4448
rect 4212 4428 4214 4448
rect 4158 4392 4214 4428
rect 4158 4140 4214 4176
rect 4158 4120 4160 4140
rect 4160 4120 4212 4140
rect 4212 4120 4214 4140
rect 4342 11192 4398 11248
rect 4526 12008 4582 12064
rect 4434 9968 4490 10024
rect 4802 13776 4858 13832
rect 5404 14170 5460 14172
rect 5484 14170 5540 14172
rect 5564 14170 5620 14172
rect 5644 14170 5700 14172
rect 5404 14118 5450 14170
rect 5450 14118 5460 14170
rect 5484 14118 5514 14170
rect 5514 14118 5526 14170
rect 5526 14118 5540 14170
rect 5564 14118 5578 14170
rect 5578 14118 5590 14170
rect 5590 14118 5620 14170
rect 5644 14118 5654 14170
rect 5654 14118 5700 14170
rect 5404 14116 5460 14118
rect 5484 14116 5540 14118
rect 5564 14116 5620 14118
rect 5644 14116 5700 14118
rect 5722 13776 5778 13832
rect 5404 13082 5460 13084
rect 5484 13082 5540 13084
rect 5564 13082 5620 13084
rect 5644 13082 5700 13084
rect 5404 13030 5450 13082
rect 5450 13030 5460 13082
rect 5484 13030 5514 13082
rect 5514 13030 5526 13082
rect 5526 13030 5540 13082
rect 5564 13030 5578 13082
rect 5578 13030 5590 13082
rect 5590 13030 5620 13082
rect 5644 13030 5654 13082
rect 5654 13030 5700 13082
rect 5404 13028 5460 13030
rect 5484 13028 5540 13030
rect 5564 13028 5620 13030
rect 5644 13028 5700 13030
rect 5404 11994 5460 11996
rect 5484 11994 5540 11996
rect 5564 11994 5620 11996
rect 5644 11994 5700 11996
rect 5404 11942 5450 11994
rect 5450 11942 5460 11994
rect 5484 11942 5514 11994
rect 5514 11942 5526 11994
rect 5526 11942 5540 11994
rect 5564 11942 5578 11994
rect 5578 11942 5590 11994
rect 5590 11942 5620 11994
rect 5644 11942 5654 11994
rect 5654 11942 5700 11994
rect 5404 11940 5460 11942
rect 5484 11940 5540 11942
rect 5564 11940 5620 11942
rect 5644 11940 5700 11942
rect 5906 13232 5962 13288
rect 6182 13932 6238 13968
rect 7102 14320 7158 14376
rect 6182 13912 6184 13932
rect 6184 13912 6236 13932
rect 6236 13912 6238 13932
rect 7010 13932 7066 13968
rect 7010 13912 7012 13932
rect 7012 13912 7064 13932
rect 7064 13912 7066 13932
rect 6366 13252 6422 13288
rect 6366 13232 6368 13252
rect 6368 13232 6420 13252
rect 6420 13232 6422 13252
rect 5814 11192 5870 11248
rect 5262 11056 5318 11112
rect 4526 7928 4582 7984
rect 4526 6316 4582 6352
rect 4526 6296 4528 6316
rect 4528 6296 4580 6316
rect 4580 6296 4582 6316
rect 5170 9580 5226 9616
rect 5170 9560 5172 9580
rect 5172 9560 5224 9580
rect 5224 9560 5226 9580
rect 4618 3440 4674 3496
rect 3054 1808 3110 1864
rect 2962 856 3018 912
rect 5404 10906 5460 10908
rect 5484 10906 5540 10908
rect 5564 10906 5620 10908
rect 5644 10906 5700 10908
rect 5404 10854 5450 10906
rect 5450 10854 5460 10906
rect 5484 10854 5514 10906
rect 5514 10854 5526 10906
rect 5526 10854 5540 10906
rect 5564 10854 5578 10906
rect 5578 10854 5590 10906
rect 5590 10854 5620 10906
rect 5644 10854 5654 10906
rect 5654 10854 5700 10906
rect 5404 10852 5460 10854
rect 5484 10852 5540 10854
rect 5564 10852 5620 10854
rect 5644 10852 5700 10854
rect 5404 9818 5460 9820
rect 5484 9818 5540 9820
rect 5564 9818 5620 9820
rect 5644 9818 5700 9820
rect 5404 9766 5450 9818
rect 5450 9766 5460 9818
rect 5484 9766 5514 9818
rect 5514 9766 5526 9818
rect 5526 9766 5540 9818
rect 5564 9766 5578 9818
rect 5578 9766 5590 9818
rect 5590 9766 5620 9818
rect 5644 9766 5654 9818
rect 5654 9766 5700 9818
rect 5404 9764 5460 9766
rect 5484 9764 5540 9766
rect 5564 9764 5620 9766
rect 5644 9764 5700 9766
rect 5906 10668 5962 10704
rect 5906 10648 5908 10668
rect 5908 10648 5960 10668
rect 5960 10648 5962 10668
rect 5722 9016 5778 9072
rect 5404 8730 5460 8732
rect 5484 8730 5540 8732
rect 5564 8730 5620 8732
rect 5644 8730 5700 8732
rect 5404 8678 5450 8730
rect 5450 8678 5460 8730
rect 5484 8678 5514 8730
rect 5514 8678 5526 8730
rect 5526 8678 5540 8730
rect 5564 8678 5578 8730
rect 5578 8678 5590 8730
rect 5590 8678 5620 8730
rect 5644 8678 5654 8730
rect 5654 8678 5700 8730
rect 5404 8676 5460 8678
rect 5484 8676 5540 8678
rect 5564 8676 5620 8678
rect 5644 8676 5700 8678
rect 5078 8472 5134 8528
rect 5262 8472 5318 8528
rect 4894 4528 4950 4584
rect 5404 7642 5460 7644
rect 5484 7642 5540 7644
rect 5564 7642 5620 7644
rect 5644 7642 5700 7644
rect 5404 7590 5450 7642
rect 5450 7590 5460 7642
rect 5484 7590 5514 7642
rect 5514 7590 5526 7642
rect 5526 7590 5540 7642
rect 5564 7590 5578 7642
rect 5578 7590 5590 7642
rect 5590 7590 5620 7642
rect 5644 7590 5654 7642
rect 5654 7590 5700 7642
rect 5404 7588 5460 7590
rect 5484 7588 5540 7590
rect 5564 7588 5620 7590
rect 5644 7588 5700 7590
rect 5404 6554 5460 6556
rect 5484 6554 5540 6556
rect 5564 6554 5620 6556
rect 5644 6554 5700 6556
rect 5404 6502 5450 6554
rect 5450 6502 5460 6554
rect 5484 6502 5514 6554
rect 5514 6502 5526 6554
rect 5526 6502 5540 6554
rect 5564 6502 5578 6554
rect 5578 6502 5590 6554
rect 5590 6502 5620 6554
rect 5644 6502 5654 6554
rect 5654 6502 5700 6554
rect 5404 6500 5460 6502
rect 5484 6500 5540 6502
rect 5564 6500 5620 6502
rect 5644 6500 5700 6502
rect 5404 5466 5460 5468
rect 5484 5466 5540 5468
rect 5564 5466 5620 5468
rect 5644 5466 5700 5468
rect 5404 5414 5450 5466
rect 5450 5414 5460 5466
rect 5484 5414 5514 5466
rect 5514 5414 5526 5466
rect 5526 5414 5540 5466
rect 5564 5414 5578 5466
rect 5578 5414 5590 5466
rect 5590 5414 5620 5466
rect 5644 5414 5654 5466
rect 5654 5414 5700 5466
rect 5404 5412 5460 5414
rect 5484 5412 5540 5414
rect 5564 5412 5620 5414
rect 5644 5412 5700 5414
rect 5906 5616 5962 5672
rect 5404 4378 5460 4380
rect 5484 4378 5540 4380
rect 5564 4378 5620 4380
rect 5644 4378 5700 4380
rect 5404 4326 5450 4378
rect 5450 4326 5460 4378
rect 5484 4326 5514 4378
rect 5514 4326 5526 4378
rect 5526 4326 5540 4378
rect 5564 4326 5578 4378
rect 5578 4326 5590 4378
rect 5590 4326 5620 4378
rect 5644 4326 5654 4378
rect 5654 4326 5700 4378
rect 5404 4324 5460 4326
rect 5484 4324 5540 4326
rect 5564 4324 5620 4326
rect 5644 4324 5700 4326
rect 5906 3576 5962 3632
rect 5078 3304 5134 3360
rect 5262 3304 5318 3360
rect 5404 3290 5460 3292
rect 5484 3290 5540 3292
rect 5564 3290 5620 3292
rect 5644 3290 5700 3292
rect 5404 3238 5450 3290
rect 5450 3238 5460 3290
rect 5484 3238 5514 3290
rect 5514 3238 5526 3290
rect 5526 3238 5540 3290
rect 5564 3238 5578 3290
rect 5578 3238 5590 3290
rect 5590 3238 5620 3290
rect 5644 3238 5654 3290
rect 5654 3238 5700 3290
rect 5404 3236 5460 3238
rect 5484 3236 5540 3238
rect 5564 3236 5620 3238
rect 5644 3236 5700 3238
rect 5906 2932 5908 2952
rect 5908 2932 5960 2952
rect 5960 2932 5962 2952
rect 5906 2896 5962 2932
rect 6550 5072 6606 5128
rect 6458 2896 6514 2952
rect 6826 9016 6882 9072
rect 6734 8744 6790 8800
rect 6826 8608 6882 8664
rect 7628 14714 7684 14716
rect 7708 14714 7764 14716
rect 7788 14714 7844 14716
rect 7868 14714 7924 14716
rect 7628 14662 7674 14714
rect 7674 14662 7684 14714
rect 7708 14662 7738 14714
rect 7738 14662 7750 14714
rect 7750 14662 7764 14714
rect 7788 14662 7802 14714
rect 7802 14662 7814 14714
rect 7814 14662 7844 14714
rect 7868 14662 7878 14714
rect 7878 14662 7924 14714
rect 7628 14660 7684 14662
rect 7708 14660 7764 14662
rect 7788 14660 7844 14662
rect 7868 14660 7924 14662
rect 7628 13626 7684 13628
rect 7708 13626 7764 13628
rect 7788 13626 7844 13628
rect 7868 13626 7924 13628
rect 7628 13574 7674 13626
rect 7674 13574 7684 13626
rect 7708 13574 7738 13626
rect 7738 13574 7750 13626
rect 7750 13574 7764 13626
rect 7788 13574 7802 13626
rect 7802 13574 7814 13626
rect 7814 13574 7844 13626
rect 7868 13574 7878 13626
rect 7878 13574 7924 13626
rect 7628 13572 7684 13574
rect 7708 13572 7764 13574
rect 7788 13572 7844 13574
rect 7868 13572 7924 13574
rect 7628 12538 7684 12540
rect 7708 12538 7764 12540
rect 7788 12538 7844 12540
rect 7868 12538 7924 12540
rect 7628 12486 7674 12538
rect 7674 12486 7684 12538
rect 7708 12486 7738 12538
rect 7738 12486 7750 12538
rect 7750 12486 7764 12538
rect 7788 12486 7802 12538
rect 7802 12486 7814 12538
rect 7814 12486 7844 12538
rect 7868 12486 7878 12538
rect 7878 12486 7924 12538
rect 7628 12484 7684 12486
rect 7708 12484 7764 12486
rect 7788 12484 7844 12486
rect 7868 12484 7924 12486
rect 7628 11450 7684 11452
rect 7708 11450 7764 11452
rect 7788 11450 7844 11452
rect 7868 11450 7924 11452
rect 7628 11398 7674 11450
rect 7674 11398 7684 11450
rect 7708 11398 7738 11450
rect 7738 11398 7750 11450
rect 7750 11398 7764 11450
rect 7788 11398 7802 11450
rect 7802 11398 7814 11450
rect 7814 11398 7844 11450
rect 7868 11398 7878 11450
rect 7878 11398 7924 11450
rect 7628 11396 7684 11398
rect 7708 11396 7764 11398
rect 7788 11396 7844 11398
rect 7868 11396 7924 11398
rect 7628 10362 7684 10364
rect 7708 10362 7764 10364
rect 7788 10362 7844 10364
rect 7868 10362 7924 10364
rect 7628 10310 7674 10362
rect 7674 10310 7684 10362
rect 7708 10310 7738 10362
rect 7738 10310 7750 10362
rect 7750 10310 7764 10362
rect 7788 10310 7802 10362
rect 7802 10310 7814 10362
rect 7814 10310 7844 10362
rect 7868 10310 7878 10362
rect 7878 10310 7924 10362
rect 7628 10308 7684 10310
rect 7708 10308 7764 10310
rect 7788 10308 7844 10310
rect 7868 10308 7924 10310
rect 7628 9274 7684 9276
rect 7708 9274 7764 9276
rect 7788 9274 7844 9276
rect 7868 9274 7924 9276
rect 7628 9222 7674 9274
rect 7674 9222 7684 9274
rect 7708 9222 7738 9274
rect 7738 9222 7750 9274
rect 7750 9222 7764 9274
rect 7788 9222 7802 9274
rect 7802 9222 7814 9274
rect 7814 9222 7844 9274
rect 7868 9222 7878 9274
rect 7878 9222 7924 9274
rect 7628 9220 7684 9222
rect 7708 9220 7764 9222
rect 7788 9220 7844 9222
rect 7868 9220 7924 9222
rect 8206 14492 8208 14512
rect 8208 14492 8260 14512
rect 8260 14492 8262 14512
rect 8206 14456 8262 14492
rect 8206 8744 8262 8800
rect 8114 8628 8170 8664
rect 8114 8608 8116 8628
rect 8116 8608 8168 8628
rect 8168 8608 8170 8628
rect 8482 11464 8538 11520
rect 8298 8608 8354 8664
rect 7628 8186 7684 8188
rect 7708 8186 7764 8188
rect 7788 8186 7844 8188
rect 7868 8186 7924 8188
rect 7628 8134 7674 8186
rect 7674 8134 7684 8186
rect 7708 8134 7738 8186
rect 7738 8134 7750 8186
rect 7750 8134 7764 8186
rect 7788 8134 7802 8186
rect 7802 8134 7814 8186
rect 7814 8134 7844 8186
rect 7868 8134 7878 8186
rect 7878 8134 7924 8186
rect 7628 8132 7684 8134
rect 7708 8132 7764 8134
rect 7788 8132 7844 8134
rect 7868 8132 7924 8134
rect 8758 8780 8760 8800
rect 8760 8780 8812 8800
rect 8812 8780 8814 8800
rect 8758 8744 8814 8780
rect 8206 7928 8262 7984
rect 7628 7098 7684 7100
rect 7708 7098 7764 7100
rect 7788 7098 7844 7100
rect 7868 7098 7924 7100
rect 7628 7046 7674 7098
rect 7674 7046 7684 7098
rect 7708 7046 7738 7098
rect 7738 7046 7750 7098
rect 7750 7046 7764 7098
rect 7788 7046 7802 7098
rect 7802 7046 7814 7098
rect 7814 7046 7844 7098
rect 7868 7046 7878 7098
rect 7878 7046 7924 7098
rect 7628 7044 7684 7046
rect 7708 7044 7764 7046
rect 7788 7044 7844 7046
rect 7868 7044 7924 7046
rect 7194 5208 7250 5264
rect 7654 6704 7710 6760
rect 7746 6296 7802 6352
rect 7470 6160 7526 6216
rect 7628 6010 7684 6012
rect 7708 6010 7764 6012
rect 7788 6010 7844 6012
rect 7868 6010 7924 6012
rect 7628 5958 7674 6010
rect 7674 5958 7684 6010
rect 7708 5958 7738 6010
rect 7738 5958 7750 6010
rect 7750 5958 7764 6010
rect 7788 5958 7802 6010
rect 7802 5958 7814 6010
rect 7814 5958 7844 6010
rect 7868 5958 7878 6010
rect 7878 5958 7924 6010
rect 7628 5956 7684 5958
rect 7708 5956 7764 5958
rect 7788 5956 7844 5958
rect 7868 5956 7924 5958
rect 7654 5208 7710 5264
rect 7286 4120 7342 4176
rect 7286 3440 7342 3496
rect 7628 4922 7684 4924
rect 7708 4922 7764 4924
rect 7788 4922 7844 4924
rect 7868 4922 7924 4924
rect 7628 4870 7674 4922
rect 7674 4870 7684 4922
rect 7708 4870 7738 4922
rect 7738 4870 7750 4922
rect 7750 4870 7764 4922
rect 7788 4870 7802 4922
rect 7802 4870 7814 4922
rect 7814 4870 7844 4922
rect 7868 4870 7878 4922
rect 7878 4870 7924 4922
rect 7628 4868 7684 4870
rect 7708 4868 7764 4870
rect 7788 4868 7844 4870
rect 7868 4868 7924 4870
rect 8206 6296 8262 6352
rect 7628 3834 7684 3836
rect 7708 3834 7764 3836
rect 7788 3834 7844 3836
rect 7868 3834 7924 3836
rect 7628 3782 7674 3834
rect 7674 3782 7684 3834
rect 7708 3782 7738 3834
rect 7738 3782 7750 3834
rect 7750 3782 7764 3834
rect 7788 3782 7802 3834
rect 7802 3782 7814 3834
rect 7814 3782 7844 3834
rect 7868 3782 7878 3834
rect 7878 3782 7924 3834
rect 7628 3780 7684 3782
rect 7708 3780 7764 3782
rect 7788 3780 7844 3782
rect 7868 3780 7924 3782
rect 12076 14714 12132 14716
rect 12156 14714 12212 14716
rect 12236 14714 12292 14716
rect 12316 14714 12372 14716
rect 12076 14662 12122 14714
rect 12122 14662 12132 14714
rect 12156 14662 12186 14714
rect 12186 14662 12198 14714
rect 12198 14662 12212 14714
rect 12236 14662 12250 14714
rect 12250 14662 12262 14714
rect 12262 14662 12292 14714
rect 12316 14662 12326 14714
rect 12326 14662 12372 14714
rect 12076 14660 12132 14662
rect 12156 14660 12212 14662
rect 12236 14660 12292 14662
rect 12316 14660 12372 14662
rect 9126 9016 9182 9072
rect 9126 5480 9182 5536
rect 7628 2746 7684 2748
rect 7708 2746 7764 2748
rect 7788 2746 7844 2748
rect 7868 2746 7924 2748
rect 7628 2694 7674 2746
rect 7674 2694 7684 2746
rect 7708 2694 7738 2746
rect 7738 2694 7750 2746
rect 7750 2694 7764 2746
rect 7788 2694 7802 2746
rect 7802 2694 7814 2746
rect 7814 2694 7844 2746
rect 7868 2694 7878 2746
rect 7878 2694 7924 2746
rect 7628 2692 7684 2694
rect 7708 2692 7764 2694
rect 7788 2692 7844 2694
rect 7868 2692 7924 2694
rect 9310 8780 9312 8800
rect 9312 8780 9364 8800
rect 9364 8780 9366 8800
rect 9310 8744 9366 8780
rect 9494 8608 9550 8664
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9898 14170
rect 9898 14118 9908 14170
rect 9932 14118 9962 14170
rect 9962 14118 9974 14170
rect 9974 14118 9988 14170
rect 10012 14118 10026 14170
rect 10026 14118 10038 14170
rect 10038 14118 10068 14170
rect 10092 14118 10102 14170
rect 10102 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9898 13082
rect 9898 13030 9908 13082
rect 9932 13030 9962 13082
rect 9962 13030 9974 13082
rect 9974 13030 9988 13082
rect 10012 13030 10026 13082
rect 10026 13030 10038 13082
rect 10038 13030 10068 13082
rect 10092 13030 10102 13082
rect 10102 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9898 11994
rect 9898 11942 9908 11994
rect 9932 11942 9962 11994
rect 9962 11942 9974 11994
rect 9974 11942 9988 11994
rect 10012 11942 10026 11994
rect 10026 11942 10038 11994
rect 10038 11942 10068 11994
rect 10092 11942 10102 11994
rect 10102 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9898 10906
rect 9898 10854 9908 10906
rect 9932 10854 9962 10906
rect 9962 10854 9974 10906
rect 9974 10854 9988 10906
rect 10012 10854 10026 10906
rect 10026 10854 10038 10906
rect 10038 10854 10068 10906
rect 10092 10854 10102 10906
rect 10102 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 10414 11056 10470 11112
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9898 9818
rect 9898 9766 9908 9818
rect 9932 9766 9962 9818
rect 9962 9766 9974 9818
rect 9974 9766 9988 9818
rect 10012 9766 10026 9818
rect 10026 9766 10038 9818
rect 10038 9766 10068 9818
rect 10092 9766 10102 9818
rect 10102 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9898 8730
rect 9898 8678 9908 8730
rect 9932 8678 9962 8730
rect 9962 8678 9974 8730
rect 9974 8678 9988 8730
rect 10012 8678 10026 8730
rect 10026 8678 10038 8730
rect 10038 8678 10068 8730
rect 10092 8678 10102 8730
rect 10102 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 9678 7928 9734 7984
rect 10046 7964 10048 7984
rect 10048 7964 10100 7984
rect 10100 7964 10102 7984
rect 10046 7928 10102 7964
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9898 7642
rect 9898 7590 9908 7642
rect 9932 7590 9962 7642
rect 9962 7590 9974 7642
rect 9974 7590 9988 7642
rect 10012 7590 10026 7642
rect 10026 7590 10038 7642
rect 10038 7590 10068 7642
rect 10092 7590 10102 7642
rect 10102 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9898 6554
rect 9898 6502 9908 6554
rect 9932 6502 9962 6554
rect 9962 6502 9974 6554
rect 9974 6502 9988 6554
rect 10012 6502 10026 6554
rect 10026 6502 10038 6554
rect 10038 6502 10068 6554
rect 10092 6502 10102 6554
rect 10102 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 10414 9424 10470 9480
rect 9678 5480 9734 5536
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9898 5466
rect 9898 5414 9908 5466
rect 9932 5414 9962 5466
rect 9962 5414 9974 5466
rect 9974 5414 9988 5466
rect 10012 5414 10026 5466
rect 10026 5414 10038 5466
rect 10038 5414 10068 5466
rect 10092 5414 10102 5466
rect 10102 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9898 4378
rect 9898 4326 9908 4378
rect 9932 4326 9962 4378
rect 9962 4326 9974 4378
rect 9974 4326 9988 4378
rect 10012 4326 10026 4378
rect 10026 4326 10038 4378
rect 10038 4326 10068 4378
rect 10092 4326 10102 4378
rect 10102 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 10874 11056 10930 11112
rect 11150 11600 11206 11656
rect 11242 10648 11298 10704
rect 11150 9444 11206 9480
rect 11150 9424 11152 9444
rect 11152 9424 11204 9444
rect 11204 9424 11206 9444
rect 11610 9988 11666 10024
rect 11610 9968 11612 9988
rect 11612 9968 11664 9988
rect 11664 9968 11666 9988
rect 12076 13626 12132 13628
rect 12156 13626 12212 13628
rect 12236 13626 12292 13628
rect 12316 13626 12372 13628
rect 12076 13574 12122 13626
rect 12122 13574 12132 13626
rect 12156 13574 12186 13626
rect 12186 13574 12198 13626
rect 12198 13574 12212 13626
rect 12236 13574 12250 13626
rect 12250 13574 12262 13626
rect 12262 13574 12292 13626
rect 12316 13574 12326 13626
rect 12326 13574 12372 13626
rect 12076 13572 12132 13574
rect 12156 13572 12212 13574
rect 12236 13572 12292 13574
rect 12316 13572 12372 13574
rect 12076 12538 12132 12540
rect 12156 12538 12212 12540
rect 12236 12538 12292 12540
rect 12316 12538 12372 12540
rect 12076 12486 12122 12538
rect 12122 12486 12132 12538
rect 12156 12486 12186 12538
rect 12186 12486 12198 12538
rect 12198 12486 12212 12538
rect 12236 12486 12250 12538
rect 12250 12486 12262 12538
rect 12262 12486 12292 12538
rect 12316 12486 12326 12538
rect 12326 12486 12372 12538
rect 12076 12484 12132 12486
rect 12156 12484 12212 12486
rect 12236 12484 12292 12486
rect 12316 12484 12372 12486
rect 11518 8608 11574 8664
rect 11242 7792 11298 7848
rect 11518 6840 11574 6896
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9898 3290
rect 9898 3238 9908 3290
rect 9932 3238 9962 3290
rect 9962 3238 9974 3290
rect 9974 3238 9988 3290
rect 10012 3238 10026 3290
rect 10026 3238 10038 3290
rect 10038 3238 10068 3290
rect 10092 3238 10102 3290
rect 10102 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 5404 2202 5460 2204
rect 5484 2202 5540 2204
rect 5564 2202 5620 2204
rect 5644 2202 5700 2204
rect 5404 2150 5450 2202
rect 5450 2150 5460 2202
rect 5484 2150 5514 2202
rect 5514 2150 5526 2202
rect 5526 2150 5540 2202
rect 5564 2150 5578 2202
rect 5578 2150 5590 2202
rect 5590 2150 5620 2202
rect 5644 2150 5654 2202
rect 5654 2150 5700 2202
rect 5404 2148 5460 2150
rect 5484 2148 5540 2150
rect 5564 2148 5620 2150
rect 5644 2148 5700 2150
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9898 2202
rect 9898 2150 9908 2202
rect 9932 2150 9962 2202
rect 9962 2150 9974 2202
rect 9974 2150 9988 2202
rect 10012 2150 10026 2202
rect 10026 2150 10038 2202
rect 10038 2150 10068 2202
rect 10092 2150 10102 2202
rect 10102 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 11058 4664 11114 4720
rect 10874 4120 10930 4176
rect 11242 4528 11298 4584
rect 11518 4020 11520 4040
rect 11520 4020 11572 4040
rect 11572 4020 11574 4040
rect 11518 3984 11574 4020
rect 14300 14170 14356 14172
rect 14380 14170 14436 14172
rect 14460 14170 14516 14172
rect 14540 14170 14596 14172
rect 14300 14118 14346 14170
rect 14346 14118 14356 14170
rect 14380 14118 14410 14170
rect 14410 14118 14422 14170
rect 14422 14118 14436 14170
rect 14460 14118 14474 14170
rect 14474 14118 14486 14170
rect 14486 14118 14516 14170
rect 14540 14118 14550 14170
rect 14550 14118 14596 14170
rect 14300 14116 14356 14118
rect 14380 14116 14436 14118
rect 14460 14116 14516 14118
rect 14540 14116 14596 14118
rect 14094 13368 14150 13424
rect 12076 11450 12132 11452
rect 12156 11450 12212 11452
rect 12236 11450 12292 11452
rect 12316 11450 12372 11452
rect 12076 11398 12122 11450
rect 12122 11398 12132 11450
rect 12156 11398 12186 11450
rect 12186 11398 12198 11450
rect 12198 11398 12212 11450
rect 12236 11398 12250 11450
rect 12250 11398 12262 11450
rect 12262 11398 12292 11450
rect 12316 11398 12326 11450
rect 12326 11398 12372 11450
rect 12076 11396 12132 11398
rect 12156 11396 12212 11398
rect 12236 11396 12292 11398
rect 12316 11396 12372 11398
rect 12076 10362 12132 10364
rect 12156 10362 12212 10364
rect 12236 10362 12292 10364
rect 12316 10362 12372 10364
rect 12076 10310 12122 10362
rect 12122 10310 12132 10362
rect 12156 10310 12186 10362
rect 12186 10310 12198 10362
rect 12198 10310 12212 10362
rect 12236 10310 12250 10362
rect 12250 10310 12262 10362
rect 12262 10310 12292 10362
rect 12316 10310 12326 10362
rect 12326 10310 12372 10362
rect 12076 10308 12132 10310
rect 12156 10308 12212 10310
rect 12236 10308 12292 10310
rect 12316 10308 12372 10310
rect 12076 9274 12132 9276
rect 12156 9274 12212 9276
rect 12236 9274 12292 9276
rect 12316 9274 12372 9276
rect 12076 9222 12122 9274
rect 12122 9222 12132 9274
rect 12156 9222 12186 9274
rect 12186 9222 12198 9274
rect 12198 9222 12212 9274
rect 12236 9222 12250 9274
rect 12250 9222 12262 9274
rect 12262 9222 12292 9274
rect 12316 9222 12326 9274
rect 12326 9222 12372 9274
rect 12076 9220 12132 9222
rect 12156 9220 12212 9222
rect 12236 9220 12292 9222
rect 12316 9220 12372 9222
rect 12530 9172 12586 9208
rect 12806 9324 12808 9344
rect 12808 9324 12860 9344
rect 12860 9324 12862 9344
rect 12806 9288 12862 9324
rect 12530 9152 12532 9172
rect 12532 9152 12584 9172
rect 12584 9152 12586 9172
rect 12898 9152 12954 9208
rect 11978 8744 12034 8800
rect 11978 8492 12034 8528
rect 11978 8472 11980 8492
rect 11980 8472 12032 8492
rect 12032 8472 12034 8492
rect 12076 8186 12132 8188
rect 12156 8186 12212 8188
rect 12236 8186 12292 8188
rect 12316 8186 12372 8188
rect 12076 8134 12122 8186
rect 12122 8134 12132 8186
rect 12156 8134 12186 8186
rect 12186 8134 12198 8186
rect 12198 8134 12212 8186
rect 12236 8134 12250 8186
rect 12250 8134 12262 8186
rect 12262 8134 12292 8186
rect 12316 8134 12326 8186
rect 12326 8134 12372 8186
rect 12076 8132 12132 8134
rect 12156 8132 12212 8134
rect 12236 8132 12292 8134
rect 12316 8132 12372 8134
rect 11978 7792 12034 7848
rect 12076 7098 12132 7100
rect 12156 7098 12212 7100
rect 12236 7098 12292 7100
rect 12316 7098 12372 7100
rect 12076 7046 12122 7098
rect 12122 7046 12132 7098
rect 12156 7046 12186 7098
rect 12186 7046 12198 7098
rect 12198 7046 12212 7098
rect 12236 7046 12250 7098
rect 12250 7046 12262 7098
rect 12262 7046 12292 7098
rect 12316 7046 12326 7098
rect 12326 7046 12372 7098
rect 12076 7044 12132 7046
rect 12156 7044 12212 7046
rect 12236 7044 12292 7046
rect 12316 7044 12372 7046
rect 12076 6010 12132 6012
rect 12156 6010 12212 6012
rect 12236 6010 12292 6012
rect 12316 6010 12372 6012
rect 12076 5958 12122 6010
rect 12122 5958 12132 6010
rect 12156 5958 12186 6010
rect 12186 5958 12198 6010
rect 12198 5958 12212 6010
rect 12236 5958 12250 6010
rect 12250 5958 12262 6010
rect 12262 5958 12292 6010
rect 12316 5958 12326 6010
rect 12326 5958 12372 6010
rect 12076 5956 12132 5958
rect 12156 5956 12212 5958
rect 12236 5956 12292 5958
rect 12316 5956 12372 5958
rect 13358 9968 13414 10024
rect 13542 9152 13598 9208
rect 13726 8744 13782 8800
rect 13818 8608 13874 8664
rect 13358 7928 13414 7984
rect 13266 7248 13322 7304
rect 13082 5616 13138 5672
rect 12076 4922 12132 4924
rect 12156 4922 12212 4924
rect 12236 4922 12292 4924
rect 12316 4922 12372 4924
rect 12076 4870 12122 4922
rect 12122 4870 12132 4922
rect 12156 4870 12186 4922
rect 12186 4870 12198 4922
rect 12198 4870 12212 4922
rect 12236 4870 12250 4922
rect 12250 4870 12262 4922
rect 12262 4870 12292 4922
rect 12316 4870 12326 4922
rect 12326 4870 12372 4922
rect 12076 4868 12132 4870
rect 12156 4868 12212 4870
rect 12236 4868 12292 4870
rect 12316 4868 12372 4870
rect 11978 4256 12034 4312
rect 12990 5072 13046 5128
rect 12076 3834 12132 3836
rect 12156 3834 12212 3836
rect 12236 3834 12292 3836
rect 12316 3834 12372 3836
rect 12076 3782 12122 3834
rect 12122 3782 12132 3834
rect 12156 3782 12186 3834
rect 12186 3782 12198 3834
rect 12198 3782 12212 3834
rect 12236 3782 12250 3834
rect 12250 3782 12262 3834
rect 12262 3782 12292 3834
rect 12316 3782 12326 3834
rect 12326 3782 12372 3834
rect 12076 3780 12132 3782
rect 12156 3780 12212 3782
rect 12236 3780 12292 3782
rect 12316 3780 12372 3782
rect 12438 3304 12494 3360
rect 12076 2746 12132 2748
rect 12156 2746 12212 2748
rect 12236 2746 12292 2748
rect 12316 2746 12372 2748
rect 12076 2694 12122 2746
rect 12122 2694 12132 2746
rect 12156 2694 12186 2746
rect 12186 2694 12198 2746
rect 12198 2694 12212 2746
rect 12236 2694 12250 2746
rect 12250 2694 12262 2746
rect 12262 2694 12292 2746
rect 12316 2694 12326 2746
rect 12326 2694 12372 2746
rect 12076 2692 12132 2694
rect 12156 2692 12212 2694
rect 12236 2692 12292 2694
rect 12316 2692 12372 2694
rect 12714 3984 12770 4040
rect 12714 3884 12716 3904
rect 12716 3884 12768 3904
rect 12768 3884 12770 3904
rect 12714 3848 12770 3884
rect 13450 5480 13506 5536
rect 13726 6840 13782 6896
rect 14300 13082 14356 13084
rect 14380 13082 14436 13084
rect 14460 13082 14516 13084
rect 14540 13082 14596 13084
rect 14300 13030 14346 13082
rect 14346 13030 14356 13082
rect 14380 13030 14410 13082
rect 14410 13030 14422 13082
rect 14422 13030 14436 13082
rect 14460 13030 14474 13082
rect 14474 13030 14486 13082
rect 14486 13030 14516 13082
rect 14540 13030 14550 13082
rect 14550 13030 14596 13082
rect 14300 13028 14356 13030
rect 14380 13028 14436 13030
rect 14460 13028 14516 13030
rect 14540 13028 14596 13030
rect 14300 11994 14356 11996
rect 14380 11994 14436 11996
rect 14460 11994 14516 11996
rect 14540 11994 14596 11996
rect 14300 11942 14346 11994
rect 14346 11942 14356 11994
rect 14380 11942 14410 11994
rect 14410 11942 14422 11994
rect 14422 11942 14436 11994
rect 14460 11942 14474 11994
rect 14474 11942 14486 11994
rect 14486 11942 14516 11994
rect 14540 11942 14550 11994
rect 14550 11942 14596 11994
rect 14300 11940 14356 11942
rect 14380 11940 14436 11942
rect 14460 11940 14516 11942
rect 14540 11940 14596 11942
rect 13726 5752 13782 5808
rect 13358 3984 13414 4040
rect 13726 4256 13782 4312
rect 13634 3984 13690 4040
rect 13634 3712 13690 3768
rect 14300 10906 14356 10908
rect 14380 10906 14436 10908
rect 14460 10906 14516 10908
rect 14540 10906 14596 10908
rect 14300 10854 14346 10906
rect 14346 10854 14356 10906
rect 14380 10854 14410 10906
rect 14410 10854 14422 10906
rect 14422 10854 14436 10906
rect 14460 10854 14474 10906
rect 14474 10854 14486 10906
rect 14486 10854 14516 10906
rect 14540 10854 14550 10906
rect 14550 10854 14596 10906
rect 14300 10852 14356 10854
rect 14380 10852 14436 10854
rect 14460 10852 14516 10854
rect 14540 10852 14596 10854
rect 14300 9818 14356 9820
rect 14380 9818 14436 9820
rect 14460 9818 14516 9820
rect 14540 9818 14596 9820
rect 14300 9766 14346 9818
rect 14346 9766 14356 9818
rect 14380 9766 14410 9818
rect 14410 9766 14422 9818
rect 14422 9766 14436 9818
rect 14460 9766 14474 9818
rect 14474 9766 14486 9818
rect 14486 9766 14516 9818
rect 14540 9766 14550 9818
rect 14550 9766 14596 9818
rect 14300 9764 14356 9766
rect 14380 9764 14436 9766
rect 14460 9764 14516 9766
rect 14540 9764 14596 9766
rect 14300 8730 14356 8732
rect 14380 8730 14436 8732
rect 14460 8730 14516 8732
rect 14540 8730 14596 8732
rect 14300 8678 14346 8730
rect 14346 8678 14356 8730
rect 14380 8678 14410 8730
rect 14410 8678 14422 8730
rect 14422 8678 14436 8730
rect 14460 8678 14474 8730
rect 14474 8678 14486 8730
rect 14486 8678 14516 8730
rect 14540 8678 14550 8730
rect 14550 8678 14596 8730
rect 14300 8676 14356 8678
rect 14380 8676 14436 8678
rect 14460 8676 14516 8678
rect 14540 8676 14596 8678
rect 14554 7928 14610 7984
rect 14300 7642 14356 7644
rect 14380 7642 14436 7644
rect 14460 7642 14516 7644
rect 14540 7642 14596 7644
rect 14300 7590 14346 7642
rect 14346 7590 14356 7642
rect 14380 7590 14410 7642
rect 14410 7590 14422 7642
rect 14422 7590 14436 7642
rect 14460 7590 14474 7642
rect 14474 7590 14486 7642
rect 14486 7590 14516 7642
rect 14540 7590 14550 7642
rect 14550 7590 14596 7642
rect 14300 7588 14356 7590
rect 14380 7588 14436 7590
rect 14460 7588 14516 7590
rect 14540 7588 14596 7590
rect 14300 6554 14356 6556
rect 14380 6554 14436 6556
rect 14460 6554 14516 6556
rect 14540 6554 14596 6556
rect 14300 6502 14346 6554
rect 14346 6502 14356 6554
rect 14380 6502 14410 6554
rect 14410 6502 14422 6554
rect 14422 6502 14436 6554
rect 14460 6502 14474 6554
rect 14474 6502 14486 6554
rect 14486 6502 14516 6554
rect 14540 6502 14550 6554
rect 14550 6502 14596 6554
rect 14300 6500 14356 6502
rect 14380 6500 14436 6502
rect 14460 6500 14516 6502
rect 14540 6500 14596 6502
rect 14300 5466 14356 5468
rect 14380 5466 14436 5468
rect 14460 5466 14516 5468
rect 14540 5466 14596 5468
rect 14300 5414 14346 5466
rect 14346 5414 14356 5466
rect 14380 5414 14410 5466
rect 14410 5414 14422 5466
rect 14422 5414 14436 5466
rect 14460 5414 14474 5466
rect 14474 5414 14486 5466
rect 14486 5414 14516 5466
rect 14540 5414 14550 5466
rect 14550 5414 14596 5466
rect 14300 5412 14356 5414
rect 14380 5412 14436 5414
rect 14460 5412 14516 5414
rect 14540 5412 14596 5414
rect 13818 3848 13874 3904
rect 13542 3476 13544 3496
rect 13544 3476 13596 3496
rect 13596 3476 13598 3496
rect 13542 3440 13598 3476
rect 14300 4378 14356 4380
rect 14380 4378 14436 4380
rect 14460 4378 14516 4380
rect 14540 4378 14596 4380
rect 14300 4326 14346 4378
rect 14346 4326 14356 4378
rect 14380 4326 14410 4378
rect 14410 4326 14422 4378
rect 14422 4326 14436 4378
rect 14460 4326 14474 4378
rect 14474 4326 14486 4378
rect 14486 4326 14516 4378
rect 14540 4326 14550 4378
rect 14550 4326 14596 4378
rect 14300 4324 14356 4326
rect 14380 4324 14436 4326
rect 14460 4324 14516 4326
rect 14540 4324 14596 4326
rect 14830 8200 14886 8256
rect 14830 7928 14886 7984
rect 14094 3984 14150 4040
rect 14300 3290 14356 3292
rect 14380 3290 14436 3292
rect 14460 3290 14516 3292
rect 14540 3290 14596 3292
rect 14300 3238 14346 3290
rect 14346 3238 14356 3290
rect 14380 3238 14410 3290
rect 14410 3238 14422 3290
rect 14422 3238 14436 3290
rect 14460 3238 14474 3290
rect 14474 3238 14486 3290
rect 14486 3238 14516 3290
rect 14540 3238 14550 3290
rect 14550 3238 14596 3290
rect 14300 3236 14356 3238
rect 14380 3236 14436 3238
rect 14460 3236 14516 3238
rect 14540 3236 14596 3238
rect 14300 2202 14356 2204
rect 14380 2202 14436 2204
rect 14460 2202 14516 2204
rect 14540 2202 14596 2204
rect 14300 2150 14346 2202
rect 14346 2150 14356 2202
rect 14380 2150 14410 2202
rect 14410 2150 14422 2202
rect 14422 2150 14436 2202
rect 14460 2150 14474 2202
rect 14474 2150 14486 2202
rect 14486 2150 14516 2202
rect 14540 2150 14550 2202
rect 14550 2150 14596 2202
rect 14300 2148 14356 2150
rect 14380 2148 14436 2150
rect 14460 2148 14516 2150
rect 14540 2148 14596 2150
rect 3882 176 3938 232
rect 15106 12416 15162 12472
rect 15198 10648 15254 10704
rect 15198 10532 15254 10568
rect 15198 10512 15200 10532
rect 15200 10512 15252 10532
rect 15252 10512 15254 10532
rect 15198 8880 15254 8936
rect 15290 7792 15346 7848
rect 15106 3984 15162 4040
rect 15290 6160 15346 6216
rect 16118 16768 16174 16824
rect 16302 16360 16358 16416
rect 16118 15544 16174 15600
rect 16210 15136 16266 15192
rect 15474 9288 15530 9344
rect 15566 8880 15622 8936
rect 15934 11056 15990 11112
rect 15842 9016 15898 9072
rect 15934 8744 15990 8800
rect 15750 7792 15806 7848
rect 15382 5344 15438 5400
rect 15566 3984 15622 4040
rect 15750 3032 15806 3088
rect 15934 5208 15990 5264
rect 16394 15952 16450 16008
rect 16524 14714 16580 14716
rect 16604 14714 16660 14716
rect 16684 14714 16740 14716
rect 16764 14714 16820 14716
rect 16524 14662 16570 14714
rect 16570 14662 16580 14714
rect 16604 14662 16634 14714
rect 16634 14662 16646 14714
rect 16646 14662 16660 14714
rect 16684 14662 16698 14714
rect 16698 14662 16710 14714
rect 16710 14662 16740 14714
rect 16764 14662 16774 14714
rect 16774 14662 16820 14714
rect 16524 14660 16580 14662
rect 16604 14660 16660 14662
rect 16684 14660 16740 14662
rect 16764 14660 16820 14662
rect 16524 13626 16580 13628
rect 16604 13626 16660 13628
rect 16684 13626 16740 13628
rect 16764 13626 16820 13628
rect 16524 13574 16570 13626
rect 16570 13574 16580 13626
rect 16604 13574 16634 13626
rect 16634 13574 16646 13626
rect 16646 13574 16660 13626
rect 16684 13574 16698 13626
rect 16698 13574 16710 13626
rect 16710 13574 16740 13626
rect 16764 13574 16774 13626
rect 16774 13574 16820 13626
rect 16524 13572 16580 13574
rect 16604 13572 16660 13574
rect 16684 13572 16740 13574
rect 16764 13572 16820 13574
rect 17038 13812 17040 13832
rect 17040 13812 17092 13832
rect 17092 13812 17094 13832
rect 17038 13776 17094 13812
rect 16524 12538 16580 12540
rect 16604 12538 16660 12540
rect 16684 12538 16740 12540
rect 16764 12538 16820 12540
rect 16524 12486 16570 12538
rect 16570 12486 16580 12538
rect 16604 12486 16634 12538
rect 16634 12486 16646 12538
rect 16646 12486 16660 12538
rect 16684 12486 16698 12538
rect 16698 12486 16710 12538
rect 16710 12486 16740 12538
rect 16764 12486 16774 12538
rect 16774 12486 16820 12538
rect 16524 12484 16580 12486
rect 16604 12484 16660 12486
rect 16684 12484 16740 12486
rect 16764 12484 16820 12486
rect 16524 11450 16580 11452
rect 16604 11450 16660 11452
rect 16684 11450 16740 11452
rect 16764 11450 16820 11452
rect 16524 11398 16570 11450
rect 16570 11398 16580 11450
rect 16604 11398 16634 11450
rect 16634 11398 16646 11450
rect 16646 11398 16660 11450
rect 16684 11398 16698 11450
rect 16698 11398 16710 11450
rect 16710 11398 16740 11450
rect 16764 11398 16774 11450
rect 16774 11398 16820 11450
rect 16524 11396 16580 11398
rect 16604 11396 16660 11398
rect 16684 11396 16740 11398
rect 16764 11396 16820 11398
rect 16118 8608 16174 8664
rect 17406 14728 17462 14784
rect 17498 13776 17554 13832
rect 17314 12688 17370 12744
rect 17682 14184 17738 14240
rect 17682 13368 17738 13424
rect 17682 12960 17738 13016
rect 17682 12552 17738 12608
rect 16670 10956 16672 10976
rect 16672 10956 16724 10976
rect 16724 10956 16726 10976
rect 16670 10920 16726 10956
rect 17130 10784 17186 10840
rect 16524 10362 16580 10364
rect 16604 10362 16660 10364
rect 16684 10362 16740 10364
rect 16764 10362 16820 10364
rect 16524 10310 16570 10362
rect 16570 10310 16580 10362
rect 16604 10310 16634 10362
rect 16634 10310 16646 10362
rect 16646 10310 16660 10362
rect 16684 10310 16698 10362
rect 16698 10310 16710 10362
rect 16710 10310 16740 10362
rect 16764 10310 16774 10362
rect 16774 10310 16820 10362
rect 16524 10308 16580 10310
rect 16604 10308 16660 10310
rect 16684 10308 16740 10310
rect 16764 10308 16820 10310
rect 16394 9560 16450 9616
rect 16302 9424 16358 9480
rect 16524 9274 16580 9276
rect 16604 9274 16660 9276
rect 16684 9274 16740 9276
rect 16764 9274 16820 9276
rect 16524 9222 16570 9274
rect 16570 9222 16580 9274
rect 16604 9222 16634 9274
rect 16634 9222 16646 9274
rect 16646 9222 16660 9274
rect 16684 9222 16698 9274
rect 16698 9222 16710 9274
rect 16710 9222 16740 9274
rect 16764 9222 16774 9274
rect 16774 9222 16820 9274
rect 16524 9220 16580 9222
rect 16604 9220 16660 9222
rect 16684 9220 16740 9222
rect 16764 9220 16820 9222
rect 16670 8780 16672 8800
rect 16672 8780 16724 8800
rect 16724 8780 16726 8800
rect 16670 8744 16726 8780
rect 16524 8186 16580 8188
rect 16604 8186 16660 8188
rect 16684 8186 16740 8188
rect 16764 8186 16820 8188
rect 16524 8134 16570 8186
rect 16570 8134 16580 8186
rect 16604 8134 16634 8186
rect 16634 8134 16646 8186
rect 16646 8134 16660 8186
rect 16684 8134 16698 8186
rect 16698 8134 16710 8186
rect 16710 8134 16740 8186
rect 16764 8134 16774 8186
rect 16774 8134 16820 8186
rect 16524 8132 16580 8134
rect 16604 8132 16660 8134
rect 16684 8132 16740 8134
rect 16764 8132 16820 8134
rect 16118 6704 16174 6760
rect 17774 12144 17830 12200
rect 17682 11736 17738 11792
rect 17406 11500 17408 11520
rect 17408 11500 17460 11520
rect 17460 11500 17462 11520
rect 17406 11464 17462 11500
rect 17498 11192 17554 11248
rect 17682 10784 17738 10840
rect 17682 10376 17738 10432
rect 16210 5480 16266 5536
rect 16118 4528 16174 4584
rect 16524 7098 16580 7100
rect 16604 7098 16660 7100
rect 16684 7098 16740 7100
rect 16764 7098 16820 7100
rect 16524 7046 16570 7098
rect 16570 7046 16580 7098
rect 16604 7046 16634 7098
rect 16634 7046 16646 7098
rect 16646 7046 16660 7098
rect 16684 7046 16698 7098
rect 16698 7046 16710 7098
rect 16710 7046 16740 7098
rect 16764 7046 16774 7098
rect 16774 7046 16820 7098
rect 16524 7044 16580 7046
rect 16604 7044 16660 7046
rect 16684 7044 16740 7046
rect 16764 7044 16820 7046
rect 16670 6860 16726 6896
rect 16670 6840 16672 6860
rect 16672 6840 16724 6860
rect 16724 6840 16726 6860
rect 16762 6296 16818 6352
rect 16486 6196 16488 6216
rect 16488 6196 16540 6216
rect 16540 6196 16542 6216
rect 16486 6160 16542 6196
rect 16524 6010 16580 6012
rect 16604 6010 16660 6012
rect 16684 6010 16740 6012
rect 16764 6010 16820 6012
rect 16524 5958 16570 6010
rect 16570 5958 16580 6010
rect 16604 5958 16634 6010
rect 16634 5958 16646 6010
rect 16646 5958 16660 6010
rect 16684 5958 16698 6010
rect 16698 5958 16710 6010
rect 16710 5958 16740 6010
rect 16764 5958 16774 6010
rect 16774 5958 16820 6010
rect 16524 5956 16580 5958
rect 16604 5956 16660 5958
rect 16684 5956 16740 5958
rect 16764 5956 16820 5958
rect 16578 5616 16634 5672
rect 16854 5344 16910 5400
rect 16524 4922 16580 4924
rect 16604 4922 16660 4924
rect 16684 4922 16740 4924
rect 16764 4922 16820 4924
rect 16524 4870 16570 4922
rect 16570 4870 16580 4922
rect 16604 4870 16634 4922
rect 16634 4870 16646 4922
rect 16646 4870 16660 4922
rect 16684 4870 16698 4922
rect 16698 4870 16710 4922
rect 16710 4870 16740 4922
rect 16764 4870 16774 4922
rect 16774 4870 16820 4922
rect 16524 4868 16580 4870
rect 16604 4868 16660 4870
rect 16684 4868 16740 4870
rect 16764 4868 16820 4870
rect 16854 4256 16910 4312
rect 16670 4020 16672 4040
rect 16672 4020 16724 4040
rect 16724 4020 16726 4040
rect 16670 3984 16726 4020
rect 15934 3168 15990 3224
rect 16524 3834 16580 3836
rect 16604 3834 16660 3836
rect 16684 3834 16740 3836
rect 16764 3834 16820 3836
rect 16524 3782 16570 3834
rect 16570 3782 16580 3834
rect 16604 3782 16634 3834
rect 16634 3782 16646 3834
rect 16646 3782 16660 3834
rect 16684 3782 16698 3834
rect 16698 3782 16710 3834
rect 16710 3782 16740 3834
rect 16764 3782 16774 3834
rect 16774 3782 16820 3834
rect 16524 3780 16580 3782
rect 16604 3780 16660 3782
rect 16684 3780 16740 3782
rect 16764 3780 16820 3782
rect 17774 9288 17830 9344
rect 18786 13232 18842 13288
rect 17958 9968 18014 10024
rect 18418 10004 18420 10024
rect 18420 10004 18472 10024
rect 18472 10004 18474 10024
rect 18418 9968 18474 10004
rect 17590 8744 17646 8800
rect 17866 9016 17922 9072
rect 17222 7692 17224 7712
rect 17224 7692 17276 7712
rect 17276 7692 17278 7712
rect 17222 7656 17278 7692
rect 17406 7248 17462 7304
rect 17406 6432 17462 6488
rect 17130 5480 17186 5536
rect 16302 2896 16358 2952
rect 16524 2746 16580 2748
rect 16604 2746 16660 2748
rect 16684 2746 16740 2748
rect 16764 2746 16820 2748
rect 16524 2694 16570 2746
rect 16570 2694 16580 2746
rect 16604 2694 16634 2746
rect 16634 2694 16646 2746
rect 16646 2694 16660 2746
rect 16684 2694 16698 2746
rect 16698 2694 16710 2746
rect 16710 2694 16740 2746
rect 16764 2694 16774 2746
rect 16774 2694 16820 2746
rect 16524 2692 16580 2694
rect 16604 2692 16660 2694
rect 16684 2692 16740 2694
rect 16764 2692 16820 2694
rect 15198 176 15254 232
rect 17130 3460 17186 3496
rect 17130 3440 17132 3460
rect 17132 3440 17184 3460
rect 17184 3440 17186 3460
rect 17130 3052 17186 3088
rect 17130 3032 17132 3052
rect 17132 3032 17184 3052
rect 17184 3032 17186 3052
rect 16946 1400 17002 1456
rect 17958 7828 17960 7848
rect 17960 7828 18012 7848
rect 18012 7828 18014 7848
rect 17958 7792 18014 7828
rect 17958 7384 18014 7440
rect 17774 4800 17830 4856
rect 17498 4120 17554 4176
rect 17866 4392 17922 4448
rect 17682 3576 17738 3632
rect 17866 3168 17922 3224
rect 18050 6160 18106 6216
rect 18510 8608 18566 8664
rect 18418 8200 18474 8256
rect 18418 7792 18474 7848
rect 18418 6996 18474 7032
rect 18418 6976 18420 6996
rect 18420 6976 18472 6996
rect 18472 6976 18474 6996
rect 18418 6568 18474 6624
rect 18418 5616 18474 5672
rect 18050 5108 18052 5128
rect 18052 5108 18104 5128
rect 18104 5108 18106 5128
rect 18050 5072 18106 5108
rect 18786 7520 18842 7576
rect 18050 3168 18106 3224
rect 18418 3984 18474 4040
rect 17590 1808 17646 1864
rect 17314 992 17370 1048
rect 18418 2624 18474 2680
rect 17866 2216 17922 2272
rect 17774 856 17830 912
<< metal3 >>
rect 0 16826 800 16856
rect 3785 16826 3851 16829
rect 0 16824 3851 16826
rect 0 16768 3790 16824
rect 3846 16768 3851 16824
rect 0 16766 3851 16768
rect 0 16736 800 16766
rect 3785 16763 3851 16766
rect 16113 16826 16179 16829
rect 19200 16826 20000 16856
rect 16113 16824 20000 16826
rect 16113 16768 16118 16824
rect 16174 16768 20000 16824
rect 16113 16766 20000 16768
rect 16113 16763 16179 16766
rect 19200 16736 20000 16766
rect 0 16418 800 16448
rect 3877 16418 3943 16421
rect 0 16416 3943 16418
rect 0 16360 3882 16416
rect 3938 16360 3943 16416
rect 0 16358 3943 16360
rect 0 16328 800 16358
rect 3877 16355 3943 16358
rect 16297 16418 16363 16421
rect 19200 16418 20000 16448
rect 16297 16416 20000 16418
rect 16297 16360 16302 16416
rect 16358 16360 20000 16416
rect 16297 16358 20000 16360
rect 16297 16355 16363 16358
rect 19200 16328 20000 16358
rect 0 16010 800 16040
rect 3049 16010 3115 16013
rect 0 16008 3115 16010
rect 0 15952 3054 16008
rect 3110 15952 3115 16008
rect 0 15950 3115 15952
rect 0 15920 800 15950
rect 3049 15947 3115 15950
rect 16389 16010 16455 16013
rect 19200 16010 20000 16040
rect 16389 16008 20000 16010
rect 16389 15952 16394 16008
rect 16450 15952 20000 16008
rect 16389 15950 20000 15952
rect 16389 15947 16455 15950
rect 19200 15920 20000 15950
rect 0 15602 800 15632
rect 4153 15602 4219 15605
rect 0 15600 4219 15602
rect 0 15544 4158 15600
rect 4214 15544 4219 15600
rect 0 15542 4219 15544
rect 0 15512 800 15542
rect 4153 15539 4219 15542
rect 16113 15602 16179 15605
rect 19200 15602 20000 15632
rect 16113 15600 20000 15602
rect 16113 15544 16118 15600
rect 16174 15544 20000 15600
rect 16113 15542 20000 15544
rect 16113 15539 16179 15542
rect 19200 15512 20000 15542
rect 0 15194 800 15224
rect 3601 15194 3667 15197
rect 0 15192 3667 15194
rect 0 15136 3606 15192
rect 3662 15136 3667 15192
rect 0 15134 3667 15136
rect 0 15104 800 15134
rect 3601 15131 3667 15134
rect 16205 15194 16271 15197
rect 19200 15194 20000 15224
rect 16205 15192 20000 15194
rect 16205 15136 16210 15192
rect 16266 15136 20000 15192
rect 16205 15134 20000 15136
rect 16205 15131 16271 15134
rect 19200 15104 20000 15134
rect 0 14786 800 14816
rect 2957 14786 3023 14789
rect 0 14784 3023 14786
rect 0 14728 2962 14784
rect 3018 14728 3023 14784
rect 0 14726 3023 14728
rect 0 14696 800 14726
rect 2957 14723 3023 14726
rect 17401 14786 17467 14789
rect 19200 14786 20000 14816
rect 17401 14784 20000 14786
rect 17401 14728 17406 14784
rect 17462 14728 20000 14784
rect 17401 14726 20000 14728
rect 17401 14723 17467 14726
rect 3168 14720 3488 14721
rect 3168 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3488 14720
rect 3168 14655 3488 14656
rect 7616 14720 7936 14721
rect 7616 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7936 14720
rect 7616 14655 7936 14656
rect 12064 14720 12384 14721
rect 12064 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12384 14720
rect 12064 14655 12384 14656
rect 16512 14720 16832 14721
rect 16512 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16832 14720
rect 19200 14696 20000 14726
rect 16512 14655 16832 14656
rect 2221 14514 2287 14517
rect 8201 14514 8267 14517
rect 2221 14512 8267 14514
rect 2221 14456 2226 14512
rect 2282 14456 8206 14512
rect 8262 14456 8267 14512
rect 2221 14454 8267 14456
rect 2221 14451 2287 14454
rect 8201 14451 8267 14454
rect 0 14378 800 14408
rect 3049 14378 3115 14381
rect 0 14376 3115 14378
rect 0 14320 3054 14376
rect 3110 14320 3115 14376
rect 0 14318 3115 14320
rect 0 14288 800 14318
rect 3049 14315 3115 14318
rect 3417 14378 3483 14381
rect 7097 14378 7163 14381
rect 3417 14376 7163 14378
rect 3417 14320 3422 14376
rect 3478 14320 7102 14376
rect 7158 14320 7163 14376
rect 3417 14318 7163 14320
rect 3417 14315 3483 14318
rect 7097 14315 7163 14318
rect 17677 14242 17743 14245
rect 19200 14242 20000 14272
rect 17677 14240 20000 14242
rect 17677 14184 17682 14240
rect 17738 14184 20000 14240
rect 17677 14182 20000 14184
rect 17677 14179 17743 14182
rect 5392 14176 5712 14177
rect 5392 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5712 14176
rect 5392 14111 5712 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 14288 14176 14608 14177
rect 14288 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14608 14176
rect 19200 14152 20000 14182
rect 14288 14111 14608 14112
rect 0 13970 800 14000
rect 2221 13970 2287 13973
rect 0 13968 2287 13970
rect 0 13912 2226 13968
rect 2282 13912 2287 13968
rect 0 13910 2287 13912
rect 0 13880 800 13910
rect 2221 13907 2287 13910
rect 6177 13970 6243 13973
rect 7005 13970 7071 13973
rect 6177 13968 7071 13970
rect 6177 13912 6182 13968
rect 6238 13912 7010 13968
rect 7066 13912 7071 13968
rect 6177 13910 7071 13912
rect 6177 13907 6243 13910
rect 7005 13907 7071 13910
rect 4797 13834 4863 13837
rect 5717 13834 5783 13837
rect 4797 13832 5783 13834
rect 4797 13776 4802 13832
rect 4858 13776 5722 13832
rect 5778 13776 5783 13832
rect 4797 13774 5783 13776
rect 4797 13771 4863 13774
rect 5717 13771 5783 13774
rect 16246 13772 16252 13836
rect 16316 13834 16322 13836
rect 17033 13834 17099 13837
rect 16316 13832 17099 13834
rect 16316 13776 17038 13832
rect 17094 13776 17099 13832
rect 16316 13774 17099 13776
rect 16316 13772 16322 13774
rect 17033 13771 17099 13774
rect 17493 13834 17559 13837
rect 19200 13834 20000 13864
rect 17493 13832 20000 13834
rect 17493 13776 17498 13832
rect 17554 13776 20000 13832
rect 17493 13774 20000 13776
rect 17493 13771 17559 13774
rect 19200 13744 20000 13774
rect 3168 13632 3488 13633
rect 0 13562 800 13592
rect 3168 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3488 13632
rect 3168 13567 3488 13568
rect 7616 13632 7936 13633
rect 7616 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7936 13632
rect 7616 13567 7936 13568
rect 12064 13632 12384 13633
rect 12064 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12384 13632
rect 12064 13567 12384 13568
rect 16512 13632 16832 13633
rect 16512 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16832 13632
rect 16512 13567 16832 13568
rect 2773 13562 2839 13565
rect 0 13560 2839 13562
rect 0 13504 2778 13560
rect 2834 13504 2839 13560
rect 0 13502 2839 13504
rect 0 13472 800 13502
rect 2773 13499 2839 13502
rect 2957 13426 3023 13429
rect 14089 13426 14155 13429
rect 2822 13424 14155 13426
rect 2822 13368 2962 13424
rect 3018 13368 14094 13424
rect 14150 13368 14155 13424
rect 2822 13366 14155 13368
rect 2822 13293 2882 13366
rect 2957 13363 3023 13366
rect 14089 13363 14155 13366
rect 17677 13426 17743 13429
rect 19200 13426 20000 13456
rect 17677 13424 20000 13426
rect 17677 13368 17682 13424
rect 17738 13368 20000 13424
rect 17677 13366 20000 13368
rect 17677 13363 17743 13366
rect 19200 13336 20000 13366
rect 2773 13288 2882 13293
rect 2773 13232 2778 13288
rect 2834 13232 2882 13288
rect 2773 13230 2882 13232
rect 3509 13290 3575 13293
rect 5901 13290 5967 13293
rect 3509 13288 5967 13290
rect 3509 13232 3514 13288
rect 3570 13232 5906 13288
rect 5962 13232 5967 13288
rect 3509 13230 5967 13232
rect 2773 13227 2839 13230
rect 3509 13227 3575 13230
rect 5901 13227 5967 13230
rect 6361 13290 6427 13293
rect 18781 13290 18847 13293
rect 6361 13288 18847 13290
rect 6361 13232 6366 13288
rect 6422 13232 18786 13288
rect 18842 13232 18847 13288
rect 6361 13230 18847 13232
rect 6361 13227 6427 13230
rect 18781 13227 18847 13230
rect 0 13154 800 13184
rect 2221 13154 2287 13157
rect 0 13152 2287 13154
rect 0 13096 2226 13152
rect 2282 13096 2287 13152
rect 0 13094 2287 13096
rect 0 13064 800 13094
rect 2221 13091 2287 13094
rect 5392 13088 5712 13089
rect 5392 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5712 13088
rect 5392 13023 5712 13024
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 14288 13088 14608 13089
rect 14288 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14608 13088
rect 14288 13023 14608 13024
rect 17677 13018 17743 13021
rect 19200 13018 20000 13048
rect 17677 13016 20000 13018
rect 17677 12960 17682 13016
rect 17738 12960 20000 13016
rect 17677 12958 20000 12960
rect 17677 12955 17743 12958
rect 19200 12928 20000 12958
rect 1945 12882 2011 12885
rect 3734 12882 3740 12884
rect 1945 12880 3740 12882
rect 1945 12824 1950 12880
rect 2006 12824 3740 12880
rect 1945 12822 3740 12824
rect 1945 12819 2011 12822
rect 3734 12820 3740 12822
rect 3804 12820 3810 12884
rect 0 12746 800 12776
rect 2221 12746 2287 12749
rect 0 12744 2287 12746
rect 0 12688 2226 12744
rect 2282 12688 2287 12744
rect 0 12686 2287 12688
rect 0 12656 800 12686
rect 2221 12683 2287 12686
rect 12566 12684 12572 12748
rect 12636 12746 12642 12748
rect 17309 12746 17375 12749
rect 12636 12744 17375 12746
rect 12636 12688 17314 12744
rect 17370 12688 17375 12744
rect 12636 12686 17375 12688
rect 12636 12684 12642 12686
rect 17309 12683 17375 12686
rect 17677 12610 17743 12613
rect 19200 12610 20000 12640
rect 17677 12608 20000 12610
rect 17677 12552 17682 12608
rect 17738 12552 20000 12608
rect 17677 12550 20000 12552
rect 17677 12547 17743 12550
rect 3168 12544 3488 12545
rect 3168 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3488 12544
rect 3168 12479 3488 12480
rect 7616 12544 7936 12545
rect 7616 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7936 12544
rect 7616 12479 7936 12480
rect 12064 12544 12384 12545
rect 12064 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12384 12544
rect 12064 12479 12384 12480
rect 16512 12544 16832 12545
rect 16512 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16832 12544
rect 19200 12520 20000 12550
rect 16512 12479 16832 12480
rect 15101 12474 15167 12477
rect 15694 12474 15700 12476
rect 15101 12472 15700 12474
rect 15101 12416 15106 12472
rect 15162 12416 15700 12472
rect 15101 12414 15700 12416
rect 15101 12411 15167 12414
rect 15694 12412 15700 12414
rect 15764 12412 15770 12476
rect 0 12338 800 12368
rect 3233 12338 3299 12341
rect 0 12336 3299 12338
rect 0 12280 3238 12336
rect 3294 12280 3299 12336
rect 0 12278 3299 12280
rect 0 12248 800 12278
rect 3233 12275 3299 12278
rect 17769 12202 17835 12205
rect 19200 12202 20000 12232
rect 17769 12200 20000 12202
rect 17769 12144 17774 12200
rect 17830 12144 20000 12200
rect 17769 12142 20000 12144
rect 17769 12139 17835 12142
rect 19200 12112 20000 12142
rect 2957 12066 3023 12069
rect 4521 12066 4587 12069
rect 2957 12064 4587 12066
rect 2957 12008 2962 12064
rect 3018 12008 4526 12064
rect 4582 12008 4587 12064
rect 2957 12006 4587 12008
rect 2957 12003 3023 12006
rect 4521 12003 4587 12006
rect 5392 12000 5712 12001
rect 0 11930 800 11960
rect 5392 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5712 12000
rect 5392 11935 5712 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 14288 12000 14608 12001
rect 14288 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14608 12000
rect 14288 11935 14608 11936
rect 2773 11930 2839 11933
rect 0 11928 2839 11930
rect 0 11872 2778 11928
rect 2834 11872 2839 11928
rect 0 11870 2839 11872
rect 0 11840 800 11870
rect 2773 11867 2839 11870
rect 3693 11794 3759 11797
rect 12566 11794 12572 11796
rect 3693 11792 12572 11794
rect 3693 11736 3698 11792
rect 3754 11736 12572 11792
rect 3693 11734 12572 11736
rect 3693 11731 3759 11734
rect 12566 11732 12572 11734
rect 12636 11732 12642 11796
rect 17677 11794 17743 11797
rect 19200 11794 20000 11824
rect 17677 11792 20000 11794
rect 17677 11736 17682 11792
rect 17738 11736 20000 11792
rect 17677 11734 20000 11736
rect 17677 11731 17743 11734
rect 19200 11704 20000 11734
rect 3969 11658 4035 11661
rect 11145 11658 11211 11661
rect 3969 11656 11211 11658
rect 3969 11600 3974 11656
rect 4030 11600 11150 11656
rect 11206 11600 11211 11656
rect 3969 11598 11211 11600
rect 3969 11595 4035 11598
rect 11145 11595 11211 11598
rect 11286 11598 17234 11658
rect 8477 11522 8543 11525
rect 11286 11522 11346 11598
rect 17174 11524 17234 11598
rect 8477 11520 11346 11522
rect 8477 11464 8482 11520
rect 8538 11464 11346 11520
rect 8477 11462 11346 11464
rect 8477 11459 8543 11462
rect 17166 11460 17172 11524
rect 17236 11522 17242 11524
rect 17401 11522 17467 11525
rect 17236 11520 17467 11522
rect 17236 11464 17406 11520
rect 17462 11464 17467 11520
rect 17236 11462 17467 11464
rect 17236 11460 17242 11462
rect 17401 11459 17467 11462
rect 3168 11456 3488 11457
rect 0 11386 800 11416
rect 3168 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3488 11456
rect 3168 11391 3488 11392
rect 7616 11456 7936 11457
rect 7616 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7936 11456
rect 7616 11391 7936 11392
rect 12064 11456 12384 11457
rect 12064 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12384 11456
rect 12064 11391 12384 11392
rect 16512 11456 16832 11457
rect 16512 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16832 11456
rect 16512 11391 16832 11392
rect 2221 11386 2287 11389
rect 0 11384 2330 11386
rect 0 11328 2226 11384
rect 2282 11328 2330 11384
rect 0 11326 2330 11328
rect 0 11296 800 11326
rect 2221 11323 2330 11326
rect 2270 11250 2330 11323
rect 3417 11250 3483 11253
rect 2270 11248 3483 11250
rect 2270 11192 3422 11248
rect 3478 11192 3483 11248
rect 2270 11190 3483 11192
rect 3417 11187 3483 11190
rect 4061 11250 4127 11253
rect 4337 11250 4403 11253
rect 5809 11250 5875 11253
rect 15326 11250 15332 11252
rect 4061 11248 5642 11250
rect 4061 11192 4066 11248
rect 4122 11192 4342 11248
rect 4398 11192 5642 11248
rect 4061 11190 5642 11192
rect 4061 11187 4127 11190
rect 4337 11187 4403 11190
rect 1945 11114 2011 11117
rect 5257 11114 5323 11117
rect 1945 11112 5323 11114
rect 1945 11056 1950 11112
rect 2006 11056 5262 11112
rect 5318 11056 5323 11112
rect 1945 11054 5323 11056
rect 5582 11114 5642 11190
rect 5809 11248 15332 11250
rect 5809 11192 5814 11248
rect 5870 11192 15332 11248
rect 5809 11190 15332 11192
rect 5809 11187 5875 11190
rect 15326 11188 15332 11190
rect 15396 11188 15402 11252
rect 17493 11250 17559 11253
rect 19200 11250 20000 11280
rect 17493 11248 20000 11250
rect 17493 11192 17498 11248
rect 17554 11192 20000 11248
rect 17493 11190 20000 11192
rect 17493 11187 17559 11190
rect 19200 11160 20000 11190
rect 10409 11114 10475 11117
rect 5582 11112 10475 11114
rect 5582 11056 10414 11112
rect 10470 11056 10475 11112
rect 5582 11054 10475 11056
rect 1945 11051 2011 11054
rect 5257 11051 5323 11054
rect 10409 11051 10475 11054
rect 10869 11114 10935 11117
rect 13854 11114 13860 11116
rect 10869 11112 13860 11114
rect 10869 11056 10874 11112
rect 10930 11056 13860 11112
rect 10869 11054 13860 11056
rect 10869 11051 10935 11054
rect 13854 11052 13860 11054
rect 13924 11052 13930 11116
rect 15929 11114 15995 11117
rect 16982 11114 16988 11116
rect 15929 11112 16988 11114
rect 15929 11056 15934 11112
rect 15990 11056 16988 11112
rect 15929 11054 16988 11056
rect 15929 11051 15995 11054
rect 16982 11052 16988 11054
rect 17052 11052 17058 11116
rect 0 10978 800 11008
rect 2221 10978 2287 10981
rect 0 10976 2287 10978
rect 0 10920 2226 10976
rect 2282 10920 2287 10976
rect 0 10918 2287 10920
rect 0 10888 800 10918
rect 2221 10915 2287 10918
rect 16665 10978 16731 10981
rect 17350 10978 17356 10980
rect 16665 10976 17356 10978
rect 16665 10920 16670 10976
rect 16726 10920 17356 10976
rect 16665 10918 17356 10920
rect 16665 10915 16731 10918
rect 17350 10916 17356 10918
rect 17420 10916 17426 10980
rect 5392 10912 5712 10913
rect 5392 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5712 10912
rect 5392 10847 5712 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 14288 10912 14608 10913
rect 14288 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14608 10912
rect 14288 10847 14608 10848
rect 17125 10842 17191 10845
rect 14966 10840 17191 10842
rect 14966 10784 17130 10840
rect 17186 10784 17191 10840
rect 14966 10782 17191 10784
rect 1577 10706 1643 10709
rect 5901 10706 5967 10709
rect 1577 10704 5967 10706
rect 1577 10648 1582 10704
rect 1638 10648 5906 10704
rect 5962 10648 5967 10704
rect 1577 10646 5967 10648
rect 1577 10643 1643 10646
rect 5901 10643 5967 10646
rect 11237 10706 11303 10709
rect 14966 10706 15026 10782
rect 17125 10779 17191 10782
rect 17677 10842 17743 10845
rect 19200 10842 20000 10872
rect 17677 10840 20000 10842
rect 17677 10784 17682 10840
rect 17738 10784 20000 10840
rect 17677 10782 20000 10784
rect 17677 10779 17743 10782
rect 19200 10752 20000 10782
rect 15193 10708 15259 10709
rect 11237 10704 15026 10706
rect 11237 10648 11242 10704
rect 11298 10648 15026 10704
rect 11237 10646 15026 10648
rect 11237 10643 11303 10646
rect 15142 10644 15148 10708
rect 15212 10706 15259 10708
rect 15212 10704 15304 10706
rect 15254 10648 15304 10704
rect 15212 10646 15304 10648
rect 15212 10644 15259 10646
rect 15193 10643 15259 10644
rect 0 10570 800 10600
rect 1485 10570 1551 10573
rect 0 10568 1551 10570
rect 0 10512 1490 10568
rect 1546 10512 1551 10568
rect 0 10510 1551 10512
rect 0 10480 800 10510
rect 1485 10507 1551 10510
rect 6862 10508 6868 10572
rect 6932 10570 6938 10572
rect 15193 10570 15259 10573
rect 6932 10568 15259 10570
rect 6932 10512 15198 10568
rect 15254 10512 15259 10568
rect 6932 10510 15259 10512
rect 6932 10508 6938 10510
rect 15193 10507 15259 10510
rect 17677 10434 17743 10437
rect 19200 10434 20000 10464
rect 17677 10432 20000 10434
rect 17677 10376 17682 10432
rect 17738 10376 20000 10432
rect 17677 10374 20000 10376
rect 17677 10371 17743 10374
rect 3168 10368 3488 10369
rect 3168 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3488 10368
rect 3168 10303 3488 10304
rect 7616 10368 7936 10369
rect 7616 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7936 10368
rect 7616 10303 7936 10304
rect 12064 10368 12384 10369
rect 12064 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12384 10368
rect 12064 10303 12384 10304
rect 16512 10368 16832 10369
rect 16512 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16832 10368
rect 19200 10344 20000 10374
rect 16512 10303 16832 10304
rect 0 10162 800 10192
rect 1853 10162 1919 10165
rect 0 10160 1919 10162
rect 0 10104 1858 10160
rect 1914 10104 1919 10160
rect 0 10102 1919 10104
rect 0 10072 800 10102
rect 1853 10099 1919 10102
rect 3550 10100 3556 10164
rect 3620 10162 3626 10164
rect 3693 10162 3759 10165
rect 3620 10160 3759 10162
rect 3620 10104 3698 10160
rect 3754 10104 3759 10160
rect 3620 10102 3759 10104
rect 3620 10100 3626 10102
rect 3693 10099 3759 10102
rect 2313 10026 2379 10029
rect 4429 10026 4495 10029
rect 11605 10026 11671 10029
rect 2313 10024 11671 10026
rect 2313 9968 2318 10024
rect 2374 9968 4434 10024
rect 4490 9968 11610 10024
rect 11666 9968 11671 10024
rect 2313 9966 11671 9968
rect 2313 9963 2379 9966
rect 4429 9963 4495 9966
rect 11605 9963 11671 9966
rect 13353 10026 13419 10029
rect 17953 10026 18019 10029
rect 13353 10024 18019 10026
rect 13353 9968 13358 10024
rect 13414 9968 17958 10024
rect 18014 9968 18019 10024
rect 13353 9966 18019 9968
rect 13353 9963 13419 9966
rect 17953 9963 18019 9966
rect 18413 10026 18479 10029
rect 19200 10026 20000 10056
rect 18413 10024 20000 10026
rect 18413 9968 18418 10024
rect 18474 9968 20000 10024
rect 18413 9966 20000 9968
rect 18413 9963 18479 9966
rect 19200 9936 20000 9966
rect 5392 9824 5712 9825
rect 0 9754 800 9784
rect 5392 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5712 9824
rect 5392 9759 5712 9760
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 14288 9824 14608 9825
rect 14288 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14608 9824
rect 14288 9759 14608 9760
rect 2405 9754 2471 9757
rect 0 9752 2471 9754
rect 0 9696 2410 9752
rect 2466 9696 2471 9752
rect 0 9694 2471 9696
rect 0 9664 800 9694
rect 2405 9691 2471 9694
rect 2589 9618 2655 9621
rect 5165 9618 5231 9621
rect 2589 9616 5231 9618
rect 2589 9560 2594 9616
rect 2650 9560 5170 9616
rect 5226 9560 5231 9616
rect 2589 9558 5231 9560
rect 2589 9555 2655 9558
rect 5165 9555 5231 9558
rect 16389 9618 16455 9621
rect 19200 9618 20000 9648
rect 16389 9616 20000 9618
rect 16389 9560 16394 9616
rect 16450 9560 20000 9616
rect 16389 9558 20000 9560
rect 16389 9555 16455 9558
rect 19200 9528 20000 9558
rect 3601 9482 3667 9485
rect 10409 9482 10475 9485
rect 3601 9480 10475 9482
rect 3601 9424 3606 9480
rect 3662 9424 10414 9480
rect 10470 9424 10475 9480
rect 3601 9422 10475 9424
rect 3601 9419 3667 9422
rect 10409 9419 10475 9422
rect 11145 9482 11211 9485
rect 11145 9480 12588 9482
rect 11145 9424 11150 9480
rect 11206 9424 12588 9480
rect 11145 9422 12588 9424
rect 11145 9419 11211 9422
rect 0 9346 800 9376
rect 1301 9346 1367 9349
rect 0 9344 1367 9346
rect 0 9288 1306 9344
rect 1362 9288 1367 9344
rect 0 9286 1367 9288
rect 12528 9346 12588 9422
rect 15326 9420 15332 9484
rect 15396 9482 15402 9484
rect 16297 9482 16363 9485
rect 15396 9480 16363 9482
rect 15396 9424 16302 9480
rect 16358 9424 16363 9480
rect 15396 9422 16363 9424
rect 15396 9420 15402 9422
rect 16297 9419 16363 9422
rect 12801 9346 12867 9349
rect 15469 9346 15535 9349
rect 12528 9344 15535 9346
rect 12528 9288 12806 9344
rect 12862 9288 15474 9344
rect 15530 9288 15535 9344
rect 12528 9286 15535 9288
rect 0 9256 800 9286
rect 1301 9283 1367 9286
rect 12801 9283 12867 9286
rect 15469 9283 15535 9286
rect 17769 9346 17835 9349
rect 17769 9344 17970 9346
rect 17769 9288 17774 9344
rect 17830 9288 17970 9344
rect 17769 9286 17970 9288
rect 17769 9283 17835 9286
rect 3168 9280 3488 9281
rect 3168 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3488 9280
rect 3168 9215 3488 9216
rect 7616 9280 7936 9281
rect 7616 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7936 9280
rect 7616 9215 7936 9216
rect 12064 9280 12384 9281
rect 12064 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12384 9280
rect 12064 9215 12384 9216
rect 16512 9280 16832 9281
rect 16512 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16832 9280
rect 16512 9215 16832 9216
rect 12525 9210 12591 9213
rect 12893 9210 12959 9213
rect 13537 9210 13603 9213
rect 12525 9208 13603 9210
rect 12525 9152 12530 9208
rect 12586 9152 12898 9208
rect 12954 9152 13542 9208
rect 13598 9152 13603 9208
rect 12525 9150 13603 9152
rect 17910 9210 17970 9286
rect 19200 9210 20000 9240
rect 17910 9150 20000 9210
rect 12525 9147 12591 9150
rect 12893 9147 12959 9150
rect 13537 9147 13603 9150
rect 19200 9120 20000 9150
rect 2405 9074 2471 9077
rect 5717 9074 5783 9077
rect 2405 9072 5783 9074
rect 2405 9016 2410 9072
rect 2466 9016 5722 9072
rect 5778 9016 5783 9072
rect 2405 9014 5783 9016
rect 2405 9011 2471 9014
rect 5717 9011 5783 9014
rect 6821 9074 6887 9077
rect 9121 9074 9187 9077
rect 15837 9074 15903 9077
rect 17861 9074 17927 9077
rect 6821 9072 17927 9074
rect 6821 9016 6826 9072
rect 6882 9016 9126 9072
rect 9182 9016 15842 9072
rect 15898 9016 17866 9072
rect 17922 9016 17927 9072
rect 6821 9014 17927 9016
rect 6821 9011 6887 9014
rect 9121 9011 9187 9014
rect 15837 9011 15903 9014
rect 17861 9011 17927 9014
rect 0 8938 800 8968
rect 3049 8938 3115 8941
rect 0 8936 3115 8938
rect 0 8880 3054 8936
rect 3110 8880 3115 8936
rect 0 8878 3115 8880
rect 0 8848 800 8878
rect 3049 8875 3115 8878
rect 3417 8938 3483 8941
rect 3693 8938 3759 8941
rect 15193 8938 15259 8941
rect 15561 8938 15627 8941
rect 3417 8936 15627 8938
rect 3417 8880 3422 8936
rect 3478 8880 3698 8936
rect 3754 8880 15198 8936
rect 15254 8880 15566 8936
rect 15622 8880 15627 8936
rect 3417 8878 15627 8880
rect 3417 8875 3483 8878
rect 3693 8875 3759 8878
rect 15193 8875 15259 8878
rect 15561 8875 15627 8878
rect 6729 8802 6795 8805
rect 8201 8802 8267 8805
rect 6729 8800 8267 8802
rect 6729 8744 6734 8800
rect 6790 8744 8206 8800
rect 8262 8744 8267 8800
rect 6729 8742 8267 8744
rect 6729 8739 6795 8742
rect 8201 8739 8267 8742
rect 8753 8802 8819 8805
rect 9305 8802 9371 8805
rect 8753 8800 9371 8802
rect 8753 8744 8758 8800
rect 8814 8744 9310 8800
rect 9366 8744 9371 8800
rect 8753 8742 9371 8744
rect 8753 8739 8819 8742
rect 9305 8739 9371 8742
rect 11973 8802 12039 8805
rect 13721 8802 13787 8805
rect 11973 8800 13787 8802
rect 11973 8744 11978 8800
rect 12034 8744 13726 8800
rect 13782 8744 13787 8800
rect 11973 8742 13787 8744
rect 11973 8739 12039 8742
rect 13721 8739 13787 8742
rect 15929 8802 15995 8805
rect 16062 8802 16068 8804
rect 15929 8800 16068 8802
rect 15929 8744 15934 8800
rect 15990 8744 16068 8800
rect 15929 8742 16068 8744
rect 15929 8739 15995 8742
rect 16062 8740 16068 8742
rect 16132 8802 16138 8804
rect 16665 8802 16731 8805
rect 16132 8800 16731 8802
rect 16132 8744 16670 8800
rect 16726 8744 16731 8800
rect 16132 8742 16731 8744
rect 16132 8740 16138 8742
rect 16665 8739 16731 8742
rect 17585 8802 17651 8805
rect 19200 8802 20000 8832
rect 17585 8800 20000 8802
rect 17585 8744 17590 8800
rect 17646 8744 20000 8800
rect 17585 8742 20000 8744
rect 17585 8739 17651 8742
rect 5392 8736 5712 8737
rect 5392 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5712 8736
rect 5392 8671 5712 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 14288 8736 14608 8737
rect 14288 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14608 8736
rect 19200 8712 20000 8742
rect 14288 8671 14608 8672
rect 6821 8666 6887 8669
rect 8109 8666 8175 8669
rect 6821 8664 8175 8666
rect 6821 8608 6826 8664
rect 6882 8608 8114 8664
rect 8170 8608 8175 8664
rect 6821 8606 8175 8608
rect 6821 8603 6887 8606
rect 8109 8603 8175 8606
rect 8293 8666 8359 8669
rect 9489 8666 9555 8669
rect 8293 8664 9555 8666
rect 8293 8608 8298 8664
rect 8354 8608 9494 8664
rect 9550 8608 9555 8664
rect 8293 8606 9555 8608
rect 8293 8603 8359 8606
rect 9489 8603 9555 8606
rect 11513 8666 11579 8669
rect 13813 8666 13879 8669
rect 11513 8664 13879 8666
rect 11513 8608 11518 8664
rect 11574 8608 13818 8664
rect 13874 8608 13879 8664
rect 11513 8606 13879 8608
rect 11513 8603 11579 8606
rect 13813 8603 13879 8606
rect 16113 8666 16179 8669
rect 18505 8666 18571 8669
rect 16113 8664 18571 8666
rect 16113 8608 16118 8664
rect 16174 8608 18510 8664
rect 18566 8608 18571 8664
rect 16113 8606 18571 8608
rect 16113 8603 16179 8606
rect 18505 8603 18571 8606
rect 0 8530 800 8560
rect 1669 8530 1735 8533
rect 0 8528 1735 8530
rect 0 8472 1674 8528
rect 1730 8472 1735 8528
rect 0 8470 1735 8472
rect 0 8440 800 8470
rect 1669 8467 1735 8470
rect 2129 8530 2195 8533
rect 5073 8530 5139 8533
rect 2129 8528 5139 8530
rect 2129 8472 2134 8528
rect 2190 8472 5078 8528
rect 5134 8472 5139 8528
rect 2129 8470 5139 8472
rect 2129 8467 2195 8470
rect 5073 8467 5139 8470
rect 5257 8530 5323 8533
rect 11973 8530 12039 8533
rect 5257 8528 12039 8530
rect 5257 8472 5262 8528
rect 5318 8472 11978 8528
rect 12034 8472 12039 8528
rect 5257 8470 12039 8472
rect 13816 8530 13876 8603
rect 17350 8530 17356 8532
rect 13816 8470 17356 8530
rect 5257 8467 5323 8470
rect 11973 8467 12039 8470
rect 17350 8468 17356 8470
rect 17420 8468 17426 8532
rect 3877 8394 3943 8397
rect 16062 8394 16068 8396
rect 3877 8392 16068 8394
rect 3877 8336 3882 8392
rect 3938 8336 16068 8392
rect 3877 8334 16068 8336
rect 3877 8331 3943 8334
rect 16062 8332 16068 8334
rect 16132 8332 16138 8396
rect 14825 8258 14891 8261
rect 14958 8258 14964 8260
rect 14825 8256 14964 8258
rect 14825 8200 14830 8256
rect 14886 8200 14964 8256
rect 14825 8198 14964 8200
rect 14825 8195 14891 8198
rect 14958 8196 14964 8198
rect 15028 8196 15034 8260
rect 18413 8258 18479 8261
rect 19200 8258 20000 8288
rect 18413 8256 20000 8258
rect 18413 8200 18418 8256
rect 18474 8200 20000 8256
rect 18413 8198 20000 8200
rect 18413 8195 18479 8198
rect 3168 8192 3488 8193
rect 0 8122 800 8152
rect 3168 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3488 8192
rect 3168 8127 3488 8128
rect 7616 8192 7936 8193
rect 7616 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7936 8192
rect 7616 8127 7936 8128
rect 12064 8192 12384 8193
rect 12064 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12384 8192
rect 12064 8127 12384 8128
rect 16512 8192 16832 8193
rect 16512 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16832 8192
rect 19200 8168 20000 8198
rect 16512 8127 16832 8128
rect 1853 8122 1919 8125
rect 0 8120 1919 8122
rect 0 8064 1858 8120
rect 1914 8064 1919 8120
rect 0 8062 1919 8064
rect 0 8032 800 8062
rect 1853 8059 1919 8062
rect 2221 7986 2287 7989
rect 4521 7986 4587 7989
rect 8201 7986 8267 7989
rect 2221 7984 8267 7986
rect 2221 7928 2226 7984
rect 2282 7928 4526 7984
rect 4582 7928 8206 7984
rect 8262 7928 8267 7984
rect 2221 7926 8267 7928
rect 2221 7923 2287 7926
rect 4521 7923 4587 7926
rect 8201 7923 8267 7926
rect 9673 7986 9739 7989
rect 10041 7986 10107 7989
rect 13353 7986 13419 7989
rect 9673 7984 13419 7986
rect 9673 7928 9678 7984
rect 9734 7928 10046 7984
rect 10102 7928 13358 7984
rect 13414 7928 13419 7984
rect 9673 7926 13419 7928
rect 9673 7923 9739 7926
rect 10041 7923 10107 7926
rect 13353 7923 13419 7926
rect 14549 7986 14615 7989
rect 14825 7986 14891 7989
rect 14549 7984 14891 7986
rect 14549 7928 14554 7984
rect 14610 7928 14830 7984
rect 14886 7928 14891 7984
rect 14549 7926 14891 7928
rect 14549 7923 14615 7926
rect 14825 7923 14891 7926
rect 1945 7850 2011 7853
rect 3141 7850 3207 7853
rect 11237 7850 11303 7853
rect 1945 7848 11303 7850
rect 1945 7792 1950 7848
rect 2006 7792 3146 7848
rect 3202 7792 11242 7848
rect 11298 7792 11303 7848
rect 1945 7790 11303 7792
rect 1945 7787 2011 7790
rect 3141 7787 3207 7790
rect 11237 7787 11303 7790
rect 11973 7850 12039 7853
rect 15285 7850 15351 7853
rect 11973 7848 15351 7850
rect 11973 7792 11978 7848
rect 12034 7792 15290 7848
rect 15346 7792 15351 7848
rect 11973 7790 15351 7792
rect 11973 7787 12039 7790
rect 15285 7787 15351 7790
rect 15745 7850 15811 7853
rect 17953 7850 18019 7853
rect 15745 7848 18019 7850
rect 15745 7792 15750 7848
rect 15806 7792 17958 7848
rect 18014 7792 18019 7848
rect 15745 7790 18019 7792
rect 15745 7787 15811 7790
rect 17953 7787 18019 7790
rect 18413 7850 18479 7853
rect 19200 7850 20000 7880
rect 18413 7848 20000 7850
rect 18413 7792 18418 7848
rect 18474 7792 20000 7848
rect 18413 7790 20000 7792
rect 18413 7787 18479 7790
rect 19200 7760 20000 7790
rect 0 7714 800 7744
rect 1485 7714 1551 7717
rect 0 7712 1551 7714
rect 0 7656 1490 7712
rect 1546 7656 1551 7712
rect 0 7654 1551 7656
rect 0 7624 800 7654
rect 1485 7651 1551 7654
rect 17217 7714 17283 7717
rect 17350 7714 17356 7716
rect 17217 7712 17356 7714
rect 17217 7656 17222 7712
rect 17278 7656 17356 7712
rect 17217 7654 17356 7656
rect 17217 7651 17283 7654
rect 17350 7652 17356 7654
rect 17420 7652 17426 7716
rect 5392 7648 5712 7649
rect 5392 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5712 7648
rect 5392 7583 5712 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 14288 7648 14608 7649
rect 14288 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14608 7648
rect 14288 7583 14608 7584
rect 18781 7578 18847 7581
rect 16438 7576 18847 7578
rect 16438 7520 18786 7576
rect 18842 7520 18847 7576
rect 16438 7518 18847 7520
rect 3141 7442 3207 7445
rect 16438 7442 16498 7518
rect 18781 7515 18847 7518
rect 3141 7440 16498 7442
rect 3141 7384 3146 7440
rect 3202 7384 16498 7440
rect 3141 7382 16498 7384
rect 17953 7442 18019 7445
rect 19200 7442 20000 7472
rect 17953 7440 20000 7442
rect 17953 7384 17958 7440
rect 18014 7384 20000 7440
rect 17953 7382 20000 7384
rect 3141 7379 3207 7382
rect 17953 7379 18019 7382
rect 19200 7352 20000 7382
rect 0 7306 800 7336
rect 2221 7306 2287 7309
rect 0 7304 2287 7306
rect 0 7248 2226 7304
rect 2282 7248 2287 7304
rect 0 7246 2287 7248
rect 0 7216 800 7246
rect 2221 7243 2287 7246
rect 13261 7306 13327 7309
rect 17401 7306 17467 7309
rect 13261 7304 17467 7306
rect 13261 7248 13266 7304
rect 13322 7248 17406 7304
rect 17462 7248 17467 7304
rect 13261 7246 17467 7248
rect 13261 7243 13327 7246
rect 17401 7243 17467 7246
rect 3168 7104 3488 7105
rect 3168 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3488 7104
rect 3168 7039 3488 7040
rect 7616 7104 7936 7105
rect 7616 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7936 7104
rect 7616 7039 7936 7040
rect 12064 7104 12384 7105
rect 12064 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12384 7104
rect 12064 7039 12384 7040
rect 16512 7104 16832 7105
rect 16512 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16832 7104
rect 16512 7039 16832 7040
rect 18413 7034 18479 7037
rect 19200 7034 20000 7064
rect 18413 7032 20000 7034
rect 18413 6976 18418 7032
rect 18474 6976 20000 7032
rect 18413 6974 20000 6976
rect 18413 6971 18479 6974
rect 19200 6944 20000 6974
rect 0 6898 800 6928
rect 2313 6898 2379 6901
rect 0 6896 2379 6898
rect 0 6840 2318 6896
rect 2374 6840 2379 6896
rect 0 6838 2379 6840
rect 0 6808 800 6838
rect 2313 6835 2379 6838
rect 11513 6898 11579 6901
rect 13721 6898 13787 6901
rect 16665 6898 16731 6901
rect 11513 6896 16731 6898
rect 11513 6840 11518 6896
rect 11574 6840 13726 6896
rect 13782 6840 16670 6896
rect 16726 6840 16731 6896
rect 11513 6838 16731 6840
rect 11513 6835 11579 6838
rect 13721 6835 13787 6838
rect 16665 6835 16731 6838
rect 7649 6762 7715 6765
rect 16113 6762 16179 6765
rect 7649 6760 16179 6762
rect 7649 6704 7654 6760
rect 7710 6704 16118 6760
rect 16174 6704 16179 6760
rect 7649 6702 16179 6704
rect 7649 6699 7715 6702
rect 16113 6699 16179 6702
rect 18413 6626 18479 6629
rect 19200 6626 20000 6656
rect 18413 6624 20000 6626
rect 18413 6568 18418 6624
rect 18474 6568 20000 6624
rect 18413 6566 20000 6568
rect 18413 6563 18479 6566
rect 5392 6560 5712 6561
rect 0 6490 800 6520
rect 5392 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5712 6560
rect 5392 6495 5712 6496
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 14288 6560 14608 6561
rect 14288 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14608 6560
rect 19200 6536 20000 6566
rect 14288 6495 14608 6496
rect 1853 6490 1919 6493
rect 17401 6490 17467 6493
rect 0 6488 1919 6490
rect 0 6432 1858 6488
rect 1914 6432 1919 6488
rect 0 6430 1919 6432
rect 0 6400 800 6430
rect 1853 6427 1919 6430
rect 14966 6488 17467 6490
rect 14966 6432 17406 6488
rect 17462 6432 17467 6488
rect 14966 6430 17467 6432
rect 4521 6354 4587 6357
rect 7741 6354 7807 6357
rect 4521 6352 7807 6354
rect 4521 6296 4526 6352
rect 4582 6296 7746 6352
rect 7802 6296 7807 6352
rect 4521 6294 7807 6296
rect 4521 6291 4587 6294
rect 7741 6291 7807 6294
rect 8201 6354 8267 6357
rect 14966 6354 15026 6430
rect 17401 6427 17467 6430
rect 16757 6354 16823 6357
rect 8201 6352 15026 6354
rect 8201 6296 8206 6352
rect 8262 6296 15026 6352
rect 8201 6294 15026 6296
rect 15150 6352 16823 6354
rect 15150 6296 16762 6352
rect 16818 6296 16823 6352
rect 15150 6294 16823 6296
rect 8201 6291 8267 6294
rect 1853 6218 1919 6221
rect 7465 6218 7531 6221
rect 15150 6218 15210 6294
rect 16757 6291 16823 6294
rect 1853 6216 2790 6218
rect 1853 6160 1858 6216
rect 1914 6160 2790 6216
rect 1853 6158 2790 6160
rect 1853 6155 1919 6158
rect 0 6082 800 6112
rect 1485 6082 1551 6085
rect 0 6080 1551 6082
rect 0 6024 1490 6080
rect 1546 6024 1551 6080
rect 0 6022 1551 6024
rect 0 5992 800 6022
rect 1485 6019 1551 6022
rect 2730 5810 2790 6158
rect 7465 6216 15210 6218
rect 7465 6160 7470 6216
rect 7526 6160 15210 6216
rect 7465 6158 15210 6160
rect 15285 6218 15351 6221
rect 16246 6218 16252 6220
rect 15285 6216 16252 6218
rect 15285 6160 15290 6216
rect 15346 6160 16252 6216
rect 15285 6158 16252 6160
rect 7465 6155 7531 6158
rect 15285 6155 15351 6158
rect 16246 6156 16252 6158
rect 16316 6218 16322 6220
rect 16481 6218 16547 6221
rect 16316 6216 16547 6218
rect 16316 6160 16486 6216
rect 16542 6160 16547 6216
rect 16316 6158 16547 6160
rect 16316 6156 16322 6158
rect 16481 6155 16547 6158
rect 18045 6218 18111 6221
rect 19200 6218 20000 6248
rect 18045 6216 20000 6218
rect 18045 6160 18050 6216
rect 18106 6160 20000 6216
rect 18045 6158 20000 6160
rect 18045 6155 18111 6158
rect 19200 6128 20000 6158
rect 3168 6016 3488 6017
rect 3168 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3488 6016
rect 3168 5951 3488 5952
rect 7616 6016 7936 6017
rect 7616 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7936 6016
rect 7616 5951 7936 5952
rect 12064 6016 12384 6017
rect 12064 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12384 6016
rect 12064 5951 12384 5952
rect 16512 6016 16832 6017
rect 16512 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16832 6016
rect 16512 5951 16832 5952
rect 13721 5810 13787 5813
rect 2730 5808 13787 5810
rect 2730 5752 13726 5808
rect 13782 5752 13787 5808
rect 2730 5750 13787 5752
rect 1761 5674 1827 5677
rect 3049 5674 3115 5677
rect 1761 5672 3115 5674
rect 1761 5616 1766 5672
rect 1822 5616 3054 5672
rect 3110 5616 3115 5672
rect 1761 5614 3115 5616
rect 1761 5611 1827 5614
rect 3049 5611 3115 5614
rect 0 5538 800 5568
rect 3742 5541 3802 5750
rect 13721 5747 13787 5750
rect 4061 5674 4127 5677
rect 5901 5674 5967 5677
rect 4061 5672 5967 5674
rect 4061 5616 4066 5672
rect 4122 5616 5906 5672
rect 5962 5616 5967 5672
rect 4061 5614 5967 5616
rect 4061 5611 4127 5614
rect 5901 5611 5967 5614
rect 13077 5674 13143 5677
rect 16573 5674 16639 5677
rect 13077 5672 16639 5674
rect 13077 5616 13082 5672
rect 13138 5616 16578 5672
rect 16634 5616 16639 5672
rect 13077 5614 16639 5616
rect 13077 5611 13143 5614
rect 13494 5541 13554 5614
rect 16573 5611 16639 5614
rect 18413 5674 18479 5677
rect 19200 5674 20000 5704
rect 18413 5672 20000 5674
rect 18413 5616 18418 5672
rect 18474 5616 20000 5672
rect 18413 5614 20000 5616
rect 18413 5611 18479 5614
rect 19200 5584 20000 5614
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 3693 5536 3802 5541
rect 3693 5480 3698 5536
rect 3754 5480 3802 5536
rect 3693 5478 3802 5480
rect 9121 5538 9187 5541
rect 9673 5538 9739 5541
rect 9121 5536 9739 5538
rect 9121 5480 9126 5536
rect 9182 5480 9678 5536
rect 9734 5480 9739 5536
rect 9121 5478 9739 5480
rect 3693 5475 3759 5478
rect 9121 5475 9187 5478
rect 9673 5475 9739 5478
rect 13445 5536 13554 5541
rect 13445 5480 13450 5536
rect 13506 5480 13554 5536
rect 13445 5478 13554 5480
rect 13445 5475 13511 5478
rect 16062 5476 16068 5540
rect 16132 5538 16138 5540
rect 16205 5538 16271 5541
rect 16132 5536 16271 5538
rect 16132 5480 16210 5536
rect 16266 5480 16271 5536
rect 16132 5478 16271 5480
rect 16132 5476 16138 5478
rect 16205 5475 16271 5478
rect 17125 5540 17191 5541
rect 17125 5536 17172 5540
rect 17236 5538 17242 5540
rect 17125 5480 17130 5536
rect 17125 5476 17172 5480
rect 17236 5478 17282 5538
rect 17236 5476 17242 5478
rect 17125 5475 17191 5476
rect 5392 5472 5712 5473
rect 5392 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5712 5472
rect 5392 5407 5712 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 14288 5472 14608 5473
rect 14288 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14608 5472
rect 14288 5407 14608 5408
rect 15377 5402 15443 5405
rect 16849 5402 16915 5405
rect 15377 5400 16915 5402
rect 15377 5344 15382 5400
rect 15438 5344 16854 5400
rect 16910 5344 16915 5400
rect 15377 5342 16915 5344
rect 15377 5339 15443 5342
rect 16849 5339 16915 5342
rect 7189 5266 7255 5269
rect 7649 5266 7715 5269
rect 7189 5264 7715 5266
rect 7189 5208 7194 5264
rect 7250 5208 7654 5264
rect 7710 5208 7715 5264
rect 7189 5206 7715 5208
rect 7189 5203 7255 5206
rect 7649 5203 7715 5206
rect 15929 5266 15995 5269
rect 19200 5266 20000 5296
rect 15929 5264 20000 5266
rect 15929 5208 15934 5264
rect 15990 5208 20000 5264
rect 15929 5206 20000 5208
rect 15929 5203 15995 5206
rect 19200 5176 20000 5206
rect 0 5130 800 5160
rect 1485 5130 1551 5133
rect 0 5128 1551 5130
rect 0 5072 1490 5128
rect 1546 5072 1551 5128
rect 0 5070 1551 5072
rect 0 5040 800 5070
rect 1485 5067 1551 5070
rect 2221 5130 2287 5133
rect 6545 5130 6611 5133
rect 2221 5128 6611 5130
rect 2221 5072 2226 5128
rect 2282 5072 6550 5128
rect 6606 5072 6611 5128
rect 2221 5070 6611 5072
rect 2221 5067 2287 5070
rect 6545 5067 6611 5070
rect 12985 5130 13051 5133
rect 18045 5130 18111 5133
rect 12985 5128 18111 5130
rect 12985 5072 12990 5128
rect 13046 5072 18050 5128
rect 18106 5072 18111 5128
rect 12985 5070 18111 5072
rect 12985 5067 13051 5070
rect 18045 5067 18111 5070
rect 3168 4928 3488 4929
rect 3168 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3488 4928
rect 3168 4863 3488 4864
rect 7616 4928 7936 4929
rect 7616 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7936 4928
rect 7616 4863 7936 4864
rect 12064 4928 12384 4929
rect 12064 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12384 4928
rect 12064 4863 12384 4864
rect 16512 4928 16832 4929
rect 16512 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16832 4928
rect 16512 4863 16832 4864
rect 17769 4858 17835 4861
rect 19200 4858 20000 4888
rect 17769 4856 20000 4858
rect 17769 4800 17774 4856
rect 17830 4800 20000 4856
rect 17769 4798 20000 4800
rect 17769 4795 17835 4798
rect 19200 4768 20000 4798
rect 0 4722 800 4752
rect 1853 4722 1919 4725
rect 0 4720 1919 4722
rect 0 4664 1858 4720
rect 1914 4664 1919 4720
rect 0 4662 1919 4664
rect 0 4632 800 4662
rect 1853 4659 1919 4662
rect 11053 4722 11119 4725
rect 14958 4722 14964 4724
rect 11053 4720 14964 4722
rect 11053 4664 11058 4720
rect 11114 4664 14964 4720
rect 11053 4662 14964 4664
rect 11053 4659 11119 4662
rect 14958 4660 14964 4662
rect 15028 4660 15034 4724
rect 2037 4586 2103 4589
rect 2405 4586 2471 4589
rect 4889 4586 4955 4589
rect 2037 4584 4955 4586
rect 2037 4528 2042 4584
rect 2098 4528 2410 4584
rect 2466 4528 4894 4584
rect 4950 4528 4955 4584
rect 2037 4526 4955 4528
rect 2037 4523 2103 4526
rect 2405 4523 2471 4526
rect 4889 4523 4955 4526
rect 11237 4586 11303 4589
rect 16113 4586 16179 4589
rect 11237 4584 16179 4586
rect 11237 4528 11242 4584
rect 11298 4528 16118 4584
rect 16174 4528 16179 4584
rect 11237 4526 16179 4528
rect 11237 4523 11303 4526
rect 16113 4523 16179 4526
rect 3734 4388 3740 4452
rect 3804 4450 3810 4452
rect 4153 4450 4219 4453
rect 3804 4448 4219 4450
rect 3804 4392 4158 4448
rect 4214 4392 4219 4448
rect 3804 4390 4219 4392
rect 3804 4388 3810 4390
rect 4153 4387 4219 4390
rect 17861 4450 17927 4453
rect 19200 4450 20000 4480
rect 17861 4448 20000 4450
rect 17861 4392 17866 4448
rect 17922 4392 20000 4448
rect 17861 4390 20000 4392
rect 17861 4387 17927 4390
rect 5392 4384 5712 4385
rect 0 4314 800 4344
rect 5392 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5712 4384
rect 5392 4319 5712 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 14288 4384 14608 4385
rect 14288 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14608 4384
rect 19200 4360 20000 4390
rect 14288 4319 14608 4320
rect 1485 4314 1551 4317
rect 0 4312 1551 4314
rect 0 4256 1490 4312
rect 1546 4256 1551 4312
rect 0 4254 1551 4256
rect 0 4224 800 4254
rect 1485 4251 1551 4254
rect 2497 4314 2563 4317
rect 11973 4314 12039 4317
rect 13721 4314 13787 4317
rect 2497 4312 2790 4314
rect 2497 4256 2502 4312
rect 2558 4256 2790 4312
rect 2497 4254 2790 4256
rect 2497 4251 2563 4254
rect 2730 4042 2790 4254
rect 11973 4312 13787 4314
rect 11973 4256 11978 4312
rect 12034 4256 13726 4312
rect 13782 4256 13787 4312
rect 11973 4254 13787 4256
rect 11973 4251 12039 4254
rect 13721 4251 13787 4254
rect 14958 4252 14964 4316
rect 15028 4314 15034 4316
rect 16849 4314 16915 4317
rect 15028 4312 16915 4314
rect 15028 4256 16854 4312
rect 16910 4256 16915 4312
rect 15028 4254 16915 4256
rect 15028 4252 15034 4254
rect 16849 4251 16915 4254
rect 4153 4178 4219 4181
rect 7281 4178 7347 4181
rect 4153 4176 7347 4178
rect 4153 4120 4158 4176
rect 4214 4120 7286 4176
rect 7342 4120 7347 4176
rect 4153 4118 7347 4120
rect 4153 4115 4219 4118
rect 7281 4115 7347 4118
rect 10869 4178 10935 4181
rect 17493 4178 17559 4181
rect 10869 4176 17559 4178
rect 10869 4120 10874 4176
rect 10930 4120 17498 4176
rect 17554 4120 17559 4176
rect 10869 4118 17559 4120
rect 10869 4115 10935 4118
rect 17493 4115 17559 4118
rect 3785 4042 3851 4045
rect 2730 4040 3851 4042
rect 2730 3984 3790 4040
rect 3846 3984 3851 4040
rect 2730 3982 3851 3984
rect 3785 3979 3851 3982
rect 11513 4042 11579 4045
rect 12709 4042 12775 4045
rect 11513 4040 12775 4042
rect 11513 3984 11518 4040
rect 11574 3984 12714 4040
rect 12770 3984 12775 4040
rect 11513 3982 12775 3984
rect 11513 3979 11579 3982
rect 12709 3979 12775 3982
rect 13353 4042 13419 4045
rect 13629 4042 13695 4045
rect 13353 4040 13695 4042
rect 13353 3984 13358 4040
rect 13414 3984 13634 4040
rect 13690 3984 13695 4040
rect 13353 3982 13695 3984
rect 13353 3979 13419 3982
rect 13629 3979 13695 3982
rect 13854 3980 13860 4044
rect 13924 4042 13930 4044
rect 14089 4042 14155 4045
rect 13924 4040 14155 4042
rect 13924 3984 14094 4040
rect 14150 3984 14155 4040
rect 13924 3982 14155 3984
rect 13924 3980 13930 3982
rect 14089 3979 14155 3982
rect 15101 4044 15167 4045
rect 15101 4040 15148 4044
rect 15212 4042 15218 4044
rect 15561 4042 15627 4045
rect 15694 4042 15700 4044
rect 15101 3984 15106 4040
rect 15101 3980 15148 3984
rect 15212 3982 15258 4042
rect 15561 4040 15700 4042
rect 15561 3984 15566 4040
rect 15622 3984 15700 4040
rect 15561 3982 15700 3984
rect 15212 3980 15218 3982
rect 15101 3979 15167 3980
rect 15561 3979 15627 3982
rect 15694 3980 15700 3982
rect 15764 3980 15770 4044
rect 16665 4042 16731 4045
rect 15886 4040 16731 4042
rect 15886 3984 16670 4040
rect 16726 3984 16731 4040
rect 15886 3982 16731 3984
rect 0 3906 800 3936
rect 1485 3906 1551 3909
rect 0 3904 1551 3906
rect 0 3848 1490 3904
rect 1546 3848 1551 3904
rect 0 3846 1551 3848
rect 0 3816 800 3846
rect 1485 3843 1551 3846
rect 12709 3906 12775 3909
rect 13813 3906 13879 3909
rect 12709 3904 13879 3906
rect 12709 3848 12714 3904
rect 12770 3848 13818 3904
rect 13874 3848 13879 3904
rect 12709 3846 13879 3848
rect 12709 3843 12775 3846
rect 13813 3843 13879 3846
rect 3168 3840 3488 3841
rect 3168 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3488 3840
rect 3168 3775 3488 3776
rect 7616 3840 7936 3841
rect 7616 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7936 3840
rect 7616 3775 7936 3776
rect 12064 3840 12384 3841
rect 12064 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12384 3840
rect 12064 3775 12384 3776
rect 13629 3770 13695 3773
rect 15886 3770 15946 3982
rect 16665 3979 16731 3982
rect 18413 4042 18479 4045
rect 19200 4042 20000 4072
rect 18413 4040 20000 4042
rect 18413 3984 18418 4040
rect 18474 3984 20000 4040
rect 18413 3982 20000 3984
rect 18413 3979 18479 3982
rect 19200 3952 20000 3982
rect 16512 3840 16832 3841
rect 16512 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16832 3840
rect 16512 3775 16832 3776
rect 13629 3768 15946 3770
rect 13629 3712 13634 3768
rect 13690 3712 15946 3768
rect 13629 3710 15946 3712
rect 13629 3707 13695 3710
rect 2773 3634 2839 3637
rect 5901 3634 5967 3637
rect 2773 3632 5967 3634
rect 2773 3576 2778 3632
rect 2834 3576 5906 3632
rect 5962 3576 5967 3632
rect 2773 3574 5967 3576
rect 2773 3571 2839 3574
rect 5901 3571 5967 3574
rect 17677 3634 17743 3637
rect 19200 3634 20000 3664
rect 17677 3632 20000 3634
rect 17677 3576 17682 3632
rect 17738 3576 20000 3632
rect 17677 3574 20000 3576
rect 17677 3571 17743 3574
rect 19200 3544 20000 3574
rect 0 3498 800 3528
rect 1485 3498 1551 3501
rect 0 3496 1551 3498
rect 0 3440 1490 3496
rect 1546 3440 1551 3496
rect 0 3438 1551 3440
rect 0 3408 800 3438
rect 1485 3435 1551 3438
rect 1853 3498 1919 3501
rect 3233 3498 3299 3501
rect 1853 3496 3299 3498
rect 1853 3440 1858 3496
rect 1914 3440 3238 3496
rect 3294 3440 3299 3496
rect 1853 3438 3299 3440
rect 1853 3435 1919 3438
rect 3233 3435 3299 3438
rect 3417 3498 3483 3501
rect 3550 3498 3556 3500
rect 3417 3496 3556 3498
rect 3417 3440 3422 3496
rect 3478 3440 3556 3496
rect 3417 3438 3556 3440
rect 3417 3435 3483 3438
rect 3550 3436 3556 3438
rect 3620 3436 3626 3500
rect 4613 3498 4679 3501
rect 6862 3498 6868 3500
rect 4613 3496 6868 3498
rect 4613 3440 4618 3496
rect 4674 3440 6868 3496
rect 4613 3438 6868 3440
rect 4613 3435 4679 3438
rect 6862 3436 6868 3438
rect 6932 3436 6938 3500
rect 7281 3498 7347 3501
rect 13537 3498 13603 3501
rect 7281 3496 13603 3498
rect 7281 3440 7286 3496
rect 7342 3440 13542 3496
rect 13598 3440 13603 3496
rect 7281 3438 13603 3440
rect 7281 3435 7347 3438
rect 13537 3435 13603 3438
rect 16982 3436 16988 3500
rect 17052 3498 17058 3500
rect 17125 3498 17191 3501
rect 17052 3496 17191 3498
rect 17052 3440 17130 3496
rect 17186 3440 17191 3496
rect 17052 3438 17191 3440
rect 17052 3436 17058 3438
rect 17125 3435 17191 3438
rect 2129 3362 2195 3365
rect 5073 3362 5139 3365
rect 5257 3362 5323 3365
rect 2129 3360 5323 3362
rect 2129 3304 2134 3360
rect 2190 3304 5078 3360
rect 5134 3304 5262 3360
rect 5318 3304 5323 3360
rect 2129 3302 5323 3304
rect 2129 3299 2195 3302
rect 5073 3299 5139 3302
rect 5257 3299 5323 3302
rect 12433 3362 12499 3365
rect 12566 3362 12572 3364
rect 12433 3360 12572 3362
rect 12433 3304 12438 3360
rect 12494 3304 12572 3360
rect 12433 3302 12572 3304
rect 12433 3299 12499 3302
rect 12566 3300 12572 3302
rect 12636 3300 12642 3364
rect 5392 3296 5712 3297
rect 5392 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5712 3296
rect 5392 3231 5712 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 14288 3296 14608 3297
rect 14288 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14608 3296
rect 14288 3231 14608 3232
rect 15929 3226 15995 3229
rect 17861 3226 17927 3229
rect 15929 3224 17927 3226
rect 15929 3168 15934 3224
rect 15990 3168 17866 3224
rect 17922 3168 17927 3224
rect 15929 3166 17927 3168
rect 15929 3163 15995 3166
rect 17861 3163 17927 3166
rect 18045 3226 18111 3229
rect 19200 3226 20000 3256
rect 18045 3224 20000 3226
rect 18045 3168 18050 3224
rect 18106 3168 20000 3224
rect 18045 3166 20000 3168
rect 18045 3163 18111 3166
rect 19200 3136 20000 3166
rect 0 3090 800 3120
rect 1853 3090 1919 3093
rect 0 3088 1919 3090
rect 0 3032 1858 3088
rect 1914 3032 1919 3088
rect 0 3030 1919 3032
rect 0 3000 800 3030
rect 1853 3027 1919 3030
rect 15745 3090 15811 3093
rect 17125 3090 17191 3093
rect 15745 3088 17191 3090
rect 15745 3032 15750 3088
rect 15806 3032 17130 3088
rect 17186 3032 17191 3088
rect 15745 3030 17191 3032
rect 15745 3027 15811 3030
rect 17125 3027 17191 3030
rect 5901 2954 5967 2957
rect 6453 2954 6519 2957
rect 16297 2954 16363 2957
rect 5901 2952 16363 2954
rect 5901 2896 5906 2952
rect 5962 2896 6458 2952
rect 6514 2896 16302 2952
rect 16358 2896 16363 2952
rect 5901 2894 16363 2896
rect 5901 2891 5967 2894
rect 6453 2891 6519 2894
rect 16297 2891 16363 2894
rect 3168 2752 3488 2753
rect 0 2682 800 2712
rect 3168 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3488 2752
rect 3168 2687 3488 2688
rect 7616 2752 7936 2753
rect 7616 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7936 2752
rect 7616 2687 7936 2688
rect 12064 2752 12384 2753
rect 12064 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12384 2752
rect 12064 2687 12384 2688
rect 16512 2752 16832 2753
rect 16512 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16832 2752
rect 16512 2687 16832 2688
rect 1485 2682 1551 2685
rect 0 2680 1551 2682
rect 0 2624 1490 2680
rect 1546 2624 1551 2680
rect 0 2622 1551 2624
rect 0 2592 800 2622
rect 1485 2619 1551 2622
rect 18413 2682 18479 2685
rect 19200 2682 20000 2712
rect 18413 2680 20000 2682
rect 18413 2624 18418 2680
rect 18474 2624 20000 2680
rect 18413 2622 20000 2624
rect 18413 2619 18479 2622
rect 19200 2592 20000 2622
rect 0 2274 800 2304
rect 1485 2274 1551 2277
rect 0 2272 1551 2274
rect 0 2216 1490 2272
rect 1546 2216 1551 2272
rect 0 2214 1551 2216
rect 0 2184 800 2214
rect 1485 2211 1551 2214
rect 17861 2274 17927 2277
rect 19200 2274 20000 2304
rect 17861 2272 20000 2274
rect 17861 2216 17866 2272
rect 17922 2216 20000 2272
rect 17861 2214 20000 2216
rect 17861 2211 17927 2214
rect 5392 2208 5712 2209
rect 5392 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5712 2208
rect 5392 2143 5712 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 14288 2208 14608 2209
rect 14288 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14608 2208
rect 19200 2184 20000 2214
rect 14288 2143 14608 2144
rect 0 1866 800 1896
rect 3049 1866 3115 1869
rect 0 1864 3115 1866
rect 0 1808 3054 1864
rect 3110 1808 3115 1864
rect 0 1806 3115 1808
rect 0 1776 800 1806
rect 3049 1803 3115 1806
rect 17585 1866 17651 1869
rect 19200 1866 20000 1896
rect 17585 1864 20000 1866
rect 17585 1808 17590 1864
rect 17646 1808 20000 1864
rect 17585 1806 20000 1808
rect 17585 1803 17651 1806
rect 19200 1776 20000 1806
rect 0 1458 800 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 800 1398
rect 2773 1395 2839 1398
rect 16941 1458 17007 1461
rect 19200 1458 20000 1488
rect 16941 1456 20000 1458
rect 16941 1400 16946 1456
rect 17002 1400 20000 1456
rect 16941 1398 20000 1400
rect 16941 1395 17007 1398
rect 19200 1368 20000 1398
rect 0 1050 800 1080
rect 1577 1050 1643 1053
rect 0 1048 1643 1050
rect 0 992 1582 1048
rect 1638 992 1643 1048
rect 0 990 1643 992
rect 0 960 800 990
rect 1577 987 1643 990
rect 17309 1050 17375 1053
rect 19200 1050 20000 1080
rect 17309 1048 20000 1050
rect 17309 992 17314 1048
rect 17370 992 20000 1048
rect 17309 990 20000 992
rect 17309 987 17375 990
rect 19200 960 20000 990
rect 2957 914 3023 917
rect 1534 912 3023 914
rect 1534 856 2962 912
rect 3018 856 3023 912
rect 1534 854 3023 856
rect 0 642 800 672
rect 1534 642 1594 854
rect 2957 851 3023 854
rect 17769 914 17835 917
rect 17769 912 17970 914
rect 17769 856 17774 912
rect 17830 856 17970 912
rect 17769 854 17970 856
rect 17769 851 17835 854
rect 0 582 1594 642
rect 17910 642 17970 854
rect 19200 642 20000 672
rect 17910 582 20000 642
rect 0 552 800 582
rect 19200 552 20000 582
rect 0 234 800 264
rect 3877 234 3943 237
rect 0 232 3943 234
rect 0 176 3882 232
rect 3938 176 3943 232
rect 0 174 3943 176
rect 0 144 800 174
rect 3877 171 3943 174
rect 15193 234 15259 237
rect 19200 234 20000 264
rect 15193 232 20000 234
rect 15193 176 15198 232
rect 15254 176 20000 232
rect 15193 174 20000 176
rect 15193 171 15259 174
rect 19200 144 20000 174
<< via3 >>
rect 3176 14716 3240 14720
rect 3176 14660 3180 14716
rect 3180 14660 3236 14716
rect 3236 14660 3240 14716
rect 3176 14656 3240 14660
rect 3256 14716 3320 14720
rect 3256 14660 3260 14716
rect 3260 14660 3316 14716
rect 3316 14660 3320 14716
rect 3256 14656 3320 14660
rect 3336 14716 3400 14720
rect 3336 14660 3340 14716
rect 3340 14660 3396 14716
rect 3396 14660 3400 14716
rect 3336 14656 3400 14660
rect 3416 14716 3480 14720
rect 3416 14660 3420 14716
rect 3420 14660 3476 14716
rect 3476 14660 3480 14716
rect 3416 14656 3480 14660
rect 7624 14716 7688 14720
rect 7624 14660 7628 14716
rect 7628 14660 7684 14716
rect 7684 14660 7688 14716
rect 7624 14656 7688 14660
rect 7704 14716 7768 14720
rect 7704 14660 7708 14716
rect 7708 14660 7764 14716
rect 7764 14660 7768 14716
rect 7704 14656 7768 14660
rect 7784 14716 7848 14720
rect 7784 14660 7788 14716
rect 7788 14660 7844 14716
rect 7844 14660 7848 14716
rect 7784 14656 7848 14660
rect 7864 14716 7928 14720
rect 7864 14660 7868 14716
rect 7868 14660 7924 14716
rect 7924 14660 7928 14716
rect 7864 14656 7928 14660
rect 12072 14716 12136 14720
rect 12072 14660 12076 14716
rect 12076 14660 12132 14716
rect 12132 14660 12136 14716
rect 12072 14656 12136 14660
rect 12152 14716 12216 14720
rect 12152 14660 12156 14716
rect 12156 14660 12212 14716
rect 12212 14660 12216 14716
rect 12152 14656 12216 14660
rect 12232 14716 12296 14720
rect 12232 14660 12236 14716
rect 12236 14660 12292 14716
rect 12292 14660 12296 14716
rect 12232 14656 12296 14660
rect 12312 14716 12376 14720
rect 12312 14660 12316 14716
rect 12316 14660 12372 14716
rect 12372 14660 12376 14716
rect 12312 14656 12376 14660
rect 16520 14716 16584 14720
rect 16520 14660 16524 14716
rect 16524 14660 16580 14716
rect 16580 14660 16584 14716
rect 16520 14656 16584 14660
rect 16600 14716 16664 14720
rect 16600 14660 16604 14716
rect 16604 14660 16660 14716
rect 16660 14660 16664 14716
rect 16600 14656 16664 14660
rect 16680 14716 16744 14720
rect 16680 14660 16684 14716
rect 16684 14660 16740 14716
rect 16740 14660 16744 14716
rect 16680 14656 16744 14660
rect 16760 14716 16824 14720
rect 16760 14660 16764 14716
rect 16764 14660 16820 14716
rect 16820 14660 16824 14716
rect 16760 14656 16824 14660
rect 5400 14172 5464 14176
rect 5400 14116 5404 14172
rect 5404 14116 5460 14172
rect 5460 14116 5464 14172
rect 5400 14112 5464 14116
rect 5480 14172 5544 14176
rect 5480 14116 5484 14172
rect 5484 14116 5540 14172
rect 5540 14116 5544 14172
rect 5480 14112 5544 14116
rect 5560 14172 5624 14176
rect 5560 14116 5564 14172
rect 5564 14116 5620 14172
rect 5620 14116 5624 14172
rect 5560 14112 5624 14116
rect 5640 14172 5704 14176
rect 5640 14116 5644 14172
rect 5644 14116 5700 14172
rect 5700 14116 5704 14172
rect 5640 14112 5704 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 14296 14172 14360 14176
rect 14296 14116 14300 14172
rect 14300 14116 14356 14172
rect 14356 14116 14360 14172
rect 14296 14112 14360 14116
rect 14376 14172 14440 14176
rect 14376 14116 14380 14172
rect 14380 14116 14436 14172
rect 14436 14116 14440 14172
rect 14376 14112 14440 14116
rect 14456 14172 14520 14176
rect 14456 14116 14460 14172
rect 14460 14116 14516 14172
rect 14516 14116 14520 14172
rect 14456 14112 14520 14116
rect 14536 14172 14600 14176
rect 14536 14116 14540 14172
rect 14540 14116 14596 14172
rect 14596 14116 14600 14172
rect 14536 14112 14600 14116
rect 16252 13772 16316 13836
rect 3176 13628 3240 13632
rect 3176 13572 3180 13628
rect 3180 13572 3236 13628
rect 3236 13572 3240 13628
rect 3176 13568 3240 13572
rect 3256 13628 3320 13632
rect 3256 13572 3260 13628
rect 3260 13572 3316 13628
rect 3316 13572 3320 13628
rect 3256 13568 3320 13572
rect 3336 13628 3400 13632
rect 3336 13572 3340 13628
rect 3340 13572 3396 13628
rect 3396 13572 3400 13628
rect 3336 13568 3400 13572
rect 3416 13628 3480 13632
rect 3416 13572 3420 13628
rect 3420 13572 3476 13628
rect 3476 13572 3480 13628
rect 3416 13568 3480 13572
rect 7624 13628 7688 13632
rect 7624 13572 7628 13628
rect 7628 13572 7684 13628
rect 7684 13572 7688 13628
rect 7624 13568 7688 13572
rect 7704 13628 7768 13632
rect 7704 13572 7708 13628
rect 7708 13572 7764 13628
rect 7764 13572 7768 13628
rect 7704 13568 7768 13572
rect 7784 13628 7848 13632
rect 7784 13572 7788 13628
rect 7788 13572 7844 13628
rect 7844 13572 7848 13628
rect 7784 13568 7848 13572
rect 7864 13628 7928 13632
rect 7864 13572 7868 13628
rect 7868 13572 7924 13628
rect 7924 13572 7928 13628
rect 7864 13568 7928 13572
rect 12072 13628 12136 13632
rect 12072 13572 12076 13628
rect 12076 13572 12132 13628
rect 12132 13572 12136 13628
rect 12072 13568 12136 13572
rect 12152 13628 12216 13632
rect 12152 13572 12156 13628
rect 12156 13572 12212 13628
rect 12212 13572 12216 13628
rect 12152 13568 12216 13572
rect 12232 13628 12296 13632
rect 12232 13572 12236 13628
rect 12236 13572 12292 13628
rect 12292 13572 12296 13628
rect 12232 13568 12296 13572
rect 12312 13628 12376 13632
rect 12312 13572 12316 13628
rect 12316 13572 12372 13628
rect 12372 13572 12376 13628
rect 12312 13568 12376 13572
rect 16520 13628 16584 13632
rect 16520 13572 16524 13628
rect 16524 13572 16580 13628
rect 16580 13572 16584 13628
rect 16520 13568 16584 13572
rect 16600 13628 16664 13632
rect 16600 13572 16604 13628
rect 16604 13572 16660 13628
rect 16660 13572 16664 13628
rect 16600 13568 16664 13572
rect 16680 13628 16744 13632
rect 16680 13572 16684 13628
rect 16684 13572 16740 13628
rect 16740 13572 16744 13628
rect 16680 13568 16744 13572
rect 16760 13628 16824 13632
rect 16760 13572 16764 13628
rect 16764 13572 16820 13628
rect 16820 13572 16824 13628
rect 16760 13568 16824 13572
rect 5400 13084 5464 13088
rect 5400 13028 5404 13084
rect 5404 13028 5460 13084
rect 5460 13028 5464 13084
rect 5400 13024 5464 13028
rect 5480 13084 5544 13088
rect 5480 13028 5484 13084
rect 5484 13028 5540 13084
rect 5540 13028 5544 13084
rect 5480 13024 5544 13028
rect 5560 13084 5624 13088
rect 5560 13028 5564 13084
rect 5564 13028 5620 13084
rect 5620 13028 5624 13084
rect 5560 13024 5624 13028
rect 5640 13084 5704 13088
rect 5640 13028 5644 13084
rect 5644 13028 5700 13084
rect 5700 13028 5704 13084
rect 5640 13024 5704 13028
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 14296 13084 14360 13088
rect 14296 13028 14300 13084
rect 14300 13028 14356 13084
rect 14356 13028 14360 13084
rect 14296 13024 14360 13028
rect 14376 13084 14440 13088
rect 14376 13028 14380 13084
rect 14380 13028 14436 13084
rect 14436 13028 14440 13084
rect 14376 13024 14440 13028
rect 14456 13084 14520 13088
rect 14456 13028 14460 13084
rect 14460 13028 14516 13084
rect 14516 13028 14520 13084
rect 14456 13024 14520 13028
rect 14536 13084 14600 13088
rect 14536 13028 14540 13084
rect 14540 13028 14596 13084
rect 14596 13028 14600 13084
rect 14536 13024 14600 13028
rect 3740 12820 3804 12884
rect 12572 12684 12636 12748
rect 3176 12540 3240 12544
rect 3176 12484 3180 12540
rect 3180 12484 3236 12540
rect 3236 12484 3240 12540
rect 3176 12480 3240 12484
rect 3256 12540 3320 12544
rect 3256 12484 3260 12540
rect 3260 12484 3316 12540
rect 3316 12484 3320 12540
rect 3256 12480 3320 12484
rect 3336 12540 3400 12544
rect 3336 12484 3340 12540
rect 3340 12484 3396 12540
rect 3396 12484 3400 12540
rect 3336 12480 3400 12484
rect 3416 12540 3480 12544
rect 3416 12484 3420 12540
rect 3420 12484 3476 12540
rect 3476 12484 3480 12540
rect 3416 12480 3480 12484
rect 7624 12540 7688 12544
rect 7624 12484 7628 12540
rect 7628 12484 7684 12540
rect 7684 12484 7688 12540
rect 7624 12480 7688 12484
rect 7704 12540 7768 12544
rect 7704 12484 7708 12540
rect 7708 12484 7764 12540
rect 7764 12484 7768 12540
rect 7704 12480 7768 12484
rect 7784 12540 7848 12544
rect 7784 12484 7788 12540
rect 7788 12484 7844 12540
rect 7844 12484 7848 12540
rect 7784 12480 7848 12484
rect 7864 12540 7928 12544
rect 7864 12484 7868 12540
rect 7868 12484 7924 12540
rect 7924 12484 7928 12540
rect 7864 12480 7928 12484
rect 12072 12540 12136 12544
rect 12072 12484 12076 12540
rect 12076 12484 12132 12540
rect 12132 12484 12136 12540
rect 12072 12480 12136 12484
rect 12152 12540 12216 12544
rect 12152 12484 12156 12540
rect 12156 12484 12212 12540
rect 12212 12484 12216 12540
rect 12152 12480 12216 12484
rect 12232 12540 12296 12544
rect 12232 12484 12236 12540
rect 12236 12484 12292 12540
rect 12292 12484 12296 12540
rect 12232 12480 12296 12484
rect 12312 12540 12376 12544
rect 12312 12484 12316 12540
rect 12316 12484 12372 12540
rect 12372 12484 12376 12540
rect 12312 12480 12376 12484
rect 16520 12540 16584 12544
rect 16520 12484 16524 12540
rect 16524 12484 16580 12540
rect 16580 12484 16584 12540
rect 16520 12480 16584 12484
rect 16600 12540 16664 12544
rect 16600 12484 16604 12540
rect 16604 12484 16660 12540
rect 16660 12484 16664 12540
rect 16600 12480 16664 12484
rect 16680 12540 16744 12544
rect 16680 12484 16684 12540
rect 16684 12484 16740 12540
rect 16740 12484 16744 12540
rect 16680 12480 16744 12484
rect 16760 12540 16824 12544
rect 16760 12484 16764 12540
rect 16764 12484 16820 12540
rect 16820 12484 16824 12540
rect 16760 12480 16824 12484
rect 15700 12412 15764 12476
rect 5400 11996 5464 12000
rect 5400 11940 5404 11996
rect 5404 11940 5460 11996
rect 5460 11940 5464 11996
rect 5400 11936 5464 11940
rect 5480 11996 5544 12000
rect 5480 11940 5484 11996
rect 5484 11940 5540 11996
rect 5540 11940 5544 11996
rect 5480 11936 5544 11940
rect 5560 11996 5624 12000
rect 5560 11940 5564 11996
rect 5564 11940 5620 11996
rect 5620 11940 5624 11996
rect 5560 11936 5624 11940
rect 5640 11996 5704 12000
rect 5640 11940 5644 11996
rect 5644 11940 5700 11996
rect 5700 11940 5704 11996
rect 5640 11936 5704 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 14296 11996 14360 12000
rect 14296 11940 14300 11996
rect 14300 11940 14356 11996
rect 14356 11940 14360 11996
rect 14296 11936 14360 11940
rect 14376 11996 14440 12000
rect 14376 11940 14380 11996
rect 14380 11940 14436 11996
rect 14436 11940 14440 11996
rect 14376 11936 14440 11940
rect 14456 11996 14520 12000
rect 14456 11940 14460 11996
rect 14460 11940 14516 11996
rect 14516 11940 14520 11996
rect 14456 11936 14520 11940
rect 14536 11996 14600 12000
rect 14536 11940 14540 11996
rect 14540 11940 14596 11996
rect 14596 11940 14600 11996
rect 14536 11936 14600 11940
rect 12572 11732 12636 11796
rect 17172 11460 17236 11524
rect 3176 11452 3240 11456
rect 3176 11396 3180 11452
rect 3180 11396 3236 11452
rect 3236 11396 3240 11452
rect 3176 11392 3240 11396
rect 3256 11452 3320 11456
rect 3256 11396 3260 11452
rect 3260 11396 3316 11452
rect 3316 11396 3320 11452
rect 3256 11392 3320 11396
rect 3336 11452 3400 11456
rect 3336 11396 3340 11452
rect 3340 11396 3396 11452
rect 3396 11396 3400 11452
rect 3336 11392 3400 11396
rect 3416 11452 3480 11456
rect 3416 11396 3420 11452
rect 3420 11396 3476 11452
rect 3476 11396 3480 11452
rect 3416 11392 3480 11396
rect 7624 11452 7688 11456
rect 7624 11396 7628 11452
rect 7628 11396 7684 11452
rect 7684 11396 7688 11452
rect 7624 11392 7688 11396
rect 7704 11452 7768 11456
rect 7704 11396 7708 11452
rect 7708 11396 7764 11452
rect 7764 11396 7768 11452
rect 7704 11392 7768 11396
rect 7784 11452 7848 11456
rect 7784 11396 7788 11452
rect 7788 11396 7844 11452
rect 7844 11396 7848 11452
rect 7784 11392 7848 11396
rect 7864 11452 7928 11456
rect 7864 11396 7868 11452
rect 7868 11396 7924 11452
rect 7924 11396 7928 11452
rect 7864 11392 7928 11396
rect 12072 11452 12136 11456
rect 12072 11396 12076 11452
rect 12076 11396 12132 11452
rect 12132 11396 12136 11452
rect 12072 11392 12136 11396
rect 12152 11452 12216 11456
rect 12152 11396 12156 11452
rect 12156 11396 12212 11452
rect 12212 11396 12216 11452
rect 12152 11392 12216 11396
rect 12232 11452 12296 11456
rect 12232 11396 12236 11452
rect 12236 11396 12292 11452
rect 12292 11396 12296 11452
rect 12232 11392 12296 11396
rect 12312 11452 12376 11456
rect 12312 11396 12316 11452
rect 12316 11396 12372 11452
rect 12372 11396 12376 11452
rect 12312 11392 12376 11396
rect 16520 11452 16584 11456
rect 16520 11396 16524 11452
rect 16524 11396 16580 11452
rect 16580 11396 16584 11452
rect 16520 11392 16584 11396
rect 16600 11452 16664 11456
rect 16600 11396 16604 11452
rect 16604 11396 16660 11452
rect 16660 11396 16664 11452
rect 16600 11392 16664 11396
rect 16680 11452 16744 11456
rect 16680 11396 16684 11452
rect 16684 11396 16740 11452
rect 16740 11396 16744 11452
rect 16680 11392 16744 11396
rect 16760 11452 16824 11456
rect 16760 11396 16764 11452
rect 16764 11396 16820 11452
rect 16820 11396 16824 11452
rect 16760 11392 16824 11396
rect 15332 11188 15396 11252
rect 13860 11052 13924 11116
rect 16988 11052 17052 11116
rect 17356 10916 17420 10980
rect 5400 10908 5464 10912
rect 5400 10852 5404 10908
rect 5404 10852 5460 10908
rect 5460 10852 5464 10908
rect 5400 10848 5464 10852
rect 5480 10908 5544 10912
rect 5480 10852 5484 10908
rect 5484 10852 5540 10908
rect 5540 10852 5544 10908
rect 5480 10848 5544 10852
rect 5560 10908 5624 10912
rect 5560 10852 5564 10908
rect 5564 10852 5620 10908
rect 5620 10852 5624 10908
rect 5560 10848 5624 10852
rect 5640 10908 5704 10912
rect 5640 10852 5644 10908
rect 5644 10852 5700 10908
rect 5700 10852 5704 10908
rect 5640 10848 5704 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 14296 10908 14360 10912
rect 14296 10852 14300 10908
rect 14300 10852 14356 10908
rect 14356 10852 14360 10908
rect 14296 10848 14360 10852
rect 14376 10908 14440 10912
rect 14376 10852 14380 10908
rect 14380 10852 14436 10908
rect 14436 10852 14440 10908
rect 14376 10848 14440 10852
rect 14456 10908 14520 10912
rect 14456 10852 14460 10908
rect 14460 10852 14516 10908
rect 14516 10852 14520 10908
rect 14456 10848 14520 10852
rect 14536 10908 14600 10912
rect 14536 10852 14540 10908
rect 14540 10852 14596 10908
rect 14596 10852 14600 10908
rect 14536 10848 14600 10852
rect 15148 10704 15212 10708
rect 15148 10648 15198 10704
rect 15198 10648 15212 10704
rect 15148 10644 15212 10648
rect 6868 10508 6932 10572
rect 3176 10364 3240 10368
rect 3176 10308 3180 10364
rect 3180 10308 3236 10364
rect 3236 10308 3240 10364
rect 3176 10304 3240 10308
rect 3256 10364 3320 10368
rect 3256 10308 3260 10364
rect 3260 10308 3316 10364
rect 3316 10308 3320 10364
rect 3256 10304 3320 10308
rect 3336 10364 3400 10368
rect 3336 10308 3340 10364
rect 3340 10308 3396 10364
rect 3396 10308 3400 10364
rect 3336 10304 3400 10308
rect 3416 10364 3480 10368
rect 3416 10308 3420 10364
rect 3420 10308 3476 10364
rect 3476 10308 3480 10364
rect 3416 10304 3480 10308
rect 7624 10364 7688 10368
rect 7624 10308 7628 10364
rect 7628 10308 7684 10364
rect 7684 10308 7688 10364
rect 7624 10304 7688 10308
rect 7704 10364 7768 10368
rect 7704 10308 7708 10364
rect 7708 10308 7764 10364
rect 7764 10308 7768 10364
rect 7704 10304 7768 10308
rect 7784 10364 7848 10368
rect 7784 10308 7788 10364
rect 7788 10308 7844 10364
rect 7844 10308 7848 10364
rect 7784 10304 7848 10308
rect 7864 10364 7928 10368
rect 7864 10308 7868 10364
rect 7868 10308 7924 10364
rect 7924 10308 7928 10364
rect 7864 10304 7928 10308
rect 12072 10364 12136 10368
rect 12072 10308 12076 10364
rect 12076 10308 12132 10364
rect 12132 10308 12136 10364
rect 12072 10304 12136 10308
rect 12152 10364 12216 10368
rect 12152 10308 12156 10364
rect 12156 10308 12212 10364
rect 12212 10308 12216 10364
rect 12152 10304 12216 10308
rect 12232 10364 12296 10368
rect 12232 10308 12236 10364
rect 12236 10308 12292 10364
rect 12292 10308 12296 10364
rect 12232 10304 12296 10308
rect 12312 10364 12376 10368
rect 12312 10308 12316 10364
rect 12316 10308 12372 10364
rect 12372 10308 12376 10364
rect 12312 10304 12376 10308
rect 16520 10364 16584 10368
rect 16520 10308 16524 10364
rect 16524 10308 16580 10364
rect 16580 10308 16584 10364
rect 16520 10304 16584 10308
rect 16600 10364 16664 10368
rect 16600 10308 16604 10364
rect 16604 10308 16660 10364
rect 16660 10308 16664 10364
rect 16600 10304 16664 10308
rect 16680 10364 16744 10368
rect 16680 10308 16684 10364
rect 16684 10308 16740 10364
rect 16740 10308 16744 10364
rect 16680 10304 16744 10308
rect 16760 10364 16824 10368
rect 16760 10308 16764 10364
rect 16764 10308 16820 10364
rect 16820 10308 16824 10364
rect 16760 10304 16824 10308
rect 3556 10100 3620 10164
rect 5400 9820 5464 9824
rect 5400 9764 5404 9820
rect 5404 9764 5460 9820
rect 5460 9764 5464 9820
rect 5400 9760 5464 9764
rect 5480 9820 5544 9824
rect 5480 9764 5484 9820
rect 5484 9764 5540 9820
rect 5540 9764 5544 9820
rect 5480 9760 5544 9764
rect 5560 9820 5624 9824
rect 5560 9764 5564 9820
rect 5564 9764 5620 9820
rect 5620 9764 5624 9820
rect 5560 9760 5624 9764
rect 5640 9820 5704 9824
rect 5640 9764 5644 9820
rect 5644 9764 5700 9820
rect 5700 9764 5704 9820
rect 5640 9760 5704 9764
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 14296 9820 14360 9824
rect 14296 9764 14300 9820
rect 14300 9764 14356 9820
rect 14356 9764 14360 9820
rect 14296 9760 14360 9764
rect 14376 9820 14440 9824
rect 14376 9764 14380 9820
rect 14380 9764 14436 9820
rect 14436 9764 14440 9820
rect 14376 9760 14440 9764
rect 14456 9820 14520 9824
rect 14456 9764 14460 9820
rect 14460 9764 14516 9820
rect 14516 9764 14520 9820
rect 14456 9760 14520 9764
rect 14536 9820 14600 9824
rect 14536 9764 14540 9820
rect 14540 9764 14596 9820
rect 14596 9764 14600 9820
rect 14536 9760 14600 9764
rect 15332 9420 15396 9484
rect 3176 9276 3240 9280
rect 3176 9220 3180 9276
rect 3180 9220 3236 9276
rect 3236 9220 3240 9276
rect 3176 9216 3240 9220
rect 3256 9276 3320 9280
rect 3256 9220 3260 9276
rect 3260 9220 3316 9276
rect 3316 9220 3320 9276
rect 3256 9216 3320 9220
rect 3336 9276 3400 9280
rect 3336 9220 3340 9276
rect 3340 9220 3396 9276
rect 3396 9220 3400 9276
rect 3336 9216 3400 9220
rect 3416 9276 3480 9280
rect 3416 9220 3420 9276
rect 3420 9220 3476 9276
rect 3476 9220 3480 9276
rect 3416 9216 3480 9220
rect 7624 9276 7688 9280
rect 7624 9220 7628 9276
rect 7628 9220 7684 9276
rect 7684 9220 7688 9276
rect 7624 9216 7688 9220
rect 7704 9276 7768 9280
rect 7704 9220 7708 9276
rect 7708 9220 7764 9276
rect 7764 9220 7768 9276
rect 7704 9216 7768 9220
rect 7784 9276 7848 9280
rect 7784 9220 7788 9276
rect 7788 9220 7844 9276
rect 7844 9220 7848 9276
rect 7784 9216 7848 9220
rect 7864 9276 7928 9280
rect 7864 9220 7868 9276
rect 7868 9220 7924 9276
rect 7924 9220 7928 9276
rect 7864 9216 7928 9220
rect 12072 9276 12136 9280
rect 12072 9220 12076 9276
rect 12076 9220 12132 9276
rect 12132 9220 12136 9276
rect 12072 9216 12136 9220
rect 12152 9276 12216 9280
rect 12152 9220 12156 9276
rect 12156 9220 12212 9276
rect 12212 9220 12216 9276
rect 12152 9216 12216 9220
rect 12232 9276 12296 9280
rect 12232 9220 12236 9276
rect 12236 9220 12292 9276
rect 12292 9220 12296 9276
rect 12232 9216 12296 9220
rect 12312 9276 12376 9280
rect 12312 9220 12316 9276
rect 12316 9220 12372 9276
rect 12372 9220 12376 9276
rect 12312 9216 12376 9220
rect 16520 9276 16584 9280
rect 16520 9220 16524 9276
rect 16524 9220 16580 9276
rect 16580 9220 16584 9276
rect 16520 9216 16584 9220
rect 16600 9276 16664 9280
rect 16600 9220 16604 9276
rect 16604 9220 16660 9276
rect 16660 9220 16664 9276
rect 16600 9216 16664 9220
rect 16680 9276 16744 9280
rect 16680 9220 16684 9276
rect 16684 9220 16740 9276
rect 16740 9220 16744 9276
rect 16680 9216 16744 9220
rect 16760 9276 16824 9280
rect 16760 9220 16764 9276
rect 16764 9220 16820 9276
rect 16820 9220 16824 9276
rect 16760 9216 16824 9220
rect 16068 8740 16132 8804
rect 5400 8732 5464 8736
rect 5400 8676 5404 8732
rect 5404 8676 5460 8732
rect 5460 8676 5464 8732
rect 5400 8672 5464 8676
rect 5480 8732 5544 8736
rect 5480 8676 5484 8732
rect 5484 8676 5540 8732
rect 5540 8676 5544 8732
rect 5480 8672 5544 8676
rect 5560 8732 5624 8736
rect 5560 8676 5564 8732
rect 5564 8676 5620 8732
rect 5620 8676 5624 8732
rect 5560 8672 5624 8676
rect 5640 8732 5704 8736
rect 5640 8676 5644 8732
rect 5644 8676 5700 8732
rect 5700 8676 5704 8732
rect 5640 8672 5704 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 14296 8732 14360 8736
rect 14296 8676 14300 8732
rect 14300 8676 14356 8732
rect 14356 8676 14360 8732
rect 14296 8672 14360 8676
rect 14376 8732 14440 8736
rect 14376 8676 14380 8732
rect 14380 8676 14436 8732
rect 14436 8676 14440 8732
rect 14376 8672 14440 8676
rect 14456 8732 14520 8736
rect 14456 8676 14460 8732
rect 14460 8676 14516 8732
rect 14516 8676 14520 8732
rect 14456 8672 14520 8676
rect 14536 8732 14600 8736
rect 14536 8676 14540 8732
rect 14540 8676 14596 8732
rect 14596 8676 14600 8732
rect 14536 8672 14600 8676
rect 17356 8468 17420 8532
rect 16068 8332 16132 8396
rect 14964 8196 15028 8260
rect 3176 8188 3240 8192
rect 3176 8132 3180 8188
rect 3180 8132 3236 8188
rect 3236 8132 3240 8188
rect 3176 8128 3240 8132
rect 3256 8188 3320 8192
rect 3256 8132 3260 8188
rect 3260 8132 3316 8188
rect 3316 8132 3320 8188
rect 3256 8128 3320 8132
rect 3336 8188 3400 8192
rect 3336 8132 3340 8188
rect 3340 8132 3396 8188
rect 3396 8132 3400 8188
rect 3336 8128 3400 8132
rect 3416 8188 3480 8192
rect 3416 8132 3420 8188
rect 3420 8132 3476 8188
rect 3476 8132 3480 8188
rect 3416 8128 3480 8132
rect 7624 8188 7688 8192
rect 7624 8132 7628 8188
rect 7628 8132 7684 8188
rect 7684 8132 7688 8188
rect 7624 8128 7688 8132
rect 7704 8188 7768 8192
rect 7704 8132 7708 8188
rect 7708 8132 7764 8188
rect 7764 8132 7768 8188
rect 7704 8128 7768 8132
rect 7784 8188 7848 8192
rect 7784 8132 7788 8188
rect 7788 8132 7844 8188
rect 7844 8132 7848 8188
rect 7784 8128 7848 8132
rect 7864 8188 7928 8192
rect 7864 8132 7868 8188
rect 7868 8132 7924 8188
rect 7924 8132 7928 8188
rect 7864 8128 7928 8132
rect 12072 8188 12136 8192
rect 12072 8132 12076 8188
rect 12076 8132 12132 8188
rect 12132 8132 12136 8188
rect 12072 8128 12136 8132
rect 12152 8188 12216 8192
rect 12152 8132 12156 8188
rect 12156 8132 12212 8188
rect 12212 8132 12216 8188
rect 12152 8128 12216 8132
rect 12232 8188 12296 8192
rect 12232 8132 12236 8188
rect 12236 8132 12292 8188
rect 12292 8132 12296 8188
rect 12232 8128 12296 8132
rect 12312 8188 12376 8192
rect 12312 8132 12316 8188
rect 12316 8132 12372 8188
rect 12372 8132 12376 8188
rect 12312 8128 12376 8132
rect 16520 8188 16584 8192
rect 16520 8132 16524 8188
rect 16524 8132 16580 8188
rect 16580 8132 16584 8188
rect 16520 8128 16584 8132
rect 16600 8188 16664 8192
rect 16600 8132 16604 8188
rect 16604 8132 16660 8188
rect 16660 8132 16664 8188
rect 16600 8128 16664 8132
rect 16680 8188 16744 8192
rect 16680 8132 16684 8188
rect 16684 8132 16740 8188
rect 16740 8132 16744 8188
rect 16680 8128 16744 8132
rect 16760 8188 16824 8192
rect 16760 8132 16764 8188
rect 16764 8132 16820 8188
rect 16820 8132 16824 8188
rect 16760 8128 16824 8132
rect 17356 7652 17420 7716
rect 5400 7644 5464 7648
rect 5400 7588 5404 7644
rect 5404 7588 5460 7644
rect 5460 7588 5464 7644
rect 5400 7584 5464 7588
rect 5480 7644 5544 7648
rect 5480 7588 5484 7644
rect 5484 7588 5540 7644
rect 5540 7588 5544 7644
rect 5480 7584 5544 7588
rect 5560 7644 5624 7648
rect 5560 7588 5564 7644
rect 5564 7588 5620 7644
rect 5620 7588 5624 7644
rect 5560 7584 5624 7588
rect 5640 7644 5704 7648
rect 5640 7588 5644 7644
rect 5644 7588 5700 7644
rect 5700 7588 5704 7644
rect 5640 7584 5704 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 14296 7644 14360 7648
rect 14296 7588 14300 7644
rect 14300 7588 14356 7644
rect 14356 7588 14360 7644
rect 14296 7584 14360 7588
rect 14376 7644 14440 7648
rect 14376 7588 14380 7644
rect 14380 7588 14436 7644
rect 14436 7588 14440 7644
rect 14376 7584 14440 7588
rect 14456 7644 14520 7648
rect 14456 7588 14460 7644
rect 14460 7588 14516 7644
rect 14516 7588 14520 7644
rect 14456 7584 14520 7588
rect 14536 7644 14600 7648
rect 14536 7588 14540 7644
rect 14540 7588 14596 7644
rect 14596 7588 14600 7644
rect 14536 7584 14600 7588
rect 3176 7100 3240 7104
rect 3176 7044 3180 7100
rect 3180 7044 3236 7100
rect 3236 7044 3240 7100
rect 3176 7040 3240 7044
rect 3256 7100 3320 7104
rect 3256 7044 3260 7100
rect 3260 7044 3316 7100
rect 3316 7044 3320 7100
rect 3256 7040 3320 7044
rect 3336 7100 3400 7104
rect 3336 7044 3340 7100
rect 3340 7044 3396 7100
rect 3396 7044 3400 7100
rect 3336 7040 3400 7044
rect 3416 7100 3480 7104
rect 3416 7044 3420 7100
rect 3420 7044 3476 7100
rect 3476 7044 3480 7100
rect 3416 7040 3480 7044
rect 7624 7100 7688 7104
rect 7624 7044 7628 7100
rect 7628 7044 7684 7100
rect 7684 7044 7688 7100
rect 7624 7040 7688 7044
rect 7704 7100 7768 7104
rect 7704 7044 7708 7100
rect 7708 7044 7764 7100
rect 7764 7044 7768 7100
rect 7704 7040 7768 7044
rect 7784 7100 7848 7104
rect 7784 7044 7788 7100
rect 7788 7044 7844 7100
rect 7844 7044 7848 7100
rect 7784 7040 7848 7044
rect 7864 7100 7928 7104
rect 7864 7044 7868 7100
rect 7868 7044 7924 7100
rect 7924 7044 7928 7100
rect 7864 7040 7928 7044
rect 12072 7100 12136 7104
rect 12072 7044 12076 7100
rect 12076 7044 12132 7100
rect 12132 7044 12136 7100
rect 12072 7040 12136 7044
rect 12152 7100 12216 7104
rect 12152 7044 12156 7100
rect 12156 7044 12212 7100
rect 12212 7044 12216 7100
rect 12152 7040 12216 7044
rect 12232 7100 12296 7104
rect 12232 7044 12236 7100
rect 12236 7044 12292 7100
rect 12292 7044 12296 7100
rect 12232 7040 12296 7044
rect 12312 7100 12376 7104
rect 12312 7044 12316 7100
rect 12316 7044 12372 7100
rect 12372 7044 12376 7100
rect 12312 7040 12376 7044
rect 16520 7100 16584 7104
rect 16520 7044 16524 7100
rect 16524 7044 16580 7100
rect 16580 7044 16584 7100
rect 16520 7040 16584 7044
rect 16600 7100 16664 7104
rect 16600 7044 16604 7100
rect 16604 7044 16660 7100
rect 16660 7044 16664 7100
rect 16600 7040 16664 7044
rect 16680 7100 16744 7104
rect 16680 7044 16684 7100
rect 16684 7044 16740 7100
rect 16740 7044 16744 7100
rect 16680 7040 16744 7044
rect 16760 7100 16824 7104
rect 16760 7044 16764 7100
rect 16764 7044 16820 7100
rect 16820 7044 16824 7100
rect 16760 7040 16824 7044
rect 5400 6556 5464 6560
rect 5400 6500 5404 6556
rect 5404 6500 5460 6556
rect 5460 6500 5464 6556
rect 5400 6496 5464 6500
rect 5480 6556 5544 6560
rect 5480 6500 5484 6556
rect 5484 6500 5540 6556
rect 5540 6500 5544 6556
rect 5480 6496 5544 6500
rect 5560 6556 5624 6560
rect 5560 6500 5564 6556
rect 5564 6500 5620 6556
rect 5620 6500 5624 6556
rect 5560 6496 5624 6500
rect 5640 6556 5704 6560
rect 5640 6500 5644 6556
rect 5644 6500 5700 6556
rect 5700 6500 5704 6556
rect 5640 6496 5704 6500
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 14296 6556 14360 6560
rect 14296 6500 14300 6556
rect 14300 6500 14356 6556
rect 14356 6500 14360 6556
rect 14296 6496 14360 6500
rect 14376 6556 14440 6560
rect 14376 6500 14380 6556
rect 14380 6500 14436 6556
rect 14436 6500 14440 6556
rect 14376 6496 14440 6500
rect 14456 6556 14520 6560
rect 14456 6500 14460 6556
rect 14460 6500 14516 6556
rect 14516 6500 14520 6556
rect 14456 6496 14520 6500
rect 14536 6556 14600 6560
rect 14536 6500 14540 6556
rect 14540 6500 14596 6556
rect 14596 6500 14600 6556
rect 14536 6496 14600 6500
rect 16252 6156 16316 6220
rect 3176 6012 3240 6016
rect 3176 5956 3180 6012
rect 3180 5956 3236 6012
rect 3236 5956 3240 6012
rect 3176 5952 3240 5956
rect 3256 6012 3320 6016
rect 3256 5956 3260 6012
rect 3260 5956 3316 6012
rect 3316 5956 3320 6012
rect 3256 5952 3320 5956
rect 3336 6012 3400 6016
rect 3336 5956 3340 6012
rect 3340 5956 3396 6012
rect 3396 5956 3400 6012
rect 3336 5952 3400 5956
rect 3416 6012 3480 6016
rect 3416 5956 3420 6012
rect 3420 5956 3476 6012
rect 3476 5956 3480 6012
rect 3416 5952 3480 5956
rect 7624 6012 7688 6016
rect 7624 5956 7628 6012
rect 7628 5956 7684 6012
rect 7684 5956 7688 6012
rect 7624 5952 7688 5956
rect 7704 6012 7768 6016
rect 7704 5956 7708 6012
rect 7708 5956 7764 6012
rect 7764 5956 7768 6012
rect 7704 5952 7768 5956
rect 7784 6012 7848 6016
rect 7784 5956 7788 6012
rect 7788 5956 7844 6012
rect 7844 5956 7848 6012
rect 7784 5952 7848 5956
rect 7864 6012 7928 6016
rect 7864 5956 7868 6012
rect 7868 5956 7924 6012
rect 7924 5956 7928 6012
rect 7864 5952 7928 5956
rect 12072 6012 12136 6016
rect 12072 5956 12076 6012
rect 12076 5956 12132 6012
rect 12132 5956 12136 6012
rect 12072 5952 12136 5956
rect 12152 6012 12216 6016
rect 12152 5956 12156 6012
rect 12156 5956 12212 6012
rect 12212 5956 12216 6012
rect 12152 5952 12216 5956
rect 12232 6012 12296 6016
rect 12232 5956 12236 6012
rect 12236 5956 12292 6012
rect 12292 5956 12296 6012
rect 12232 5952 12296 5956
rect 12312 6012 12376 6016
rect 12312 5956 12316 6012
rect 12316 5956 12372 6012
rect 12372 5956 12376 6012
rect 12312 5952 12376 5956
rect 16520 6012 16584 6016
rect 16520 5956 16524 6012
rect 16524 5956 16580 6012
rect 16580 5956 16584 6012
rect 16520 5952 16584 5956
rect 16600 6012 16664 6016
rect 16600 5956 16604 6012
rect 16604 5956 16660 6012
rect 16660 5956 16664 6012
rect 16600 5952 16664 5956
rect 16680 6012 16744 6016
rect 16680 5956 16684 6012
rect 16684 5956 16740 6012
rect 16740 5956 16744 6012
rect 16680 5952 16744 5956
rect 16760 6012 16824 6016
rect 16760 5956 16764 6012
rect 16764 5956 16820 6012
rect 16820 5956 16824 6012
rect 16760 5952 16824 5956
rect 16068 5476 16132 5540
rect 17172 5536 17236 5540
rect 17172 5480 17186 5536
rect 17186 5480 17236 5536
rect 17172 5476 17236 5480
rect 5400 5468 5464 5472
rect 5400 5412 5404 5468
rect 5404 5412 5460 5468
rect 5460 5412 5464 5468
rect 5400 5408 5464 5412
rect 5480 5468 5544 5472
rect 5480 5412 5484 5468
rect 5484 5412 5540 5468
rect 5540 5412 5544 5468
rect 5480 5408 5544 5412
rect 5560 5468 5624 5472
rect 5560 5412 5564 5468
rect 5564 5412 5620 5468
rect 5620 5412 5624 5468
rect 5560 5408 5624 5412
rect 5640 5468 5704 5472
rect 5640 5412 5644 5468
rect 5644 5412 5700 5468
rect 5700 5412 5704 5468
rect 5640 5408 5704 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 14296 5468 14360 5472
rect 14296 5412 14300 5468
rect 14300 5412 14356 5468
rect 14356 5412 14360 5468
rect 14296 5408 14360 5412
rect 14376 5468 14440 5472
rect 14376 5412 14380 5468
rect 14380 5412 14436 5468
rect 14436 5412 14440 5468
rect 14376 5408 14440 5412
rect 14456 5468 14520 5472
rect 14456 5412 14460 5468
rect 14460 5412 14516 5468
rect 14516 5412 14520 5468
rect 14456 5408 14520 5412
rect 14536 5468 14600 5472
rect 14536 5412 14540 5468
rect 14540 5412 14596 5468
rect 14596 5412 14600 5468
rect 14536 5408 14600 5412
rect 3176 4924 3240 4928
rect 3176 4868 3180 4924
rect 3180 4868 3236 4924
rect 3236 4868 3240 4924
rect 3176 4864 3240 4868
rect 3256 4924 3320 4928
rect 3256 4868 3260 4924
rect 3260 4868 3316 4924
rect 3316 4868 3320 4924
rect 3256 4864 3320 4868
rect 3336 4924 3400 4928
rect 3336 4868 3340 4924
rect 3340 4868 3396 4924
rect 3396 4868 3400 4924
rect 3336 4864 3400 4868
rect 3416 4924 3480 4928
rect 3416 4868 3420 4924
rect 3420 4868 3476 4924
rect 3476 4868 3480 4924
rect 3416 4864 3480 4868
rect 7624 4924 7688 4928
rect 7624 4868 7628 4924
rect 7628 4868 7684 4924
rect 7684 4868 7688 4924
rect 7624 4864 7688 4868
rect 7704 4924 7768 4928
rect 7704 4868 7708 4924
rect 7708 4868 7764 4924
rect 7764 4868 7768 4924
rect 7704 4864 7768 4868
rect 7784 4924 7848 4928
rect 7784 4868 7788 4924
rect 7788 4868 7844 4924
rect 7844 4868 7848 4924
rect 7784 4864 7848 4868
rect 7864 4924 7928 4928
rect 7864 4868 7868 4924
rect 7868 4868 7924 4924
rect 7924 4868 7928 4924
rect 7864 4864 7928 4868
rect 12072 4924 12136 4928
rect 12072 4868 12076 4924
rect 12076 4868 12132 4924
rect 12132 4868 12136 4924
rect 12072 4864 12136 4868
rect 12152 4924 12216 4928
rect 12152 4868 12156 4924
rect 12156 4868 12212 4924
rect 12212 4868 12216 4924
rect 12152 4864 12216 4868
rect 12232 4924 12296 4928
rect 12232 4868 12236 4924
rect 12236 4868 12292 4924
rect 12292 4868 12296 4924
rect 12232 4864 12296 4868
rect 12312 4924 12376 4928
rect 12312 4868 12316 4924
rect 12316 4868 12372 4924
rect 12372 4868 12376 4924
rect 12312 4864 12376 4868
rect 16520 4924 16584 4928
rect 16520 4868 16524 4924
rect 16524 4868 16580 4924
rect 16580 4868 16584 4924
rect 16520 4864 16584 4868
rect 16600 4924 16664 4928
rect 16600 4868 16604 4924
rect 16604 4868 16660 4924
rect 16660 4868 16664 4924
rect 16600 4864 16664 4868
rect 16680 4924 16744 4928
rect 16680 4868 16684 4924
rect 16684 4868 16740 4924
rect 16740 4868 16744 4924
rect 16680 4864 16744 4868
rect 16760 4924 16824 4928
rect 16760 4868 16764 4924
rect 16764 4868 16820 4924
rect 16820 4868 16824 4924
rect 16760 4864 16824 4868
rect 14964 4660 15028 4724
rect 3740 4388 3804 4452
rect 5400 4380 5464 4384
rect 5400 4324 5404 4380
rect 5404 4324 5460 4380
rect 5460 4324 5464 4380
rect 5400 4320 5464 4324
rect 5480 4380 5544 4384
rect 5480 4324 5484 4380
rect 5484 4324 5540 4380
rect 5540 4324 5544 4380
rect 5480 4320 5544 4324
rect 5560 4380 5624 4384
rect 5560 4324 5564 4380
rect 5564 4324 5620 4380
rect 5620 4324 5624 4380
rect 5560 4320 5624 4324
rect 5640 4380 5704 4384
rect 5640 4324 5644 4380
rect 5644 4324 5700 4380
rect 5700 4324 5704 4380
rect 5640 4320 5704 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 14296 4380 14360 4384
rect 14296 4324 14300 4380
rect 14300 4324 14356 4380
rect 14356 4324 14360 4380
rect 14296 4320 14360 4324
rect 14376 4380 14440 4384
rect 14376 4324 14380 4380
rect 14380 4324 14436 4380
rect 14436 4324 14440 4380
rect 14376 4320 14440 4324
rect 14456 4380 14520 4384
rect 14456 4324 14460 4380
rect 14460 4324 14516 4380
rect 14516 4324 14520 4380
rect 14456 4320 14520 4324
rect 14536 4380 14600 4384
rect 14536 4324 14540 4380
rect 14540 4324 14596 4380
rect 14596 4324 14600 4380
rect 14536 4320 14600 4324
rect 14964 4252 15028 4316
rect 13860 3980 13924 4044
rect 15148 4040 15212 4044
rect 15148 3984 15162 4040
rect 15162 3984 15212 4040
rect 15148 3980 15212 3984
rect 15700 3980 15764 4044
rect 3176 3836 3240 3840
rect 3176 3780 3180 3836
rect 3180 3780 3236 3836
rect 3236 3780 3240 3836
rect 3176 3776 3240 3780
rect 3256 3836 3320 3840
rect 3256 3780 3260 3836
rect 3260 3780 3316 3836
rect 3316 3780 3320 3836
rect 3256 3776 3320 3780
rect 3336 3836 3400 3840
rect 3336 3780 3340 3836
rect 3340 3780 3396 3836
rect 3396 3780 3400 3836
rect 3336 3776 3400 3780
rect 3416 3836 3480 3840
rect 3416 3780 3420 3836
rect 3420 3780 3476 3836
rect 3476 3780 3480 3836
rect 3416 3776 3480 3780
rect 7624 3836 7688 3840
rect 7624 3780 7628 3836
rect 7628 3780 7684 3836
rect 7684 3780 7688 3836
rect 7624 3776 7688 3780
rect 7704 3836 7768 3840
rect 7704 3780 7708 3836
rect 7708 3780 7764 3836
rect 7764 3780 7768 3836
rect 7704 3776 7768 3780
rect 7784 3836 7848 3840
rect 7784 3780 7788 3836
rect 7788 3780 7844 3836
rect 7844 3780 7848 3836
rect 7784 3776 7848 3780
rect 7864 3836 7928 3840
rect 7864 3780 7868 3836
rect 7868 3780 7924 3836
rect 7924 3780 7928 3836
rect 7864 3776 7928 3780
rect 12072 3836 12136 3840
rect 12072 3780 12076 3836
rect 12076 3780 12132 3836
rect 12132 3780 12136 3836
rect 12072 3776 12136 3780
rect 12152 3836 12216 3840
rect 12152 3780 12156 3836
rect 12156 3780 12212 3836
rect 12212 3780 12216 3836
rect 12152 3776 12216 3780
rect 12232 3836 12296 3840
rect 12232 3780 12236 3836
rect 12236 3780 12292 3836
rect 12292 3780 12296 3836
rect 12232 3776 12296 3780
rect 12312 3836 12376 3840
rect 12312 3780 12316 3836
rect 12316 3780 12372 3836
rect 12372 3780 12376 3836
rect 12312 3776 12376 3780
rect 16520 3836 16584 3840
rect 16520 3780 16524 3836
rect 16524 3780 16580 3836
rect 16580 3780 16584 3836
rect 16520 3776 16584 3780
rect 16600 3836 16664 3840
rect 16600 3780 16604 3836
rect 16604 3780 16660 3836
rect 16660 3780 16664 3836
rect 16600 3776 16664 3780
rect 16680 3836 16744 3840
rect 16680 3780 16684 3836
rect 16684 3780 16740 3836
rect 16740 3780 16744 3836
rect 16680 3776 16744 3780
rect 16760 3836 16824 3840
rect 16760 3780 16764 3836
rect 16764 3780 16820 3836
rect 16820 3780 16824 3836
rect 16760 3776 16824 3780
rect 3556 3436 3620 3500
rect 6868 3436 6932 3500
rect 16988 3436 17052 3500
rect 12572 3300 12636 3364
rect 5400 3292 5464 3296
rect 5400 3236 5404 3292
rect 5404 3236 5460 3292
rect 5460 3236 5464 3292
rect 5400 3232 5464 3236
rect 5480 3292 5544 3296
rect 5480 3236 5484 3292
rect 5484 3236 5540 3292
rect 5540 3236 5544 3292
rect 5480 3232 5544 3236
rect 5560 3292 5624 3296
rect 5560 3236 5564 3292
rect 5564 3236 5620 3292
rect 5620 3236 5624 3292
rect 5560 3232 5624 3236
rect 5640 3292 5704 3296
rect 5640 3236 5644 3292
rect 5644 3236 5700 3292
rect 5700 3236 5704 3292
rect 5640 3232 5704 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 14296 3292 14360 3296
rect 14296 3236 14300 3292
rect 14300 3236 14356 3292
rect 14356 3236 14360 3292
rect 14296 3232 14360 3236
rect 14376 3292 14440 3296
rect 14376 3236 14380 3292
rect 14380 3236 14436 3292
rect 14436 3236 14440 3292
rect 14376 3232 14440 3236
rect 14456 3292 14520 3296
rect 14456 3236 14460 3292
rect 14460 3236 14516 3292
rect 14516 3236 14520 3292
rect 14456 3232 14520 3236
rect 14536 3292 14600 3296
rect 14536 3236 14540 3292
rect 14540 3236 14596 3292
rect 14596 3236 14600 3292
rect 14536 3232 14600 3236
rect 3176 2748 3240 2752
rect 3176 2692 3180 2748
rect 3180 2692 3236 2748
rect 3236 2692 3240 2748
rect 3176 2688 3240 2692
rect 3256 2748 3320 2752
rect 3256 2692 3260 2748
rect 3260 2692 3316 2748
rect 3316 2692 3320 2748
rect 3256 2688 3320 2692
rect 3336 2748 3400 2752
rect 3336 2692 3340 2748
rect 3340 2692 3396 2748
rect 3396 2692 3400 2748
rect 3336 2688 3400 2692
rect 3416 2748 3480 2752
rect 3416 2692 3420 2748
rect 3420 2692 3476 2748
rect 3476 2692 3480 2748
rect 3416 2688 3480 2692
rect 7624 2748 7688 2752
rect 7624 2692 7628 2748
rect 7628 2692 7684 2748
rect 7684 2692 7688 2748
rect 7624 2688 7688 2692
rect 7704 2748 7768 2752
rect 7704 2692 7708 2748
rect 7708 2692 7764 2748
rect 7764 2692 7768 2748
rect 7704 2688 7768 2692
rect 7784 2748 7848 2752
rect 7784 2692 7788 2748
rect 7788 2692 7844 2748
rect 7844 2692 7848 2748
rect 7784 2688 7848 2692
rect 7864 2748 7928 2752
rect 7864 2692 7868 2748
rect 7868 2692 7924 2748
rect 7924 2692 7928 2748
rect 7864 2688 7928 2692
rect 12072 2748 12136 2752
rect 12072 2692 12076 2748
rect 12076 2692 12132 2748
rect 12132 2692 12136 2748
rect 12072 2688 12136 2692
rect 12152 2748 12216 2752
rect 12152 2692 12156 2748
rect 12156 2692 12212 2748
rect 12212 2692 12216 2748
rect 12152 2688 12216 2692
rect 12232 2748 12296 2752
rect 12232 2692 12236 2748
rect 12236 2692 12292 2748
rect 12292 2692 12296 2748
rect 12232 2688 12296 2692
rect 12312 2748 12376 2752
rect 12312 2692 12316 2748
rect 12316 2692 12372 2748
rect 12372 2692 12376 2748
rect 12312 2688 12376 2692
rect 16520 2748 16584 2752
rect 16520 2692 16524 2748
rect 16524 2692 16580 2748
rect 16580 2692 16584 2748
rect 16520 2688 16584 2692
rect 16600 2748 16664 2752
rect 16600 2692 16604 2748
rect 16604 2692 16660 2748
rect 16660 2692 16664 2748
rect 16600 2688 16664 2692
rect 16680 2748 16744 2752
rect 16680 2692 16684 2748
rect 16684 2692 16740 2748
rect 16740 2692 16744 2748
rect 16680 2688 16744 2692
rect 16760 2748 16824 2752
rect 16760 2692 16764 2748
rect 16764 2692 16820 2748
rect 16820 2692 16824 2748
rect 16760 2688 16824 2692
rect 5400 2204 5464 2208
rect 5400 2148 5404 2204
rect 5404 2148 5460 2204
rect 5460 2148 5464 2204
rect 5400 2144 5464 2148
rect 5480 2204 5544 2208
rect 5480 2148 5484 2204
rect 5484 2148 5540 2204
rect 5540 2148 5544 2204
rect 5480 2144 5544 2148
rect 5560 2204 5624 2208
rect 5560 2148 5564 2204
rect 5564 2148 5620 2204
rect 5620 2148 5624 2204
rect 5560 2144 5624 2148
rect 5640 2204 5704 2208
rect 5640 2148 5644 2204
rect 5644 2148 5700 2204
rect 5700 2148 5704 2204
rect 5640 2144 5704 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 14296 2204 14360 2208
rect 14296 2148 14300 2204
rect 14300 2148 14356 2204
rect 14356 2148 14360 2204
rect 14296 2144 14360 2148
rect 14376 2204 14440 2208
rect 14376 2148 14380 2204
rect 14380 2148 14436 2204
rect 14436 2148 14440 2204
rect 14376 2144 14440 2148
rect 14456 2204 14520 2208
rect 14456 2148 14460 2204
rect 14460 2148 14516 2204
rect 14516 2148 14520 2204
rect 14456 2144 14520 2148
rect 14536 2204 14600 2208
rect 14536 2148 14540 2204
rect 14540 2148 14596 2204
rect 14596 2148 14600 2204
rect 14536 2144 14600 2148
<< metal4 >>
rect 3168 14720 3488 14736
rect 3168 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3488 14720
rect 3168 13632 3488 14656
rect 3168 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3488 13632
rect 3168 12544 3488 13568
rect 5392 14176 5712 14736
rect 5392 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5712 14176
rect 5392 13088 5712 14112
rect 5392 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5712 13088
rect 3739 12884 3805 12885
rect 3739 12820 3740 12884
rect 3804 12820 3805 12884
rect 3739 12819 3805 12820
rect 3168 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3488 12544
rect 3168 11456 3488 12480
rect 3168 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3488 11456
rect 3168 10368 3488 11392
rect 3168 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3488 10368
rect 3168 9280 3488 10304
rect 3555 10164 3621 10165
rect 3555 10100 3556 10164
rect 3620 10100 3621 10164
rect 3555 10099 3621 10100
rect 3168 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3488 9280
rect 3168 8192 3488 9216
rect 3168 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3488 8192
rect 3168 7104 3488 8128
rect 3168 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3488 7104
rect 3168 6016 3488 7040
rect 3168 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3488 6016
rect 3168 4928 3488 5952
rect 3168 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3488 4928
rect 3168 3840 3488 4864
rect 3168 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3488 3840
rect 3168 2752 3488 3776
rect 3558 3501 3618 10099
rect 3742 4453 3802 12819
rect 5392 12000 5712 13024
rect 5392 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5712 12000
rect 5392 10912 5712 11936
rect 5392 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5712 10912
rect 5392 9824 5712 10848
rect 7616 14720 7936 14736
rect 7616 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7936 14720
rect 7616 13632 7936 14656
rect 7616 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7936 13632
rect 7616 12544 7936 13568
rect 7616 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7936 12544
rect 7616 11456 7936 12480
rect 7616 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7936 11456
rect 6867 10572 6933 10573
rect 6867 10508 6868 10572
rect 6932 10508 6933 10572
rect 6867 10507 6933 10508
rect 5392 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5712 9824
rect 5392 8736 5712 9760
rect 5392 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5712 8736
rect 5392 7648 5712 8672
rect 5392 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5712 7648
rect 5392 6560 5712 7584
rect 5392 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5712 6560
rect 5392 5472 5712 6496
rect 5392 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5712 5472
rect 3739 4452 3805 4453
rect 3739 4388 3740 4452
rect 3804 4388 3805 4452
rect 3739 4387 3805 4388
rect 5392 4384 5712 5408
rect 5392 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5712 4384
rect 3555 3500 3621 3501
rect 3555 3436 3556 3500
rect 3620 3436 3621 3500
rect 3555 3435 3621 3436
rect 3168 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3488 2752
rect 3168 2128 3488 2688
rect 5392 3296 5712 4320
rect 6870 3501 6930 10507
rect 7616 10368 7936 11392
rect 7616 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7936 10368
rect 7616 9280 7936 10304
rect 7616 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7936 9280
rect 7616 8192 7936 9216
rect 7616 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7936 8192
rect 7616 7104 7936 8128
rect 7616 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7936 7104
rect 7616 6016 7936 7040
rect 7616 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7936 6016
rect 7616 4928 7936 5952
rect 7616 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7936 4928
rect 7616 3840 7936 4864
rect 7616 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7936 3840
rect 6867 3500 6933 3501
rect 6867 3436 6868 3500
rect 6932 3436 6933 3500
rect 6867 3435 6933 3436
rect 5392 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5712 3296
rect 5392 2208 5712 3232
rect 5392 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5712 2208
rect 5392 2128 5712 2144
rect 7616 2752 7936 3776
rect 7616 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7936 2752
rect 7616 2128 7936 2688
rect 9840 14176 10160 14736
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 2208 10160 3232
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 12064 14720 12384 14736
rect 12064 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12384 14720
rect 12064 13632 12384 14656
rect 12064 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12384 13632
rect 12064 12544 12384 13568
rect 14288 14176 14608 14736
rect 14288 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14608 14176
rect 14288 13088 14608 14112
rect 16512 14720 16832 14736
rect 16512 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16832 14720
rect 16251 13836 16317 13837
rect 16251 13772 16252 13836
rect 16316 13772 16317 13836
rect 16251 13771 16317 13772
rect 14288 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14608 13088
rect 12571 12748 12637 12749
rect 12571 12684 12572 12748
rect 12636 12684 12637 12748
rect 12571 12683 12637 12684
rect 12064 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12384 12544
rect 12064 11456 12384 12480
rect 12574 11797 12634 12683
rect 14288 12000 14608 13024
rect 15699 12476 15765 12477
rect 15699 12412 15700 12476
rect 15764 12412 15765 12476
rect 15699 12411 15765 12412
rect 14288 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14608 12000
rect 12571 11796 12637 11797
rect 12571 11732 12572 11796
rect 12636 11732 12637 11796
rect 12571 11731 12637 11732
rect 12064 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12384 11456
rect 12064 10368 12384 11392
rect 12064 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12384 10368
rect 12064 9280 12384 10304
rect 12064 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12384 9280
rect 12064 8192 12384 9216
rect 12064 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12384 8192
rect 12064 7104 12384 8128
rect 12064 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12384 7104
rect 12064 6016 12384 7040
rect 12064 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12384 6016
rect 12064 4928 12384 5952
rect 12064 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12384 4928
rect 12064 3840 12384 4864
rect 12064 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12384 3840
rect 12064 2752 12384 3776
rect 12574 3365 12634 11731
rect 13859 11116 13925 11117
rect 13859 11052 13860 11116
rect 13924 11052 13925 11116
rect 13859 11051 13925 11052
rect 13862 4045 13922 11051
rect 14288 10912 14608 11936
rect 15331 11252 15397 11253
rect 15331 11188 15332 11252
rect 15396 11188 15397 11252
rect 15331 11187 15397 11188
rect 14288 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14608 10912
rect 14288 9824 14608 10848
rect 15147 10708 15213 10709
rect 15147 10644 15148 10708
rect 15212 10644 15213 10708
rect 15147 10643 15213 10644
rect 14288 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14608 9824
rect 14288 8736 14608 9760
rect 14288 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14608 8736
rect 14288 7648 14608 8672
rect 14963 8260 15029 8261
rect 14963 8196 14964 8260
rect 15028 8196 15029 8260
rect 14963 8195 15029 8196
rect 14288 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14608 7648
rect 14288 6560 14608 7584
rect 14288 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14608 6560
rect 14288 5472 14608 6496
rect 14288 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14608 5472
rect 14288 4384 14608 5408
rect 14966 4725 15026 8195
rect 14963 4724 15029 4725
rect 14963 4660 14964 4724
rect 15028 4660 15029 4724
rect 14963 4659 15029 4660
rect 14288 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14608 4384
rect 13859 4044 13925 4045
rect 13859 3980 13860 4044
rect 13924 3980 13925 4044
rect 13859 3979 13925 3980
rect 12571 3364 12637 3365
rect 12571 3300 12572 3364
rect 12636 3300 12637 3364
rect 12571 3299 12637 3300
rect 12064 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12384 2752
rect 12064 2128 12384 2688
rect 14288 3296 14608 4320
rect 14966 4317 15026 4659
rect 14963 4316 15029 4317
rect 14963 4252 14964 4316
rect 15028 4252 15029 4316
rect 14963 4251 15029 4252
rect 15150 4045 15210 10643
rect 15334 9485 15394 11187
rect 15331 9484 15397 9485
rect 15331 9420 15332 9484
rect 15396 9420 15397 9484
rect 15331 9419 15397 9420
rect 15702 4045 15762 12411
rect 16067 8804 16133 8805
rect 16067 8740 16068 8804
rect 16132 8740 16133 8804
rect 16067 8739 16133 8740
rect 16070 8397 16130 8739
rect 16067 8396 16133 8397
rect 16067 8332 16068 8396
rect 16132 8332 16133 8396
rect 16067 8331 16133 8332
rect 16070 5541 16130 8331
rect 16254 6221 16314 13771
rect 16512 13632 16832 14656
rect 16512 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16832 13632
rect 16512 12544 16832 13568
rect 16512 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16832 12544
rect 16512 11456 16832 12480
rect 17171 11524 17237 11525
rect 17171 11460 17172 11524
rect 17236 11460 17237 11524
rect 17171 11459 17237 11460
rect 16512 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16832 11456
rect 16512 10368 16832 11392
rect 16987 11116 17053 11117
rect 16987 11052 16988 11116
rect 17052 11052 17053 11116
rect 16987 11051 17053 11052
rect 16512 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16832 10368
rect 16512 9280 16832 10304
rect 16512 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16832 9280
rect 16512 8192 16832 9216
rect 16512 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16832 8192
rect 16512 7104 16832 8128
rect 16512 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16832 7104
rect 16251 6220 16317 6221
rect 16251 6156 16252 6220
rect 16316 6156 16317 6220
rect 16251 6155 16317 6156
rect 16512 6016 16832 7040
rect 16512 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16832 6016
rect 16067 5540 16133 5541
rect 16067 5476 16068 5540
rect 16132 5476 16133 5540
rect 16067 5475 16133 5476
rect 16512 4928 16832 5952
rect 16512 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16832 4928
rect 15147 4044 15213 4045
rect 15147 3980 15148 4044
rect 15212 3980 15213 4044
rect 15147 3979 15213 3980
rect 15699 4044 15765 4045
rect 15699 3980 15700 4044
rect 15764 3980 15765 4044
rect 15699 3979 15765 3980
rect 14288 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14608 3296
rect 14288 2208 14608 3232
rect 14288 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14608 2208
rect 14288 2128 14608 2144
rect 16512 3840 16832 4864
rect 16512 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16832 3840
rect 16512 2752 16832 3776
rect 16990 3501 17050 11051
rect 17174 5541 17234 11459
rect 17355 10980 17421 10981
rect 17355 10916 17356 10980
rect 17420 10916 17421 10980
rect 17355 10915 17421 10916
rect 17358 8533 17418 10915
rect 17355 8532 17421 8533
rect 17355 8468 17356 8532
rect 17420 8468 17421 8532
rect 17355 8467 17421 8468
rect 17358 7717 17418 8467
rect 17355 7716 17421 7717
rect 17355 7652 17356 7716
rect 17420 7652 17421 7716
rect 17355 7651 17421 7652
rect 17171 5540 17237 5541
rect 17171 5476 17172 5540
rect 17236 5476 17237 5540
rect 17171 5475 17237 5476
rect 16987 3500 17053 3501
rect 16987 3436 16988 3500
rect 17052 3436 17053 3500
rect 16987 3435 17053 3436
rect 16512 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16832 2752
rect 16512 2128 16832 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__18__A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__19__A
timestamp 1649977179
transform -1 0 5612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__20__A
timestamp 1649977179
transform -1 0 5428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A
timestamp 1649977179
transform -1 0 5060 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__22__A
timestamp 1649977179
transform -1 0 5980 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__23__A
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__24__A
timestamp 1649977179
transform -1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__25__A
timestamp 1649977179
transform -1 0 5796 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__26__A
timestamp 1649977179
transform -1 0 5244 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__27__A
timestamp 1649977179
transform -1 0 4048 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__28__A
timestamp 1649977179
transform -1 0 2760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__29__A
timestamp 1649977179
transform -1 0 4232 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__30__A
timestamp 1649977179
transform -1 0 3680 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__31__A
timestamp 1649977179
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__32__A
timestamp 1649977179
transform -1 0 2668 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__35__A
timestamp 1649977179
transform -1 0 11408 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A
timestamp 1649977179
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A
timestamp 1649977179
transform -1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform -1 0 16560 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform -1 0 17848 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform -1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform -1 0 15548 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform -1 0 8188 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform 1 0 15456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__47__A
timestamp 1649977179
transform 1 0 17204 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform -1 0 5980 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform 1 0 16008 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform 1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1649977179
transform 1 0 13616 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform 1 0 14628 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform 1 0 16100 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1649977179
transform 1 0 6900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1649977179
transform 1 0 6440 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__80__A
timestamp 1649977179
transform 1 0 6256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1649977179
transform 1 0 5612 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__85__A
timestamp 1649977179
transform -1 0 2576 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_0_N_in_A
timestamp 1649977179
transform 1 0 7360 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 7452 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 5704 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 7268 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 4876 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 3680 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 6532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 8372 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 4968 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 7636 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 7452 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 8188 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 5980 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 6808 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 8004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 3588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 2484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 1564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 1564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 4140 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 4324 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 4508 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 6164 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 17664 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 16192 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 15088 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 17296 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 17296 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 14720 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 16376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 16560 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 17112 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 16744 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 15272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 16928 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 16008 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 16560 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 17020 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 17296 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 17664 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 17112 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 16928 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 7728 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 13248 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 10672 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 16560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 11408 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 14996 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 12420 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 12604 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 14536 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 9384 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 10028 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 10672 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 11960 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 4508 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4140 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4232 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7912 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 8280 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4232 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 4048 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 2576 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 2668 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 3956 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 3312 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4600 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7360 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5704 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7176 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 5244 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9844 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 7728 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 6992 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14260 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 16008 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13892 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11776 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11592 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14536 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 17112 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 16928 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14996 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 17296 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 15640 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 16376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 18216 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 16008 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 16376 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 17020 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 18584 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0__A
timestamp 1649977179
transform -1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13708 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 14168 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 14168 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12144 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 10304 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2116 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22
timestamp 1649977179
transform 1 0 3128 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33
timestamp 1649977179
transform 1 0 4140 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49
timestamp 1649977179
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 1649977179
transform 1 0 7084 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_119
timestamp 1649977179
transform 1 0 12052 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_128
timestamp 1649977179
transform 1 0 12880 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_135
timestamp 1649977179
transform 1 0 13524 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_185
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_30
timestamp 1649977179
transform 1 0 3864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_47
timestamp 1649977179
transform 1 0 5428 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_50
timestamp 1649977179
transform 1 0 5704 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_80
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_104
timestamp 1649977179
transform 1 0 10672 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_149
timestamp 1649977179
transform 1 0 14812 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_53
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_91
timestamp 1649977179
transform 1 0 9476 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_98
timestamp 1649977179
transform 1 0 10120 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_108
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_159
timestamp 1649977179
transform 1 0 15732 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_177
timestamp 1649977179
transform 1 0 17388 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_16
timestamp 1649977179
transform 1 0 2576 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_67
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_108
timestamp 1649977179
transform 1 0 11040 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_159
timestamp 1649977179
transform 1 0 15732 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_7
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_38
timestamp 1649977179
transform 1 0 4600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_66
timestamp 1649977179
transform 1 0 7176 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_76
timestamp 1649977179
transform 1 0 8096 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_129
timestamp 1649977179
transform 1 0 12972 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_102
timestamp 1649977179
transform 1 0 10488 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_5
timestamp 1649977179
transform 1 0 1564 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_21
timestamp 1649977179
transform 1 0 3036 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_40
timestamp 1649977179
transform 1 0 4784 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_70 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7544 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_144
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_164
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_65 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_73
timestamp 1649977179
transform 1 0 7820 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_106 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10856 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_145
timestamp 1649977179
transform 1 0 14444 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_185
timestamp 1649977179
transform 1 0 18124 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_44
timestamp 1649977179
transform 1 0 5152 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_86 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9016 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_98
timestamp 1649977179
transform 1 0 10120 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_102
timestamp 1649977179
transform 1 0 10488 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_115 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_119
timestamp 1649977179
transform 1 0 12052 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_141
timestamp 1649977179
transform 1 0 14076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_17
timestamp 1649977179
transform 1 0 2668 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_37
timestamp 1649977179
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_67
timestamp 1649977179
transform 1 0 7268 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1649977179
transform 1 0 9476 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_101
timestamp 1649977179
transform 1 0 10396 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_185
timestamp 1649977179
transform 1 0 18124 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_33
timestamp 1649977179
transform 1 0 4140 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_37
timestamp 1649977179
transform 1 0 4508 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_63
timestamp 1649977179
transform 1 0 6900 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_80
timestamp 1649977179
transform 1 0 8464 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_15_94 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9752 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_106
timestamp 1649977179
transform 1 0 10856 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_144
timestamp 1649977179
transform 1 0 14352 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_46
timestamp 1649977179
transform 1 0 5336 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_118
timestamp 1649977179
transform 1 0 11960 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_122
timestamp 1649977179
transform 1 0 12328 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_170
timestamp 1649977179
transform 1 0 16744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_13
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_29
timestamp 1649977179
transform 1 0 3772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_46
timestamp 1649977179
transform 1 0 5336 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_73
timestamp 1649977179
transform 1 0 7820 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_87
timestamp 1649977179
transform 1 0 9108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_99
timestamp 1649977179
transform 1 0 10212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_165
timestamp 1649977179
transform 1 0 16284 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_42
timestamp 1649977179
transform 1 0 4968 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_59
timestamp 1649977179
transform 1 0 6532 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_71
timestamp 1649977179
transform 1 0 7636 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_169
timestamp 1649977179
transform 1 0 16652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_23
timestamp 1649977179
transform 1 0 3220 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_59
timestamp 1649977179
transform 1 0 6532 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_71
timestamp 1649977179
transform 1 0 7636 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_83
timestamp 1649977179
transform 1 0 8740 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_95
timestamp 1649977179
transform 1 0 9844 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_107
timestamp 1649977179
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_64
timestamp 1649977179
transform 1 0 6992 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_76
timestamp 1649977179
transform 1 0 8096 0 1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_33
timestamp 1649977179
transform 1 0 4140 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_71
timestamp 1649977179
transform 1 0 7636 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_83
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_95
timestamp 1649977179
transform 1 0 9844 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1649977179
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_133
timestamp 1649977179
transform 1 0 13340 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_139
timestamp 1649977179
transform 1 0 13892 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_21_148
timestamp 1649977179
transform 1 0 14720 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_157
timestamp 1649977179
transform 1 0 15548 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_23
timestamp 1649977179
transform 1 0 3220 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_61
timestamp 1649977179
transform 1 0 6716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_66
timestamp 1649977179
transform 1 0 7176 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_79
timestamp 1649977179
transform 1 0 8372 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_93
timestamp 1649977179
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_100
timestamp 1649977179
transform 1 0 10304 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_107
timestamp 1649977179
transform 1 0 10948 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_111
timestamp 1649977179
transform 1 0 11316 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_128
timestamp 1649977179
transform 1 0 12880 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_135
timestamp 1649977179
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_169
timestamp 1649977179
transform 1 0 16652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 16560 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _18_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1649977179
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1649977179
transform 1 0 2116 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1649977179
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1649977179
transform 1 0 2392 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1649977179
transform 1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1649977179
transform 1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1649977179
transform 1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1649977179
transform 1 0 1748 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1649977179
transform 1 0 4048 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1649977179
transform 1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1649977179
transform 1 0 4324 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1649977179
transform -1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp 1649977179
transform 1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1649977179
transform 1 0 2392 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1649977179
transform -1 0 11960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1649977179
transform -1 0 17480 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1649977179
transform -1 0 15824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1649977179
transform -1 0 16192 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1649977179
transform -1 0 15180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1649977179
transform -1 0 15548 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1649977179
transform -1 0 16100 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1649977179
transform -1 0 10120 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1649977179
transform -1 0 12512 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1649977179
transform -1 0 13892 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1649977179
transform -1 0 13984 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1649977179
transform -1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1649977179
transform -1 0 16560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1649977179
transform -1 0 16376 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1649977179
transform -1 0 17664 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1649977179
transform -1 0 13984 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1649977179
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1649977179
transform -1 0 16560 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1649977179
transform -1 0 16560 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1649977179
transform -1 0 6256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1649977179
transform -1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1649977179
transform -1 0 6900 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1649977179
transform -1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1649977179
transform -1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1649977179
transform -1 0 8740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1649977179
transform 1 0 9936 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1649977179
transform -1 0 10672 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1649977179
transform -1 0 10488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform -1 0 13616 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform -1 0 12788 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform -1 0 12236 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform -1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform -1 0 13340 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform 1 0 16468 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform -1 0 11408 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform 1 0 16192 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform 1 0 13616 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform 1 0 14444 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1649977179
transform 1 0 15272 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1649977179
transform 1 0 15732 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1649977179
transform 1 0 5980 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp 1649977179
transform -1 0 3772 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp 1649977179
transform 1 0 5704 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1649977179
transform 1 0 4600 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1649977179
transform 1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _83_
timestamp 1649977179
transform -1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _84_
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _85_
timestamp 1649977179
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _86_
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8740 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk_0_N_in
timestamp 1649977179
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk_0_N_in
timestamp 1649977179
transform -1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk_0_N_in
timestamp 1649977179
transform 1 0 5244 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1649977179
transform -1 0 9200 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1649977179
transform 1 0 7912 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1649977179
transform -1 0 7636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1649977179
transform -1 0 9660 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1649977179
transform 1 0 10304 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1649977179
transform 1 0 11592 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1649977179
transform 1 0 7912 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1649977179
transform 1 0 9016 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1649977179
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1649977179
transform 1 0 1656 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1649977179
transform 1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1649977179
transform 1 0 4600 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1649977179
transform 1 0 10672 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1649977179
transform 1 0 8372 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7452 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 6256 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 3312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1649977179
transform -1 0 2300 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform -1 0 2300 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1649977179
transform -1 0 3220 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1649977179
transform -1 0 3220 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1649977179
transform -1 0 3220 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1649977179
transform -1 0 4692 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1649977179
transform -1 0 3220 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1649977179
transform -1 0 4140 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1649977179
transform -1 0 5612 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 2668 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1649977179
transform -1 0 2300 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1649977179
transform -1 0 2300 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 3128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform -1 0 2300 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform 1 0 16192 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1649977179
transform 1 0 17664 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1649977179
transform -1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1649977179
transform 1 0 17664 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1649977179
transform 1 0 16744 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1649977179
transform 1 0 16744 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1649977179
transform -1 0 16560 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1649977179
transform -1 0 17664 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1649977179
transform -1 0 16560 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1649977179
transform -1 0 15640 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input36
timestamp 1649977179
transform 1 0 17664 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform -1 0 18584 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1649977179
transform 1 0 17664 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1649977179
transform 1 0 17664 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1649977179
transform -1 0 17664 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1649977179
transform 1 0 17664 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1649977179
transform 1 0 17664 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1649977179
transform 1 0 17664 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 11776 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1649977179
transform -1 0 11408 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1649977179
transform -1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform -1 0 13064 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform 1 0 13248 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1649977179
transform -1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform -1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1649977179
transform -1 0 15456 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform 1 0 15732 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform 1 0 11960 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform -1 0 12880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform -1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform -1 0 14352 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1649977179
transform -1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform -1 0 10304 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform -1 0 10948 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform -1 0 11776 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10672 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7820 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10672 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 9660 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 9752 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__1.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6440 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 13432 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 6900 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 12144 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__2.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5428 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 7636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__3.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6440 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 12512 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 12788 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 8924 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__4.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 12788 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 13248 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform -1 0 10304 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 12052 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__5.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8280 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform -1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 14168 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 9568 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 14720 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__6.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform 1 0 14444 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 16100 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__7.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10120 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR
timestamp 1649977179
transform -1 0 15732 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE
timestamp 1649977179
transform 1 0 15272 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE
timestamp 1649977179
transform 1 0 10672 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__ebufn_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 15548 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__8.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12236 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3956 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 5336 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 6164 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 4048 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7820 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5244 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 3036 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3956 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 3312 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 5336 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5060 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8188 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6992 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9016 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8096 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11040 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12880 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10580 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 13064 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14260 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14812 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 13800 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16192 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14536 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 14168 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13984 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11960 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10396 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4508 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4600 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4600 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4416 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3772 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_0.mux_l2_in_3__149 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2852 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5244 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4876 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4600 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2668 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_1.mux_l2_in_3__150
timestamp 1649977179
transform 1 0 3128 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2668 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2208 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2208 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3220 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4048 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3220 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2760 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2392 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 4600 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform -1 0 4600 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_2.mux_l2_in_3__151
timestamp 1649977179
transform -1 0 3496 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2300 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4784 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2484 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3220 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6440 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5612 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 5428 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_3.mux_l2_in_3__152
timestamp 1649977179
transform 1 0 6256 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5428 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4784 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4600 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4508 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9200 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9016 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform -1 0 8096 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_4.mux_l2_in_3__153
timestamp 1649977179
transform -1 0 8464 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8004 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8648 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13340 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12512 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12512 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12788 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12880 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_5.mux_l2_in_3__154
timestamp 1649977179
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 13064 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12788 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 12880 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2668 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17572 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16744 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17020 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16192 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform 1 0 17112 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_6.mux_l2_in_3__155
timestamp 1649977179
transform 1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15548 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14720 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16744 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17572 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform -1 0 17296 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform -1 0 17664 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_7.mux_l2_in_3__156
timestamp 1649977179
transform 1 0 17848 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17296 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform 1 0 17020 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform 1 0 15180 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12880 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform -1 0 12972 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 13156 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12144 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 10488 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_8.mux_l2_in_3__157
timestamp 1649977179
transform -1 0 11224 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11316 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10028 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9568 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4876 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output63 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform 1 0 6808 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 3588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 2116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 5612 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 3220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform -1 0 2116 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform -1 0 2116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 2116 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform -1 0 1748 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 2116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 2116 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform -1 0 3036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 3220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform -1 0 1748 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 2116 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 1748 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform 1 0 17848 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 16192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 17848 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform 1 0 18216 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform -1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform 1 0 18216 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform 1 0 18216 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform 1 0 17112 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform 1 0 16744 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform 1 0 17848 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform 1 0 18216 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform 1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform 1 0 17480 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform 1 0 18216 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform 1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform 1 0 7176 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1649977179
transform 1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform -1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform 1 0 9016 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform -1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform -1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform 1 0 16008 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform 1 0 18216 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform -1 0 16560 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform 1 0 15824 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform -1 0 15272 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output133
timestamp 1649977179
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1649977179
transform -1 0 3680 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1649977179
transform -1 0 4600 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1649977179
transform -1 0 5244 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1649977179
transform -1 0 5980 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1649977179
transform -1 0 5980 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1649977179
transform 1 0 6348 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1649977179
transform -1 0 5612 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1649977179
transform -1 0 5704 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1649977179
transform -1 0 3588 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7728 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2668 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  repeater143
timestamp 1649977179
transform 1 0 4140 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater144
timestamp 1649977179
transform 1 0 12972 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater145
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater146
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater147
timestamp 1649977179
transform -1 0 8924 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater148
timestamp 1649977179
transform 1 0 6992 0 1 4352
box -38 -48 314 592
<< labels >>
rlabel metal2 s 7378 16400 7434 17200 6 IO_ISOL_N
port 0 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 SC_IN_BOT
port 1 nsew signal input
rlabel metal2 s 6090 16400 6146 17200 6 SC_IN_TOP
port 2 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 SC_OUT_BOT
port 3 nsew signal tristate
rlabel metal2 s 6734 16400 6790 17200 6 SC_OUT_TOP
port 4 nsew signal tristate
rlabel metal4 s 5392 2128 5712 14736 6 VGND
port 5 nsew ground input
rlabel metal4 s 9840 2128 10160 14736 6 VGND
port 5 nsew ground input
rlabel metal4 s 14288 2128 14608 14736 6 VGND
port 5 nsew ground input
rlabel metal4 s 3168 2128 3488 14736 6 VPWR
port 6 nsew power input
rlabel metal4 s 7616 2128 7936 14736 6 VPWR
port 6 nsew power input
rlabel metal4 s 12064 2128 12384 14736 6 VPWR
port 6 nsew power input
rlabel metal4 s 16512 2128 16832 14736 6 VPWR
port 6 nsew power input
rlabel metal2 s 202 0 258 800 6 bottom_grid_pin_0_
port 7 nsew signal tristate
rlabel metal2 s 2686 0 2742 800 6 bottom_grid_pin_10_
port 8 nsew signal tristate
rlabel metal2 s 3146 0 3202 800 6 bottom_grid_pin_12_
port 9 nsew signal tristate
rlabel metal2 s 3606 0 3662 800 6 bottom_grid_pin_14_
port 10 nsew signal tristate
rlabel metal2 s 4158 0 4214 800 6 bottom_grid_pin_16_
port 11 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 bottom_grid_pin_2_
port 12 nsew signal tristate
rlabel metal2 s 1122 0 1178 800 6 bottom_grid_pin_4_
port 13 nsew signal tristate
rlabel metal2 s 1674 0 1730 800 6 bottom_grid_pin_6_
port 14 nsew signal tristate
rlabel metal2 s 2134 0 2190 800 6 bottom_grid_pin_8_
port 15 nsew signal tristate
rlabel metal2 s 4618 0 4674 800 6 ccff_head
port 16 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 ccff_tail
port 17 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 chanx_left_in[0]
port 18 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_in[10]
port 19 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 chanx_left_in[11]
port 20 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 chanx_left_in[12]
port 21 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 chanx_left_in[13]
port 22 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 chanx_left_in[14]
port 23 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 chanx_left_in[15]
port 24 nsew signal input
rlabel metal3 s 0 15512 800 15632 6 chanx_left_in[16]
port 25 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 chanx_left_in[17]
port 26 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 chanx_left_in[18]
port 27 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 chanx_left_in[19]
port 28 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 chanx_left_in[1]
port 29 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[2]
port 30 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[3]
port 31 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 chanx_left_in[4]
port 32 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[5]
port 33 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[6]
port 34 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[7]
port 35 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[8]
port 36 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[9]
port 37 nsew signal input
rlabel metal3 s 0 552 800 672 6 chanx_left_out[0]
port 38 nsew signal tristate
rlabel metal3 s 0 4632 800 4752 6 chanx_left_out[10]
port 39 nsew signal tristate
rlabel metal3 s 0 5040 800 5160 6 chanx_left_out[11]
port 40 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 chanx_left_out[12]
port 41 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 chanx_left_out[13]
port 42 nsew signal tristate
rlabel metal3 s 0 6400 800 6520 6 chanx_left_out[14]
port 43 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 chanx_left_out[15]
port 44 nsew signal tristate
rlabel metal3 s 0 7216 800 7336 6 chanx_left_out[16]
port 45 nsew signal tristate
rlabel metal3 s 0 7624 800 7744 6 chanx_left_out[17]
port 46 nsew signal tristate
rlabel metal3 s 0 8032 800 8152 6 chanx_left_out[18]
port 47 nsew signal tristate
rlabel metal3 s 0 8440 800 8560 6 chanx_left_out[19]
port 48 nsew signal tristate
rlabel metal3 s 0 960 800 1080 6 chanx_left_out[1]
port 49 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 chanx_left_out[2]
port 50 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 chanx_left_out[3]
port 51 nsew signal tristate
rlabel metal3 s 0 2184 800 2304 6 chanx_left_out[4]
port 52 nsew signal tristate
rlabel metal3 s 0 2592 800 2712 6 chanx_left_out[5]
port 53 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 chanx_left_out[6]
port 54 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 chanx_left_out[7]
port 55 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 chanx_left_out[8]
port 56 nsew signal tristate
rlabel metal3 s 0 4224 800 4344 6 chanx_left_out[9]
port 57 nsew signal tristate
rlabel metal3 s 19200 8712 20000 8832 6 chanx_right_in[0]
port 58 nsew signal input
rlabel metal3 s 19200 12928 20000 13048 6 chanx_right_in[10]
port 59 nsew signal input
rlabel metal3 s 19200 13336 20000 13456 6 chanx_right_in[11]
port 60 nsew signal input
rlabel metal3 s 19200 13744 20000 13864 6 chanx_right_in[12]
port 61 nsew signal input
rlabel metal3 s 19200 14152 20000 14272 6 chanx_right_in[13]
port 62 nsew signal input
rlabel metal3 s 19200 14696 20000 14816 6 chanx_right_in[14]
port 63 nsew signal input
rlabel metal3 s 19200 15104 20000 15224 6 chanx_right_in[15]
port 64 nsew signal input
rlabel metal3 s 19200 15512 20000 15632 6 chanx_right_in[16]
port 65 nsew signal input
rlabel metal3 s 19200 15920 20000 16040 6 chanx_right_in[17]
port 66 nsew signal input
rlabel metal3 s 19200 16328 20000 16448 6 chanx_right_in[18]
port 67 nsew signal input
rlabel metal3 s 19200 16736 20000 16856 6 chanx_right_in[19]
port 68 nsew signal input
rlabel metal3 s 19200 9120 20000 9240 6 chanx_right_in[1]
port 69 nsew signal input
rlabel metal3 s 19200 9528 20000 9648 6 chanx_right_in[2]
port 70 nsew signal input
rlabel metal3 s 19200 9936 20000 10056 6 chanx_right_in[3]
port 71 nsew signal input
rlabel metal3 s 19200 10344 20000 10464 6 chanx_right_in[4]
port 72 nsew signal input
rlabel metal3 s 19200 10752 20000 10872 6 chanx_right_in[5]
port 73 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 chanx_right_in[6]
port 74 nsew signal input
rlabel metal3 s 19200 11704 20000 11824 6 chanx_right_in[7]
port 75 nsew signal input
rlabel metal3 s 19200 12112 20000 12232 6 chanx_right_in[8]
port 76 nsew signal input
rlabel metal3 s 19200 12520 20000 12640 6 chanx_right_in[9]
port 77 nsew signal input
rlabel metal3 s 19200 144 20000 264 6 chanx_right_out[0]
port 78 nsew signal tristate
rlabel metal3 s 19200 4360 20000 4480 6 chanx_right_out[10]
port 79 nsew signal tristate
rlabel metal3 s 19200 4768 20000 4888 6 chanx_right_out[11]
port 80 nsew signal tristate
rlabel metal3 s 19200 5176 20000 5296 6 chanx_right_out[12]
port 81 nsew signal tristate
rlabel metal3 s 19200 5584 20000 5704 6 chanx_right_out[13]
port 82 nsew signal tristate
rlabel metal3 s 19200 6128 20000 6248 6 chanx_right_out[14]
port 83 nsew signal tristate
rlabel metal3 s 19200 6536 20000 6656 6 chanx_right_out[15]
port 84 nsew signal tristate
rlabel metal3 s 19200 6944 20000 7064 6 chanx_right_out[16]
port 85 nsew signal tristate
rlabel metal3 s 19200 7352 20000 7472 6 chanx_right_out[17]
port 86 nsew signal tristate
rlabel metal3 s 19200 7760 20000 7880 6 chanx_right_out[18]
port 87 nsew signal tristate
rlabel metal3 s 19200 8168 20000 8288 6 chanx_right_out[19]
port 88 nsew signal tristate
rlabel metal3 s 19200 552 20000 672 6 chanx_right_out[1]
port 89 nsew signal tristate
rlabel metal3 s 19200 960 20000 1080 6 chanx_right_out[2]
port 90 nsew signal tristate
rlabel metal3 s 19200 1368 20000 1488 6 chanx_right_out[3]
port 91 nsew signal tristate
rlabel metal3 s 19200 1776 20000 1896 6 chanx_right_out[4]
port 92 nsew signal tristate
rlabel metal3 s 19200 2184 20000 2304 6 chanx_right_out[5]
port 93 nsew signal tristate
rlabel metal3 s 19200 2592 20000 2712 6 chanx_right_out[6]
port 94 nsew signal tristate
rlabel metal3 s 19200 3136 20000 3256 6 chanx_right_out[7]
port 95 nsew signal tristate
rlabel metal3 s 19200 3544 20000 3664 6 chanx_right_out[8]
port 96 nsew signal tristate
rlabel metal3 s 19200 3952 20000 4072 6 chanx_right_out[9]
port 97 nsew signal tristate
rlabel metal2 s 6642 0 6698 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[0]
port 98 nsew signal tristate
rlabel metal2 s 7102 0 7158 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[1]
port 99 nsew signal tristate
rlabel metal2 s 7654 0 7710 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[2]
port 100 nsew signal tristate
rlabel metal2 s 8114 0 8170 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[3]
port 101 nsew signal tristate
rlabel metal2 s 8666 0 8722 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[4]
port 102 nsew signal tristate
rlabel metal2 s 9126 0 9182 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[5]
port 103 nsew signal tristate
rlabel metal2 s 9678 0 9734 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[6]
port 104 nsew signal tristate
rlabel metal2 s 10138 0 10194 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[7]
port 105 nsew signal tristate
rlabel metal2 s 10598 0 10654 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR[8]
port 106 nsew signal tristate
rlabel metal2 s 11150 0 11206 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[0]
port 107 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[1]
port 108 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[2]
port 109 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[3]
port 110 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[4]
port 111 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[5]
port 112 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[6]
port 113 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[7]
port 114 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN[8]
port 115 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[0]
port 116 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[1]
port 117 nsew signal tristate
rlabel metal2 s 16670 0 16726 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[2]
port 118 nsew signal tristate
rlabel metal2 s 17130 0 17186 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[3]
port 119 nsew signal tristate
rlabel metal2 s 17590 0 17646 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[4]
port 120 nsew signal tristate
rlabel metal2 s 18142 0 18198 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[5]
port 121 nsew signal tristate
rlabel metal2 s 18602 0 18658 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[6]
port 122 nsew signal tristate
rlabel metal2 s 19154 0 19210 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[7]
port 123 nsew signal tristate
rlabel metal2 s 19614 0 19670 800 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT[8]
port 124 nsew signal tristate
rlabel metal2 s 8022 16400 8078 17200 6 prog_clk_0_N_in
port 125 nsew signal input
rlabel metal3 s 0 144 800 264 6 prog_clk_0_W_out
port 126 nsew signal tristate
rlabel metal2 s 8666 16400 8722 17200 6 top_width_0_height_0__pin_0_
port 127 nsew signal input
rlabel metal2 s 11886 16400 11942 17200 6 top_width_0_height_0__pin_10_
port 128 nsew signal input
rlabel metal2 s 14462 16400 14518 17200 6 top_width_0_height_0__pin_11_lower
port 129 nsew signal tristate
rlabel metal2 s 3514 16400 3570 17200 6 top_width_0_height_0__pin_11_upper
port 130 nsew signal tristate
rlabel metal2 s 12530 16400 12586 17200 6 top_width_0_height_0__pin_12_
port 131 nsew signal input
rlabel metal2 s 15106 16400 15162 17200 6 top_width_0_height_0__pin_13_lower
port 132 nsew signal tristate
rlabel metal2 s 4158 16400 4214 17200 6 top_width_0_height_0__pin_13_upper
port 133 nsew signal tristate
rlabel metal2 s 13174 16400 13230 17200 6 top_width_0_height_0__pin_14_
port 134 nsew signal input
rlabel metal2 s 15750 16400 15806 17200 6 top_width_0_height_0__pin_15_lower
port 135 nsew signal tristate
rlabel metal2 s 4802 16400 4858 17200 6 top_width_0_height_0__pin_15_upper
port 136 nsew signal tristate
rlabel metal2 s 13818 16400 13874 17200 6 top_width_0_height_0__pin_16_
port 137 nsew signal input
rlabel metal2 s 16394 16400 16450 17200 6 top_width_0_height_0__pin_17_lower
port 138 nsew signal tristate
rlabel metal2 s 5446 16400 5502 17200 6 top_width_0_height_0__pin_17_upper
port 139 nsew signal tristate
rlabel metal2 s 17038 16400 17094 17200 6 top_width_0_height_0__pin_1_lower
port 140 nsew signal tristate
rlabel metal2 s 294 16400 350 17200 6 top_width_0_height_0__pin_1_upper
port 141 nsew signal tristate
rlabel metal2 s 9310 16400 9366 17200 6 top_width_0_height_0__pin_2_
port 142 nsew signal input
rlabel metal2 s 17682 16400 17738 17200 6 top_width_0_height_0__pin_3_lower
port 143 nsew signal tristate
rlabel metal2 s 938 16400 994 17200 6 top_width_0_height_0__pin_3_upper
port 144 nsew signal tristate
rlabel metal2 s 9954 16400 10010 17200 6 top_width_0_height_0__pin_4_
port 145 nsew signal input
rlabel metal2 s 18326 16400 18382 17200 6 top_width_0_height_0__pin_5_lower
port 146 nsew signal tristate
rlabel metal2 s 1582 16400 1638 17200 6 top_width_0_height_0__pin_5_upper
port 147 nsew signal tristate
rlabel metal2 s 10598 16400 10654 17200 6 top_width_0_height_0__pin_6_
port 148 nsew signal input
rlabel metal2 s 18970 16400 19026 17200 6 top_width_0_height_0__pin_7_lower
port 149 nsew signal tristate
rlabel metal2 s 2226 16400 2282 17200 6 top_width_0_height_0__pin_7_upper
port 150 nsew signal tristate
rlabel metal2 s 11242 16400 11298 17200 6 top_width_0_height_0__pin_8_
port 151 nsew signal input
rlabel metal2 s 19614 16400 19670 17200 6 top_width_0_height_0__pin_9_lower
port 152 nsew signal tristate
rlabel metal2 s 2870 16400 2926 17200 6 top_width_0_height_0__pin_9_upper
port 153 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
