* NGSPICE file created from cby_0__1_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_1 abstract view
.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_8 abstract view
.subckt sky130_fd_sc_hd__ebufn_8 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

.subckt cby_0__1_ IO_ISOL_N VGND VPWR ccff_head ccff_tail chany_bottom_in[0] chany_bottom_in[10]
+ chany_bottom_in[11] chany_bottom_in[12] chany_bottom_in[13] chany_bottom_in[14]
+ chany_bottom_in[15] chany_bottom_in[16] chany_bottom_in[17] chany_bottom_in[18]
+ chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2] chany_bottom_in[3] chany_bottom_in[4]
+ chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7] chany_bottom_in[8] chany_bottom_in[9]
+ chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11] chany_bottom_out[12]
+ chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15] chany_bottom_out[16]
+ chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19] chany_bottom_out[1]
+ chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4] chany_bottom_out[5]
+ chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8] chany_bottom_out[9]
+ chany_top_in[0] chany_top_in[10] chany_top_in[11] chany_top_in[12] chany_top_in[13]
+ chany_top_in[14] chany_top_in[15] chany_top_in[16] chany_top_in[17] chany_top_in[18]
+ chany_top_in[19] chany_top_in[1] chany_top_in[2] chany_top_in[3] chany_top_in[4]
+ chany_top_in[5] chany_top_in[6] chany_top_in[7] chany_top_in[8] chany_top_in[9]
+ chany_top_out[0] chany_top_out[10] chany_top_out[11] chany_top_out[12] chany_top_out[13]
+ chany_top_out[14] chany_top_out[15] chany_top_out[16] chany_top_out[17] chany_top_out[18]
+ chany_top_out[19] chany_top_out[1] chany_top_out[2] chany_top_out[3] chany_top_out[4]
+ chany_top_out[5] chany_top_out[6] chany_top_out[7] chany_top_out[8] chany_top_out[9]
+ gfpga_pad_EMBEDDED_IO_HD_SOC_DIR gfpga_pad_EMBEDDED_IO_HD_SOC_IN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
+ left_grid_pin_0_ prog_clk_0_E_in right_width_0_height_0__pin_0_ right_width_0_height_0__pin_1_lower
+ right_width_0_height_0__pin_1_upper
XFILLER_22_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input18_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput75 _19_/X VGND VGND VPWR VPWR chany_top_out[18] sky130_fd_sc_hd__buf_2
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput53 _38_/X VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
Xoutput64 _30_/X VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
Xoutput86 output86/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_DIR sky130_fd_sc_hd__buf_2
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput76 _20_/X VGND VGND VPWR VPWR chany_top_out[19] sky130_fd_sc_hd__buf_2
XANTENNA_input30_A chany_top_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput54 _39_/X VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
Xoutput65 _31_/X VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
Xoutput87 output87/A VGND VGND VPWR VPWR left_grid_pin_0_ sky130_fd_sc_hd__buf_2
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_87 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_68 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput88 _21_/X VGND VGND VPWR VPWR right_width_0_height_0__pin_1_upper sky130_fd_sc_hd__buf_2
XANTENNA_input23_A chany_top_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput66 _42_/X VGND VGND VPWR VPWR chany_top_out[0] sky130_fd_sc_hd__buf_2
Xoutput77 _02_/X VGND VGND VPWR VPWR chany_top_out[1] sky130_fd_sc_hd__buf_2
XFILLER_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput55 _40_/X VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xprog_clk_0_FTB00 prog_clk_0_E_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
X_29_ _29_/A VGND VGND VPWR VPWR _29_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput67 _11_/X VGND VGND VPWR VPWR chany_top_out[10] sky130_fd_sc_hd__buf_2
Xoutput78 _03_/X VGND VGND VPWR VPWR chany_top_out[2] sky130_fd_sc_hd__buf_2
Xoutput45 output45/A VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_2
XFILLER_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput56 _41_/X VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input16_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input8_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_28_ _28_/A VGND VGND VPWR VPWR _28_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput46 _22_/X VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
Xoutput57 _23_/X VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
Xoutput68 _12_/X VGND VGND VPWR VPWR chany_top_out[11] sky130_fd_sc_hd__buf_2
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput79 _04_/X VGND VGND VPWR VPWR chany_top_out[3] sky130_fd_sc_hd__buf_2
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input39_A chany_top_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_27_ _27_/A VGND VGND VPWR VPWR _27_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput69 _13_/X VGND VGND VPWR VPWR chany_top_out[12] sky130_fd_sc_hd__buf_2
Xoutput47 _32_/X VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
Xoutput58 _24_/X VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input21_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_49 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_40 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_26_ _26_/A VGND VGND VPWR VPWR _26_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_09_ _09_/A VGND VGND VPWR VPWR _09_/X sky130_fd_sc_hd__clkbuf_1
Xoutput48 _33_/X VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
Xoutput59 _25_/X VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input14_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_ mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_right_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_input6_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR output86/A
+ VGND VGND VPWR VPWR logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y
+ sky130_fd_sc_hd__inv_1
XFILLER_23_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_42_ _42_/A VGND VGND VPWR VPWR _42_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25_ _25_/A VGND VGND VPWR VPWR _25_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input44_A right_width_0_height_0__pin_0_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_08_ _08_/A VGND VGND VPWR VPWR _08_/X sky130_fd_sc_hd__clkbuf_1
Xoutput49 _34_/X VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_ mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_right_ipin_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l3_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_41_ _41_/A VGND VGND VPWR VPWR _41_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24_ _24_/A VGND VGND VPWR VPWR _24_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input37_A chany_top_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_ipin_0.mux_l2_in_3__89 VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_3_/A0
+ mux_right_ipin_0.mux_l2_in_3__89/LO sky130_fd_sc_hd__conb_1
X_07_ _07_/A VGND VGND VPWR VPWR _07_/X sky130_fd_sc_hd__clkbuf_1
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_ mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK
+ mux_right_ipin_0.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_3_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_12_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_40_ _40_/A VGND VGND VPWR VPWR _40_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_23_ _23_/A VGND VGND VPWR VPWR _23_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_06_ _06_/A VGND VGND VPWR VPWR _06_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK
+ input2/X VGND VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_27_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input12_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_96 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input4_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_22_ _22_/A VGND VGND VPWR VPWR _22_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_05_ _05_/A VGND VGND VPWR VPWR _05_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE input43/X
+ logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR/Y VGND
+ VGND VPWR VPWR right_width_0_height_0__pin_1_lower sky130_fd_sc_hd__ebufn_8
XANTENNA_input42_A chany_top_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_21_ right_width_0_height_0__pin_1_lower VGND VGND VPWR VPWR _21_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_04_ _04_/A VGND VGND VPWR VPWR _04_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input35_A chany_top_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_20_ _20_/A VGND VGND VPWR VPWR _20_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput1 IO_ISOL_N VGND VGND VPWR VPWR input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_03_ _03_/A VGND VGND VPWR VPWR _03_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input28_A chany_top_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input10_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input2_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput2 ccff_head VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__clkbuf_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_02_ _02_/A VGND VGND VPWR VPWR _02_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_24_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input40_A chany_top_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_ mux_right_ipin_0.mux_l4_in_0_/X VGND VGND
+ VPWR VPWR output87/A sky130_fd_sc_hd__clkbuf_1
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 chany_bottom_in[0] VGND VGND VPWR VPWR _42_/A sky130_fd_sc_hd__clkbuf_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_8 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_E_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input33_A chany_top_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_24 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_16 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 chany_bottom_in[10] VGND VGND VPWR VPWR _11_/A sky130_fd_sc_hd__clkbuf_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput40 chany_top_in[7] VGND VGND VPWR VPWR _29_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_21_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input26_A chany_top_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__21__A right_width_0_height_0__pin_1_lower VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_0.mux_l2_in_3_ mux_right_ipin_0.mux_l2_in_3_/A0 _38_/A mux_right_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_3_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_36 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_28 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput5 chany_bottom_in[11] VGND VGND VPWR VPWR _12_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_right_ipin_0.mux_l4_in_0_ mux_right_ipin_0.mux_l3_in_1_/X mux_right_ipin_0.mux_l3_in_0_/X
+ hold1/A VGND VGND VPWR VPWR mux_right_ipin_0.mux_l4_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_27 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput30 chany_top_in[16] VGND VGND VPWR VPWR _38_/A sky130_fd_sc_hd__clkbuf_1
Xinput41 chany_top_in[8] VGND VGND VPWR VPWR _30_/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_0.mux_l3_in_1_ mux_right_ipin_0.mux_l2_in_3_/X mux_right_ipin_0.mux_l2_in_2_/X
+ mux_right_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l3_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_12_106 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input19_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_right_ipin_0.mux_l2_in_2_ _17_/A _32_/A mux_right_ipin_0.mux_l2_in_3_/S VGND
+ VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_1_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_19_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 chany_bottom_in[12] VGND VGND VPWR VPWR _13_/A sky130_fd_sc_hd__clkbuf_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput31 chany_top_in[17] VGND VGND VPWR VPWR _39_/A sky130_fd_sc_hd__clkbuf_1
Xmux_right_ipin_0.mux_l3_in_0_ mux_right_ipin_0.mux_l2_in_1_/X mux_right_ipin_0.mux_l2_in_0_/X
+ mux_right_ipin_0.mux_l3_in_1_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l3_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xinput20 chany_bottom_in[7] VGND VGND VPWR VPWR _08_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_7_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput42 chany_top_in[9] VGND VGND VPWR VPWR _31_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_118 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input31_A chany_top_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_ipin_0.mux_l2_in_1_ _11_/A mux_right_ipin_0.mux_l1_in_2_/X mux_right_ipin_0.mux_l2_in_3_/S
+ VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_right_ipin_0.mux_l1_in_2_ _26_/A _05_/A mux_right_ipin_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xclkbuf_1_0__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ VGND VGND VPWR VPWR mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 chany_bottom_in[13] VGND VGND VPWR VPWR _14_/A sky130_fd_sc_hd__clkbuf_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput32 chany_top_in[18] VGND VGND VPWR VPWR _40_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput43 gfpga_pad_EMBEDDED_IO_HD_SOC_IN VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput21 chany_bottom_in[8] VGND VGND VPWR VPWR _09_/A sky130_fd_sc_hd__clkbuf_1
Xinput10 chany_bottom_in[16] VGND VGND VPWR VPWR _17_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE input44/X
+ output86/A VGND VGND VPWR VPWR gfpga_pad_EMBEDDED_IO_HD_SOC_OUT sky130_fd_sc_hd__ebufn_8
XFILLER_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_0.mux_l2_in_0_ mux_right_ipin_0.mux_l1_in_1_/X mux_right_ipin_0.mux_l1_in_0_/X
+ mux_right_ipin_0.mux_l2_in_3_/S VGND VGND VPWR VPWR mux_right_ipin_0.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input24_A chany_top_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_right_ipin_0.mux_l1_in_1_ _24_/A _03_/A mux_right_ipin_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 chany_bottom_in[14] VGND VGND VPWR VPWR _15_/A sky130_fd_sc_hd__clkbuf_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_39 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput33 chany_top_in[19] VGND VGND VPWR VPWR _41_/A sky130_fd_sc_hd__clkbuf_1
X_39_ _39_/A VGND VGND VPWR VPWR _39_/X sky130_fd_sc_hd__clkbuf_1
Xinput22 chany_bottom_in[9] VGND VGND VPWR VPWR _10_/A sky130_fd_sc_hd__clkbuf_1
Xinput44 right_width_0_height_0__pin_0_ VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_1
Xinput11 chany_bottom_in[17] VGND VGND VPWR VPWR _18_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input17_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input9_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_right_ipin_0.mux_l1_in_0_ _22_/A _42_/A mux_right_ipin_0.mux_l1_in_2_/S VGND
+ VGND VPWR VPWR mux_right_ipin_0.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 chany_bottom_in[15] VGND VGND VPWR VPWR _16_/A sky130_fd_sc_hd__clkbuf_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput34 chany_top_in[1] VGND VGND VPWR VPWR _23_/A sky130_fd_sc_hd__clkbuf_1
Xinput23 chany_top_in[0] VGND VGND VPWR VPWR _22_/A sky130_fd_sc_hd__clkbuf_1
Xinput12 chany_bottom_in[18] VGND VGND VPWR VPWR _19_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_38_ _38_/A VGND VGND VPWR VPWR _38_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput24 chany_top_in[10] VGND VGND VPWR VPWR _32_/A sky130_fd_sc_hd__clkbuf_1
Xinput35 chany_top_in[2] VGND VGND VPWR VPWR _24_/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_14_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput13 chany_bottom_in[19] VGND VGND VPWR VPWR _20_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_37_ _37_/A VGND VGND VPWR VPWR _37_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_7_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input22_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput25 chany_top_in[11] VGND VGND VPWR VPWR _33_/A sky130_fd_sc_hd__clkbuf_1
Xinput36 chany_top_in[3] VGND VGND VPWR VPWR _25_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput14 chany_bottom_in[1] VGND VGND VPWR VPWR _02_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_31 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_36_ _36_/A VGND VGND VPWR VPWR _36_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_22_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_19_ _19_/A VGND VGND VPWR VPWR _19_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input15_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input7_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_43 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput26 chany_top_in[12] VGND VGND VPWR VPWR _34_/A sky130_fd_sc_hd__clkbuf_1
Xinput37 chany_top_in[4] VGND VGND VPWR VPWR _26_/A sky130_fd_sc_hd__clkbuf_1
X_35_ _35_/A VGND VGND VPWR VPWR _35_/X sky130_fd_sc_hd__clkbuf_1
Xinput15 chany_bottom_in[2] VGND VGND VPWR VPWR _03_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
+ mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_/CLK hold1/X VGND VGND VPWR VPWR output45/A
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_18_ _18_/A VGND VGND VPWR VPWR _18_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_4_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_20 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_20 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput27 chany_top_in[13] VGND VGND VPWR VPWR _35_/A sky130_fd_sc_hd__clkbuf_1
Xinput38 chany_top_in[5] VGND VGND VPWR VPWR _27_/A sky130_fd_sc_hd__clkbuf_1
X_34_ _34_/A VGND VGND VPWR VPWR _34_/X sky130_fd_sc_hd__clkbuf_1
Xinput16 chany_bottom_in[3] VGND VGND VPWR VPWR _04_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA_input38_A chany_top_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_17_ _17_/A VGND VGND VPWR VPWR _17_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_17_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input20_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_32 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
+ clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk/X
+ VGND VGND VPWR VPWR mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_7 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput28 chany_top_in[14] VGND VGND VPWR VPWR _36_/A sky130_fd_sc_hd__clkbuf_1
Xinput39 chany_top_in[6] VGND VGND VPWR VPWR _28_/A sky130_fd_sc_hd__clkbuf_1
X_33_ _33_/A VGND VGND VPWR VPWR _33_/X sky130_fd_sc_hd__clkbuf_1
Xinput17 chany_bottom_in[4] VGND VGND VPWR VPWR _05_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_16_ _16_/A VGND VGND VPWR VPWR _16_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_77 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input13_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_44 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input5_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput29 chany_top_in[15] VGND VGND VPWR VPWR _37_/A sky130_fd_sc_hd__clkbuf_1
Xinput18 chany_bottom_in[5] VGND VGND VPWR VPWR _06_/A sky130_fd_sc_hd__clkbuf_1
X_32_ _32_/A VGND VGND VPWR VPWR _32_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_15_ _15_/A VGND VGND VPWR VPWR _15_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_89 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input43_A gfpga_pad_EMBEDDED_IO_HD_SOC_IN VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput19 chany_bottom_in[6] VGND VGND VPWR VPWR _07_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_31_ _31_/A VGND VGND VPWR VPWR _31_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_14_ _14_/A VGND VGND VPWR VPWR _14_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input36_A chany_top_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_91 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_30_ _30_/A VGND VGND VPWR VPWR _30_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13_ _13_/A VGND VGND VPWR VPWR _13_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input29_A chany_top_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input11_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input3_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_15 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_12_ _12_/A VGND VGND VPWR VPWR _12_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_3_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input41_A chany_top_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput80 _05_/X VGND VGND VPWR VPWR chany_top_out[4] sky130_fd_sc_hd__buf_2
XFILLER_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_11_ _11_/A VGND VGND VPWR VPWR _11_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_8_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input34_A chany_top_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput70 _14_/X VGND VGND VPWR VPWR chany_top_out[13] sky130_fd_sc_hd__buf_2
Xoutput81 _06_/X VGND VGND VPWR VPWR chany_top_out[5] sky130_fd_sc_hd__buf_2
XFILLER_7_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xlogical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE output45/A
+ input1/X VGND VGND VPWR VPWR output86/A sky130_fd_sc_hd__or2b_2
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_10_ _10_/A VGND VGND VPWR VPWR _10_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_94 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input27_A chany_top_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_61 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput71 _15_/X VGND VGND VPWR VPWR chany_top_out[14] sky130_fd_sc_hd__buf_2
Xoutput82 _07_/X VGND VGND VPWR VPWR chany_top_out[6] sky130_fd_sc_hd__buf_2
Xoutput60 _26_/X VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_11_19 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_29 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input1_A IO_ISOL_N VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_53 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput72 _16_/X VGND VGND VPWR VPWR chany_top_out[15] sky130_fd_sc_hd__buf_2
Xoutput83 _08_/X VGND VGND VPWR VPWR chany_top_out[7] sky130_fd_sc_hd__buf_2
XFILLER_15_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput50 _35_/X VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
Xoutput61 _27_/X VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input32_A chany_top_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_65 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput73 _17_/X VGND VGND VPWR VPWR chany_top_out[16] sky130_fd_sc_hd__buf_2
Xoutput84 _09_/X VGND VGND VPWR VPWR chany_top_out[8] sky130_fd_sc_hd__buf_2
Xoutput51 _36_/X VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
Xoutput62 _28_/X VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_8 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input25_A chany_top_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_3 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput52 _37_/X VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
Xoutput74 _18_/X VGND VGND VPWR VPWR chany_top_out[17] sky130_fd_sc_hd__buf_2
Xoutput85 _10_/X VGND VGND VPWR VPWR chany_top_out[9] sky130_fd_sc_hd__buf_2
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput63 _29_/X VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
.ends

