magic
tech sky130A
magscale 1 2
timestamp 1650894746
<< viali >>
rect 2237 22185 2271 22219
rect 11345 22185 11379 22219
rect 17877 22185 17911 22219
rect 19257 22185 19291 22219
rect 13185 22117 13219 22151
rect 22017 22117 22051 22151
rect 10977 22049 11011 22083
rect 20085 22049 20119 22083
rect 1685 21981 1719 22015
rect 1777 21981 1811 22015
rect 2329 21981 2363 22015
rect 2697 21981 2731 22015
rect 3249 21981 3283 22015
rect 3341 21981 3375 22015
rect 4077 21981 4111 22015
rect 4445 21981 4479 22015
rect 5457 21981 5491 22015
rect 6193 21981 6227 22015
rect 8217 21981 8251 22015
rect 8309 21981 8343 22015
rect 8585 21981 8619 22015
rect 8953 21981 8987 22015
rect 10333 21981 10367 22015
rect 11621 21981 11655 22015
rect 11897 21981 11931 22015
rect 12173 21981 12207 22015
rect 12633 21981 12667 22015
rect 12817 21981 12851 22015
rect 13921 21981 13955 22015
rect 14105 21981 14139 22015
rect 15577 21981 15611 22015
rect 16313 21981 16347 22015
rect 16865 21981 16899 22015
rect 17601 21981 17635 22015
rect 17693 21981 17727 22015
rect 18061 21981 18095 22015
rect 18797 21981 18831 22015
rect 19441 21981 19475 22015
rect 20637 21981 20671 22015
rect 20913 21981 20947 22015
rect 21649 21981 21683 22015
rect 21833 21981 21867 22015
rect 22385 21981 22419 22015
rect 23121 21981 23155 22015
rect 3985 21913 4019 21947
rect 6561 21913 6595 21947
rect 7972 21913 8006 21947
rect 9597 21913 9631 21947
rect 10793 21913 10827 21947
rect 13001 21913 13035 21947
rect 19993 21913 20027 21947
rect 1501 21845 1535 21879
rect 1961 21845 1995 21879
rect 2513 21845 2547 21879
rect 2881 21845 2915 21879
rect 3065 21845 3099 21879
rect 3525 21845 3559 21879
rect 4261 21845 4295 21879
rect 4629 21845 4663 21879
rect 4813 21845 4847 21879
rect 5549 21845 5583 21879
rect 6469 21845 6503 21879
rect 6837 21845 6871 21879
rect 8493 21845 8527 21879
rect 8769 21845 8803 21879
rect 9689 21845 9723 21879
rect 10425 21845 10459 21879
rect 10885 21845 10919 21879
rect 11805 21845 11839 21879
rect 12081 21845 12115 21879
rect 12357 21845 12391 21879
rect 13277 21845 13311 21879
rect 14749 21845 14783 21879
rect 14933 21845 14967 21879
rect 15669 21845 15703 21879
rect 16405 21845 16439 21879
rect 16681 21845 16715 21879
rect 16957 21845 16991 21879
rect 18705 21845 18739 21879
rect 18981 21845 19015 21879
rect 19533 21845 19567 21879
rect 19901 21845 19935 21879
rect 20453 21845 20487 21879
rect 20729 21845 20763 21879
rect 21005 21845 21039 21879
rect 22201 21845 22235 21879
rect 22477 21845 22511 21879
rect 1501 21641 1535 21675
rect 4813 21641 4847 21675
rect 6837 21641 6871 21675
rect 9413 21641 9447 21675
rect 9965 21641 9999 21675
rect 12449 21641 12483 21675
rect 18061 21641 18095 21675
rect 21281 21641 21315 21675
rect 22753 21641 22787 21675
rect 4997 21573 5031 21607
rect 5181 21573 5215 21607
rect 7542 21573 7576 21607
rect 11100 21573 11134 21607
rect 11529 21573 11563 21607
rect 16948 21573 16982 21607
rect 18420 21573 18454 21607
rect 1685 21505 1719 21539
rect 1777 21505 1811 21539
rect 2881 21505 2915 21539
rect 3700 21505 3734 21539
rect 5365 21505 5399 21539
rect 6193 21505 6227 21539
rect 7297 21505 7331 21539
rect 8861 21505 8895 21539
rect 9321 21505 9355 21539
rect 9597 21505 9631 21539
rect 9689 21505 9723 21539
rect 12173 21505 12207 21539
rect 12265 21505 12299 21539
rect 13185 21505 13219 21539
rect 13645 21505 13679 21539
rect 14289 21505 14323 21539
rect 14556 21505 14590 21539
rect 15761 21505 15795 21539
rect 20749 21505 20783 21539
rect 21097 21505 21131 21539
rect 21649 21505 21683 21539
rect 22477 21505 22511 21539
rect 22569 21505 22603 21539
rect 23121 21505 23155 21539
rect 2605 21437 2639 21471
rect 2789 21437 2823 21471
rect 3433 21437 3467 21471
rect 6561 21437 6595 21471
rect 6745 21437 6779 21471
rect 11345 21437 11379 21471
rect 13369 21437 13403 21471
rect 13553 21437 13587 21471
rect 16681 21437 16715 21471
rect 18153 21437 18187 21471
rect 21005 21437 21039 21471
rect 9045 21369 9079 21403
rect 14105 21369 14139 21403
rect 16405 21369 16439 21403
rect 2421 21301 2455 21335
rect 3249 21301 3283 21335
rect 5549 21301 5583 21335
rect 7205 21301 7239 21335
rect 8677 21301 8711 21335
rect 9137 21301 9171 21335
rect 9873 21301 9907 21335
rect 12541 21301 12575 21335
rect 14013 21301 14047 21335
rect 15669 21301 15703 21335
rect 19533 21301 19567 21335
rect 19625 21301 19659 21335
rect 21465 21301 21499 21335
rect 21833 21301 21867 21335
rect 22937 21301 22971 21335
rect 4261 21097 4295 21131
rect 9597 21097 9631 21131
rect 11437 21097 11471 21131
rect 14105 21097 14139 21131
rect 18981 21097 19015 21131
rect 21373 21097 21407 21131
rect 5733 21029 5767 21063
rect 16957 21029 16991 21063
rect 1593 20961 1627 20995
rect 1685 20961 1719 20995
rect 10057 20961 10091 20995
rect 11529 20961 11563 20995
rect 12541 20961 12575 20995
rect 15485 20961 15519 20995
rect 15577 20961 15611 20995
rect 17233 20961 17267 20995
rect 18061 20961 18095 20995
rect 2237 20893 2271 20927
rect 3801 20893 3835 20927
rect 4353 20893 4387 20927
rect 5917 20893 5951 20927
rect 7297 20893 7331 20927
rect 8769 20893 8803 20927
rect 8953 20893 8987 20927
rect 11805 20893 11839 20927
rect 12808 20893 12842 20927
rect 15844 20893 15878 20927
rect 18245 20893 18279 20927
rect 18797 20893 18831 20927
rect 19901 20893 19935 20927
rect 19993 20893 20027 20927
rect 21465 20893 21499 20927
rect 1777 20825 1811 20859
rect 2493 20825 2527 20859
rect 3985 20825 4019 20859
rect 4620 20825 4654 20859
rect 8502 20825 8536 20859
rect 9689 20825 9723 20859
rect 10302 20825 10336 20859
rect 15240 20825 15274 20859
rect 20238 20825 20272 20859
rect 21710 20825 21744 20859
rect 22937 20825 22971 20859
rect 2145 20757 2179 20791
rect 3617 20757 3651 20791
rect 6561 20757 6595 20791
rect 6653 20757 6687 20791
rect 7389 20757 7423 20791
rect 12449 20757 12483 20791
rect 13921 20757 13955 20791
rect 17325 20757 17359 20791
rect 17417 20757 17451 20791
rect 17785 20757 17819 20791
rect 18153 20757 18187 20791
rect 18613 20757 18647 20791
rect 19257 20757 19291 20791
rect 22845 20757 22879 20791
rect 1777 20553 1811 20587
rect 3709 20553 3743 20587
rect 6193 20553 6227 20587
rect 7757 20553 7791 20587
rect 8217 20553 8251 20587
rect 8769 20553 8803 20587
rect 11897 20553 11931 20587
rect 13553 20553 13587 20587
rect 14013 20553 14047 20587
rect 14565 20553 14599 20587
rect 14933 20553 14967 20587
rect 15669 20553 15703 20587
rect 19349 20553 19383 20587
rect 19717 20553 19751 20587
rect 19993 20553 20027 20587
rect 22845 20553 22879 20587
rect 4721 20485 4755 20519
rect 6622 20485 6656 20519
rect 9229 20485 9263 20519
rect 11161 20485 11195 20519
rect 16865 20485 16899 20519
rect 17049 20485 17083 20519
rect 18245 20485 18279 20519
rect 20514 20485 20548 20519
rect 1501 20417 1535 20451
rect 2890 20417 2924 20451
rect 3157 20417 3191 20451
rect 3617 20417 3651 20451
rect 4077 20417 4111 20451
rect 4813 20417 4847 20451
rect 5080 20417 5114 20451
rect 6377 20417 6411 20451
rect 9689 20417 9723 20451
rect 9956 20417 9990 20451
rect 11713 20417 11747 20451
rect 12081 20417 12115 20451
rect 12173 20417 12207 20451
rect 12440 20417 12474 20451
rect 13829 20417 13863 20451
rect 15025 20417 15059 20451
rect 16129 20417 16163 20451
rect 17233 20417 17267 20451
rect 18889 20417 18923 20451
rect 19809 20417 19843 20451
rect 22201 20417 22235 20451
rect 22661 20417 22695 20451
rect 3893 20349 3927 20383
rect 8309 20349 8343 20383
rect 8401 20349 8435 20383
rect 9321 20349 9355 20383
rect 9505 20349 9539 20383
rect 14381 20349 14415 20383
rect 14473 20349 14507 20383
rect 15945 20349 15979 20383
rect 16037 20349 16071 20383
rect 17509 20349 17543 20383
rect 19165 20349 19199 20383
rect 19257 20349 19291 20383
rect 20269 20349 20303 20383
rect 21925 20349 21959 20383
rect 22109 20349 22143 20383
rect 11529 20281 11563 20315
rect 13645 20281 13679 20315
rect 21649 20281 21683 20315
rect 1685 20213 1719 20247
rect 3249 20213 3283 20247
rect 7849 20213 7883 20247
rect 8861 20213 8895 20247
rect 11069 20213 11103 20247
rect 16497 20213 16531 20247
rect 16681 20213 16715 20247
rect 22569 20213 22603 20247
rect 23029 20213 23063 20247
rect 4445 20009 4479 20043
rect 7205 20009 7239 20043
rect 8033 20009 8067 20043
rect 9781 20009 9815 20043
rect 11345 20009 11379 20043
rect 13737 20009 13771 20043
rect 14105 20009 14139 20043
rect 14933 20009 14967 20043
rect 22661 20009 22695 20043
rect 5089 19941 5123 19975
rect 6745 19941 6779 19975
rect 9873 19941 9907 19975
rect 5273 19873 5307 19907
rect 6101 19873 6135 19907
rect 6837 19873 6871 19907
rect 7757 19873 7791 19907
rect 8677 19873 8711 19907
rect 11253 19873 11287 19907
rect 11897 19873 11931 19907
rect 13093 19873 13127 19907
rect 14565 19873 14599 19907
rect 14657 19873 14691 19907
rect 18705 19873 18739 19907
rect 18889 19873 18923 19907
rect 19720 19873 19754 19907
rect 1501 19805 1535 19839
rect 3617 19805 3651 19839
rect 3801 19805 3835 19839
rect 4629 19805 4663 19839
rect 4905 19805 4939 19839
rect 5457 19805 5491 19839
rect 9137 19805 9171 19839
rect 12817 19805 12851 19839
rect 13369 19805 13403 19839
rect 14473 19805 14507 19839
rect 15577 19805 15611 19839
rect 15669 19805 15703 19839
rect 16405 19805 16439 19839
rect 18153 19805 18187 19839
rect 19257 19805 19291 19839
rect 19993 19805 20027 19839
rect 21189 19805 21223 19839
rect 21445 19805 21479 19839
rect 22845 19805 22879 19839
rect 1768 19737 1802 19771
rect 2973 19737 3007 19771
rect 5549 19737 5583 19771
rect 7021 19737 7055 19771
rect 7665 19737 7699 19771
rect 8493 19737 8527 19771
rect 10986 19737 11020 19771
rect 13277 19737 13311 19771
rect 17908 19737 17942 19771
rect 2881 19669 2915 19703
rect 4813 19669 4847 19703
rect 5917 19669 5951 19703
rect 6285 19669 6319 19703
rect 6377 19669 6411 19703
rect 7573 19669 7607 19703
rect 8401 19669 8435 19703
rect 9045 19669 9079 19703
rect 11713 19669 11747 19703
rect 11805 19669 11839 19703
rect 12173 19669 12207 19703
rect 13921 19669 13955 19703
rect 16313 19669 16347 19703
rect 16589 19669 16623 19703
rect 16773 19669 16807 19703
rect 18245 19669 18279 19703
rect 18613 19669 18647 19703
rect 19723 19669 19757 19703
rect 21097 19669 21131 19703
rect 22569 19669 22603 19703
rect 23029 19669 23063 19703
rect 1593 19465 1627 19499
rect 3065 19465 3099 19499
rect 4813 19465 4847 19499
rect 4905 19465 4939 19499
rect 6377 19465 6411 19499
rect 6929 19465 6963 19499
rect 9137 19465 9171 19499
rect 10057 19465 10091 19499
rect 10333 19465 10367 19499
rect 11345 19465 11379 19499
rect 11989 19465 12023 19499
rect 14381 19465 14415 19499
rect 16957 19465 16991 19499
rect 18981 19465 19015 19499
rect 21833 19465 21867 19499
rect 22293 19465 22327 19499
rect 23029 19465 23063 19499
rect 4353 19397 4387 19431
rect 5273 19397 5307 19431
rect 10701 19397 10735 19431
rect 13216 19397 13250 19431
rect 15301 19397 15335 19431
rect 16129 19397 16163 19431
rect 1409 19329 1443 19363
rect 1685 19329 1719 19363
rect 1952 19329 1986 19363
rect 3341 19329 3375 19363
rect 3985 19329 4019 19363
rect 4445 19329 4479 19363
rect 6009 19329 6043 19363
rect 6745 19329 6779 19363
rect 7297 19329 7331 19363
rect 7620 19329 7654 19363
rect 9229 19329 9263 19363
rect 9689 19329 9723 19363
rect 9965 19329 9999 19363
rect 10241 19329 10275 19363
rect 11161 19329 11195 19363
rect 11529 19329 11563 19363
rect 11805 19329 11839 19363
rect 13461 19329 13495 19363
rect 14013 19329 14047 19363
rect 14841 19329 14875 19363
rect 14933 19329 14967 19363
rect 15945 19329 15979 19363
rect 16773 19329 16807 19363
rect 19073 19329 19107 19363
rect 19993 19329 20027 19363
rect 20913 19329 20947 19363
rect 21005 19329 21039 19363
rect 21649 19329 21683 19363
rect 22201 19329 22235 19363
rect 22845 19329 22879 19363
rect 4169 19261 4203 19295
rect 5365 19261 5399 19295
rect 5457 19261 5491 19295
rect 7205 19261 7239 19295
rect 7760 19261 7794 19295
rect 7987 19261 8021 19295
rect 10793 19261 10827 19295
rect 10885 19261 10919 19295
rect 13737 19261 13771 19295
rect 13921 19261 13955 19295
rect 15025 19261 15059 19295
rect 16405 19261 16439 19295
rect 17141 19261 17175 19295
rect 17464 19261 17498 19295
rect 17604 19261 17638 19295
rect 17877 19261 17911 19295
rect 22385 19261 22419 19295
rect 22661 19261 22695 19295
rect 3249 19193 3283 19227
rect 9505 19193 9539 19227
rect 19809 19193 19843 19227
rect 5825 19125 5859 19159
rect 6193 19125 6227 19159
rect 9413 19125 9447 19159
rect 9781 19125 9815 19159
rect 11713 19125 11747 19159
rect 12081 19125 12115 19159
rect 14473 19125 14507 19159
rect 16221 19125 16255 19159
rect 19717 19125 19751 19159
rect 20269 19125 20303 19159
rect 4813 18921 4847 18955
rect 12817 18921 12851 18955
rect 13921 18921 13955 18955
rect 14105 18921 14139 18955
rect 15577 18921 15611 18955
rect 17325 18921 17359 18955
rect 20545 18921 20579 18955
rect 23029 18921 23063 18955
rect 7205 18853 7239 18887
rect 17233 18853 17267 18887
rect 18889 18853 18923 18887
rect 4445 18785 4479 18819
rect 5457 18785 5491 18819
rect 10241 18785 10275 18819
rect 11023 18785 11057 18819
rect 17877 18785 17911 18819
rect 1501 18717 1535 18751
rect 2145 18717 2179 18751
rect 2881 18717 2915 18751
rect 3617 18717 3651 18751
rect 5181 18717 5215 18751
rect 6285 18717 6319 18751
rect 7021 18717 7055 18751
rect 7941 18717 7975 18751
rect 8677 18717 8711 18751
rect 9597 18717 9631 18751
rect 10517 18717 10551 18751
rect 11253 18717 11287 18751
rect 12633 18717 12667 18751
rect 12909 18717 12943 18751
rect 13737 18717 13771 18751
rect 15485 18717 15519 18751
rect 16957 18717 16991 18751
rect 17049 18717 17083 18751
rect 17785 18717 17819 18751
rect 18797 18717 18831 18751
rect 19073 18717 19107 18751
rect 19349 18717 19383 18751
rect 19441 18717 19475 18751
rect 21925 18717 21959 18751
rect 22661 18717 22695 18751
rect 22845 18717 22879 18751
rect 4721 18649 4755 18683
rect 8953 18649 8987 18683
rect 15240 18649 15274 18683
rect 16712 18649 16746 18683
rect 20177 18649 20211 18683
rect 21680 18649 21714 18683
rect 2237 18581 2271 18615
rect 2973 18581 3007 18615
rect 3801 18581 3835 18615
rect 4169 18581 4203 18615
rect 4261 18581 4295 18615
rect 5273 18581 5307 18615
rect 5641 18581 5675 18615
rect 6377 18581 6411 18615
rect 7297 18581 7331 18615
rect 8033 18581 8067 18615
rect 9689 18581 9723 18615
rect 10057 18581 10091 18615
rect 10149 18581 10183 18615
rect 10983 18581 11017 18615
rect 12357 18581 12391 18615
rect 12541 18581 12575 18615
rect 13553 18581 13587 18615
rect 17693 18581 17727 18615
rect 18153 18581 18187 18615
rect 22017 18581 22051 18615
rect 1685 18377 1719 18411
rect 4905 18377 4939 18411
rect 5733 18377 5767 18411
rect 9419 18377 9453 18411
rect 10885 18377 10919 18411
rect 11529 18377 11563 18411
rect 12817 18377 12851 18411
rect 14565 18377 14599 18411
rect 16681 18377 16715 18411
rect 17049 18377 17083 18411
rect 18245 18377 18279 18411
rect 18613 18377 18647 18411
rect 19165 18377 19199 18411
rect 21557 18377 21591 18411
rect 22293 18377 22327 18411
rect 22753 18377 22787 18411
rect 3770 18309 3804 18343
rect 5365 18309 5399 18343
rect 6193 18309 6227 18343
rect 7542 18309 7576 18343
rect 8769 18309 8803 18343
rect 18153 18309 18187 18343
rect 19892 18309 19926 18343
rect 22201 18309 22235 18343
rect 1501 18241 1535 18275
rect 1777 18241 1811 18275
rect 2053 18241 2087 18275
rect 2320 18241 2354 18275
rect 3525 18241 3559 18275
rect 6009 18241 6043 18275
rect 7021 18241 7055 18275
rect 7297 18241 7331 18275
rect 11161 18241 11195 18275
rect 11897 18241 11931 18275
rect 11989 18241 12023 18275
rect 12909 18241 12943 18275
rect 14013 18241 14047 18275
rect 14473 18241 14507 18275
rect 15117 18241 15151 18275
rect 15384 18241 15418 18275
rect 17509 18241 17543 18275
rect 18429 18241 18463 18275
rect 21281 18241 21315 18275
rect 21373 18241 21407 18275
rect 22845 18241 22879 18275
rect 5089 18173 5123 18207
rect 5273 18173 5307 18207
rect 8953 18173 8987 18207
rect 9416 18173 9450 18207
rect 9689 18173 9723 18207
rect 12081 18173 12115 18207
rect 12725 18173 12759 18207
rect 14289 18173 14323 18207
rect 17141 18173 17175 18207
rect 17233 18173 17267 18207
rect 18889 18173 18923 18207
rect 19073 18173 19107 18207
rect 19625 18173 19659 18207
rect 22477 18173 22511 18207
rect 1961 18105 1995 18139
rect 10793 18105 10827 18139
rect 12449 18105 12483 18139
rect 16497 18105 16531 18139
rect 21005 18105 21039 18139
rect 3433 18037 3467 18071
rect 6377 18037 6411 18071
rect 8677 18037 8711 18071
rect 11345 18037 11379 18071
rect 13277 18037 13311 18071
rect 13369 18037 13403 18071
rect 14933 18037 14967 18071
rect 19533 18037 19567 18071
rect 21097 18037 21131 18071
rect 21833 18037 21867 18071
rect 23029 18037 23063 18071
rect 1685 17833 1719 17867
rect 3157 17833 3191 17867
rect 3985 17833 4019 17867
rect 6469 17833 6503 17867
rect 6745 17833 6779 17867
rect 11437 17833 11471 17867
rect 12909 17833 12943 17867
rect 14105 17833 14139 17867
rect 17325 17833 17359 17867
rect 19257 17833 19291 17867
rect 22845 17833 22879 17867
rect 3341 17765 3375 17799
rect 8677 17765 8711 17799
rect 13001 17765 13035 17799
rect 16313 17765 16347 17799
rect 17601 17765 17635 17799
rect 21373 17765 21407 17799
rect 1777 17697 1811 17731
rect 8122 17697 8156 17731
rect 9689 17697 9723 17731
rect 10057 17697 10091 17731
rect 13461 17697 13495 17731
rect 13553 17697 13587 17731
rect 14657 17697 14691 17731
rect 16037 17697 16071 17731
rect 16865 17697 16899 17731
rect 21465 17697 21499 17731
rect 1501 17629 1535 17663
rect 2044 17629 2078 17663
rect 3433 17629 3467 17663
rect 3801 17629 3835 17663
rect 4077 17629 4111 17663
rect 5089 17629 5123 17663
rect 6561 17629 6595 17663
rect 7849 17629 7883 17663
rect 8585 17629 8619 17663
rect 11529 17629 11563 17663
rect 11796 17629 11830 17663
rect 14473 17629 14507 17663
rect 15117 17629 15151 17663
rect 17141 17629 17175 17663
rect 17417 17629 17451 17663
rect 17693 17629 17727 17663
rect 20637 17629 20671 17663
rect 20729 17629 20763 17663
rect 21721 17629 21755 17663
rect 23121 17629 23155 17663
rect 4813 17561 4847 17595
rect 5356 17561 5390 17595
rect 8953 17561 8987 17595
rect 10324 17561 10358 17595
rect 13921 17561 13955 17595
rect 15301 17561 15335 17595
rect 16773 17561 16807 17595
rect 17960 17561 17994 17595
rect 20392 17561 20426 17595
rect 3617 17493 3651 17527
rect 8118 17493 8152 17527
rect 13369 17493 13403 17527
rect 14565 17493 14599 17527
rect 14933 17493 14967 17527
rect 16681 17493 16715 17527
rect 19073 17493 19107 17527
rect 22937 17493 22971 17527
rect 1501 17289 1535 17323
rect 3249 17289 3283 17323
rect 3341 17289 3375 17323
rect 4537 17289 4571 17323
rect 4721 17289 4755 17323
rect 6377 17289 6411 17323
rect 8861 17289 8895 17323
rect 9689 17289 9723 17323
rect 13461 17289 13495 17323
rect 13921 17289 13955 17323
rect 14289 17289 14323 17323
rect 16497 17289 16531 17323
rect 17417 17289 17451 17323
rect 19257 17289 19291 17323
rect 20085 17289 20119 17323
rect 20821 17289 20855 17323
rect 21189 17289 21223 17323
rect 21833 17289 21867 17323
rect 22201 17289 22235 17323
rect 22293 17289 22327 17323
rect 9229 17221 9263 17255
rect 10824 17221 10858 17255
rect 11345 17221 11379 17255
rect 12256 17221 12290 17255
rect 21281 17221 21315 17255
rect 22845 17221 22879 17255
rect 2614 17153 2648 17187
rect 2881 17153 2915 17187
rect 4169 17153 4203 17187
rect 5080 17153 5114 17187
rect 6745 17153 6779 17187
rect 8318 17153 8352 17187
rect 8585 17153 8619 17187
rect 11069 17153 11103 17187
rect 11713 17153 11747 17187
rect 13829 17153 13863 17187
rect 14657 17153 14691 17187
rect 15117 17153 15151 17187
rect 15384 17153 15418 17187
rect 16681 17153 16715 17187
rect 18541 17153 18575 17187
rect 18797 17153 18831 17187
rect 20729 17153 20763 17187
rect 3157 17085 3191 17119
rect 3893 17085 3927 17119
rect 4077 17085 4111 17119
rect 4813 17085 4847 17119
rect 6837 17085 6871 17119
rect 6929 17085 6963 17119
rect 9321 17085 9355 17119
rect 9413 17085 9447 17119
rect 11989 17085 12023 17119
rect 14105 17085 14139 17119
rect 14749 17085 14783 17119
rect 14841 17085 14875 17119
rect 19073 17085 19107 17119
rect 19165 17085 19199 17119
rect 20177 17085 20211 17119
rect 20361 17085 20395 17119
rect 21465 17085 21499 17119
rect 22477 17085 22511 17119
rect 3709 17017 3743 17051
rect 6193 17017 6227 17051
rect 19625 17017 19659 17051
rect 22661 17017 22695 17051
rect 7205 16949 7239 16983
rect 8769 16949 8803 16983
rect 11621 16949 11655 16983
rect 11897 16949 11931 16983
rect 13369 16949 13403 16983
rect 17325 16949 17359 16983
rect 19717 16949 19751 16983
rect 20545 16949 20579 16983
rect 23121 16949 23155 16983
rect 3801 16745 3835 16779
rect 6009 16745 6043 16779
rect 6929 16745 6963 16779
rect 8125 16745 8159 16779
rect 16313 16745 16347 16779
rect 18797 16745 18831 16779
rect 18613 16677 18647 16711
rect 19901 16677 19935 16711
rect 2697 16609 2731 16643
rect 4445 16609 4479 16643
rect 4629 16609 4663 16643
rect 6561 16609 6595 16643
rect 6653 16609 6687 16643
rect 7573 16609 7607 16643
rect 7665 16609 7699 16643
rect 9045 16609 9079 16643
rect 9229 16609 9263 16643
rect 13829 16609 13863 16643
rect 14841 16609 14875 16643
rect 17233 16609 17267 16643
rect 20453 16609 20487 16643
rect 21465 16609 21499 16643
rect 1501 16541 1535 16575
rect 2421 16541 2455 16575
rect 2881 16541 2915 16575
rect 3617 16541 3651 16575
rect 4896 16541 4930 16575
rect 6469 16541 6503 16575
rect 7757 16541 7791 16575
rect 8401 16541 8435 16575
rect 8493 16541 8527 16575
rect 11161 16541 11195 16575
rect 12357 16541 12391 16575
rect 13562 16541 13596 16575
rect 14749 16541 14783 16575
rect 16957 16541 16991 16575
rect 17489 16541 17523 16575
rect 18889 16541 18923 16575
rect 19257 16541 19291 16575
rect 19993 16541 20027 16575
rect 20729 16541 20763 16575
rect 23121 16541 23155 16575
rect 4261 16473 4295 16507
rect 10916 16473 10950 16507
rect 15108 16473 15142 16507
rect 17141 16473 17175 16507
rect 20637 16473 20671 16507
rect 21189 16473 21223 16507
rect 21732 16473 21766 16507
rect 1685 16405 1719 16439
rect 1777 16405 1811 16439
rect 2789 16405 2823 16439
rect 3249 16405 3283 16439
rect 3433 16405 3467 16439
rect 4169 16405 4203 16439
rect 6101 16405 6135 16439
rect 7113 16405 7147 16439
rect 8217 16405 8251 16439
rect 9321 16405 9355 16439
rect 9689 16405 9723 16439
rect 9781 16405 9815 16439
rect 11437 16405 11471 16439
rect 11713 16405 11747 16439
rect 12449 16405 12483 16439
rect 14105 16405 14139 16439
rect 16221 16405 16255 16439
rect 19073 16405 19107 16439
rect 20177 16405 20211 16439
rect 21097 16405 21131 16439
rect 22845 16405 22879 16439
rect 22937 16405 22971 16439
rect 2881 16201 2915 16235
rect 3709 16201 3743 16235
rect 5181 16201 5215 16235
rect 5457 16201 5491 16235
rect 8033 16201 8067 16235
rect 9505 16201 9539 16235
rect 9965 16201 9999 16235
rect 12173 16201 12207 16235
rect 13645 16201 13679 16235
rect 15117 16201 15151 16235
rect 16221 16201 16255 16235
rect 3341 16133 3375 16167
rect 14004 16133 14038 16167
rect 18092 16133 18126 16167
rect 19901 16133 19935 16167
rect 22753 16133 22787 16167
rect 1768 16065 1802 16099
rect 4068 16065 4102 16099
rect 5273 16065 5307 16099
rect 5549 16065 5583 16099
rect 6193 16065 6227 16099
rect 7205 16065 7239 16099
rect 7297 16065 7331 16099
rect 9146 16065 9180 16099
rect 9413 16065 9447 16099
rect 11078 16065 11112 16099
rect 11345 16065 11379 16099
rect 11529 16065 11563 16099
rect 12265 16065 12299 16099
rect 12521 16065 12555 16099
rect 13737 16065 13771 16099
rect 15209 16065 15243 16099
rect 16037 16065 16071 16099
rect 16313 16065 16347 16099
rect 16681 16065 16715 16099
rect 18337 16065 18371 16099
rect 18797 16065 18831 16099
rect 19257 16065 19291 16099
rect 19993 16065 20027 16099
rect 21373 16065 21407 16099
rect 21649 16065 21683 16099
rect 22477 16065 22511 16099
rect 22569 16065 22603 16099
rect 1501 15997 1535 16031
rect 3065 15997 3099 16031
rect 3249 15997 3283 16031
rect 3801 15997 3835 16031
rect 6377 15997 6411 16031
rect 18521 15997 18555 16031
rect 18705 15997 18739 16031
rect 22937 15997 22971 16031
rect 6561 15929 6595 15963
rect 16497 15929 16531 15963
rect 16865 15929 16899 15963
rect 20729 15929 20763 15963
rect 7941 15861 7975 15895
rect 15853 15861 15887 15895
rect 16957 15861 16991 15895
rect 19165 15861 19199 15895
rect 20637 15861 20671 15895
rect 21465 15861 21499 15895
rect 21833 15861 21867 15895
rect 23121 15861 23155 15895
rect 2053 15657 2087 15691
rect 3525 15657 3559 15691
rect 4169 15657 4203 15691
rect 5641 15657 5675 15691
rect 8953 15657 8987 15691
rect 10517 15657 10551 15691
rect 12357 15657 12391 15691
rect 13461 15657 13495 15691
rect 13645 15657 13679 15691
rect 13921 15657 13955 15691
rect 15761 15657 15795 15691
rect 18705 15657 18739 15691
rect 19993 15657 20027 15691
rect 21097 15657 21131 15691
rect 22845 15657 22879 15691
rect 3801 15589 3835 15623
rect 10425 15589 10459 15623
rect 11529 15589 11563 15623
rect 17877 15589 17911 15623
rect 2145 15521 2179 15555
rect 6469 15521 6503 15555
rect 6653 15521 6687 15555
rect 9873 15521 9907 15555
rect 9965 15521 9999 15555
rect 11161 15521 11195 15555
rect 14289 15521 14323 15555
rect 18061 15521 18095 15555
rect 18245 15521 18279 15555
rect 19441 15521 19475 15555
rect 20177 15521 20211 15555
rect 20361 15521 20395 15555
rect 21465 15521 21499 15555
rect 1409 15453 1443 15487
rect 3985 15453 4019 15487
rect 4261 15453 4295 15487
rect 4997 15453 5031 15487
rect 5917 15453 5951 15487
rect 7205 15453 7239 15487
rect 9597 15453 9631 15487
rect 10057 15453 10091 15487
rect 10977 15453 11011 15487
rect 11345 15453 11379 15487
rect 11713 15453 11747 15487
rect 13737 15453 13771 15487
rect 14556 15453 14590 15487
rect 16405 15453 16439 15487
rect 16497 15453 16531 15487
rect 18889 15453 18923 15487
rect 20913 15453 20947 15487
rect 21181 15453 21215 15487
rect 23121 15453 23155 15487
rect 2390 15385 2424 15419
rect 7472 15385 7506 15419
rect 14197 15385 14231 15419
rect 16764 15385 16798 15419
rect 18337 15385 18371 15419
rect 20453 15385 20487 15419
rect 21732 15385 21766 15419
rect 4905 15317 4939 15351
rect 5733 15317 5767 15351
rect 6009 15317 6043 15351
rect 6561 15317 6595 15351
rect 7039 15317 7073 15351
rect 8585 15317 8619 15351
rect 10885 15317 10919 15351
rect 15669 15317 15703 15351
rect 19073 15317 19107 15351
rect 19533 15317 19567 15351
rect 19625 15317 19659 15351
rect 20821 15317 20855 15351
rect 21373 15317 21407 15351
rect 22937 15317 22971 15351
rect 1409 15113 1443 15147
rect 4261 15113 4295 15147
rect 5825 15113 5859 15147
rect 8033 15113 8067 15147
rect 9406 15113 9440 15147
rect 11621 15113 11655 15147
rect 16681 15113 16715 15147
rect 18429 15113 18463 15147
rect 18889 15113 18923 15147
rect 19349 15113 19383 15147
rect 19809 15113 19843 15147
rect 20913 15113 20947 15147
rect 21373 15113 21407 15147
rect 22201 15113 22235 15147
rect 22661 15113 22695 15147
rect 2544 15045 2578 15079
rect 4353 15045 4387 15079
rect 5089 15045 5123 15079
rect 10793 15045 10827 15079
rect 14105 15045 14139 15079
rect 14565 15045 14599 15079
rect 22109 15045 22143 15079
rect 2789 14977 2823 15011
rect 2881 14977 2915 15011
rect 3137 14977 3171 15011
rect 5733 14977 5767 15011
rect 7490 14977 7524 15011
rect 9965 14977 9999 15011
rect 11345 14977 11379 15011
rect 12745 14977 12779 15011
rect 13001 14977 13035 15011
rect 14381 14977 14415 15011
rect 15761 14977 15795 15011
rect 16497 14977 16531 15011
rect 17805 14977 17839 15011
rect 18061 14977 18095 15011
rect 18521 14977 18555 15011
rect 19441 14977 19475 15011
rect 19901 14977 19935 15011
rect 21281 14977 21315 15011
rect 22845 14977 22879 15011
rect 23121 14977 23155 15011
rect 6009 14909 6043 14943
rect 7757 14909 7791 14943
rect 9137 14909 9171 14943
rect 9410 14909 9444 14943
rect 9873 14909 9907 14943
rect 15301 14909 15335 14943
rect 18337 14909 18371 14943
rect 19165 14909 19199 14943
rect 20729 14909 20763 14943
rect 21465 14909 21499 14943
rect 22017 14909 22051 14943
rect 6377 14841 6411 14875
rect 14197 14841 14231 14875
rect 22937 14841 22971 14875
rect 5365 14773 5399 14807
rect 11069 14773 11103 14807
rect 11161 14773 11195 14807
rect 13921 14773 13955 14807
rect 15577 14773 15611 14807
rect 15853 14773 15887 14807
rect 22569 14773 22603 14807
rect 1593 14569 1627 14603
rect 2053 14569 2087 14603
rect 2421 14569 2455 14603
rect 2697 14569 2731 14603
rect 2973 14569 3007 14603
rect 4169 14569 4203 14603
rect 8953 14569 8987 14603
rect 10149 14569 10183 14603
rect 10425 14569 10459 14603
rect 13553 14569 13587 14603
rect 15945 14569 15979 14603
rect 17601 14569 17635 14603
rect 19073 14569 19107 14603
rect 21005 14569 21039 14603
rect 22569 14569 22603 14603
rect 1777 14501 1811 14535
rect 10517 14501 10551 14535
rect 17509 14501 17543 14535
rect 4629 14433 4663 14467
rect 4813 14433 4847 14467
rect 4997 14433 5031 14467
rect 7573 14433 7607 14467
rect 7803 14433 7837 14467
rect 9505 14433 9539 14467
rect 11161 14433 11195 14467
rect 16129 14433 16163 14467
rect 18429 14433 18463 14467
rect 21189 14433 21223 14467
rect 1409 14365 1443 14399
rect 1961 14365 1995 14399
rect 2237 14365 2271 14399
rect 2605 14365 2639 14399
rect 2881 14365 2915 14399
rect 3617 14365 3651 14399
rect 3985 14365 4019 14399
rect 8309 14365 8343 14399
rect 9965 14365 9999 14399
rect 10241 14365 10275 14399
rect 10885 14365 10919 14399
rect 12081 14365 12115 14399
rect 12173 14365 12207 14399
rect 12909 14365 12943 14399
rect 14749 14365 14783 14399
rect 15485 14365 15519 14399
rect 16385 14365 16419 14399
rect 18245 14365 18279 14399
rect 18705 14365 18739 14399
rect 20370 14365 20404 14399
rect 20637 14365 20671 14399
rect 20913 14365 20947 14399
rect 21456 14365 21490 14399
rect 23121 14365 23155 14399
rect 5264 14297 5298 14331
rect 9321 14297 9355 14331
rect 9873 14297 9907 14331
rect 10977 14297 11011 14331
rect 15577 14297 15611 14331
rect 15761 14297 15795 14331
rect 4537 14229 4571 14263
rect 6377 14229 6411 14263
rect 6469 14229 6503 14263
rect 7842 14229 7876 14263
rect 9413 14229 9447 14263
rect 11437 14229 11471 14263
rect 12817 14229 12851 14263
rect 14105 14229 14139 14263
rect 14841 14229 14875 14263
rect 18613 14229 18647 14263
rect 19257 14229 19291 14263
rect 20729 14229 20763 14263
rect 22661 14229 22695 14263
rect 22937 14229 22971 14263
rect 2789 14025 2823 14059
rect 5733 14025 5767 14059
rect 6653 14025 6687 14059
rect 7113 14025 7147 14059
rect 8309 14025 8343 14059
rect 9229 14025 9263 14059
rect 10885 14025 10919 14059
rect 14565 14025 14599 14059
rect 16129 14025 16163 14059
rect 19901 14025 19935 14059
rect 21373 14025 21407 14059
rect 21649 14025 21683 14059
rect 22109 14025 22143 14059
rect 22201 14025 22235 14059
rect 9321 13957 9355 13991
rect 10425 13957 10459 13991
rect 11774 13957 11808 13991
rect 16497 13957 16531 13991
rect 2605 13889 2639 13923
rect 3148 13889 3182 13923
rect 4353 13889 4387 13923
rect 4620 13889 4654 13923
rect 6009 13889 6043 13923
rect 7021 13889 7055 13923
rect 7481 13889 7515 13923
rect 8401 13889 8435 13923
rect 8585 13889 8619 13923
rect 9965 13889 9999 13923
rect 10517 13889 10551 13923
rect 11161 13889 11195 13923
rect 11529 13889 11563 13923
rect 13185 13889 13219 13923
rect 13452 13889 13486 13923
rect 14657 13889 14691 13923
rect 14924 13889 14958 13923
rect 16313 13889 16347 13923
rect 16681 13889 16715 13923
rect 17601 13889 17635 13923
rect 17785 13889 17819 13923
rect 18521 13889 18555 13923
rect 18788 13889 18822 13923
rect 19993 13889 20027 13923
rect 20249 13889 20283 13923
rect 21465 13889 21499 13923
rect 22845 13889 22879 13923
rect 23121 13889 23155 13923
rect 2881 13821 2915 13855
rect 6101 13821 6135 13855
rect 7205 13821 7239 13855
rect 8125 13821 8159 13855
rect 10333 13821 10367 13855
rect 10977 13821 11011 13855
rect 17325 13821 17359 13855
rect 18429 13821 18463 13855
rect 21925 13821 21959 13855
rect 4261 13753 4295 13787
rect 17417 13753 17451 13787
rect 1961 13685 1995 13719
rect 5825 13685 5859 13719
rect 12909 13685 12943 13719
rect 16037 13685 16071 13719
rect 22569 13685 22603 13719
rect 22661 13685 22695 13719
rect 22937 13685 22971 13719
rect 5641 13481 5675 13515
rect 7021 13481 7055 13515
rect 9321 13481 9355 13515
rect 11897 13481 11931 13515
rect 13921 13481 13955 13515
rect 16129 13481 16163 13515
rect 19349 13481 19383 13515
rect 22661 13481 22695 13515
rect 22845 13481 22879 13515
rect 3525 13413 3559 13447
rect 4537 13413 4571 13447
rect 8493 13413 8527 13447
rect 10149 13413 10183 13447
rect 12357 13413 12391 13447
rect 22937 13413 22971 13447
rect 3893 13345 3927 13379
rect 5181 13345 5215 13379
rect 9505 13345 9539 13379
rect 18797 13345 18831 13379
rect 19073 13345 19107 13379
rect 21097 13345 21131 13379
rect 21281 13345 21315 13379
rect 1409 13277 1443 13311
rect 2145 13277 2179 13311
rect 4169 13277 4203 13311
rect 5089 13277 5123 13311
rect 6285 13277 6319 13311
rect 6377 13277 6411 13311
rect 7113 13277 7147 13311
rect 7369 13277 7403 13311
rect 8769 13277 8803 13311
rect 9137 13277 9171 13311
rect 10241 13277 10275 13311
rect 10517 13277 10551 13311
rect 11989 13277 12023 13311
rect 12173 13277 12207 13311
rect 12541 13277 12575 13311
rect 14749 13277 14783 13311
rect 15016 13277 15050 13311
rect 16865 13277 16899 13311
rect 17049 13277 17083 13311
rect 17785 13277 17819 13311
rect 19993 13277 20027 13311
rect 20361 13277 20395 13311
rect 20821 13277 20855 13311
rect 23121 13277 23155 13311
rect 2390 13209 2424 13243
rect 4077 13209 4111 13243
rect 10762 13209 10796 13243
rect 12808 13209 12842 13243
rect 21526 13209 21560 13243
rect 2053 13141 2087 13175
rect 4629 13141 4663 13175
rect 4997 13141 5031 13175
rect 8585 13141 8619 13175
rect 9689 13141 9723 13175
rect 9781 13141 9815 13175
rect 10425 13141 10459 13175
rect 16221 13141 16255 13175
rect 17693 13141 17727 13175
rect 18429 13141 18463 13175
rect 20177 13141 20211 13175
rect 20453 13141 20487 13175
rect 20913 13141 20947 13175
rect 1869 12937 1903 12971
rect 3525 12937 3559 12971
rect 5457 12937 5491 12971
rect 6101 12937 6135 12971
rect 8769 12937 8803 12971
rect 9321 12937 9355 12971
rect 9781 12937 9815 12971
rect 10149 12937 10183 12971
rect 10517 12937 10551 12971
rect 11529 12937 11563 12971
rect 11897 12937 11931 12971
rect 18889 12937 18923 12971
rect 19625 12937 19659 12971
rect 20269 12937 20303 12971
rect 21833 12937 21867 12971
rect 22661 12937 22695 12971
rect 5641 12869 5675 12903
rect 5806 12869 5840 12903
rect 10609 12869 10643 12903
rect 13676 12869 13710 12903
rect 14381 12869 14415 12903
rect 15209 12869 15243 12903
rect 2993 12801 3027 12835
rect 3249 12801 3283 12835
rect 4169 12801 4203 12835
rect 4813 12801 4847 12835
rect 5917 12801 5951 12835
rect 6377 12801 6411 12835
rect 6837 12801 6871 12835
rect 8134 12801 8168 12835
rect 8401 12801 8435 12835
rect 8861 12801 8895 12835
rect 9689 12801 9723 12835
rect 11161 12801 11195 12835
rect 13921 12801 13955 12835
rect 15301 12801 15335 12835
rect 16497 12801 16531 12835
rect 17049 12801 17083 12835
rect 17509 12801 17543 12835
rect 17776 12801 17810 12835
rect 18981 12801 19015 12835
rect 19809 12801 19843 12835
rect 21393 12801 21427 12835
rect 21649 12801 21683 12835
rect 22201 12801 22235 12835
rect 23121 12801 23155 12835
rect 4905 12733 4939 12767
rect 5089 12733 5123 12767
rect 8677 12733 8711 12767
rect 9873 12733 9907 12767
rect 10793 12733 10827 12767
rect 10977 12733 11011 12767
rect 11989 12733 12023 12767
rect 12081 12733 12115 12767
rect 14197 12733 14231 12767
rect 14289 12733 14323 12767
rect 15393 12733 15427 12767
rect 16865 12733 16899 12767
rect 16957 12733 16991 12767
rect 22293 12733 22327 12767
rect 22477 12733 22511 12767
rect 6653 12665 6687 12699
rect 12541 12665 12575 12699
rect 4445 12597 4479 12631
rect 6561 12597 6595 12631
rect 7021 12597 7055 12631
rect 9229 12597 9263 12631
rect 14749 12597 14783 12631
rect 14841 12597 14875 12631
rect 15853 12597 15887 12631
rect 17417 12597 17451 12631
rect 19993 12597 20027 12631
rect 20177 12597 20211 12631
rect 22937 12597 22971 12631
rect 3801 12393 3835 12427
rect 9137 12393 9171 12427
rect 10149 12393 10183 12427
rect 14933 12393 14967 12427
rect 17049 12393 17083 12427
rect 19625 12393 19659 12427
rect 21557 12393 21591 12427
rect 3433 12325 3467 12359
rect 8769 12325 8803 12359
rect 2053 12257 2087 12291
rect 13921 12257 13955 12291
rect 14197 12257 14231 12291
rect 14381 12257 14415 12291
rect 15669 12257 15703 12291
rect 18521 12257 18555 12291
rect 20223 12257 20257 12291
rect 21741 12257 21775 12291
rect 2309 12189 2343 12223
rect 4445 12189 4479 12223
rect 4537 12189 4571 12223
rect 5457 12189 5491 12223
rect 5641 12189 5675 12223
rect 6653 12189 6687 12223
rect 7869 12189 7903 12223
rect 8125 12189 8159 12223
rect 8585 12189 8619 12223
rect 8953 12189 8987 12223
rect 10057 12189 10091 12223
rect 11529 12189 11563 12223
rect 14473 12189 14507 12223
rect 15577 12189 15611 12223
rect 15936 12189 15970 12223
rect 18254 12189 18288 12223
rect 19073 12189 19107 12223
rect 19717 12189 19751 12223
rect 20453 12189 20487 12223
rect 9413 12121 9447 12155
rect 11262 12121 11296 12155
rect 12173 12121 12207 12155
rect 22008 12121 22042 12155
rect 5181 12053 5215 12087
rect 6009 12053 6043 12087
rect 6745 12053 6779 12087
rect 14841 12053 14875 12087
rect 17141 12053 17175 12087
rect 18613 12053 18647 12087
rect 19441 12053 19475 12087
rect 20183 12053 20217 12087
rect 23121 12053 23155 12087
rect 1777 11849 1811 11883
rect 3617 11849 3651 11883
rect 3709 11849 3743 11883
rect 4261 11849 4295 11883
rect 5365 11849 5399 11883
rect 8125 11849 8159 11883
rect 8493 11849 8527 11883
rect 8953 11849 8987 11883
rect 11345 11849 11379 11883
rect 11989 11849 12023 11883
rect 14749 11849 14783 11883
rect 15209 11849 15243 11883
rect 18521 11849 18555 11883
rect 20453 11849 20487 11883
rect 20821 11849 20855 11883
rect 21373 11849 21407 11883
rect 21833 11849 21867 11883
rect 22293 11849 22327 11883
rect 2912 11781 2946 11815
rect 6990 11781 7024 11815
rect 8585 11781 8619 11815
rect 14013 11781 14047 11815
rect 17408 11781 17442 11815
rect 18858 11781 18892 11815
rect 21281 11781 21315 11815
rect 22661 11781 22695 11815
rect 4077 11713 4111 11747
rect 4537 11713 4571 11747
rect 4997 11713 5031 11747
rect 6101 11713 6135 11747
rect 6561 11713 6595 11747
rect 9045 11713 9079 11747
rect 9965 11713 9999 11747
rect 10221 11713 10255 11747
rect 13369 11713 13403 11747
rect 15393 11713 15427 11747
rect 15669 11713 15703 11747
rect 16129 11713 16163 11747
rect 16865 11713 16899 11747
rect 22201 11713 22235 11747
rect 23121 11713 23155 11747
rect 3157 11645 3191 11679
rect 3893 11645 3927 11679
rect 4721 11645 4755 11679
rect 4905 11645 4939 11679
rect 6745 11645 6779 11679
rect 8401 11645 8435 11679
rect 12081 11645 12115 11679
rect 12173 11645 12207 11679
rect 13185 11645 13219 11679
rect 13277 11645 13311 11679
rect 14565 11645 14599 11679
rect 14657 11645 14691 11679
rect 15945 11645 15979 11679
rect 16037 11645 16071 11679
rect 17141 11645 17175 11679
rect 18613 11645 18647 11679
rect 20177 11645 20211 11679
rect 20361 11645 20395 11679
rect 21465 11645 21499 11679
rect 22385 11645 22419 11679
rect 6377 11577 6411 11611
rect 11621 11577 11655 11611
rect 15485 11577 15519 11611
rect 16681 11577 16715 11611
rect 3249 11509 3283 11543
rect 4353 11509 4387 11543
rect 5457 11509 5491 11543
rect 9689 11509 9723 11543
rect 13737 11509 13771 11543
rect 13921 11509 13955 11543
rect 15117 11509 15151 11543
rect 16497 11509 16531 11543
rect 19993 11509 20027 11543
rect 20913 11509 20947 11543
rect 22937 11509 22971 11543
rect 3157 11305 3191 11339
rect 3985 11305 4019 11339
rect 4261 11305 4295 11339
rect 9137 11305 9171 11339
rect 9229 11305 9263 11339
rect 11437 11305 11471 11339
rect 13737 11305 13771 11339
rect 14841 11305 14875 11339
rect 15669 11305 15703 11339
rect 17601 11305 17635 11339
rect 18705 11305 18739 11339
rect 21005 11305 21039 11339
rect 3617 11237 3651 11271
rect 9965 11237 9999 11271
rect 15945 11237 15979 11271
rect 17509 11237 17543 11271
rect 18981 11237 19015 11271
rect 20637 11237 20671 11271
rect 20821 11237 20855 11271
rect 22477 11237 22511 11271
rect 22753 11237 22787 11271
rect 22937 11237 22971 11271
rect 4997 11169 5031 11203
rect 5825 11169 5859 11203
rect 6285 11169 6319 11203
rect 11345 11169 11379 11203
rect 14289 11169 14323 11203
rect 15117 11169 15151 11203
rect 16957 11169 16991 11203
rect 17049 11169 17083 11203
rect 18061 11169 18095 11203
rect 19257 11169 19291 11203
rect 1777 11101 1811 11135
rect 3433 11101 3467 11135
rect 3801 11101 3835 11135
rect 4077 11101 4111 11135
rect 5549 11101 5583 11135
rect 6929 11101 6963 11135
rect 8401 11101 8435 11135
rect 8953 11101 8987 11135
rect 9873 11101 9907 11135
rect 12081 11101 12115 11135
rect 12357 11101 12391 11135
rect 12624 11101 12658 11135
rect 14473 11101 14507 11135
rect 15761 11101 15795 11135
rect 16681 11101 16715 11135
rect 17141 11101 17175 11135
rect 17785 11101 17819 11135
rect 18337 11101 18371 11135
rect 21097 11101 21131 11135
rect 21353 11101 21387 11135
rect 22569 11101 22603 11135
rect 23121 11101 23155 11135
rect 2044 11033 2078 11067
rect 4721 11033 4755 11067
rect 8156 11033 8190 11067
rect 11078 11033 11112 11067
rect 15209 11033 15243 11067
rect 16037 11033 16071 11067
rect 18245 11033 18279 11067
rect 18889 11033 18923 11067
rect 19502 11033 19536 11067
rect 4353 10965 4387 10999
rect 4813 10965 4847 10999
rect 5181 10965 5215 10999
rect 5641 10965 5675 10999
rect 7021 10965 7055 10999
rect 14381 10965 14415 10999
rect 15301 10965 15335 10999
rect 3985 10761 4019 10795
rect 4353 10761 4387 10795
rect 7389 10761 7423 10795
rect 7849 10761 7883 10795
rect 8217 10761 8251 10795
rect 8677 10761 8711 10795
rect 8769 10761 8803 10795
rect 9137 10761 9171 10795
rect 10609 10761 10643 10795
rect 11069 10761 11103 10795
rect 14013 10761 14047 10795
rect 14381 10761 14415 10795
rect 15117 10761 15151 10795
rect 16957 10761 16991 10795
rect 22477 10761 22511 10795
rect 23121 10761 23155 10795
rect 5948 10693 5982 10727
rect 9229 10693 9263 10727
rect 10425 10693 10459 10727
rect 15853 10693 15887 10727
rect 20085 10693 20119 10727
rect 2033 10625 2067 10659
rect 3893 10625 3927 10659
rect 6193 10625 6227 10659
rect 7021 10625 7055 10659
rect 7481 10625 7515 10659
rect 8309 10625 8343 10659
rect 9597 10625 9631 10659
rect 10977 10625 11011 10659
rect 12173 10625 12207 10659
rect 12440 10625 12474 10659
rect 14473 10625 14507 10659
rect 15209 10625 15243 10659
rect 17049 10625 17083 10659
rect 17601 10625 17635 10659
rect 17969 10625 18003 10659
rect 20269 10625 20303 10659
rect 20525 10625 20559 10659
rect 21833 10625 21867 10659
rect 22937 10625 22971 10659
rect 1777 10557 1811 10591
rect 4445 10557 4479 10591
rect 4629 10557 4663 10591
rect 7205 10557 7239 10591
rect 8125 10557 8159 10591
rect 9321 10557 9355 10591
rect 11161 10557 11195 10591
rect 13737 10557 13771 10591
rect 13921 10557 13955 10591
rect 16497 10557 16531 10591
rect 16865 10557 16899 10591
rect 18292 10557 18326 10591
rect 18432 10557 18466 10591
rect 18705 10557 18739 10591
rect 22569 10557 22603 10591
rect 3157 10489 3191 10523
rect 13553 10489 13587 10523
rect 17785 10489 17819 10523
rect 3249 10421 3283 10455
rect 4813 10421 4847 10455
rect 6377 10421 6411 10455
rect 11529 10421 11563 10455
rect 17417 10421 17451 10455
rect 19809 10421 19843 10455
rect 21649 10421 21683 10455
rect 6193 10217 6227 10251
rect 7205 10217 7239 10251
rect 8953 10217 8987 10251
rect 11989 10217 12023 10251
rect 13645 10217 13679 10251
rect 14289 10217 14323 10251
rect 17325 10217 17359 10251
rect 19901 10217 19935 10251
rect 21833 10217 21867 10251
rect 22937 10217 22971 10251
rect 3617 10149 3651 10183
rect 6101 10149 6135 10183
rect 22845 10149 22879 10183
rect 3157 10081 3191 10115
rect 4261 10081 4295 10115
rect 4445 10081 4479 10115
rect 6745 10081 6779 10115
rect 9505 10081 9539 10115
rect 20499 10081 20533 10115
rect 22385 10081 22419 10115
rect 22477 10081 22511 10115
rect 3433 10013 3467 10047
rect 4721 10013 4755 10047
rect 8318 10013 8352 10047
rect 8585 10013 8619 10047
rect 9873 10013 9907 10047
rect 13369 10013 13403 10047
rect 13461 10013 13495 10047
rect 14105 10013 14139 10047
rect 15761 10013 15795 10047
rect 15853 10013 15887 10047
rect 18705 10013 18739 10047
rect 19073 10013 19107 10047
rect 19257 10013 19291 10047
rect 19993 10013 20027 10047
rect 20729 10013 20763 10047
rect 23121 10013 23155 10047
rect 2912 9945 2946 9979
rect 4169 9945 4203 9979
rect 4966 9945 5000 9979
rect 10118 9945 10152 9979
rect 13124 9945 13158 9979
rect 15516 9945 15550 9979
rect 16120 9945 16154 9979
rect 18460 9945 18494 9979
rect 18889 9945 18923 9979
rect 22293 9945 22327 9979
rect 1777 9877 1811 9911
rect 3801 9877 3835 9911
rect 6561 9877 6595 9911
rect 6653 9877 6687 9911
rect 9321 9877 9355 9911
rect 9413 9877 9447 9911
rect 11253 9877 11287 9911
rect 14381 9877 14415 9911
rect 17233 9877 17267 9911
rect 20459 9877 20493 9911
rect 21925 9877 21959 9911
rect 2973 9673 3007 9707
rect 4813 9673 4847 9707
rect 8769 9673 8803 9707
rect 10977 9673 11011 9707
rect 17147 9673 17181 9707
rect 18521 9673 18555 9707
rect 21833 9673 21867 9707
rect 22201 9673 22235 9707
rect 3065 9605 3099 9639
rect 3985 9605 4019 9639
rect 8861 9605 8895 9639
rect 12725 9605 12759 9639
rect 14841 9605 14875 9639
rect 15669 9605 15703 9639
rect 21189 9605 21223 9639
rect 22293 9605 22327 9639
rect 23121 9605 23155 9639
rect 1409 9537 1443 9571
rect 1685 9537 1719 9571
rect 2605 9537 2639 9571
rect 3525 9537 3559 9571
rect 4721 9537 4755 9571
rect 5937 9537 5971 9571
rect 6193 9537 6227 9571
rect 7297 9537 7331 9571
rect 7389 9537 7423 9571
rect 7645 9537 7679 9571
rect 9505 9537 9539 9571
rect 9597 9537 9631 9571
rect 9864 9537 9898 9571
rect 12081 9537 12115 9571
rect 13277 9537 13311 9571
rect 14381 9537 14415 9571
rect 15853 9537 15887 9571
rect 17417 9537 17451 9571
rect 18613 9537 18647 9571
rect 19349 9537 19383 9571
rect 19616 9537 19650 9571
rect 22845 9537 22879 9571
rect 2881 9469 2915 9503
rect 14473 9469 14507 9503
rect 14565 9469 14599 9503
rect 16497 9469 16531 9503
rect 16681 9469 16715 9503
rect 17187 9469 17221 9503
rect 19257 9469 19291 9503
rect 21281 9469 21315 9503
rect 21465 9469 21499 9503
rect 22477 9469 22511 9503
rect 3433 9401 3467 9435
rect 3709 9401 3743 9435
rect 14013 9401 14047 9435
rect 20729 9401 20763 9435
rect 22661 9401 22695 9435
rect 1593 9333 1627 9367
rect 1961 9333 1995 9367
rect 6653 9333 6687 9367
rect 13921 9333 13955 9367
rect 20821 9333 20855 9367
rect 3617 9129 3651 9163
rect 4537 9129 4571 9163
rect 5457 9129 5491 9163
rect 13461 9129 13495 9163
rect 14197 9129 14231 9163
rect 18981 9129 19015 9163
rect 21557 9129 21591 9163
rect 3801 9061 3835 9095
rect 8769 9061 8803 9095
rect 17417 9061 17451 9095
rect 1409 8993 1443 9027
rect 3065 8993 3099 9027
rect 5089 8993 5123 9027
rect 5549 8993 5583 9027
rect 11253 8993 11287 9027
rect 12909 8993 12943 9027
rect 16773 8993 16807 9027
rect 16957 8993 16991 9027
rect 18061 8993 18095 9027
rect 20637 8993 20671 9027
rect 21741 8993 21775 9027
rect 1665 8925 1699 8959
rect 4445 8925 4479 8959
rect 7389 8925 7423 8959
rect 9137 8925 9171 8959
rect 14381 8925 14415 8959
rect 15853 8925 15887 8959
rect 17049 8925 17083 8959
rect 18337 8925 18371 8959
rect 19717 8925 19751 8959
rect 20913 8925 20947 8959
rect 3157 8857 3191 8891
rect 5816 8857 5850 8891
rect 7634 8857 7668 8891
rect 9382 8857 9416 8891
rect 11498 8857 11532 8891
rect 14648 8857 14682 8891
rect 19441 8857 19475 8891
rect 19901 8857 19935 8891
rect 21986 8857 22020 8891
rect 2789 8789 2823 8823
rect 3249 8789 3283 8823
rect 4905 8789 4939 8823
rect 4997 8789 5031 8823
rect 6929 8789 6963 8823
rect 10517 8789 10551 8823
rect 12633 8789 12667 8823
rect 13001 8789 13035 8823
rect 13093 8789 13127 8823
rect 15761 8789 15795 8823
rect 16497 8789 16531 8823
rect 23121 8789 23155 8823
rect 3525 8585 3559 8619
rect 3893 8585 3927 8619
rect 4353 8585 4387 8619
rect 5365 8585 5399 8619
rect 7021 8585 7055 8619
rect 9781 8585 9815 8619
rect 10149 8585 10183 8619
rect 10701 8585 10735 8619
rect 13369 8585 13403 8619
rect 14933 8585 14967 8619
rect 16221 8585 16255 8619
rect 17325 8585 17359 8619
rect 18337 8585 18371 8619
rect 20177 8585 20211 8619
rect 20637 8585 20671 8619
rect 4813 8517 4847 8551
rect 7573 8517 7607 8551
rect 8554 8517 8588 8551
rect 13728 8517 13762 8551
rect 15301 8517 15335 8551
rect 18696 8517 18730 8551
rect 2053 8449 2087 8483
rect 2320 8449 2354 8483
rect 4721 8449 4755 8483
rect 5733 8449 5767 8483
rect 6377 8449 6411 8483
rect 8217 8449 8251 8483
rect 8309 8449 8343 8483
rect 11345 8449 11379 8483
rect 11989 8449 12023 8483
rect 12245 8449 12279 8483
rect 13461 8449 13495 8483
rect 16129 8449 16163 8483
rect 16681 8449 16715 8483
rect 17417 8449 17451 8483
rect 18429 8449 18463 8483
rect 20269 8449 20303 8483
rect 21373 8449 21407 8483
rect 21833 8449 21867 8483
rect 22569 8449 22603 8483
rect 3985 8381 4019 8415
rect 4169 8381 4203 8415
rect 4997 8381 5031 8415
rect 5825 8381 5859 8415
rect 6009 8381 6043 8415
rect 10241 8381 10275 8415
rect 10425 8381 10459 8415
rect 15393 8381 15427 8415
rect 15485 8381 15519 8415
rect 16313 8381 16347 8415
rect 20085 8381 20119 8415
rect 20729 8381 20763 8415
rect 21465 8381 21499 8415
rect 22477 8381 22511 8415
rect 22753 8381 22787 8415
rect 3433 8313 3467 8347
rect 9689 8313 9723 8347
rect 15761 8313 15795 8347
rect 18061 8313 18095 8347
rect 14841 8245 14875 8279
rect 19809 8245 19843 8279
rect 4629 8041 4663 8075
rect 5457 8041 5491 8075
rect 7573 8041 7607 8075
rect 8125 8041 8159 8075
rect 9505 8041 9539 8075
rect 13185 8041 13219 8075
rect 21373 8041 21407 8075
rect 22937 8041 22971 8075
rect 3893 7973 3927 8007
rect 19073 7973 19107 8007
rect 2237 7905 2271 7939
rect 5181 7905 5215 7939
rect 10241 7905 10275 7939
rect 13093 7905 13127 7939
rect 13645 7905 13679 7939
rect 13737 7905 13771 7939
rect 15485 7905 15519 7939
rect 18521 7905 18555 7939
rect 19720 7905 19754 7939
rect 19993 7905 20027 7939
rect 2145 7837 2179 7871
rect 2504 7837 2538 7871
rect 4537 7837 4571 7871
rect 6837 7837 6871 7871
rect 6929 7837 6963 7871
rect 8769 7837 8803 7871
rect 10149 7837 10183 7871
rect 12837 7837 12871 7871
rect 16037 7837 16071 7871
rect 17509 7837 17543 7871
rect 18705 7837 18739 7871
rect 19247 7837 19281 7871
rect 21189 7837 21223 7871
rect 21465 7837 21499 7871
rect 23121 7837 23155 7871
rect 1501 7769 1535 7803
rect 6592 7769 6626 7803
rect 9321 7769 9355 7803
rect 10508 7769 10542 7803
rect 15218 7769 15252 7803
rect 16304 7769 16338 7803
rect 18153 7769 18187 7803
rect 21732 7769 21766 7803
rect 3617 7701 3651 7735
rect 4997 7701 5031 7735
rect 5089 7701 5123 7735
rect 9229 7701 9263 7735
rect 11621 7701 11655 7735
rect 11713 7701 11747 7735
rect 13553 7701 13587 7735
rect 14105 7701 14139 7735
rect 17417 7701 17451 7735
rect 18613 7701 18647 7735
rect 19723 7701 19757 7735
rect 21097 7701 21131 7735
rect 22845 7701 22879 7735
rect 1409 7497 1443 7531
rect 3249 7497 3283 7531
rect 6469 7497 6503 7531
rect 11529 7497 11563 7531
rect 11805 7497 11839 7531
rect 12633 7497 12667 7531
rect 14565 7497 14599 7531
rect 15301 7497 15335 7531
rect 16129 7497 16163 7531
rect 19717 7497 19751 7531
rect 20085 7497 20119 7531
rect 20821 7497 20855 7531
rect 21925 7497 21959 7531
rect 10701 7429 10735 7463
rect 14473 7429 14507 7463
rect 17794 7429 17828 7463
rect 22293 7429 22327 7463
rect 1593 7361 1627 7395
rect 2798 7361 2832 7395
rect 4362 7361 4396 7395
rect 5069 7361 5103 7395
rect 6745 7361 6779 7395
rect 9054 7361 9088 7395
rect 9321 7361 9355 7395
rect 9413 7361 9447 7395
rect 10609 7361 10643 7395
rect 11345 7361 11379 7395
rect 12265 7361 12299 7395
rect 15209 7361 15243 7395
rect 15945 7361 15979 7395
rect 19369 7361 19403 7395
rect 19636 7361 19670 7395
rect 20913 7361 20947 7395
rect 21465 7361 21499 7395
rect 23029 7361 23063 7395
rect 3065 7293 3099 7327
rect 4629 7293 4663 7327
rect 4813 7293 4847 7327
rect 7297 7293 7331 7327
rect 10149 7293 10183 7327
rect 11989 7293 12023 7327
rect 12173 7293 12207 7327
rect 18061 7293 18095 7327
rect 20177 7293 20211 7327
rect 20361 7293 20395 7327
rect 20729 7293 20763 7327
rect 22385 7293 22419 7327
rect 22569 7293 22603 7327
rect 6193 7225 6227 7259
rect 16221 7225 16255 7259
rect 16681 7225 16715 7259
rect 21649 7225 21683 7259
rect 22845 7225 22879 7259
rect 1685 7157 1719 7191
rect 7573 7157 7607 7191
rect 7941 7157 7975 7191
rect 10425 7157 10459 7191
rect 13001 7157 13035 7191
rect 16497 7157 16531 7191
rect 18245 7157 18279 7191
rect 21281 7157 21315 7191
rect 1685 6953 1719 6987
rect 12173 6953 12207 6987
rect 17969 6953 18003 6987
rect 19073 6953 19107 6987
rect 22569 6953 22603 6987
rect 22477 6885 22511 6919
rect 1869 6817 1903 6851
rect 3985 6817 4019 6851
rect 6193 6817 6227 6851
rect 7297 6817 7331 6851
rect 8585 6817 8619 6851
rect 12265 6817 12299 6851
rect 14749 6817 14783 6851
rect 17509 6817 17543 6851
rect 17601 6817 17635 6851
rect 18429 6817 18463 6851
rect 19349 6817 19383 6851
rect 21097 6817 21131 6851
rect 2513 6749 2547 6783
rect 3617 6749 3651 6783
rect 4252 6749 4286 6783
rect 5457 6749 5491 6783
rect 7205 6749 7239 6783
rect 7941 6749 7975 6783
rect 10333 6749 10367 6783
rect 10793 6749 10827 6783
rect 12909 6749 12943 6783
rect 13012 6749 13046 6783
rect 14105 6749 14139 6783
rect 15485 6749 15519 6783
rect 16957 6749 16991 6783
rect 20453 6749 20487 6783
rect 20821 6749 20855 6783
rect 22753 6749 22787 6783
rect 22845 6749 22879 6783
rect 2973 6681 3007 6715
rect 8493 6681 8527 6715
rect 10088 6681 10122 6715
rect 10609 6681 10643 6715
rect 11060 6681 11094 6715
rect 13737 6681 13771 6715
rect 16690 6681 16724 6715
rect 17417 6681 17451 6715
rect 18153 6681 18187 6715
rect 19717 6681 19751 6715
rect 21364 6681 21398 6715
rect 5365 6613 5399 6647
rect 6561 6613 6595 6647
rect 8033 6613 8067 6647
rect 8401 6613 8435 6647
rect 8953 6613 8987 6647
rect 10517 6613 10551 6647
rect 13645 6613 13679 6647
rect 14841 6613 14875 6647
rect 15577 6613 15611 6647
rect 17049 6613 17083 6647
rect 18613 6613 18647 6647
rect 18705 6613 18739 6647
rect 19625 6613 19659 6647
rect 21005 6613 21039 6647
rect 23029 6613 23063 6647
rect 2421 6409 2455 6443
rect 2789 6409 2823 6443
rect 4813 6409 4847 6443
rect 7021 6409 7055 6443
rect 7481 6409 7515 6443
rect 11897 6409 11931 6443
rect 14933 6409 14967 6443
rect 16957 6409 16991 6443
rect 20183 6409 20217 6443
rect 22569 6409 22603 6443
rect 5948 6341 5982 6375
rect 8278 6341 8312 6375
rect 9597 6341 9631 6375
rect 12449 6341 12483 6375
rect 15362 6341 15396 6375
rect 18153 6341 18187 6375
rect 22661 6341 22695 6375
rect 1777 6273 1811 6307
rect 3433 6273 3467 6307
rect 4721 6273 4755 6307
rect 6193 6273 6227 6307
rect 6377 6273 6411 6307
rect 7573 6273 7607 6307
rect 8033 6273 8067 6307
rect 9965 6273 9999 6307
rect 10232 6273 10266 6307
rect 12633 6273 12667 6307
rect 12817 6273 12851 6307
rect 15117 6273 15151 6307
rect 17049 6273 17083 6307
rect 17509 6273 17543 6307
rect 18245 6273 18279 6307
rect 18501 6273 18535 6307
rect 20453 6273 20487 6307
rect 22201 6273 22235 6307
rect 22845 6273 22879 6307
rect 7389 6205 7423 6239
rect 11989 6205 12023 6239
rect 12173 6205 12207 6239
rect 13140 6205 13174 6239
rect 13280 6205 13314 6239
rect 13553 6205 13587 6239
rect 16865 6205 16899 6239
rect 19717 6205 19751 6239
rect 20180 6205 20214 6239
rect 21925 6205 21959 6239
rect 22109 6205 22143 6239
rect 4077 6137 4111 6171
rect 9413 6137 9447 6171
rect 11345 6137 11379 6171
rect 7941 6069 7975 6103
rect 9689 6069 9723 6103
rect 11529 6069 11563 6103
rect 14657 6069 14691 6103
rect 16497 6069 16531 6103
rect 17417 6069 17451 6103
rect 19625 6069 19659 6103
rect 21557 6069 21591 6103
rect 23029 6069 23063 6103
rect 4445 5865 4479 5899
rect 4629 5865 4663 5899
rect 6929 5865 6963 5899
rect 13553 5865 13587 5899
rect 13921 5865 13955 5899
rect 16681 5797 16715 5831
rect 19901 5797 19935 5831
rect 5464 5729 5498 5763
rect 8309 5729 8343 5763
rect 11437 5729 11471 5763
rect 11900 5729 11934 5763
rect 17049 5729 17083 5763
rect 19257 5729 19291 5763
rect 22937 5729 22971 5763
rect 3617 5661 3651 5695
rect 3801 5661 3835 5695
rect 5365 5661 5399 5695
rect 8585 5661 8619 5695
rect 12173 5661 12207 5695
rect 14105 5661 14139 5695
rect 16497 5661 16531 5695
rect 17417 5661 17451 5695
rect 17693 5661 17727 5695
rect 19533 5661 19567 5695
rect 21281 5661 21315 5695
rect 21465 5661 21499 5695
rect 21721 5661 21755 5695
rect 5713 5593 5747 5627
rect 8042 5593 8076 5627
rect 9597 5593 9631 5627
rect 11345 5593 11379 5627
rect 13737 5593 13771 5627
rect 14372 5593 14406 5627
rect 15761 5593 15795 5627
rect 17233 5593 17267 5627
rect 17960 5593 17994 5627
rect 21036 5593 21070 5627
rect 2973 5525 3007 5559
rect 4721 5525 4755 5559
rect 6837 5525 6871 5559
rect 8769 5525 8803 5559
rect 11903 5525 11937 5559
rect 13277 5525 13311 5559
rect 15485 5525 15519 5559
rect 17141 5525 17175 5559
rect 17601 5525 17635 5559
rect 19073 5525 19107 5559
rect 19717 5525 19751 5559
rect 22845 5525 22879 5559
rect 3249 5321 3283 5355
rect 6193 5321 6227 5355
rect 6745 5321 6779 5355
rect 7113 5321 7147 5355
rect 7665 5321 7699 5355
rect 8125 5321 8159 5355
rect 8493 5321 8527 5355
rect 8953 5321 8987 5355
rect 10701 5321 10735 5355
rect 12081 5321 12115 5355
rect 12449 5321 12483 5355
rect 16957 5321 16991 5355
rect 17417 5321 17451 5355
rect 17785 5321 17819 5355
rect 18613 5321 18647 5355
rect 19441 5321 19475 5355
rect 20269 5321 20303 5355
rect 21005 5321 21039 5355
rect 22201 5321 22235 5355
rect 3985 5253 4019 5287
rect 5080 5253 5114 5287
rect 6653 5253 6687 5287
rect 8585 5253 8619 5287
rect 10793 5253 10827 5287
rect 12541 5253 12575 5287
rect 13001 5253 13035 5287
rect 22293 5253 22327 5287
rect 22661 5253 22695 5287
rect 3341 5185 3375 5219
rect 4077 5185 4111 5219
rect 4813 5185 4847 5219
rect 7573 5185 7607 5219
rect 10066 5185 10100 5219
rect 10333 5185 10367 5219
rect 11529 5185 11563 5219
rect 15965 5185 15999 5219
rect 16313 5185 16347 5219
rect 17049 5185 17083 5219
rect 17877 5185 17911 5219
rect 18337 5185 18371 5219
rect 18981 5185 19015 5219
rect 19809 5185 19843 5219
rect 20913 5185 20947 5219
rect 21649 5185 21683 5219
rect 22845 5185 22879 5219
rect 6469 5117 6503 5151
rect 7757 5117 7791 5151
rect 8677 5117 8711 5151
rect 10517 5117 10551 5151
rect 11989 5117 12023 5151
rect 12725 5117 12759 5151
rect 14749 5117 14783 5151
rect 16221 5117 16255 5151
rect 16865 5117 16899 5151
rect 17601 5117 17635 5151
rect 19073 5117 19107 5151
rect 19165 5117 19199 5151
rect 19901 5117 19935 5151
rect 20085 5117 20119 5151
rect 22385 5117 22419 5151
rect 16497 5049 16531 5083
rect 18521 5049 18555 5083
rect 4721 4981 4755 5015
rect 7205 4981 7239 5015
rect 11161 4981 11195 5015
rect 11713 4981 11747 5015
rect 14841 4981 14875 5015
rect 18245 4981 18279 5015
rect 21833 4981 21867 5015
rect 23029 4981 23063 5015
rect 3893 4777 3927 4811
rect 5457 4777 5491 4811
rect 6929 4777 6963 4811
rect 8125 4777 8159 4811
rect 10425 4777 10459 4811
rect 10609 4777 10643 4811
rect 10977 4777 11011 4811
rect 12265 4777 12299 4811
rect 14841 4777 14875 4811
rect 18061 4777 18095 4811
rect 19073 4777 19107 4811
rect 19257 4777 19291 4811
rect 19441 4777 19475 4811
rect 21557 4777 21591 4811
rect 4721 4709 4755 4743
rect 10885 4709 10919 4743
rect 15025 4709 15059 4743
rect 20269 4709 20303 4743
rect 6377 4641 6411 4675
rect 7665 4641 7699 4675
rect 9137 4641 9171 4675
rect 11529 4641 11563 4675
rect 14289 4641 14323 4675
rect 16773 4641 16807 4675
rect 19993 4641 20027 4675
rect 20729 4641 20763 4675
rect 21741 4641 21775 4675
rect 2881 4573 2915 4607
rect 3617 4573 3651 4607
rect 4629 4573 4663 4607
rect 5365 4573 5399 4607
rect 6101 4573 6135 4607
rect 6561 4573 6595 4607
rect 7849 4573 7883 4607
rect 8769 4573 8803 4607
rect 9781 4573 9815 4607
rect 10701 4573 10735 4607
rect 11805 4573 11839 4607
rect 12173 4573 12207 4607
rect 13093 4573 13127 4607
rect 13921 4573 13955 4607
rect 16497 4573 16531 4607
rect 17417 4573 17451 4607
rect 18153 4573 18187 4607
rect 18889 4573 18923 4607
rect 20453 4573 20487 4607
rect 20821 4573 20855 4607
rect 21373 4573 21407 4607
rect 21997 4573 22031 4607
rect 2973 4505 3007 4539
rect 7481 4505 7515 4539
rect 9321 4505 9355 4539
rect 11989 4505 12023 4539
rect 14473 4505 14507 4539
rect 16252 4505 16286 4539
rect 18797 4505 18831 4539
rect 2237 4437 2271 4471
rect 3985 4437 4019 4471
rect 6469 4437 6503 4471
rect 7021 4437 7055 4471
rect 7389 4437 7423 4471
rect 8033 4437 8067 4471
rect 9229 4437 9263 4471
rect 9689 4437 9723 4471
rect 11345 4437 11379 4471
rect 11437 4437 11471 4471
rect 12449 4437 12483 4471
rect 13277 4437 13311 4471
rect 14381 4437 14415 4471
rect 15117 4437 15151 4471
rect 16865 4437 16899 4471
rect 16957 4437 16991 4471
rect 17325 4437 17359 4471
rect 19809 4437 19843 4471
rect 19901 4437 19935 4471
rect 20913 4437 20947 4471
rect 21281 4437 21315 4471
rect 23121 4437 23155 4471
rect 2973 4233 3007 4267
rect 6929 4233 6963 4267
rect 7297 4233 7331 4267
rect 7757 4233 7791 4267
rect 10241 4233 10275 4267
rect 10977 4233 11011 4267
rect 13461 4233 13495 4267
rect 16681 4233 16715 4267
rect 17049 4233 17083 4267
rect 17693 4233 17727 4267
rect 19165 4233 19199 4267
rect 19717 4233 19751 4267
rect 22937 4233 22971 4267
rect 5058 4165 5092 4199
rect 8125 4165 8159 4199
rect 17141 4165 17175 4199
rect 20514 4165 20548 4199
rect 22753 4165 22787 4199
rect 3341 4097 3375 4131
rect 4721 4097 4755 4131
rect 7481 4097 7515 4131
rect 8585 4097 8619 4131
rect 8841 4097 8875 4131
rect 10057 4097 10091 4131
rect 10517 4097 10551 4131
rect 12642 4097 12676 4131
rect 13369 4097 13403 4131
rect 13921 4097 13955 4131
rect 15373 4097 15407 4131
rect 17509 4097 17543 4131
rect 17785 4097 17819 4131
rect 18429 4097 18463 4131
rect 18797 4097 18831 4131
rect 19257 4097 19291 4131
rect 20177 4097 20211 4131
rect 21833 4097 21867 4131
rect 23121 4097 23155 4131
rect 4813 4029 4847 4063
rect 6745 4029 6779 4063
rect 6837 4029 6871 4063
rect 8217 4029 8251 4063
rect 8309 4029 8343 4063
rect 10701 4029 10735 4063
rect 10885 4029 10919 4063
rect 12909 4029 12943 4063
rect 13277 4029 13311 4063
rect 14657 4029 14691 4063
rect 15117 4029 15151 4063
rect 17325 4029 17359 4063
rect 19073 4029 19107 4063
rect 20269 4029 20303 4063
rect 3985 3961 4019 3995
rect 6193 3961 6227 3995
rect 7665 3961 7699 3995
rect 10333 3961 10367 3995
rect 16497 3961 16531 3995
rect 19993 3961 20027 3995
rect 22569 3961 22603 3995
rect 3249 3893 3283 3927
rect 4077 3893 4111 3927
rect 9965 3893 9999 3927
rect 11345 3893 11379 3927
rect 11529 3893 11563 3927
rect 13829 3893 13863 3927
rect 14565 3893 14599 3927
rect 14933 3893 14967 3927
rect 18613 3893 18647 3927
rect 19625 3893 19659 3927
rect 21649 3893 21683 3927
rect 22477 3893 22511 3927
rect 13921 3689 13955 3723
rect 15485 3689 15519 3723
rect 17049 3689 17083 3723
rect 20177 3689 20211 3723
rect 23121 3689 23155 3723
rect 6929 3621 6963 3655
rect 10977 3621 11011 3655
rect 12449 3621 12483 3655
rect 18613 3621 18647 3655
rect 2237 3553 2271 3587
rect 4629 3553 4663 3587
rect 5549 3553 5583 3587
rect 9597 3553 9631 3587
rect 17693 3553 17727 3587
rect 18061 3553 18095 3587
rect 19441 3553 19475 3587
rect 19533 3553 19567 3587
rect 20269 3553 20303 3587
rect 1593 3485 1627 3519
rect 2881 3485 2915 3519
rect 3617 3485 3651 3519
rect 3801 3485 3835 3519
rect 7113 3485 7147 3519
rect 7389 3485 7423 3519
rect 9321 3485 9355 3519
rect 11069 3485 11103 3519
rect 12541 3485 12575 3519
rect 14105 3485 14139 3519
rect 15577 3485 15611 3519
rect 17509 3485 17543 3519
rect 18889 3485 18923 3519
rect 19625 3485 19659 3519
rect 21741 3485 21775 3519
rect 5794 3417 5828 3451
rect 7634 3417 7668 3451
rect 9864 3417 9898 3451
rect 11336 3417 11370 3451
rect 12808 3417 12842 3451
rect 14372 3417 14406 3451
rect 15844 3417 15878 3451
rect 18705 3417 18739 3451
rect 20536 3417 20570 3451
rect 21986 3417 22020 3451
rect 1409 3349 1443 3383
rect 2973 3349 3007 3383
rect 7297 3349 7331 3383
rect 8769 3349 8803 3383
rect 9505 3349 9539 3383
rect 16957 3349 16991 3383
rect 17417 3349 17451 3383
rect 18153 3349 18187 3383
rect 18245 3349 18279 3383
rect 19993 3349 20027 3383
rect 21649 3349 21683 3383
rect 2513 3145 2547 3179
rect 3249 3145 3283 3179
rect 4077 3145 4111 3179
rect 6193 3145 6227 3179
rect 6377 3145 6411 3179
rect 11345 3145 11379 3179
rect 12173 3145 12207 3179
rect 13921 3145 13955 3179
rect 14565 3145 14599 3179
rect 21833 3145 21867 3179
rect 2053 3077 2087 3111
rect 7358 3077 7392 3111
rect 8953 3077 8987 3111
rect 13829 3077 13863 3111
rect 14105 3077 14139 3111
rect 16926 3077 16960 3111
rect 22293 3077 22327 3111
rect 1501 3009 1535 3043
rect 1593 3009 1627 3043
rect 2329 3009 2363 3043
rect 2605 3009 2639 3043
rect 3985 3009 4019 3043
rect 4721 3009 4755 3043
rect 4813 3009 4847 3043
rect 5080 3009 5114 3043
rect 7021 3009 7055 3043
rect 10342 3009 10376 3043
rect 10609 3009 10643 3043
rect 10701 3009 10735 3043
rect 11529 3009 11563 3043
rect 12265 3009 12299 3043
rect 12532 3009 12566 3043
rect 14841 3009 14875 3043
rect 16230 3009 16264 3043
rect 16497 3009 16531 3043
rect 16681 3009 16715 3043
rect 18153 3009 18187 3043
rect 18420 3009 18454 3043
rect 20738 3009 20772 3043
rect 21005 3009 21039 3043
rect 21281 3009 21315 3043
rect 21373 3009 21407 3043
rect 22201 3009 22235 3043
rect 22661 3009 22695 3043
rect 7113 2941 7147 2975
rect 9137 2941 9171 2975
rect 14933 2941 14967 2975
rect 22477 2941 22511 2975
rect 22845 2941 22879 2975
rect 8585 2873 8619 2907
rect 13645 2873 13679 2907
rect 18061 2873 18095 2907
rect 1777 2805 1811 2839
rect 3341 2805 3375 2839
rect 8493 2805 8527 2839
rect 9229 2805 9263 2839
rect 14381 2805 14415 2839
rect 15117 2805 15151 2839
rect 19533 2805 19567 2839
rect 19625 2805 19659 2839
rect 21097 2805 21131 2839
rect 21557 2805 21591 2839
rect 7757 2601 7791 2635
rect 8033 2601 8067 2635
rect 9413 2601 9447 2635
rect 10885 2601 10919 2635
rect 12173 2601 12207 2635
rect 13001 2601 13035 2635
rect 14749 2601 14783 2635
rect 15025 2601 15059 2635
rect 6193 2533 6227 2567
rect 11069 2533 11103 2567
rect 13277 2533 13311 2567
rect 15301 2533 15335 2567
rect 16129 2533 16163 2567
rect 16405 2533 16439 2567
rect 20729 2533 20763 2567
rect 20821 2533 20855 2567
rect 22477 2533 22511 2567
rect 22753 2533 22787 2567
rect 5641 2465 5675 2499
rect 5733 2465 5767 2499
rect 6377 2465 6411 2499
rect 8493 2465 8527 2499
rect 8677 2465 8711 2499
rect 9873 2465 9907 2499
rect 9965 2465 9999 2499
rect 12357 2465 12391 2499
rect 12541 2465 12575 2499
rect 16773 2465 16807 2499
rect 19349 2465 19383 2499
rect 21465 2465 21499 2499
rect 1869 2397 1903 2431
rect 2881 2397 2915 2431
rect 3617 2397 3651 2431
rect 4629 2397 4663 2431
rect 5365 2397 5399 2431
rect 8401 2397 8435 2431
rect 9781 2397 9815 2431
rect 10241 2397 10275 2431
rect 11253 2397 11287 2431
rect 11529 2397 11563 2431
rect 12633 2397 12667 2431
rect 13921 2397 13955 2431
rect 14105 2397 14139 2431
rect 14841 2397 14875 2431
rect 15117 2397 15151 2431
rect 15485 2397 15519 2431
rect 16221 2397 16255 2431
rect 18245 2397 18279 2431
rect 21833 2397 21867 2431
rect 22569 2397 22603 2431
rect 23121 2397 23155 2431
rect 2973 2329 3007 2363
rect 4721 2329 4755 2363
rect 5825 2329 5859 2363
rect 6622 2329 6656 2363
rect 9137 2329 9171 2363
rect 17040 2329 17074 2363
rect 19594 2329 19628 2363
rect 21281 2329 21315 2363
rect 2053 2261 2087 2295
rect 2237 2261 2271 2295
rect 3801 2261 3835 2295
rect 3985 2261 4019 2295
rect 9321 2261 9355 2295
rect 13093 2261 13127 2295
rect 18153 2261 18187 2295
rect 18889 2261 18923 2295
rect 18981 2261 19015 2295
rect 21189 2261 21223 2295
rect 22937 2261 22971 2295
<< metal1 >>
rect 5994 22924 6000 22976
rect 6052 22964 6058 22976
rect 6730 22964 6736 22976
rect 6052 22936 6736 22964
rect 6052 22924 6058 22936
rect 6730 22924 6736 22936
rect 6788 22924 6794 22976
rect 20254 22380 20260 22432
rect 20312 22420 20318 22432
rect 21910 22420 21916 22432
rect 20312 22392 21916 22420
rect 20312 22380 20318 22392
rect 21910 22380 21916 22392
rect 21968 22380 21974 22432
rect 1104 22330 23460 22352
rect 1104 22278 3749 22330
rect 3801 22278 3813 22330
rect 3865 22278 3877 22330
rect 3929 22278 3941 22330
rect 3993 22278 4005 22330
rect 4057 22278 9347 22330
rect 9399 22278 9411 22330
rect 9463 22278 9475 22330
rect 9527 22278 9539 22330
rect 9591 22278 9603 22330
rect 9655 22278 14945 22330
rect 14997 22278 15009 22330
rect 15061 22278 15073 22330
rect 15125 22278 15137 22330
rect 15189 22278 15201 22330
rect 15253 22278 20543 22330
rect 20595 22278 20607 22330
rect 20659 22278 20671 22330
rect 20723 22278 20735 22330
rect 20787 22278 20799 22330
rect 20851 22278 23460 22330
rect 1104 22256 23460 22278
rect 2225 22219 2283 22225
rect 2225 22185 2237 22219
rect 2271 22216 2283 22219
rect 8478 22216 8484 22228
rect 2271 22188 8484 22216
rect 2271 22185 2283 22188
rect 2225 22179 2283 22185
rect 8478 22176 8484 22188
rect 8536 22176 8542 22228
rect 11333 22219 11391 22225
rect 11333 22185 11345 22219
rect 11379 22216 11391 22219
rect 12526 22216 12532 22228
rect 11379 22188 12532 22216
rect 11379 22185 11391 22188
rect 11333 22179 11391 22185
rect 1946 22080 1952 22092
rect 1688 22052 1952 22080
rect 1688 22021 1716 22052
rect 1946 22040 1952 22052
rect 2004 22040 2010 22092
rect 4982 22080 4988 22092
rect 2700 22052 4988 22080
rect 1673 22015 1731 22021
rect 1673 21981 1685 22015
rect 1719 21981 1731 22015
rect 1673 21975 1731 21981
rect 1765 22015 1823 22021
rect 1765 21981 1777 22015
rect 1811 21981 1823 22015
rect 1765 21975 1823 21981
rect 1780 21944 1808 21975
rect 1854 21972 1860 22024
rect 1912 22012 1918 22024
rect 2700 22021 2728 22052
rect 4982 22040 4988 22052
rect 5040 22040 5046 22092
rect 10965 22083 11023 22089
rect 8312 22052 9168 22080
rect 2317 22015 2375 22021
rect 2317 22012 2329 22015
rect 1912 21984 2329 22012
rect 1912 21972 1918 21984
rect 2317 21981 2329 21984
rect 2363 21981 2375 22015
rect 2317 21975 2375 21981
rect 2685 22015 2743 22021
rect 2685 21981 2697 22015
rect 2731 21981 2743 22015
rect 2685 21975 2743 21981
rect 3050 21972 3056 22024
rect 3108 22012 3114 22024
rect 3237 22015 3295 22021
rect 3237 22012 3249 22015
rect 3108 21984 3249 22012
rect 3108 21972 3114 21984
rect 3237 21981 3249 21984
rect 3283 21981 3295 22015
rect 3237 21975 3295 21981
rect 3326 21972 3332 22024
rect 3384 22012 3390 22024
rect 4062 22012 4068 22024
rect 3384 21984 3429 22012
rect 4023 21984 4068 22012
rect 3384 21972 3390 21984
rect 4062 21972 4068 21984
rect 4120 21972 4126 22024
rect 4433 22015 4491 22021
rect 4433 21981 4445 22015
rect 4479 22012 4491 22015
rect 4522 22012 4528 22024
rect 4479 21984 4528 22012
rect 4479 21981 4491 21984
rect 4433 21975 4491 21981
rect 4522 21972 4528 21984
rect 4580 21972 4586 22024
rect 5166 21972 5172 22024
rect 5224 22012 5230 22024
rect 5445 22015 5503 22021
rect 5445 22012 5457 22015
rect 5224 21984 5457 22012
rect 5224 21972 5230 21984
rect 5445 21981 5457 21984
rect 5491 21981 5503 22015
rect 5445 21975 5503 21981
rect 6181 22015 6239 22021
rect 6181 21981 6193 22015
rect 6227 22012 6239 22015
rect 6454 22012 6460 22024
rect 6227 21984 6460 22012
rect 6227 21981 6239 21984
rect 6181 21975 6239 21981
rect 6454 21972 6460 21984
rect 6512 22012 6518 22024
rect 6512 21984 6868 22012
rect 6512 21972 6518 21984
rect 2038 21944 2044 21956
rect 1780 21916 2044 21944
rect 2038 21904 2044 21916
rect 2096 21904 2102 21956
rect 3973 21947 4031 21953
rect 3973 21913 3985 21947
rect 4019 21944 4031 21947
rect 6362 21944 6368 21956
rect 4019 21916 6368 21944
rect 4019 21913 4031 21916
rect 3973 21907 4031 21913
rect 6362 21904 6368 21916
rect 6420 21904 6426 21956
rect 6549 21947 6607 21953
rect 6549 21913 6561 21947
rect 6595 21944 6607 21947
rect 6730 21944 6736 21956
rect 6595 21916 6736 21944
rect 6595 21913 6607 21916
rect 6549 21907 6607 21913
rect 6730 21904 6736 21916
rect 6788 21904 6794 21956
rect 290 21836 296 21888
rect 348 21876 354 21888
rect 1489 21879 1547 21885
rect 1489 21876 1501 21879
rect 348 21848 1501 21876
rect 348 21836 354 21848
rect 1489 21845 1501 21848
rect 1535 21845 1547 21879
rect 1489 21839 1547 21845
rect 1578 21836 1584 21888
rect 1636 21876 1642 21888
rect 1949 21879 2007 21885
rect 1949 21876 1961 21879
rect 1636 21848 1961 21876
rect 1636 21836 1642 21848
rect 1949 21845 1961 21848
rect 1995 21845 2007 21879
rect 1949 21839 2007 21845
rect 2222 21836 2228 21888
rect 2280 21876 2286 21888
rect 2501 21879 2559 21885
rect 2501 21876 2513 21879
rect 2280 21848 2513 21876
rect 2280 21836 2286 21848
rect 2501 21845 2513 21848
rect 2547 21845 2559 21879
rect 2866 21876 2872 21888
rect 2827 21848 2872 21876
rect 2501 21839 2559 21845
rect 2866 21836 2872 21848
rect 2924 21836 2930 21888
rect 2958 21836 2964 21888
rect 3016 21876 3022 21888
rect 3053 21879 3111 21885
rect 3053 21876 3065 21879
rect 3016 21848 3065 21876
rect 3016 21836 3022 21848
rect 3053 21845 3065 21848
rect 3099 21845 3111 21879
rect 3510 21876 3516 21888
rect 3471 21848 3516 21876
rect 3053 21839 3111 21845
rect 3510 21836 3516 21848
rect 3568 21836 3574 21888
rect 4154 21836 4160 21888
rect 4212 21876 4218 21888
rect 4249 21879 4307 21885
rect 4249 21876 4261 21879
rect 4212 21848 4261 21876
rect 4212 21836 4218 21848
rect 4249 21845 4261 21848
rect 4295 21845 4307 21879
rect 4249 21839 4307 21845
rect 4617 21879 4675 21885
rect 4617 21845 4629 21879
rect 4663 21876 4675 21879
rect 4706 21876 4712 21888
rect 4663 21848 4712 21876
rect 4663 21845 4675 21848
rect 4617 21839 4675 21845
rect 4706 21836 4712 21848
rect 4764 21836 4770 21888
rect 4798 21836 4804 21888
rect 4856 21876 4862 21888
rect 5534 21876 5540 21888
rect 4856 21848 4901 21876
rect 5495 21848 5540 21876
rect 4856 21836 4862 21848
rect 5534 21836 5540 21848
rect 5592 21836 5598 21888
rect 5626 21836 5632 21888
rect 5684 21876 5690 21888
rect 6840 21885 6868 21984
rect 7374 21972 7380 22024
rect 7432 22012 7438 22024
rect 8312 22021 8340 22052
rect 9140 22024 9168 22052
rect 10965 22049 10977 22083
rect 11011 22049 11023 22083
rect 10965 22043 11023 22049
rect 8205 22015 8263 22021
rect 8205 22012 8217 22015
rect 7432 21984 8217 22012
rect 7432 21972 7438 21984
rect 8205 21981 8217 21984
rect 8251 21981 8263 22015
rect 8205 21975 8263 21981
rect 8297 22015 8355 22021
rect 8297 21981 8309 22015
rect 8343 21981 8355 22015
rect 8297 21975 8355 21981
rect 8478 21972 8484 22024
rect 8536 22012 8542 22024
rect 8573 22015 8631 22021
rect 8573 22012 8585 22015
rect 8536 21984 8585 22012
rect 8536 21972 8542 21984
rect 8573 21981 8585 21984
rect 8619 21981 8631 22015
rect 8573 21975 8631 21981
rect 8662 21972 8668 22024
rect 8720 22012 8726 22024
rect 8941 22015 8999 22021
rect 8941 22012 8953 22015
rect 8720 21984 8953 22012
rect 8720 21972 8726 21984
rect 8941 21981 8953 21984
rect 8987 21981 8999 22015
rect 8941 21975 8999 21981
rect 9122 21972 9128 22024
rect 9180 21972 9186 22024
rect 10318 22012 10324 22024
rect 10279 21984 10324 22012
rect 10318 21972 10324 21984
rect 10376 22012 10382 22024
rect 10980 22012 11008 22043
rect 11624 22021 11652 22188
rect 12526 22176 12532 22188
rect 12584 22176 12590 22228
rect 17678 22176 17684 22228
rect 17736 22216 17742 22228
rect 17865 22219 17923 22225
rect 17865 22216 17877 22219
rect 17736 22188 17877 22216
rect 17736 22176 17742 22188
rect 17865 22185 17877 22188
rect 17911 22185 17923 22219
rect 19245 22219 19303 22225
rect 19245 22216 19257 22219
rect 17865 22179 17923 22185
rect 17972 22188 19257 22216
rect 13078 22148 13084 22160
rect 11900 22120 13084 22148
rect 11900 22021 11928 22120
rect 13078 22108 13084 22120
rect 13136 22148 13142 22160
rect 13173 22151 13231 22157
rect 13173 22148 13185 22151
rect 13136 22120 13185 22148
rect 13136 22108 13142 22120
rect 13173 22117 13185 22120
rect 13219 22117 13231 22151
rect 13173 22111 13231 22117
rect 17972 22080 18000 22188
rect 19245 22185 19257 22188
rect 19291 22185 19303 22219
rect 22554 22216 22560 22228
rect 19245 22179 19303 22185
rect 19536 22188 22560 22216
rect 12636 22052 18000 22080
rect 10376 21984 11008 22012
rect 11609 22015 11667 22021
rect 10376 21972 10382 21984
rect 11609 21981 11621 22015
rect 11655 21981 11667 22015
rect 11609 21975 11667 21981
rect 11885 22015 11943 22021
rect 11885 21981 11897 22015
rect 11931 21981 11943 22015
rect 12158 22012 12164 22024
rect 12119 21984 12164 22012
rect 11885 21975 11943 21981
rect 12158 21972 12164 21984
rect 12216 21972 12222 22024
rect 12636 22021 12664 22052
rect 12621 22015 12679 22021
rect 12621 21981 12633 22015
rect 12667 21981 12679 22015
rect 12621 21975 12679 21981
rect 12805 22015 12863 22021
rect 12805 21981 12817 22015
rect 12851 22012 12863 22015
rect 13354 22012 13360 22024
rect 12851 21984 13360 22012
rect 12851 21981 12863 21984
rect 12805 21975 12863 21981
rect 13354 21972 13360 21984
rect 13412 21972 13418 22024
rect 13906 22012 13912 22024
rect 13867 21984 13912 22012
rect 13906 21972 13912 21984
rect 13964 21972 13970 22024
rect 14093 22015 14151 22021
rect 14093 21981 14105 22015
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 15565 22015 15623 22021
rect 15565 21981 15577 22015
rect 15611 22012 15623 22015
rect 15654 22012 15660 22024
rect 15611 21984 15660 22012
rect 15611 21981 15623 21984
rect 15565 21975 15623 21981
rect 7960 21947 8018 21953
rect 7960 21913 7972 21947
rect 8006 21944 8018 21947
rect 8110 21944 8116 21956
rect 8006 21916 8116 21944
rect 8006 21913 8018 21916
rect 7960 21907 8018 21913
rect 8110 21904 8116 21916
rect 8168 21904 8174 21956
rect 8386 21904 8392 21956
rect 8444 21944 8450 21956
rect 9585 21947 9643 21953
rect 9585 21944 9597 21947
rect 8444 21916 9597 21944
rect 8444 21904 8450 21916
rect 9585 21913 9597 21916
rect 9631 21913 9643 21947
rect 9585 21907 9643 21913
rect 10781 21947 10839 21953
rect 10781 21913 10793 21947
rect 10827 21944 10839 21947
rect 11514 21944 11520 21956
rect 10827 21916 11520 21944
rect 10827 21913 10839 21916
rect 10781 21907 10839 21913
rect 11514 21904 11520 21916
rect 11572 21904 11578 21956
rect 12434 21944 12440 21956
rect 12360 21916 12440 21944
rect 6457 21879 6515 21885
rect 6457 21876 6469 21879
rect 5684 21848 6469 21876
rect 5684 21836 5690 21848
rect 6457 21845 6469 21848
rect 6503 21845 6515 21879
rect 6457 21839 6515 21845
rect 6825 21879 6883 21885
rect 6825 21845 6837 21879
rect 6871 21845 6883 21879
rect 8478 21876 8484 21888
rect 8439 21848 8484 21876
rect 6825 21839 6883 21845
rect 8478 21836 8484 21848
rect 8536 21836 8542 21888
rect 8754 21876 8760 21888
rect 8715 21848 8760 21876
rect 8754 21836 8760 21848
rect 8812 21836 8818 21888
rect 9677 21879 9735 21885
rect 9677 21845 9689 21879
rect 9723 21876 9735 21879
rect 9950 21876 9956 21888
rect 9723 21848 9956 21876
rect 9723 21845 9735 21848
rect 9677 21839 9735 21845
rect 9950 21836 9956 21848
rect 10008 21836 10014 21888
rect 10413 21879 10471 21885
rect 10413 21845 10425 21879
rect 10459 21876 10471 21879
rect 10502 21876 10508 21888
rect 10459 21848 10508 21876
rect 10459 21845 10471 21848
rect 10413 21839 10471 21845
rect 10502 21836 10508 21848
rect 10560 21836 10566 21888
rect 10873 21879 10931 21885
rect 10873 21845 10885 21879
rect 10919 21876 10931 21879
rect 11054 21876 11060 21888
rect 10919 21848 11060 21876
rect 10919 21845 10931 21848
rect 10873 21839 10931 21845
rect 11054 21836 11060 21848
rect 11112 21836 11118 21888
rect 11790 21876 11796 21888
rect 11751 21848 11796 21876
rect 11790 21836 11796 21848
rect 11848 21836 11854 21888
rect 12066 21876 12072 21888
rect 12027 21848 12072 21876
rect 12066 21836 12072 21848
rect 12124 21836 12130 21888
rect 12360 21885 12388 21916
rect 12434 21904 12440 21916
rect 12492 21904 12498 21956
rect 12986 21944 12992 21956
rect 12947 21916 12992 21944
rect 12986 21904 12992 21916
rect 13044 21904 13050 21956
rect 13630 21904 13636 21956
rect 13688 21944 13694 21956
rect 14108 21944 14136 21975
rect 15654 21972 15660 21984
rect 15712 21972 15718 22024
rect 16298 22012 16304 22024
rect 16259 21984 16304 22012
rect 16298 21972 16304 21984
rect 16356 21972 16362 22024
rect 16853 22015 16911 22021
rect 16853 21981 16865 22015
rect 16899 21981 16911 22015
rect 16853 21975 16911 21981
rect 16574 21944 16580 21956
rect 13688 21916 14136 21944
rect 14568 21916 16580 21944
rect 13688 21904 13694 21916
rect 12345 21879 12403 21885
rect 12345 21845 12357 21879
rect 12391 21845 12403 21879
rect 12345 21839 12403 21845
rect 13265 21879 13323 21885
rect 13265 21845 13277 21879
rect 13311 21876 13323 21879
rect 13722 21876 13728 21888
rect 13311 21848 13728 21876
rect 13311 21845 13323 21848
rect 13265 21839 13323 21845
rect 13722 21836 13728 21848
rect 13780 21836 13786 21888
rect 13814 21836 13820 21888
rect 13872 21876 13878 21888
rect 14568 21876 14596 21916
rect 16574 21904 16580 21916
rect 16632 21904 16638 21956
rect 16868 21944 16896 21975
rect 17218 21972 17224 22024
rect 17276 22012 17282 22024
rect 17589 22015 17647 22021
rect 17589 22012 17601 22015
rect 17276 21984 17601 22012
rect 17276 21972 17282 21984
rect 17589 21981 17601 21984
rect 17635 21981 17647 22015
rect 17589 21975 17647 21981
rect 17678 21972 17684 22024
rect 17736 22012 17742 22024
rect 18049 22015 18107 22021
rect 17736 21984 17781 22012
rect 17736 21972 17742 21984
rect 18049 21981 18061 22015
rect 18095 22012 18107 22015
rect 18138 22012 18144 22024
rect 18095 21984 18144 22012
rect 18095 21981 18107 21984
rect 18049 21975 18107 21981
rect 18138 21972 18144 21984
rect 18196 21972 18202 22024
rect 18506 21972 18512 22024
rect 18564 22012 18570 22024
rect 18785 22015 18843 22021
rect 18785 22012 18797 22015
rect 18564 21984 18797 22012
rect 18564 21972 18570 21984
rect 18785 21981 18797 21984
rect 18831 22012 18843 22015
rect 19242 22012 19248 22024
rect 18831 21984 19248 22012
rect 18831 21981 18843 21984
rect 18785 21975 18843 21981
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 19426 21972 19432 22024
rect 19484 22012 19490 22024
rect 19536 22012 19564 22188
rect 22554 22176 22560 22188
rect 22612 22176 22618 22228
rect 21910 22108 21916 22160
rect 21968 22148 21974 22160
rect 22005 22151 22063 22157
rect 22005 22148 22017 22151
rect 21968 22120 22017 22148
rect 21968 22108 21974 22120
rect 22005 22117 22017 22120
rect 22051 22117 22063 22151
rect 22005 22111 22063 22117
rect 19978 22040 19984 22092
rect 20036 22080 20042 22092
rect 20073 22083 20131 22089
rect 20073 22080 20085 22083
rect 20036 22052 20085 22080
rect 20036 22040 20042 22052
rect 20073 22049 20085 22052
rect 20119 22049 20131 22083
rect 22186 22080 22192 22092
rect 20073 22043 20131 22049
rect 21652 22052 22192 22080
rect 19484 21984 19577 22012
rect 19628 21984 20576 22012
rect 19484 21972 19490 21984
rect 19628 21944 19656 21984
rect 16868 21916 19656 21944
rect 19702 21904 19708 21956
rect 19760 21944 19766 21956
rect 19981 21947 20039 21953
rect 19981 21944 19993 21947
rect 19760 21916 19993 21944
rect 19760 21904 19766 21916
rect 19981 21913 19993 21916
rect 20027 21913 20039 21947
rect 19981 21907 20039 21913
rect 14734 21876 14740 21888
rect 13872 21848 14596 21876
rect 14695 21848 14740 21876
rect 13872 21836 13878 21848
rect 14734 21836 14740 21848
rect 14792 21836 14798 21888
rect 14826 21836 14832 21888
rect 14884 21876 14890 21888
rect 14921 21879 14979 21885
rect 14921 21876 14933 21879
rect 14884 21848 14933 21876
rect 14884 21836 14890 21848
rect 14921 21845 14933 21848
rect 14967 21845 14979 21879
rect 14921 21839 14979 21845
rect 15657 21879 15715 21885
rect 15657 21845 15669 21879
rect 15703 21876 15715 21879
rect 15838 21876 15844 21888
rect 15703 21848 15844 21876
rect 15703 21845 15715 21848
rect 15657 21839 15715 21845
rect 15838 21836 15844 21848
rect 15896 21836 15902 21888
rect 16390 21876 16396 21888
rect 16351 21848 16396 21876
rect 16390 21836 16396 21848
rect 16448 21836 16454 21888
rect 16666 21876 16672 21888
rect 16627 21848 16672 21876
rect 16666 21836 16672 21848
rect 16724 21836 16730 21888
rect 16942 21876 16948 21888
rect 16903 21848 16948 21876
rect 16942 21836 16948 21848
rect 17000 21836 17006 21888
rect 18690 21876 18696 21888
rect 18651 21848 18696 21876
rect 18690 21836 18696 21848
rect 18748 21836 18754 21888
rect 18969 21879 19027 21885
rect 18969 21845 18981 21879
rect 19015 21876 19027 21879
rect 19058 21876 19064 21888
rect 19015 21848 19064 21876
rect 19015 21845 19027 21848
rect 18969 21839 19027 21845
rect 19058 21836 19064 21848
rect 19116 21836 19122 21888
rect 19242 21836 19248 21888
rect 19300 21876 19306 21888
rect 19521 21879 19579 21885
rect 19521 21876 19533 21879
rect 19300 21848 19533 21876
rect 19300 21836 19306 21848
rect 19521 21845 19533 21848
rect 19567 21845 19579 21879
rect 19886 21876 19892 21888
rect 19847 21848 19892 21876
rect 19521 21839 19579 21845
rect 19886 21836 19892 21848
rect 19944 21836 19950 21888
rect 20438 21876 20444 21888
rect 20399 21848 20444 21876
rect 20438 21836 20444 21848
rect 20496 21836 20502 21888
rect 20548 21876 20576 21984
rect 20622 21972 20628 22024
rect 20680 22012 20686 22024
rect 20898 22012 20904 22024
rect 20680 21984 20725 22012
rect 20859 21984 20904 22012
rect 20680 21972 20686 21984
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 21652 22021 21680 22052
rect 22186 22040 22192 22052
rect 22244 22040 22250 22092
rect 21637 22015 21695 22021
rect 21637 21981 21649 22015
rect 21683 21981 21695 22015
rect 21818 22012 21824 22024
rect 21779 21984 21824 22012
rect 21637 21975 21695 21981
rect 21818 21972 21824 21984
rect 21876 21972 21882 22024
rect 22094 21972 22100 22024
rect 22152 22012 22158 22024
rect 22373 22015 22431 22021
rect 22373 22012 22385 22015
rect 22152 21984 22385 22012
rect 22152 21972 22158 21984
rect 22373 21981 22385 21984
rect 22419 21981 22431 22015
rect 22373 21975 22431 21981
rect 22738 21972 22744 22024
rect 22796 22012 22802 22024
rect 23109 22015 23167 22021
rect 23109 22012 23121 22015
rect 22796 21984 23121 22012
rect 22796 21972 22802 21984
rect 23109 21981 23121 21984
rect 23155 21981 23167 22015
rect 23109 21975 23167 21981
rect 22922 21944 22928 21956
rect 22204 21916 22928 21944
rect 20717 21879 20775 21885
rect 20717 21876 20729 21879
rect 20548 21848 20729 21876
rect 20717 21845 20729 21848
rect 20763 21845 20775 21879
rect 20717 21839 20775 21845
rect 20993 21879 21051 21885
rect 20993 21845 21005 21879
rect 21039 21876 21051 21879
rect 21726 21876 21732 21888
rect 21039 21848 21732 21876
rect 21039 21845 21051 21848
rect 20993 21839 21051 21845
rect 21726 21836 21732 21848
rect 21784 21836 21790 21888
rect 22204 21885 22232 21916
rect 22922 21904 22928 21916
rect 22980 21904 22986 21956
rect 22189 21879 22247 21885
rect 22189 21845 22201 21879
rect 22235 21845 22247 21879
rect 22189 21839 22247 21845
rect 22370 21836 22376 21888
rect 22428 21876 22434 21888
rect 22465 21879 22523 21885
rect 22465 21876 22477 21879
rect 22428 21848 22477 21876
rect 22428 21836 22434 21848
rect 22465 21845 22477 21848
rect 22511 21845 22523 21879
rect 22465 21839 22523 21845
rect 1104 21786 23460 21808
rect 1104 21734 6548 21786
rect 6600 21734 6612 21786
rect 6664 21734 6676 21786
rect 6728 21734 6740 21786
rect 6792 21734 6804 21786
rect 6856 21734 12146 21786
rect 12198 21734 12210 21786
rect 12262 21734 12274 21786
rect 12326 21734 12338 21786
rect 12390 21734 12402 21786
rect 12454 21734 17744 21786
rect 17796 21734 17808 21786
rect 17860 21734 17872 21786
rect 17924 21734 17936 21786
rect 17988 21734 18000 21786
rect 18052 21734 23460 21786
rect 1104 21712 23460 21734
rect 934 21632 940 21684
rect 992 21672 998 21684
rect 1489 21675 1547 21681
rect 1489 21672 1501 21675
rect 992 21644 1501 21672
rect 992 21632 998 21644
rect 1489 21641 1501 21644
rect 1535 21641 1547 21675
rect 1489 21635 1547 21641
rect 2866 21632 2872 21684
rect 2924 21672 2930 21684
rect 4246 21672 4252 21684
rect 2924 21644 4252 21672
rect 2924 21632 2930 21644
rect 4246 21632 4252 21644
rect 4304 21632 4310 21684
rect 4801 21675 4859 21681
rect 4801 21641 4813 21675
rect 4847 21672 4859 21675
rect 5626 21672 5632 21684
rect 4847 21644 5212 21672
rect 4847 21641 4859 21644
rect 4801 21635 4859 21641
rect 5184 21616 5212 21644
rect 5276 21644 5632 21672
rect 2498 21564 2504 21616
rect 2556 21604 2562 21616
rect 4062 21604 4068 21616
rect 2556 21576 4068 21604
rect 2556 21564 2562 21576
rect 4062 21564 4068 21576
rect 4120 21564 4126 21616
rect 4982 21604 4988 21616
rect 4943 21576 4988 21604
rect 4982 21564 4988 21576
rect 5040 21564 5046 21616
rect 5166 21604 5172 21616
rect 5127 21576 5172 21604
rect 5166 21564 5172 21576
rect 5224 21564 5230 21616
rect 1673 21539 1731 21545
rect 1673 21505 1685 21539
rect 1719 21505 1731 21539
rect 1673 21499 1731 21505
rect 1688 21400 1716 21499
rect 1762 21496 1768 21548
rect 1820 21536 1826 21548
rect 2869 21539 2927 21545
rect 1820 21508 1865 21536
rect 1820 21496 1826 21508
rect 2869 21505 2881 21539
rect 2915 21536 2927 21539
rect 2958 21536 2964 21548
rect 2915 21508 2964 21536
rect 2915 21505 2927 21508
rect 2869 21499 2927 21505
rect 2958 21496 2964 21508
rect 3016 21496 3022 21548
rect 3688 21539 3746 21545
rect 3688 21505 3700 21539
rect 3734 21536 3746 21539
rect 4706 21536 4712 21548
rect 3734 21508 4712 21536
rect 3734 21505 3746 21508
rect 3688 21499 3746 21505
rect 4706 21496 4712 21508
rect 4764 21496 4770 21548
rect 2590 21468 2596 21480
rect 2551 21440 2596 21468
rect 2590 21428 2596 21440
rect 2648 21428 2654 21480
rect 2774 21428 2780 21480
rect 2832 21468 2838 21480
rect 3418 21468 3424 21480
rect 2832 21440 2877 21468
rect 3379 21440 3424 21468
rect 2832 21428 2838 21440
rect 3418 21428 3424 21440
rect 3476 21428 3482 21480
rect 4430 21428 4436 21480
rect 4488 21468 4494 21480
rect 5276 21468 5304 21644
rect 5626 21632 5632 21644
rect 5684 21632 5690 21684
rect 6362 21632 6368 21684
rect 6420 21672 6426 21684
rect 6825 21675 6883 21681
rect 6825 21672 6837 21675
rect 6420 21644 6837 21672
rect 6420 21632 6426 21644
rect 6825 21641 6837 21644
rect 6871 21641 6883 21675
rect 6825 21635 6883 21641
rect 6914 21632 6920 21684
rect 6972 21672 6978 21684
rect 6972 21644 8064 21672
rect 6972 21632 6978 21644
rect 5534 21564 5540 21616
rect 5592 21604 5598 21616
rect 7530 21607 7588 21613
rect 7530 21604 7542 21607
rect 5592 21576 7542 21604
rect 5592 21564 5598 21576
rect 7530 21573 7542 21576
rect 7576 21573 7588 21607
rect 7530 21567 7588 21573
rect 5353 21539 5411 21545
rect 5353 21505 5365 21539
rect 5399 21536 5411 21539
rect 5399 21508 5672 21536
rect 5399 21505 5411 21508
rect 5353 21499 5411 21505
rect 4488 21440 5304 21468
rect 4488 21428 4494 21440
rect 2682 21400 2688 21412
rect 1688 21372 2688 21400
rect 2682 21360 2688 21372
rect 2740 21360 2746 21412
rect 5644 21400 5672 21508
rect 5718 21496 5724 21548
rect 5776 21536 5782 21548
rect 6181 21539 6239 21545
rect 6181 21536 6193 21539
rect 5776 21508 6193 21536
rect 5776 21496 5782 21508
rect 6181 21505 6193 21508
rect 6227 21505 6239 21539
rect 6181 21499 6239 21505
rect 7285 21539 7343 21545
rect 7285 21505 7297 21539
rect 7331 21536 7343 21539
rect 7374 21536 7380 21548
rect 7331 21508 7380 21536
rect 7331 21505 7343 21508
rect 7285 21499 7343 21505
rect 7374 21496 7380 21508
rect 7432 21496 7438 21548
rect 8036 21536 8064 21644
rect 8938 21632 8944 21684
rect 8996 21672 9002 21684
rect 9401 21675 9459 21681
rect 9401 21672 9413 21675
rect 8996 21644 9413 21672
rect 8996 21632 9002 21644
rect 9401 21641 9413 21644
rect 9447 21641 9459 21675
rect 9858 21672 9864 21684
rect 9401 21635 9459 21641
rect 9508 21644 9864 21672
rect 8110 21564 8116 21616
rect 8168 21604 8174 21616
rect 9214 21604 9220 21616
rect 8168 21576 9220 21604
rect 8168 21564 8174 21576
rect 9214 21564 9220 21576
rect 9272 21564 9278 21616
rect 8849 21539 8907 21545
rect 8036 21508 8800 21536
rect 6454 21428 6460 21480
rect 6512 21468 6518 21480
rect 6549 21471 6607 21477
rect 6549 21468 6561 21471
rect 6512 21440 6561 21468
rect 6512 21428 6518 21440
rect 6549 21437 6561 21440
rect 6595 21437 6607 21471
rect 6549 21431 6607 21437
rect 6733 21471 6791 21477
rect 6733 21437 6745 21471
rect 6779 21468 6791 21471
rect 7190 21468 7196 21480
rect 6779 21440 7196 21468
rect 6779 21437 6791 21440
rect 6733 21431 6791 21437
rect 7190 21428 7196 21440
rect 7248 21428 7254 21480
rect 8772 21468 8800 21508
rect 8849 21505 8861 21539
rect 8895 21536 8907 21539
rect 9030 21536 9036 21548
rect 8895 21508 9036 21536
rect 8895 21505 8907 21508
rect 8849 21499 8907 21505
rect 9030 21496 9036 21508
rect 9088 21496 9094 21548
rect 9122 21496 9128 21548
rect 9180 21536 9186 21548
rect 9309 21539 9367 21545
rect 9309 21536 9321 21539
rect 9180 21508 9321 21536
rect 9180 21496 9186 21508
rect 9309 21505 9321 21508
rect 9355 21536 9367 21539
rect 9508 21536 9536 21644
rect 9858 21632 9864 21644
rect 9916 21632 9922 21684
rect 9953 21675 10011 21681
rect 9953 21641 9965 21675
rect 9999 21672 10011 21675
rect 10318 21672 10324 21684
rect 9999 21644 10324 21672
rect 9999 21641 10011 21644
rect 9953 21635 10011 21641
rect 10318 21632 10324 21644
rect 10376 21632 10382 21684
rect 12437 21675 12495 21681
rect 12437 21641 12449 21675
rect 12483 21672 12495 21675
rect 12986 21672 12992 21684
rect 12483 21644 12992 21672
rect 12483 21641 12495 21644
rect 12437 21635 12495 21641
rect 12986 21632 12992 21644
rect 13044 21632 13050 21684
rect 14182 21632 14188 21684
rect 14240 21672 14246 21684
rect 14240 21644 15700 21672
rect 14240 21632 14246 21644
rect 10226 21604 10232 21616
rect 9600 21576 10232 21604
rect 9600 21545 9628 21576
rect 10226 21564 10232 21576
rect 10284 21604 10290 21616
rect 10594 21604 10600 21616
rect 10284 21576 10600 21604
rect 10284 21564 10290 21576
rect 10594 21564 10600 21576
rect 10652 21564 10658 21616
rect 11088 21607 11146 21613
rect 11088 21573 11100 21607
rect 11134 21604 11146 21607
rect 11517 21607 11575 21613
rect 11517 21604 11529 21607
rect 11134 21576 11529 21604
rect 11134 21573 11146 21576
rect 11088 21567 11146 21573
rect 11517 21573 11529 21576
rect 11563 21573 11575 21607
rect 11517 21567 11575 21573
rect 12526 21564 12532 21616
rect 12584 21604 12590 21616
rect 12584 21576 15608 21604
rect 12584 21564 12590 21576
rect 9355 21508 9536 21536
rect 9585 21539 9643 21545
rect 9355 21505 9367 21508
rect 9309 21499 9367 21505
rect 9585 21505 9597 21539
rect 9631 21505 9643 21539
rect 9585 21499 9643 21505
rect 9674 21496 9680 21548
rect 9732 21536 9738 21548
rect 11238 21536 11244 21548
rect 9732 21508 11244 21536
rect 9732 21496 9738 21508
rect 11238 21496 11244 21508
rect 11296 21496 11302 21548
rect 12158 21536 12164 21548
rect 12119 21508 12164 21536
rect 12158 21496 12164 21508
rect 12216 21496 12222 21548
rect 12253 21539 12311 21545
rect 12253 21505 12265 21539
rect 12299 21536 12311 21539
rect 13173 21539 13231 21545
rect 12299 21508 13124 21536
rect 12299 21505 12311 21508
rect 12253 21499 12311 21505
rect 10042 21468 10048 21480
rect 8772 21440 10048 21468
rect 10042 21428 10048 21440
rect 10100 21428 10106 21480
rect 11330 21468 11336 21480
rect 11291 21440 11336 21468
rect 11330 21428 11336 21440
rect 11388 21428 11394 21480
rect 9033 21403 9091 21409
rect 5644 21372 7328 21400
rect 2314 21292 2320 21344
rect 2372 21332 2378 21344
rect 2409 21335 2467 21341
rect 2409 21332 2421 21335
rect 2372 21304 2421 21332
rect 2372 21292 2378 21304
rect 2409 21301 2421 21304
rect 2455 21301 2467 21335
rect 3234 21332 3240 21344
rect 3195 21304 3240 21332
rect 2409 21295 2467 21301
rect 3234 21292 3240 21304
rect 3292 21292 3298 21344
rect 5074 21292 5080 21344
rect 5132 21332 5138 21344
rect 5537 21335 5595 21341
rect 5537 21332 5549 21335
rect 5132 21304 5549 21332
rect 5132 21292 5138 21304
rect 5537 21301 5549 21304
rect 5583 21301 5595 21335
rect 5537 21295 5595 21301
rect 7098 21292 7104 21344
rect 7156 21332 7162 21344
rect 7193 21335 7251 21341
rect 7193 21332 7205 21335
rect 7156 21304 7205 21332
rect 7156 21292 7162 21304
rect 7193 21301 7205 21304
rect 7239 21301 7251 21335
rect 7300 21332 7328 21372
rect 8220 21372 8800 21400
rect 8220 21332 8248 21372
rect 8662 21332 8668 21344
rect 7300 21304 8248 21332
rect 8623 21304 8668 21332
rect 7193 21295 7251 21301
rect 8662 21292 8668 21304
rect 8720 21292 8726 21344
rect 8772 21332 8800 21372
rect 9033 21369 9045 21403
rect 9079 21400 9091 21403
rect 9766 21400 9772 21412
rect 9079 21372 9772 21400
rect 9079 21369 9091 21372
rect 9033 21363 9091 21369
rect 9766 21360 9772 21372
rect 9824 21360 9830 21412
rect 12066 21360 12072 21412
rect 12124 21400 12130 21412
rect 12894 21400 12900 21412
rect 12124 21372 12900 21400
rect 12124 21360 12130 21372
rect 12894 21360 12900 21372
rect 12952 21360 12958 21412
rect 13096 21400 13124 21508
rect 13173 21505 13185 21539
rect 13219 21536 13231 21539
rect 13262 21536 13268 21548
rect 13219 21508 13268 21536
rect 13219 21505 13231 21508
rect 13173 21499 13231 21505
rect 13262 21496 13268 21508
rect 13320 21496 13326 21548
rect 13633 21539 13691 21545
rect 13633 21505 13645 21539
rect 13679 21536 13691 21539
rect 14090 21536 14096 21548
rect 13679 21508 14096 21536
rect 13679 21505 13691 21508
rect 13633 21499 13691 21505
rect 14090 21496 14096 21508
rect 14148 21496 14154 21548
rect 14292 21545 14320 21576
rect 14277 21539 14335 21545
rect 14277 21505 14289 21539
rect 14323 21505 14335 21539
rect 14277 21499 14335 21505
rect 14544 21539 14602 21545
rect 14544 21505 14556 21539
rect 14590 21536 14602 21539
rect 14590 21508 15516 21536
rect 14590 21505 14602 21508
rect 14544 21499 14602 21505
rect 13354 21468 13360 21480
rect 13315 21440 13360 21468
rect 13354 21428 13360 21440
rect 13412 21428 13418 21480
rect 13538 21468 13544 21480
rect 13499 21440 13544 21468
rect 13538 21428 13544 21440
rect 13596 21428 13602 21480
rect 13722 21428 13728 21480
rect 13780 21468 13786 21480
rect 13780 21440 14320 21468
rect 13780 21428 13786 21440
rect 13170 21400 13176 21412
rect 13083 21372 13176 21400
rect 13170 21360 13176 21372
rect 13228 21400 13234 21412
rect 14093 21403 14151 21409
rect 14093 21400 14105 21403
rect 13228 21372 14105 21400
rect 13228 21360 13234 21372
rect 14093 21369 14105 21372
rect 14139 21369 14151 21403
rect 14093 21363 14151 21369
rect 9125 21335 9183 21341
rect 9125 21332 9137 21335
rect 8772 21304 9137 21332
rect 9125 21301 9137 21304
rect 9171 21301 9183 21335
rect 9125 21295 9183 21301
rect 9861 21335 9919 21341
rect 9861 21301 9873 21335
rect 9907 21332 9919 21335
rect 10410 21332 10416 21344
rect 9907 21304 10416 21332
rect 9907 21301 9919 21304
rect 9861 21295 9919 21301
rect 10410 21292 10416 21304
rect 10468 21292 10474 21344
rect 12529 21335 12587 21341
rect 12529 21301 12541 21335
rect 12575 21332 12587 21335
rect 13722 21332 13728 21344
rect 12575 21304 13728 21332
rect 12575 21301 12587 21304
rect 12529 21295 12587 21301
rect 13722 21292 13728 21304
rect 13780 21292 13786 21344
rect 13814 21292 13820 21344
rect 13872 21332 13878 21344
rect 14001 21335 14059 21341
rect 14001 21332 14013 21335
rect 13872 21304 14013 21332
rect 13872 21292 13878 21304
rect 14001 21301 14013 21304
rect 14047 21301 14059 21335
rect 14292 21332 14320 21440
rect 15488 21400 15516 21508
rect 15580 21480 15608 21576
rect 15672 21536 15700 21644
rect 16574 21632 16580 21684
rect 16632 21672 16638 21684
rect 18049 21675 18107 21681
rect 16632 21644 18000 21672
rect 16632 21632 16638 21644
rect 16942 21613 16948 21616
rect 16936 21604 16948 21613
rect 16903 21576 16948 21604
rect 16936 21567 16948 21576
rect 16942 21564 16948 21567
rect 17000 21564 17006 21616
rect 17972 21604 18000 21644
rect 18049 21641 18061 21675
rect 18095 21672 18107 21675
rect 18138 21672 18144 21684
rect 18095 21644 18144 21672
rect 18095 21641 18107 21644
rect 18049 21635 18107 21641
rect 18138 21632 18144 21644
rect 18196 21632 18202 21684
rect 19426 21672 19432 21684
rect 18340 21644 19432 21672
rect 18340 21604 18368 21644
rect 19426 21632 19432 21644
rect 19484 21632 19490 21684
rect 19610 21632 19616 21684
rect 19668 21672 19674 21684
rect 21269 21675 21327 21681
rect 21269 21672 21281 21675
rect 19668 21644 21281 21672
rect 19668 21632 19674 21644
rect 21269 21641 21281 21644
rect 21315 21641 21327 21675
rect 21269 21635 21327 21641
rect 22002 21632 22008 21684
rect 22060 21672 22066 21684
rect 22741 21675 22799 21681
rect 22741 21672 22753 21675
rect 22060 21644 22753 21672
rect 22060 21632 22066 21644
rect 22741 21641 22753 21644
rect 22787 21641 22799 21675
rect 22741 21635 22799 21641
rect 17972 21576 18368 21604
rect 18408 21607 18466 21613
rect 18408 21573 18420 21607
rect 18454 21604 18466 21607
rect 18690 21604 18696 21616
rect 18454 21576 18696 21604
rect 18454 21573 18466 21576
rect 18408 21567 18466 21573
rect 18690 21564 18696 21576
rect 18748 21564 18754 21616
rect 19058 21564 19064 21616
rect 19116 21604 19122 21616
rect 24118 21604 24124 21616
rect 19116 21576 24124 21604
rect 19116 21564 19122 21576
rect 24118 21564 24124 21576
rect 24176 21564 24182 21616
rect 15749 21539 15807 21545
rect 15749 21536 15761 21539
rect 15672 21508 15761 21536
rect 15749 21505 15761 21508
rect 15795 21505 15807 21539
rect 15749 21499 15807 21505
rect 15930 21496 15936 21548
rect 15988 21536 15994 21548
rect 20346 21536 20352 21548
rect 15988 21508 20352 21536
rect 15988 21496 15994 21508
rect 20346 21496 20352 21508
rect 20404 21496 20410 21548
rect 20737 21539 20795 21545
rect 20737 21505 20749 21539
rect 20783 21536 20795 21539
rect 20898 21536 20904 21548
rect 20783 21508 20904 21536
rect 20783 21505 20795 21508
rect 20737 21499 20795 21505
rect 20898 21496 20904 21508
rect 20956 21496 20962 21548
rect 21082 21536 21088 21548
rect 21043 21508 21088 21536
rect 21082 21496 21088 21508
rect 21140 21496 21146 21548
rect 21634 21536 21640 21548
rect 21595 21508 21640 21536
rect 21634 21496 21640 21508
rect 21692 21496 21698 21548
rect 22462 21536 22468 21548
rect 22423 21508 22468 21536
rect 22462 21496 22468 21508
rect 22520 21496 22526 21548
rect 22557 21539 22615 21545
rect 22557 21505 22569 21539
rect 22603 21505 22615 21539
rect 22557 21499 22615 21505
rect 15562 21428 15568 21480
rect 15620 21468 15626 21480
rect 16669 21471 16727 21477
rect 16669 21468 16681 21471
rect 15620 21440 16681 21468
rect 15620 21428 15626 21440
rect 16669 21437 16681 21440
rect 16715 21437 16727 21471
rect 18138 21468 18144 21480
rect 18099 21440 18144 21468
rect 16669 21431 16727 21437
rect 18138 21428 18144 21440
rect 18196 21428 18202 21480
rect 20990 21468 20996 21480
rect 20951 21440 20996 21468
rect 20990 21428 20996 21440
rect 21048 21428 21054 21480
rect 21358 21428 21364 21480
rect 21416 21468 21422 21480
rect 21818 21468 21824 21480
rect 21416 21440 21824 21468
rect 21416 21428 21422 21440
rect 21818 21428 21824 21440
rect 21876 21428 21882 21480
rect 22572 21468 22600 21499
rect 22646 21496 22652 21548
rect 22704 21536 22710 21548
rect 23109 21539 23167 21545
rect 23109 21536 23121 21539
rect 22704 21508 23121 21536
rect 22704 21496 22710 21508
rect 23109 21505 23121 21508
rect 23155 21505 23167 21539
rect 23109 21499 23167 21505
rect 23474 21468 23480 21480
rect 22572 21440 23480 21468
rect 23474 21428 23480 21440
rect 23532 21428 23538 21480
rect 16393 21403 16451 21409
rect 16393 21400 16405 21403
rect 15488 21372 16405 21400
rect 16393 21369 16405 21372
rect 16439 21369 16451 21403
rect 19978 21400 19984 21412
rect 16393 21363 16451 21369
rect 19628 21372 19984 21400
rect 19628 21344 19656 21372
rect 19978 21360 19984 21372
rect 20036 21360 20042 21412
rect 15378 21332 15384 21344
rect 14292 21304 15384 21332
rect 14001 21295 14059 21301
rect 15378 21292 15384 21304
rect 15436 21292 15442 21344
rect 15657 21335 15715 21341
rect 15657 21301 15669 21335
rect 15703 21332 15715 21335
rect 15746 21332 15752 21344
rect 15703 21304 15752 21332
rect 15703 21301 15715 21304
rect 15657 21295 15715 21301
rect 15746 21292 15752 21304
rect 15804 21292 15810 21344
rect 15930 21292 15936 21344
rect 15988 21332 15994 21344
rect 19242 21332 19248 21344
rect 15988 21304 19248 21332
rect 15988 21292 15994 21304
rect 19242 21292 19248 21304
rect 19300 21292 19306 21344
rect 19518 21332 19524 21344
rect 19479 21304 19524 21332
rect 19518 21292 19524 21304
rect 19576 21292 19582 21344
rect 19610 21292 19616 21344
rect 19668 21332 19674 21344
rect 19668 21304 19713 21332
rect 19668 21292 19674 21304
rect 19794 21292 19800 21344
rect 19852 21332 19858 21344
rect 21453 21335 21511 21341
rect 21453 21332 21465 21335
rect 19852 21304 21465 21332
rect 19852 21292 19858 21304
rect 21453 21301 21465 21304
rect 21499 21301 21511 21335
rect 21818 21332 21824 21344
rect 21779 21304 21824 21332
rect 21453 21295 21511 21301
rect 21818 21292 21824 21304
rect 21876 21292 21882 21344
rect 22830 21292 22836 21344
rect 22888 21332 22894 21344
rect 22925 21335 22983 21341
rect 22925 21332 22937 21335
rect 22888 21304 22937 21332
rect 22888 21292 22894 21304
rect 22925 21301 22937 21304
rect 22971 21301 22983 21335
rect 22925 21295 22983 21301
rect 1104 21242 23460 21264
rect 1104 21190 3749 21242
rect 3801 21190 3813 21242
rect 3865 21190 3877 21242
rect 3929 21190 3941 21242
rect 3993 21190 4005 21242
rect 4057 21190 9347 21242
rect 9399 21190 9411 21242
rect 9463 21190 9475 21242
rect 9527 21190 9539 21242
rect 9591 21190 9603 21242
rect 9655 21190 14945 21242
rect 14997 21190 15009 21242
rect 15061 21190 15073 21242
rect 15125 21190 15137 21242
rect 15189 21190 15201 21242
rect 15253 21190 20543 21242
rect 20595 21190 20607 21242
rect 20659 21190 20671 21242
rect 20723 21190 20735 21242
rect 20787 21190 20799 21242
rect 20851 21190 23460 21242
rect 1104 21168 23460 21190
rect 2590 21128 2596 21140
rect 1688 21100 2596 21128
rect 1688 21060 1716 21100
rect 2590 21088 2596 21100
rect 2648 21088 2654 21140
rect 4249 21131 4307 21137
rect 4249 21097 4261 21131
rect 4295 21128 4307 21131
rect 7650 21128 7656 21140
rect 4295 21100 7656 21128
rect 4295 21097 4307 21100
rect 4249 21091 4307 21097
rect 7650 21088 7656 21100
rect 7708 21088 7714 21140
rect 7742 21088 7748 21140
rect 7800 21128 7806 21140
rect 7800 21100 8800 21128
rect 7800 21088 7806 21100
rect 1596 21032 1716 21060
rect 1596 21001 1624 21032
rect 5350 21020 5356 21072
rect 5408 21060 5414 21072
rect 5718 21060 5724 21072
rect 5408 21032 5724 21060
rect 5408 21020 5414 21032
rect 5718 21020 5724 21032
rect 5776 21020 5782 21072
rect 1581 20995 1639 21001
rect 1581 20961 1593 20995
rect 1627 20961 1639 20995
rect 1581 20955 1639 20961
rect 1673 20995 1731 21001
rect 1673 20961 1685 20995
rect 1719 20992 1731 20995
rect 1762 20992 1768 21004
rect 1719 20964 1768 20992
rect 1719 20961 1731 20964
rect 1673 20955 1731 20961
rect 1762 20952 1768 20964
rect 1820 20952 1826 21004
rect 7098 20952 7104 21004
rect 7156 20992 7162 21004
rect 7650 20992 7656 21004
rect 7156 20964 7656 20992
rect 7156 20952 7162 20964
rect 7650 20952 7656 20964
rect 7708 20952 7714 21004
rect 8772 20992 8800 21100
rect 9214 21088 9220 21140
rect 9272 21128 9278 21140
rect 9585 21131 9643 21137
rect 9585 21128 9597 21131
rect 9272 21100 9597 21128
rect 9272 21088 9278 21100
rect 9585 21097 9597 21100
rect 9631 21097 9643 21131
rect 11330 21128 11336 21140
rect 9585 21091 9643 21097
rect 10060 21100 11336 21128
rect 9398 21020 9404 21072
rect 9456 21060 9462 21072
rect 9674 21060 9680 21072
rect 9456 21032 9680 21060
rect 9456 21020 9462 21032
rect 9674 21020 9680 21032
rect 9732 21060 9738 21072
rect 10060 21060 10088 21100
rect 11330 21088 11336 21100
rect 11388 21088 11394 21140
rect 11425 21131 11483 21137
rect 11425 21097 11437 21131
rect 11471 21128 11483 21131
rect 11882 21128 11888 21140
rect 11471 21100 11888 21128
rect 11471 21097 11483 21100
rect 11425 21091 11483 21097
rect 11882 21088 11888 21100
rect 11940 21128 11946 21140
rect 12158 21128 12164 21140
rect 11940 21100 12164 21128
rect 11940 21088 11946 21100
rect 12158 21088 12164 21100
rect 12216 21088 12222 21140
rect 12894 21088 12900 21140
rect 12952 21128 12958 21140
rect 13998 21128 14004 21140
rect 12952 21100 14004 21128
rect 12952 21088 12958 21100
rect 13998 21088 14004 21100
rect 14056 21088 14062 21140
rect 14093 21131 14151 21137
rect 14093 21097 14105 21131
rect 14139 21128 14151 21131
rect 14182 21128 14188 21140
rect 14139 21100 14188 21128
rect 14139 21097 14151 21100
rect 14093 21091 14151 21097
rect 14182 21088 14188 21100
rect 14240 21088 14246 21140
rect 18969 21131 19027 21137
rect 14568 21100 18920 21128
rect 9732 21032 10088 21060
rect 9732 21020 9738 21032
rect 10060 21001 10088 21032
rect 13906 21020 13912 21072
rect 13964 21060 13970 21072
rect 14568 21060 14596 21100
rect 13964 21032 14596 21060
rect 16945 21063 17003 21069
rect 13964 21020 13970 21032
rect 16945 21029 16957 21063
rect 16991 21029 17003 21063
rect 18892 21060 18920 21100
rect 18969 21097 18981 21131
rect 19015 21128 19027 21131
rect 19150 21128 19156 21140
rect 19015 21100 19156 21128
rect 19015 21097 19027 21100
rect 18969 21091 19027 21097
rect 19150 21088 19156 21100
rect 19208 21088 19214 21140
rect 19242 21088 19248 21140
rect 19300 21128 19306 21140
rect 20162 21128 20168 21140
rect 19300 21100 20168 21128
rect 19300 21088 19306 21100
rect 20162 21088 20168 21100
rect 20220 21088 20226 21140
rect 20346 21088 20352 21140
rect 20404 21128 20410 21140
rect 21361 21131 21419 21137
rect 21361 21128 21373 21131
rect 20404 21100 21373 21128
rect 20404 21088 20410 21100
rect 21361 21097 21373 21100
rect 21407 21128 21419 21131
rect 21634 21128 21640 21140
rect 21407 21100 21640 21128
rect 21407 21097 21419 21100
rect 21361 21091 21419 21097
rect 21634 21088 21640 21100
rect 21692 21088 21698 21140
rect 19610 21060 19616 21072
rect 18892 21032 19616 21060
rect 16945 21023 17003 21029
rect 10045 20995 10103 21001
rect 8772 20964 8984 20992
rect 2222 20924 2228 20936
rect 2183 20896 2228 20924
rect 2222 20884 2228 20896
rect 2280 20884 2286 20936
rect 2314 20884 2320 20936
rect 2372 20924 2378 20936
rect 2372 20896 2452 20924
rect 2372 20884 2378 20896
rect 1765 20859 1823 20865
rect 1765 20825 1777 20859
rect 1811 20856 1823 20859
rect 2424 20856 2452 20896
rect 3602 20884 3608 20936
rect 3660 20924 3666 20936
rect 3789 20927 3847 20933
rect 3789 20924 3801 20927
rect 3660 20896 3801 20924
rect 3660 20884 3666 20896
rect 3789 20893 3801 20896
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 4062 20884 4068 20936
rect 4120 20924 4126 20936
rect 4341 20927 4399 20933
rect 4341 20924 4353 20927
rect 4120 20896 4353 20924
rect 4120 20884 4126 20896
rect 4341 20893 4353 20896
rect 4387 20893 4399 20927
rect 5902 20924 5908 20936
rect 5863 20896 5908 20924
rect 4341 20887 4399 20893
rect 5902 20884 5908 20896
rect 5960 20884 5966 20936
rect 7285 20927 7343 20933
rect 7285 20893 7297 20927
rect 7331 20893 7343 20927
rect 7285 20887 7343 20893
rect 2481 20859 2539 20865
rect 2481 20856 2493 20859
rect 1811 20828 2360 20856
rect 2424 20828 2493 20856
rect 1811 20825 1823 20828
rect 1765 20819 1823 20825
rect 2130 20788 2136 20800
rect 2091 20760 2136 20788
rect 2130 20748 2136 20760
rect 2188 20748 2194 20800
rect 2332 20788 2360 20828
rect 2481 20825 2493 20828
rect 2527 20825 2539 20859
rect 2481 20819 2539 20825
rect 2590 20816 2596 20868
rect 2648 20856 2654 20868
rect 3973 20859 4031 20865
rect 3973 20856 3985 20859
rect 2648 20828 3985 20856
rect 2648 20816 2654 20828
rect 3973 20825 3985 20828
rect 4019 20856 4031 20859
rect 4608 20859 4666 20865
rect 4019 20828 4568 20856
rect 4019 20825 4031 20828
rect 3973 20819 4031 20825
rect 3605 20791 3663 20797
rect 3605 20788 3617 20791
rect 2332 20760 3617 20788
rect 3605 20757 3617 20760
rect 3651 20788 3663 20791
rect 3694 20788 3700 20800
rect 3651 20760 3700 20788
rect 3651 20757 3663 20760
rect 3605 20751 3663 20757
rect 3694 20748 3700 20760
rect 3752 20748 3758 20800
rect 4540 20788 4568 20828
rect 4608 20825 4620 20859
rect 4654 20856 4666 20859
rect 4798 20856 4804 20868
rect 4654 20828 4804 20856
rect 4654 20825 4666 20828
rect 4608 20819 4666 20825
rect 4798 20816 4804 20828
rect 4856 20816 4862 20868
rect 7300 20856 7328 20887
rect 7374 20884 7380 20936
rect 7432 20924 7438 20936
rect 8956 20933 8984 20964
rect 10045 20961 10057 20995
rect 10091 20961 10103 20995
rect 11514 20992 11520 21004
rect 11475 20964 11520 20992
rect 10045 20955 10103 20961
rect 11514 20952 11520 20964
rect 11572 20952 11578 21004
rect 12526 20992 12532 21004
rect 12487 20964 12532 20992
rect 12526 20952 12532 20964
rect 12584 20952 12590 21004
rect 15473 20995 15531 21001
rect 15473 20961 15485 20995
rect 15519 20992 15531 20995
rect 15562 20992 15568 21004
rect 15519 20964 15568 20992
rect 15519 20961 15531 20964
rect 15473 20955 15531 20961
rect 15562 20952 15568 20964
rect 15620 20952 15626 21004
rect 16960 20992 16988 21023
rect 19610 21020 19616 21032
rect 19668 21020 19674 21072
rect 17218 20992 17224 21004
rect 16960 20964 17224 20992
rect 17218 20952 17224 20964
rect 17276 20952 17282 21004
rect 18046 20992 18052 21004
rect 18007 20964 18052 20992
rect 18046 20952 18052 20964
rect 18104 20952 18110 21004
rect 18874 20992 18880 21004
rect 18248 20964 18880 20992
rect 8757 20927 8815 20933
rect 8757 20924 8769 20927
rect 7432 20896 8769 20924
rect 7432 20884 7438 20896
rect 8757 20893 8769 20896
rect 8803 20893 8815 20927
rect 8757 20887 8815 20893
rect 8941 20927 8999 20933
rect 8941 20893 8953 20927
rect 8987 20893 8999 20927
rect 8941 20887 8999 20893
rect 7300 20828 7420 20856
rect 5534 20788 5540 20800
rect 4540 20760 5540 20788
rect 5534 20748 5540 20760
rect 5592 20748 5598 20800
rect 6454 20748 6460 20800
rect 6512 20788 6518 20800
rect 6549 20791 6607 20797
rect 6549 20788 6561 20791
rect 6512 20760 6561 20788
rect 6512 20748 6518 20760
rect 6549 20757 6561 20760
rect 6595 20757 6607 20791
rect 6549 20751 6607 20757
rect 6641 20791 6699 20797
rect 6641 20757 6653 20791
rect 6687 20788 6699 20791
rect 7098 20788 7104 20800
rect 6687 20760 7104 20788
rect 6687 20757 6699 20760
rect 6641 20751 6699 20757
rect 7098 20748 7104 20760
rect 7156 20748 7162 20800
rect 7392 20797 7420 20828
rect 7650 20816 7656 20868
rect 7708 20856 7714 20868
rect 8110 20856 8116 20868
rect 7708 20828 8116 20856
rect 7708 20816 7714 20828
rect 8110 20816 8116 20828
rect 8168 20816 8174 20868
rect 8386 20816 8392 20868
rect 8444 20856 8450 20868
rect 8490 20859 8548 20865
rect 8490 20856 8502 20859
rect 8444 20828 8502 20856
rect 8444 20816 8450 20828
rect 8490 20825 8502 20828
rect 8536 20825 8548 20859
rect 8490 20819 8548 20825
rect 7377 20791 7435 20797
rect 7377 20757 7389 20791
rect 7423 20788 7435 20791
rect 7466 20788 7472 20800
rect 7423 20760 7472 20788
rect 7423 20757 7435 20760
rect 7377 20751 7435 20757
rect 7466 20748 7472 20760
rect 7524 20748 7530 20800
rect 8772 20788 8800 20887
rect 9306 20884 9312 20936
rect 9364 20924 9370 20936
rect 11793 20927 11851 20933
rect 9364 20896 10456 20924
rect 9364 20884 9370 20896
rect 9490 20816 9496 20868
rect 9548 20856 9554 20868
rect 9677 20859 9735 20865
rect 9677 20856 9689 20859
rect 9548 20828 9689 20856
rect 9548 20816 9554 20828
rect 9677 20825 9689 20828
rect 9723 20825 9735 20859
rect 9677 20819 9735 20825
rect 9766 20816 9772 20868
rect 9824 20856 9830 20868
rect 10290 20859 10348 20865
rect 10290 20856 10302 20859
rect 9824 20828 10302 20856
rect 9824 20816 9830 20828
rect 10290 20825 10302 20828
rect 10336 20825 10348 20859
rect 10428 20856 10456 20896
rect 11793 20893 11805 20927
rect 11839 20924 11851 20927
rect 12066 20924 12072 20936
rect 11839 20896 12072 20924
rect 11839 20893 11851 20896
rect 11793 20887 11851 20893
rect 12066 20884 12072 20896
rect 12124 20884 12130 20936
rect 12796 20927 12854 20933
rect 12796 20893 12808 20927
rect 12842 20924 12854 20927
rect 14734 20924 14740 20936
rect 12842 20896 14740 20924
rect 12842 20893 12854 20896
rect 12796 20887 12854 20893
rect 14734 20884 14740 20896
rect 14792 20884 14798 20936
rect 15378 20884 15384 20936
rect 15436 20924 15442 20936
rect 15838 20933 15844 20936
rect 15436 20896 15792 20924
rect 15436 20884 15442 20896
rect 15228 20859 15286 20865
rect 10428 20828 14412 20856
rect 10290 20819 10348 20825
rect 9398 20788 9404 20800
rect 8772 20760 9404 20788
rect 9398 20748 9404 20760
rect 9456 20748 9462 20800
rect 12437 20791 12495 20797
rect 12437 20757 12449 20791
rect 12483 20788 12495 20791
rect 12618 20788 12624 20800
rect 12483 20760 12624 20788
rect 12483 20757 12495 20760
rect 12437 20751 12495 20757
rect 12618 20748 12624 20760
rect 12676 20748 12682 20800
rect 13906 20788 13912 20800
rect 13867 20760 13912 20788
rect 13906 20748 13912 20760
rect 13964 20748 13970 20800
rect 14384 20788 14412 20828
rect 15228 20825 15240 20859
rect 15274 20856 15286 20859
rect 15654 20856 15660 20868
rect 15274 20828 15660 20856
rect 15274 20825 15286 20828
rect 15228 20819 15286 20825
rect 15654 20816 15660 20828
rect 15712 20816 15718 20868
rect 15764 20856 15792 20896
rect 15832 20887 15844 20933
rect 15896 20924 15902 20936
rect 18248 20933 18276 20964
rect 18874 20952 18880 20964
rect 18932 20952 18938 21004
rect 18233 20927 18291 20933
rect 15896 20896 15932 20924
rect 15838 20884 15844 20887
rect 15896 20884 15902 20896
rect 18233 20893 18245 20927
rect 18279 20893 18291 20927
rect 18233 20887 18291 20893
rect 18414 20884 18420 20936
rect 18472 20924 18478 20936
rect 18785 20927 18843 20933
rect 18785 20924 18797 20927
rect 18472 20896 18797 20924
rect 18472 20884 18478 20896
rect 18785 20893 18797 20896
rect 18831 20893 18843 20927
rect 19886 20924 19892 20936
rect 19847 20896 19892 20924
rect 18785 20887 18843 20893
rect 19886 20884 19892 20896
rect 19944 20884 19950 20936
rect 19978 20884 19984 20936
rect 20036 20924 20042 20936
rect 20990 20924 20996 20936
rect 20036 20896 20996 20924
rect 20036 20884 20042 20896
rect 20990 20884 20996 20896
rect 21048 20924 21054 20936
rect 21453 20927 21511 20933
rect 21453 20924 21465 20927
rect 21048 20896 21465 20924
rect 21048 20884 21054 20896
rect 21453 20893 21465 20896
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 20226 20859 20284 20865
rect 20226 20856 20238 20859
rect 15764 20828 20238 20856
rect 20226 20825 20238 20828
rect 20272 20825 20284 20859
rect 20226 20819 20284 20825
rect 20714 20816 20720 20868
rect 20772 20856 20778 20868
rect 21698 20859 21756 20865
rect 21698 20856 21710 20859
rect 20772 20828 21710 20856
rect 20772 20816 20778 20828
rect 21698 20825 21710 20828
rect 21744 20825 21756 20859
rect 21698 20819 21756 20825
rect 21910 20816 21916 20868
rect 21968 20856 21974 20868
rect 22925 20859 22983 20865
rect 22925 20856 22937 20859
rect 21968 20828 22937 20856
rect 21968 20816 21974 20828
rect 22925 20825 22937 20828
rect 22971 20825 22983 20859
rect 22925 20819 22983 20825
rect 16390 20788 16396 20800
rect 14384 20760 16396 20788
rect 16390 20748 16396 20760
rect 16448 20748 16454 20800
rect 17310 20788 17316 20800
rect 17271 20760 17316 20788
rect 17310 20748 17316 20760
rect 17368 20748 17374 20800
rect 17402 20748 17408 20800
rect 17460 20788 17466 20800
rect 17773 20791 17831 20797
rect 17460 20760 17505 20788
rect 17460 20748 17466 20760
rect 17773 20757 17785 20791
rect 17819 20788 17831 20791
rect 18141 20791 18199 20797
rect 18141 20788 18153 20791
rect 17819 20760 18153 20788
rect 17819 20757 17831 20760
rect 17773 20751 17831 20757
rect 18141 20757 18153 20760
rect 18187 20757 18199 20791
rect 18598 20788 18604 20800
rect 18559 20760 18604 20788
rect 18141 20751 18199 20757
rect 18598 20748 18604 20760
rect 18656 20748 18662 20800
rect 19245 20791 19303 20797
rect 19245 20757 19257 20791
rect 19291 20788 19303 20791
rect 20806 20788 20812 20800
rect 19291 20760 20812 20788
rect 19291 20757 19303 20760
rect 19245 20751 19303 20757
rect 20806 20748 20812 20760
rect 20864 20748 20870 20800
rect 21450 20748 21456 20800
rect 21508 20788 21514 20800
rect 22833 20791 22891 20797
rect 22833 20788 22845 20791
rect 21508 20760 22845 20788
rect 21508 20748 21514 20760
rect 22833 20757 22845 20760
rect 22879 20757 22891 20791
rect 22833 20751 22891 20757
rect 1104 20698 23460 20720
rect 1104 20646 6548 20698
rect 6600 20646 6612 20698
rect 6664 20646 6676 20698
rect 6728 20646 6740 20698
rect 6792 20646 6804 20698
rect 6856 20646 12146 20698
rect 12198 20646 12210 20698
rect 12262 20646 12274 20698
rect 12326 20646 12338 20698
rect 12390 20646 12402 20698
rect 12454 20646 17744 20698
rect 17796 20646 17808 20698
rect 17860 20646 17872 20698
rect 17924 20646 17936 20698
rect 17988 20646 18000 20698
rect 18052 20646 23460 20698
rect 1104 20624 23460 20646
rect 1762 20584 1768 20596
rect 1723 20556 1768 20584
rect 1762 20544 1768 20556
rect 1820 20544 1826 20596
rect 2222 20544 2228 20596
rect 2280 20584 2286 20596
rect 2280 20556 3188 20584
rect 2280 20544 2286 20556
rect 2130 20476 2136 20528
rect 2188 20516 2194 20528
rect 3160 20516 3188 20556
rect 3234 20544 3240 20596
rect 3292 20584 3298 20596
rect 3697 20587 3755 20593
rect 3697 20584 3709 20587
rect 3292 20556 3709 20584
rect 3292 20544 3298 20556
rect 3697 20553 3709 20556
rect 3743 20553 3755 20587
rect 3697 20547 3755 20553
rect 4062 20544 4068 20596
rect 4120 20584 4126 20596
rect 4120 20556 4844 20584
rect 4120 20544 4126 20556
rect 3418 20516 3424 20528
rect 2188 20488 3096 20516
rect 2188 20476 2194 20488
rect 1489 20451 1547 20457
rect 1489 20417 1501 20451
rect 1535 20448 1547 20451
rect 2590 20448 2596 20460
rect 1535 20420 2596 20448
rect 1535 20417 1547 20420
rect 1489 20411 1547 20417
rect 2590 20408 2596 20420
rect 2648 20408 2654 20460
rect 2866 20448 2872 20460
rect 2924 20457 2930 20460
rect 2836 20420 2872 20448
rect 2866 20408 2872 20420
rect 2924 20411 2936 20457
rect 2924 20408 2930 20411
rect 3068 20380 3096 20488
rect 3160 20488 3424 20516
rect 3160 20457 3188 20488
rect 3418 20476 3424 20488
rect 3476 20516 3482 20528
rect 4080 20516 4108 20544
rect 4706 20516 4712 20528
rect 3476 20488 4108 20516
rect 4667 20488 4712 20516
rect 3476 20476 3482 20488
rect 4706 20476 4712 20488
rect 4764 20476 4770 20528
rect 4816 20516 4844 20556
rect 5902 20544 5908 20596
rect 5960 20584 5966 20596
rect 6181 20587 6239 20593
rect 6181 20584 6193 20587
rect 5960 20556 6193 20584
rect 5960 20544 5966 20556
rect 6181 20553 6193 20556
rect 6227 20553 6239 20587
rect 7742 20584 7748 20596
rect 7703 20556 7748 20584
rect 6181 20547 6239 20553
rect 7742 20544 7748 20556
rect 7800 20544 7806 20596
rect 8205 20587 8263 20593
rect 8205 20553 8217 20587
rect 8251 20584 8263 20587
rect 8757 20587 8815 20593
rect 8251 20556 8708 20584
rect 8251 20553 8263 20556
rect 8205 20547 8263 20553
rect 4816 20488 6408 20516
rect 3145 20451 3203 20457
rect 3145 20417 3157 20451
rect 3191 20417 3203 20451
rect 3145 20411 3203 20417
rect 3605 20451 3663 20457
rect 3605 20417 3617 20451
rect 3651 20417 3663 20451
rect 3605 20411 3663 20417
rect 3620 20380 3648 20411
rect 3694 20408 3700 20460
rect 3752 20448 3758 20460
rect 4816 20457 4844 20488
rect 5074 20457 5080 20460
rect 4065 20451 4123 20457
rect 4065 20448 4077 20451
rect 3752 20420 4077 20448
rect 3752 20408 3758 20420
rect 4065 20417 4077 20420
rect 4111 20417 4123 20451
rect 4065 20411 4123 20417
rect 4801 20451 4859 20457
rect 4801 20417 4813 20451
rect 4847 20417 4859 20451
rect 5068 20448 5080 20457
rect 5035 20420 5080 20448
rect 4801 20411 4859 20417
rect 5068 20411 5080 20420
rect 5074 20408 5080 20411
rect 5132 20408 5138 20460
rect 6380 20457 6408 20488
rect 6454 20476 6460 20528
rect 6512 20516 6518 20528
rect 6610 20519 6668 20525
rect 6610 20516 6622 20519
rect 6512 20488 6622 20516
rect 6512 20476 6518 20488
rect 6610 20485 6622 20488
rect 6656 20485 6668 20519
rect 6610 20479 6668 20485
rect 8018 20476 8024 20528
rect 8076 20516 8082 20528
rect 8570 20516 8576 20528
rect 8076 20488 8576 20516
rect 8076 20476 8082 20488
rect 8570 20476 8576 20488
rect 8628 20476 8634 20528
rect 8680 20516 8708 20556
rect 8757 20553 8769 20587
rect 8803 20584 8815 20587
rect 8846 20584 8852 20596
rect 8803 20556 8852 20584
rect 8803 20553 8815 20556
rect 8757 20547 8815 20553
rect 8846 20544 8852 20556
rect 8904 20544 8910 20596
rect 9490 20584 9496 20596
rect 8956 20556 9496 20584
rect 8956 20516 8984 20556
rect 9490 20544 9496 20556
rect 9548 20544 9554 20596
rect 11885 20587 11943 20593
rect 11885 20553 11897 20587
rect 11931 20553 11943 20587
rect 11885 20547 11943 20553
rect 13541 20587 13599 20593
rect 13541 20553 13553 20587
rect 13587 20584 13599 20587
rect 13630 20584 13636 20596
rect 13587 20556 13636 20584
rect 13587 20553 13599 20556
rect 13541 20547 13599 20553
rect 8680 20488 8984 20516
rect 9217 20519 9275 20525
rect 9217 20485 9229 20519
rect 9263 20516 9275 20519
rect 11149 20519 11207 20525
rect 11149 20516 11161 20519
rect 9263 20488 11161 20516
rect 9263 20485 9275 20488
rect 9217 20479 9275 20485
rect 11149 20485 11161 20488
rect 11195 20485 11207 20519
rect 11149 20479 11207 20485
rect 6365 20451 6423 20457
rect 6365 20417 6377 20451
rect 6411 20417 6423 20451
rect 6365 20411 6423 20417
rect 7466 20408 7472 20460
rect 7524 20448 7530 20460
rect 9674 20448 9680 20460
rect 7524 20420 8432 20448
rect 9635 20420 9680 20448
rect 7524 20408 7530 20420
rect 3068 20352 3648 20380
rect 3881 20383 3939 20389
rect 3881 20349 3893 20383
rect 3927 20380 3939 20383
rect 4430 20380 4436 20392
rect 3927 20352 4436 20380
rect 3927 20349 3939 20352
rect 3881 20343 3939 20349
rect 4430 20340 4436 20352
rect 4488 20380 4494 20392
rect 4706 20380 4712 20392
rect 4488 20352 4712 20380
rect 4488 20340 4494 20352
rect 4706 20340 4712 20352
rect 4764 20340 4770 20392
rect 8018 20340 8024 20392
rect 8076 20380 8082 20392
rect 8404 20389 8432 20420
rect 9674 20408 9680 20420
rect 9732 20408 9738 20460
rect 9950 20457 9956 20460
rect 9944 20448 9956 20457
rect 9911 20420 9956 20448
rect 9944 20411 9956 20420
rect 9950 20408 9956 20411
rect 10008 20408 10014 20460
rect 11701 20451 11759 20457
rect 11701 20417 11713 20451
rect 11747 20448 11759 20451
rect 11900 20448 11928 20547
rect 13630 20544 13636 20556
rect 13688 20544 13694 20596
rect 14001 20587 14059 20593
rect 14001 20553 14013 20587
rect 14047 20584 14059 20587
rect 14553 20587 14611 20593
rect 14553 20584 14565 20587
rect 14047 20556 14565 20584
rect 14047 20553 14059 20556
rect 14001 20547 14059 20553
rect 14553 20553 14565 20556
rect 14599 20553 14611 20587
rect 14553 20547 14611 20553
rect 14921 20587 14979 20593
rect 14921 20553 14933 20587
rect 14967 20553 14979 20587
rect 15654 20584 15660 20596
rect 15615 20556 15660 20584
rect 14921 20547 14979 20553
rect 12526 20516 12532 20528
rect 12176 20488 12532 20516
rect 11747 20420 11928 20448
rect 11747 20417 11759 20420
rect 11701 20411 11759 20417
rect 11974 20408 11980 20460
rect 12032 20448 12038 20460
rect 12176 20457 12204 20488
rect 12526 20476 12532 20488
rect 12584 20516 12590 20528
rect 13446 20516 13452 20528
rect 12584 20488 13452 20516
rect 12584 20476 12590 20488
rect 13446 20476 13452 20488
rect 13504 20476 13510 20528
rect 14936 20516 14964 20547
rect 15654 20544 15660 20556
rect 15712 20544 15718 20596
rect 18598 20544 18604 20596
rect 18656 20584 18662 20596
rect 19337 20587 19395 20593
rect 19337 20584 19349 20587
rect 18656 20556 19349 20584
rect 18656 20544 18662 20556
rect 19337 20553 19349 20556
rect 19383 20553 19395 20587
rect 19702 20584 19708 20596
rect 19663 20556 19708 20584
rect 19337 20547 19395 20553
rect 19702 20544 19708 20556
rect 19760 20544 19766 20596
rect 19981 20587 20039 20593
rect 19981 20553 19993 20587
rect 20027 20584 20039 20587
rect 20027 20556 21036 20584
rect 20027 20553 20039 20556
rect 19981 20547 20039 20553
rect 14936 20488 15700 20516
rect 12069 20451 12127 20457
rect 12069 20448 12081 20451
rect 12032 20420 12081 20448
rect 12032 20408 12038 20420
rect 12069 20417 12081 20420
rect 12115 20417 12127 20451
rect 12069 20411 12127 20417
rect 12161 20451 12219 20457
rect 12161 20417 12173 20451
rect 12207 20417 12219 20451
rect 12161 20411 12219 20417
rect 12428 20451 12486 20457
rect 12428 20417 12440 20451
rect 12474 20448 12486 20451
rect 12710 20448 12716 20460
rect 12474 20420 12716 20448
rect 12474 20417 12486 20420
rect 12428 20411 12486 20417
rect 8297 20383 8355 20389
rect 8297 20380 8309 20383
rect 8076 20352 8309 20380
rect 8076 20340 8082 20352
rect 8297 20349 8309 20352
rect 8343 20349 8355 20383
rect 8297 20343 8355 20349
rect 8389 20383 8447 20389
rect 8389 20349 8401 20383
rect 8435 20349 8447 20383
rect 8389 20343 8447 20349
rect 9309 20383 9367 20389
rect 9309 20349 9321 20383
rect 9355 20349 9367 20383
rect 9309 20343 9367 20349
rect 9493 20383 9551 20389
rect 9493 20349 9505 20383
rect 9539 20349 9551 20383
rect 9493 20343 9551 20349
rect 7558 20272 7564 20324
rect 7616 20312 7622 20324
rect 8478 20312 8484 20324
rect 7616 20284 8484 20312
rect 7616 20272 7622 20284
rect 8478 20272 8484 20284
rect 8536 20272 8542 20324
rect 1673 20247 1731 20253
rect 1673 20213 1685 20247
rect 1719 20244 1731 20247
rect 3142 20244 3148 20256
rect 1719 20216 3148 20244
rect 1719 20213 1731 20216
rect 1673 20207 1731 20213
rect 3142 20204 3148 20216
rect 3200 20204 3206 20256
rect 3234 20204 3240 20256
rect 3292 20244 3298 20256
rect 3292 20216 3337 20244
rect 3292 20204 3298 20216
rect 4154 20204 4160 20256
rect 4212 20244 4218 20256
rect 4982 20244 4988 20256
rect 4212 20216 4988 20244
rect 4212 20204 4218 20216
rect 4982 20204 4988 20216
rect 5040 20244 5046 20256
rect 5994 20244 6000 20256
rect 5040 20216 6000 20244
rect 5040 20204 5046 20216
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 7834 20244 7840 20256
rect 7795 20216 7840 20244
rect 7834 20204 7840 20216
rect 7892 20204 7898 20256
rect 8294 20204 8300 20256
rect 8352 20244 8358 20256
rect 8849 20247 8907 20253
rect 8849 20244 8861 20247
rect 8352 20216 8861 20244
rect 8352 20204 8358 20216
rect 8849 20213 8861 20216
rect 8895 20244 8907 20247
rect 9214 20244 9220 20256
rect 8895 20216 9220 20244
rect 8895 20213 8907 20216
rect 8849 20207 8907 20213
rect 9214 20204 9220 20216
rect 9272 20204 9278 20256
rect 9324 20244 9352 20343
rect 9508 20312 9536 20343
rect 9674 20312 9680 20324
rect 9508 20284 9680 20312
rect 9674 20272 9680 20284
rect 9732 20272 9738 20324
rect 11146 20272 11152 20324
rect 11204 20312 11210 20324
rect 11517 20315 11575 20321
rect 11517 20312 11529 20315
rect 11204 20284 11529 20312
rect 11204 20272 11210 20284
rect 11517 20281 11529 20284
rect 11563 20281 11575 20315
rect 11517 20275 11575 20281
rect 10318 20244 10324 20256
rect 9324 20216 10324 20244
rect 10318 20204 10324 20216
rect 10376 20204 10382 20256
rect 11057 20247 11115 20253
rect 11057 20213 11069 20247
rect 11103 20244 11115 20247
rect 11238 20244 11244 20256
rect 11103 20216 11244 20244
rect 11103 20213 11115 20216
rect 11057 20207 11115 20213
rect 11238 20204 11244 20216
rect 11296 20204 11302 20256
rect 12084 20244 12112 20411
rect 12710 20408 12716 20420
rect 12768 20408 12774 20460
rect 13814 20448 13820 20460
rect 13775 20420 13820 20448
rect 13814 20408 13820 20420
rect 13872 20408 13878 20460
rect 13906 20408 13912 20460
rect 13964 20448 13970 20460
rect 14550 20448 14556 20460
rect 13964 20420 14556 20448
rect 13964 20408 13970 20420
rect 14550 20408 14556 20420
rect 14608 20448 14614 20460
rect 15013 20451 15071 20457
rect 15013 20448 15025 20451
rect 14608 20420 15025 20448
rect 14608 20408 14614 20420
rect 15013 20417 15025 20420
rect 15059 20417 15071 20451
rect 15672 20448 15700 20488
rect 15746 20476 15752 20528
rect 15804 20516 15810 20528
rect 16298 20516 16304 20528
rect 15804 20488 16304 20516
rect 15804 20476 15810 20488
rect 16298 20476 16304 20488
rect 16356 20516 16362 20528
rect 16853 20519 16911 20525
rect 16853 20516 16865 20519
rect 16356 20488 16865 20516
rect 16356 20476 16362 20488
rect 16853 20485 16865 20488
rect 16899 20485 16911 20519
rect 16853 20479 16911 20485
rect 17037 20519 17095 20525
rect 17037 20485 17049 20519
rect 17083 20516 17095 20519
rect 17954 20516 17960 20528
rect 17083 20488 17960 20516
rect 17083 20485 17095 20488
rect 17037 20479 17095 20485
rect 17954 20476 17960 20488
rect 18012 20476 18018 20528
rect 18233 20519 18291 20525
rect 18233 20485 18245 20519
rect 18279 20516 18291 20519
rect 18279 20488 19932 20516
rect 18279 20485 18291 20488
rect 18233 20479 18291 20485
rect 16117 20451 16175 20457
rect 16117 20448 16129 20451
rect 15672 20420 16129 20448
rect 15013 20411 15071 20417
rect 16117 20417 16129 20420
rect 16163 20448 16175 20451
rect 16942 20448 16948 20460
rect 16163 20420 16948 20448
rect 16163 20417 16175 20420
rect 16117 20411 16175 20417
rect 16942 20408 16948 20420
rect 17000 20408 17006 20460
rect 17218 20448 17224 20460
rect 17179 20420 17224 20448
rect 17218 20408 17224 20420
rect 17276 20408 17282 20460
rect 18877 20451 18935 20457
rect 18877 20417 18889 20451
rect 18923 20448 18935 20451
rect 18923 20420 19196 20448
rect 18923 20417 18935 20420
rect 18877 20411 18935 20417
rect 14369 20383 14427 20389
rect 14369 20349 14381 20383
rect 14415 20349 14427 20383
rect 14369 20343 14427 20349
rect 14461 20383 14519 20389
rect 14461 20349 14473 20383
rect 14507 20380 14519 20383
rect 14734 20380 14740 20392
rect 14507 20352 14740 20380
rect 14507 20349 14519 20352
rect 14461 20343 14519 20349
rect 13633 20315 13691 20321
rect 13633 20312 13645 20315
rect 13096 20284 13645 20312
rect 13096 20244 13124 20284
rect 13633 20281 13645 20284
rect 13679 20281 13691 20315
rect 13633 20275 13691 20281
rect 12084 20216 13124 20244
rect 14274 20204 14280 20256
rect 14332 20244 14338 20256
rect 14384 20244 14412 20343
rect 14734 20340 14740 20352
rect 14792 20340 14798 20392
rect 15930 20380 15936 20392
rect 15891 20352 15936 20380
rect 15930 20340 15936 20352
rect 15988 20340 15994 20392
rect 16025 20383 16083 20389
rect 16025 20349 16037 20383
rect 16071 20380 16083 20383
rect 17126 20380 17132 20392
rect 16071 20352 17132 20380
rect 16071 20349 16083 20352
rect 16025 20343 16083 20349
rect 17126 20340 17132 20352
rect 17184 20340 17190 20392
rect 17497 20383 17555 20389
rect 17497 20349 17509 20383
rect 17543 20349 17555 20383
rect 17497 20343 17555 20349
rect 15286 20272 15292 20324
rect 15344 20312 15350 20324
rect 17512 20312 17540 20343
rect 17678 20340 17684 20392
rect 17736 20380 17742 20392
rect 19058 20380 19064 20392
rect 17736 20352 19064 20380
rect 17736 20340 17742 20352
rect 19058 20340 19064 20352
rect 19116 20340 19122 20392
rect 19168 20389 19196 20420
rect 19610 20408 19616 20460
rect 19668 20448 19674 20460
rect 19797 20451 19855 20457
rect 19797 20448 19809 20451
rect 19668 20420 19809 20448
rect 19668 20408 19674 20420
rect 19797 20417 19809 20420
rect 19843 20417 19855 20451
rect 19904 20448 19932 20488
rect 20346 20476 20352 20528
rect 20404 20516 20410 20528
rect 20502 20519 20560 20525
rect 20502 20516 20514 20519
rect 20404 20488 20514 20516
rect 20404 20476 20410 20488
rect 20502 20485 20514 20488
rect 20548 20485 20560 20519
rect 21008 20516 21036 20556
rect 21174 20544 21180 20596
rect 21232 20584 21238 20596
rect 22833 20587 22891 20593
rect 22833 20584 22845 20587
rect 21232 20556 22845 20584
rect 21232 20544 21238 20556
rect 22833 20553 22845 20556
rect 22879 20553 22891 20587
rect 22833 20547 22891 20553
rect 23382 20516 23388 20528
rect 21008 20488 23388 20516
rect 20502 20479 20560 20485
rect 23382 20476 23388 20488
rect 23440 20476 23446 20528
rect 20898 20448 20904 20460
rect 19904 20420 20904 20448
rect 19797 20411 19855 20417
rect 20898 20408 20904 20420
rect 20956 20408 20962 20460
rect 20990 20408 20996 20460
rect 21048 20448 21054 20460
rect 21048 20420 21588 20448
rect 21048 20408 21054 20420
rect 19153 20383 19211 20389
rect 19153 20349 19165 20383
rect 19199 20349 19211 20383
rect 19153 20343 19211 20349
rect 15344 20284 17540 20312
rect 19168 20312 19196 20343
rect 19242 20340 19248 20392
rect 19300 20380 19306 20392
rect 19300 20352 19345 20380
rect 19300 20340 19306 20352
rect 19978 20340 19984 20392
rect 20036 20380 20042 20392
rect 20257 20383 20315 20389
rect 20257 20380 20269 20383
rect 20036 20352 20269 20380
rect 20036 20340 20042 20352
rect 20257 20349 20269 20352
rect 20303 20349 20315 20383
rect 21560 20380 21588 20420
rect 21634 20408 21640 20460
rect 21692 20448 21698 20460
rect 22189 20451 22247 20457
rect 21692 20420 21956 20448
rect 21692 20408 21698 20420
rect 21928 20389 21956 20420
rect 22189 20417 22201 20451
rect 22235 20448 22247 20451
rect 22649 20451 22707 20457
rect 22235 20420 22324 20448
rect 22235 20417 22247 20420
rect 22189 20411 22247 20417
rect 21913 20383 21971 20389
rect 21560 20352 21772 20380
rect 20257 20343 20315 20349
rect 19518 20312 19524 20324
rect 19168 20284 19524 20312
rect 15344 20272 15350 20284
rect 19518 20272 19524 20284
rect 19576 20272 19582 20324
rect 16298 20244 16304 20256
rect 14332 20216 16304 20244
rect 14332 20204 14338 20216
rect 16298 20204 16304 20216
rect 16356 20204 16362 20256
rect 16482 20244 16488 20256
rect 16443 20216 16488 20244
rect 16482 20204 16488 20216
rect 16540 20204 16546 20256
rect 16669 20247 16727 20253
rect 16669 20213 16681 20247
rect 16715 20244 16727 20247
rect 19058 20244 19064 20256
rect 16715 20216 19064 20244
rect 16715 20213 16727 20216
rect 16669 20207 16727 20213
rect 19058 20204 19064 20216
rect 19116 20204 19122 20256
rect 20272 20244 20300 20343
rect 21634 20312 21640 20324
rect 21595 20284 21640 20312
rect 21634 20272 21640 20284
rect 21692 20272 21698 20324
rect 21744 20312 21772 20352
rect 21913 20349 21925 20383
rect 21959 20349 21971 20383
rect 21913 20343 21971 20349
rect 22094 20340 22100 20392
rect 22152 20380 22158 20392
rect 22152 20352 22197 20380
rect 22152 20340 22158 20352
rect 22296 20312 22324 20420
rect 22649 20417 22661 20451
rect 22695 20448 22707 20451
rect 23014 20448 23020 20460
rect 22695 20420 23020 20448
rect 22695 20417 22707 20420
rect 22649 20411 22707 20417
rect 23014 20408 23020 20420
rect 23072 20448 23078 20460
rect 23290 20448 23296 20460
rect 23072 20420 23296 20448
rect 23072 20408 23078 20420
rect 23290 20408 23296 20420
rect 23348 20408 23354 20460
rect 21744 20284 22324 20312
rect 21174 20244 21180 20256
rect 20272 20216 21180 20244
rect 21174 20204 21180 20216
rect 21232 20204 21238 20256
rect 21266 20204 21272 20256
rect 21324 20244 21330 20256
rect 22002 20244 22008 20256
rect 21324 20216 22008 20244
rect 21324 20204 21330 20216
rect 22002 20204 22008 20216
rect 22060 20204 22066 20256
rect 22278 20204 22284 20256
rect 22336 20244 22342 20256
rect 22557 20247 22615 20253
rect 22557 20244 22569 20247
rect 22336 20216 22569 20244
rect 22336 20204 22342 20216
rect 22557 20213 22569 20216
rect 22603 20213 22615 20247
rect 23014 20244 23020 20256
rect 22975 20216 23020 20244
rect 22557 20207 22615 20213
rect 23014 20204 23020 20216
rect 23072 20204 23078 20256
rect 1104 20154 23460 20176
rect 1104 20102 3749 20154
rect 3801 20102 3813 20154
rect 3865 20102 3877 20154
rect 3929 20102 3941 20154
rect 3993 20102 4005 20154
rect 4057 20102 9347 20154
rect 9399 20102 9411 20154
rect 9463 20102 9475 20154
rect 9527 20102 9539 20154
rect 9591 20102 9603 20154
rect 9655 20102 14945 20154
rect 14997 20102 15009 20154
rect 15061 20102 15073 20154
rect 15125 20102 15137 20154
rect 15189 20102 15201 20154
rect 15253 20102 20543 20154
rect 20595 20102 20607 20154
rect 20659 20102 20671 20154
rect 20723 20102 20735 20154
rect 20787 20102 20799 20154
rect 20851 20102 23460 20154
rect 1104 20080 23460 20102
rect 2866 20000 2872 20052
rect 2924 20040 2930 20052
rect 4433 20043 4491 20049
rect 4433 20040 4445 20043
rect 2924 20012 4445 20040
rect 2924 20000 2930 20012
rect 4433 20009 4445 20012
rect 4479 20009 4491 20043
rect 4433 20003 4491 20009
rect 4614 20000 4620 20052
rect 4672 20040 4678 20052
rect 7006 20040 7012 20052
rect 4672 20012 7012 20040
rect 4672 20000 4678 20012
rect 7006 20000 7012 20012
rect 7064 20000 7070 20052
rect 7190 20040 7196 20052
rect 7151 20012 7196 20040
rect 7190 20000 7196 20012
rect 7248 20000 7254 20052
rect 8018 20040 8024 20052
rect 7979 20012 8024 20040
rect 8018 20000 8024 20012
rect 8076 20000 8082 20052
rect 9766 20040 9772 20052
rect 9727 20012 9772 20040
rect 9766 20000 9772 20012
rect 9824 20000 9830 20052
rect 11054 20000 11060 20052
rect 11112 20040 11118 20052
rect 11333 20043 11391 20049
rect 11333 20040 11345 20043
rect 11112 20012 11345 20040
rect 11112 20000 11118 20012
rect 11333 20009 11345 20012
rect 11379 20009 11391 20043
rect 11333 20003 11391 20009
rect 13538 20000 13544 20052
rect 13596 20040 13602 20052
rect 13725 20043 13783 20049
rect 13725 20040 13737 20043
rect 13596 20012 13737 20040
rect 13596 20000 13602 20012
rect 13725 20009 13737 20012
rect 13771 20009 13783 20043
rect 14090 20040 14096 20052
rect 14051 20012 14096 20040
rect 13725 20003 13783 20009
rect 14090 20000 14096 20012
rect 14148 20000 14154 20052
rect 14826 20000 14832 20052
rect 14884 20040 14890 20052
rect 14921 20043 14979 20049
rect 14921 20040 14933 20043
rect 14884 20012 14933 20040
rect 14884 20000 14890 20012
rect 14921 20009 14933 20012
rect 14967 20009 14979 20043
rect 19150 20040 19156 20052
rect 14921 20003 14979 20009
rect 15580 20012 19156 20040
rect 2590 19932 2596 19984
rect 2648 19972 2654 19984
rect 4890 19972 4896 19984
rect 2648 19944 4896 19972
rect 2648 19932 2654 19944
rect 4890 19932 4896 19944
rect 4948 19932 4954 19984
rect 5074 19972 5080 19984
rect 5035 19944 5080 19972
rect 5074 19932 5080 19944
rect 5132 19932 5138 19984
rect 5534 19932 5540 19984
rect 5592 19972 5598 19984
rect 6733 19975 6791 19981
rect 5592 19944 6224 19972
rect 5592 19932 5598 19944
rect 3142 19864 3148 19916
rect 3200 19904 3206 19916
rect 5258 19904 5264 19916
rect 3200 19876 5028 19904
rect 5219 19876 5264 19904
rect 3200 19864 3206 19876
rect 1489 19839 1547 19845
rect 1489 19805 1501 19839
rect 1535 19836 1547 19839
rect 1578 19836 1584 19848
rect 1535 19808 1584 19836
rect 1535 19805 1547 19808
rect 1489 19799 1547 19805
rect 1578 19796 1584 19808
rect 1636 19836 1642 19848
rect 2222 19836 2228 19848
rect 1636 19808 2228 19836
rect 1636 19796 1642 19808
rect 2222 19796 2228 19808
rect 2280 19796 2286 19848
rect 2774 19796 2780 19848
rect 2832 19836 2838 19848
rect 3605 19839 3663 19845
rect 3605 19836 3617 19839
rect 2832 19808 3617 19836
rect 2832 19796 2838 19808
rect 3605 19805 3617 19808
rect 3651 19805 3663 19839
rect 3605 19799 3663 19805
rect 3789 19839 3847 19845
rect 3789 19805 3801 19839
rect 3835 19805 3847 19839
rect 4614 19836 4620 19848
rect 4575 19808 4620 19836
rect 3789 19799 3847 19805
rect 1756 19771 1814 19777
rect 1756 19737 1768 19771
rect 1802 19768 1814 19771
rect 2961 19771 3019 19777
rect 2961 19768 2973 19771
rect 1802 19740 2973 19768
rect 1802 19737 1814 19740
rect 1756 19731 1814 19737
rect 2961 19737 2973 19740
rect 3007 19737 3019 19771
rect 2961 19731 3019 19737
rect 2866 19700 2872 19712
rect 2827 19672 2872 19700
rect 2866 19660 2872 19672
rect 2924 19700 2930 19712
rect 3804 19700 3832 19799
rect 4614 19796 4620 19808
rect 4672 19796 4678 19848
rect 4798 19796 4804 19848
rect 4856 19836 4862 19848
rect 4893 19839 4951 19845
rect 4893 19836 4905 19839
rect 4856 19808 4905 19836
rect 4856 19796 4862 19808
rect 4893 19805 4905 19808
rect 4939 19805 4951 19839
rect 5000 19836 5028 19876
rect 5258 19864 5264 19876
rect 5316 19864 5322 19916
rect 5902 19864 5908 19916
rect 5960 19904 5966 19916
rect 6089 19907 6147 19913
rect 6089 19904 6101 19907
rect 5960 19876 6101 19904
rect 5960 19864 5966 19876
rect 6089 19873 6101 19876
rect 6135 19873 6147 19907
rect 6196 19904 6224 19944
rect 6733 19941 6745 19975
rect 6779 19972 6791 19975
rect 7558 19972 7564 19984
rect 6779 19944 7564 19972
rect 6779 19941 6791 19944
rect 6733 19935 6791 19941
rect 7558 19932 7564 19944
rect 7616 19932 7622 19984
rect 9674 19932 9680 19984
rect 9732 19972 9738 19984
rect 9861 19975 9919 19981
rect 9861 19972 9873 19975
rect 9732 19944 9873 19972
rect 9732 19932 9738 19944
rect 9861 19941 9873 19944
rect 9907 19941 9919 19975
rect 9861 19935 9919 19941
rect 6825 19907 6883 19913
rect 6825 19904 6837 19907
rect 6196 19876 6837 19904
rect 6089 19867 6147 19873
rect 6825 19873 6837 19876
rect 6871 19873 6883 19907
rect 6825 19867 6883 19873
rect 7190 19864 7196 19916
rect 7248 19904 7254 19916
rect 7742 19904 7748 19916
rect 7248 19876 7651 19904
rect 7703 19876 7748 19904
rect 7248 19864 7254 19876
rect 5445 19839 5503 19845
rect 5445 19836 5457 19839
rect 5000 19832 5304 19836
rect 5368 19832 5457 19836
rect 5000 19808 5457 19832
rect 4893 19799 4951 19805
rect 5276 19804 5396 19808
rect 5445 19805 5457 19808
rect 5491 19805 5503 19839
rect 5445 19799 5503 19805
rect 6178 19796 6184 19848
rect 6236 19836 6242 19848
rect 7282 19836 7288 19848
rect 6236 19808 7288 19836
rect 6236 19796 6242 19808
rect 7282 19796 7288 19808
rect 7340 19796 7346 19848
rect 7623 19836 7651 19876
rect 7742 19864 7748 19876
rect 7800 19864 7806 19916
rect 8662 19904 8668 19916
rect 8623 19876 8668 19904
rect 8662 19864 8668 19876
rect 8720 19864 8726 19916
rect 9214 19904 9220 19916
rect 8772 19876 9220 19904
rect 8772 19836 8800 19876
rect 9214 19864 9220 19876
rect 9272 19864 9278 19916
rect 7623 19808 8800 19836
rect 9125 19839 9183 19845
rect 9125 19805 9137 19839
rect 9171 19836 9183 19839
rect 9876 19836 9904 19935
rect 11514 19932 11520 19984
rect 11572 19972 11578 19984
rect 11572 19944 13952 19972
rect 11572 19932 11578 19944
rect 11241 19907 11299 19913
rect 11241 19873 11253 19907
rect 11287 19904 11299 19907
rect 11330 19904 11336 19916
rect 11287 19876 11336 19904
rect 11287 19873 11299 19876
rect 11241 19867 11299 19873
rect 11330 19864 11336 19876
rect 11388 19864 11394 19916
rect 11882 19904 11888 19916
rect 11843 19876 11888 19904
rect 11882 19864 11888 19876
rect 11940 19864 11946 19916
rect 13078 19904 13084 19916
rect 13039 19876 13084 19904
rect 13078 19864 13084 19876
rect 13136 19864 13142 19916
rect 9171 19808 9904 19836
rect 9171 19805 9183 19808
rect 9125 19799 9183 19805
rect 12066 19796 12072 19848
rect 12124 19796 12130 19848
rect 12802 19836 12808 19848
rect 12763 19808 12808 19836
rect 12802 19796 12808 19808
rect 12860 19796 12866 19848
rect 13357 19839 13415 19845
rect 13357 19805 13369 19839
rect 13403 19836 13415 19839
rect 13630 19836 13636 19848
rect 13403 19808 13636 19836
rect 13403 19805 13415 19808
rect 13357 19799 13415 19805
rect 13630 19796 13636 19808
rect 13688 19796 13694 19848
rect 5074 19728 5080 19780
rect 5132 19768 5138 19780
rect 5537 19771 5595 19777
rect 5537 19768 5549 19771
rect 5132 19740 5549 19768
rect 5132 19728 5138 19740
rect 5537 19737 5549 19740
rect 5583 19737 5595 19771
rect 7009 19771 7067 19777
rect 7009 19768 7021 19771
rect 5537 19731 5595 19737
rect 5828 19740 7021 19768
rect 5828 19712 5856 19740
rect 7009 19737 7021 19740
rect 7055 19737 7067 19771
rect 7653 19771 7711 19777
rect 7653 19768 7665 19771
rect 7009 19731 7067 19737
rect 7392 19740 7665 19768
rect 2924 19672 3832 19700
rect 4801 19703 4859 19709
rect 2924 19660 2930 19672
rect 4801 19669 4813 19703
rect 4847 19700 4859 19703
rect 5810 19700 5816 19712
rect 4847 19672 5816 19700
rect 4847 19669 4859 19672
rect 4801 19663 4859 19669
rect 5810 19660 5816 19672
rect 5868 19660 5874 19712
rect 5905 19703 5963 19709
rect 5905 19669 5917 19703
rect 5951 19700 5963 19703
rect 6273 19703 6331 19709
rect 6273 19700 6285 19703
rect 5951 19672 6285 19700
rect 5951 19669 5963 19672
rect 5905 19663 5963 19669
rect 6273 19669 6285 19672
rect 6319 19669 6331 19703
rect 6273 19663 6331 19669
rect 6362 19660 6368 19712
rect 6420 19700 6426 19712
rect 6420 19672 6465 19700
rect 6420 19660 6426 19672
rect 6914 19660 6920 19712
rect 6972 19700 6978 19712
rect 7392 19700 7420 19740
rect 7653 19737 7665 19740
rect 7699 19768 7711 19771
rect 7926 19768 7932 19780
rect 7699 19740 7932 19768
rect 7699 19737 7711 19740
rect 7653 19731 7711 19737
rect 7926 19728 7932 19740
rect 7984 19728 7990 19780
rect 8481 19771 8539 19777
rect 8481 19737 8493 19771
rect 8527 19768 8539 19771
rect 9766 19768 9772 19780
rect 8527 19740 9772 19768
rect 8527 19737 8539 19740
rect 8481 19731 8539 19737
rect 9766 19728 9772 19740
rect 9824 19728 9830 19780
rect 10134 19728 10140 19780
rect 10192 19768 10198 19780
rect 10974 19771 11032 19777
rect 10974 19768 10986 19771
rect 10192 19740 10986 19768
rect 10192 19728 10198 19740
rect 10974 19737 10986 19740
rect 11020 19737 11032 19771
rect 12084 19768 12112 19796
rect 13265 19771 13323 19777
rect 13265 19768 13277 19771
rect 12084 19740 13277 19768
rect 10974 19731 11032 19737
rect 13265 19737 13277 19740
rect 13311 19737 13323 19771
rect 13265 19731 13323 19737
rect 7558 19700 7564 19712
rect 6972 19672 7420 19700
rect 7519 19672 7564 19700
rect 6972 19660 6978 19672
rect 7558 19660 7564 19672
rect 7616 19660 7622 19712
rect 8386 19700 8392 19712
rect 8347 19672 8392 19700
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 9033 19703 9091 19709
rect 9033 19669 9045 19703
rect 9079 19700 9091 19703
rect 11146 19700 11152 19712
rect 9079 19672 11152 19700
rect 9079 19669 9091 19672
rect 9033 19663 9091 19669
rect 11146 19660 11152 19672
rect 11204 19660 11210 19712
rect 11422 19660 11428 19712
rect 11480 19700 11486 19712
rect 11701 19703 11759 19709
rect 11701 19700 11713 19703
rect 11480 19672 11713 19700
rect 11480 19660 11486 19672
rect 11701 19669 11713 19672
rect 11747 19669 11759 19703
rect 11701 19663 11759 19669
rect 11790 19660 11796 19712
rect 11848 19700 11854 19712
rect 11848 19672 11893 19700
rect 11848 19660 11854 19672
rect 12066 19660 12072 19712
rect 12124 19700 12130 19712
rect 13924 19709 13952 19944
rect 13998 19932 14004 19984
rect 14056 19972 14062 19984
rect 14056 19944 14688 19972
rect 14056 19932 14062 19944
rect 14550 19904 14556 19916
rect 14511 19876 14556 19904
rect 14550 19864 14556 19876
rect 14608 19864 14614 19916
rect 14660 19913 14688 19944
rect 14645 19907 14703 19913
rect 14645 19873 14657 19907
rect 14691 19904 14703 19907
rect 15010 19904 15016 19916
rect 14691 19876 15016 19904
rect 14691 19873 14703 19876
rect 14645 19867 14703 19873
rect 15010 19864 15016 19876
rect 15068 19864 15074 19916
rect 14182 19796 14188 19848
rect 14240 19836 14246 19848
rect 15580 19845 15608 20012
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 21450 20040 21456 20052
rect 19260 20012 21456 20040
rect 18598 19864 18604 19916
rect 18656 19904 18662 19916
rect 18693 19907 18751 19913
rect 18693 19904 18705 19907
rect 18656 19876 18705 19904
rect 18656 19864 18662 19876
rect 18693 19873 18705 19876
rect 18739 19873 18751 19907
rect 18693 19867 18751 19873
rect 18877 19907 18935 19913
rect 18877 19873 18889 19907
rect 18923 19904 18935 19907
rect 19260 19904 19288 20012
rect 21450 20000 21456 20012
rect 21508 20000 21514 20052
rect 22554 20000 22560 20052
rect 22612 20040 22618 20052
rect 22649 20043 22707 20049
rect 22649 20040 22661 20043
rect 22612 20012 22661 20040
rect 22612 20000 22618 20012
rect 22649 20009 22661 20012
rect 22695 20009 22707 20043
rect 22649 20003 22707 20009
rect 18923 19876 19288 19904
rect 18923 19873 18935 19876
rect 18877 19867 18935 19873
rect 14461 19839 14519 19845
rect 14461 19836 14473 19839
rect 14240 19808 14473 19836
rect 14240 19796 14246 19808
rect 14461 19805 14473 19808
rect 14507 19805 14519 19839
rect 14461 19799 14519 19805
rect 15565 19839 15623 19845
rect 15565 19805 15577 19839
rect 15611 19805 15623 19839
rect 15565 19799 15623 19805
rect 15654 19796 15660 19848
rect 15712 19836 15718 19848
rect 16390 19836 16396 19848
rect 15712 19808 15757 19836
rect 16351 19808 16396 19836
rect 15712 19796 15718 19808
rect 16390 19796 16396 19808
rect 16448 19796 16454 19848
rect 17126 19836 17132 19848
rect 16500 19808 17132 19836
rect 14366 19728 14372 19780
rect 14424 19768 14430 19780
rect 16500 19768 16528 19808
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 18138 19836 18144 19848
rect 18099 19808 18144 19836
rect 18138 19796 18144 19808
rect 18196 19796 18202 19848
rect 17678 19768 17684 19780
rect 14424 19740 16528 19768
rect 16592 19740 17684 19768
rect 14424 19728 14430 19740
rect 12161 19703 12219 19709
rect 12161 19700 12173 19703
rect 12124 19672 12173 19700
rect 12124 19660 12130 19672
rect 12161 19669 12173 19672
rect 12207 19669 12219 19703
rect 12161 19663 12219 19669
rect 13909 19703 13967 19709
rect 13909 19669 13921 19703
rect 13955 19700 13967 19703
rect 14182 19700 14188 19712
rect 13955 19672 14188 19700
rect 13955 19669 13967 19672
rect 13909 19663 13967 19669
rect 14182 19660 14188 19672
rect 14240 19660 14246 19712
rect 16298 19700 16304 19712
rect 16259 19672 16304 19700
rect 16298 19660 16304 19672
rect 16356 19660 16362 19712
rect 16592 19709 16620 19740
rect 17678 19728 17684 19740
rect 17736 19728 17742 19780
rect 17896 19771 17954 19777
rect 17896 19737 17908 19771
rect 17942 19768 17954 19771
rect 18892 19768 18920 19867
rect 19702 19864 19708 19916
rect 19760 19904 19766 19916
rect 20990 19904 20996 19916
rect 19760 19876 20996 19904
rect 19760 19864 19766 19876
rect 20990 19864 20996 19876
rect 21048 19864 21054 19916
rect 18966 19796 18972 19848
rect 19024 19836 19030 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 19024 19808 19257 19836
rect 19024 19796 19030 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19245 19799 19303 19805
rect 19334 19796 19340 19848
rect 19392 19836 19398 19848
rect 19981 19839 20039 19845
rect 19981 19836 19993 19839
rect 19392 19808 19993 19836
rect 19392 19796 19398 19808
rect 19981 19805 19993 19808
rect 20027 19805 20039 19839
rect 21174 19836 21180 19848
rect 21135 19808 21180 19836
rect 19981 19799 20039 19805
rect 21174 19796 21180 19808
rect 21232 19796 21238 19848
rect 21433 19839 21491 19845
rect 21433 19836 21445 19839
rect 21284 19808 21445 19836
rect 17942 19740 18920 19768
rect 17942 19737 17954 19740
rect 17896 19731 17954 19737
rect 20898 19728 20904 19780
rect 20956 19768 20962 19780
rect 21284 19768 21312 19808
rect 21433 19805 21445 19808
rect 21479 19805 21491 19839
rect 21433 19799 21491 19805
rect 22833 19839 22891 19845
rect 22833 19805 22845 19839
rect 22879 19836 22891 19839
rect 23566 19836 23572 19848
rect 22879 19808 23572 19836
rect 22879 19805 22891 19808
rect 22833 19799 22891 19805
rect 23566 19796 23572 19808
rect 23624 19796 23630 19848
rect 20956 19740 21312 19768
rect 20956 19728 20962 19740
rect 16577 19703 16635 19709
rect 16577 19669 16589 19703
rect 16623 19669 16635 19703
rect 16577 19663 16635 19669
rect 16761 19703 16819 19709
rect 16761 19669 16773 19703
rect 16807 19700 16819 19703
rect 17586 19700 17592 19712
rect 16807 19672 17592 19700
rect 16807 19669 16819 19672
rect 16761 19663 16819 19669
rect 17586 19660 17592 19672
rect 17644 19660 17650 19712
rect 18230 19700 18236 19712
rect 18191 19672 18236 19700
rect 18230 19660 18236 19672
rect 18288 19660 18294 19712
rect 18598 19700 18604 19712
rect 18559 19672 18604 19700
rect 18598 19660 18604 19672
rect 18656 19660 18662 19712
rect 19610 19660 19616 19712
rect 19668 19700 19674 19712
rect 19711 19703 19769 19709
rect 19711 19700 19723 19703
rect 19668 19672 19723 19700
rect 19668 19660 19674 19672
rect 19711 19669 19723 19672
rect 19757 19669 19769 19703
rect 21082 19700 21088 19712
rect 21043 19672 21088 19700
rect 19711 19663 19769 19669
rect 21082 19660 21088 19672
rect 21140 19700 21146 19712
rect 22094 19700 22100 19712
rect 21140 19672 22100 19700
rect 21140 19660 21146 19672
rect 22094 19660 22100 19672
rect 22152 19660 22158 19712
rect 22554 19700 22560 19712
rect 22515 19672 22560 19700
rect 22554 19660 22560 19672
rect 22612 19660 22618 19712
rect 23014 19700 23020 19712
rect 22975 19672 23020 19700
rect 23014 19660 23020 19672
rect 23072 19660 23078 19712
rect 1104 19610 23460 19632
rect 1104 19558 6548 19610
rect 6600 19558 6612 19610
rect 6664 19558 6676 19610
rect 6728 19558 6740 19610
rect 6792 19558 6804 19610
rect 6856 19558 12146 19610
rect 12198 19558 12210 19610
rect 12262 19558 12274 19610
rect 12326 19558 12338 19610
rect 12390 19558 12402 19610
rect 12454 19558 17744 19610
rect 17796 19558 17808 19610
rect 17860 19558 17872 19610
rect 17924 19558 17936 19610
rect 17988 19558 18000 19610
rect 18052 19558 23460 19610
rect 1104 19536 23460 19558
rect 1486 19456 1492 19508
rect 1544 19496 1550 19508
rect 1581 19499 1639 19505
rect 1581 19496 1593 19499
rect 1544 19468 1593 19496
rect 1544 19456 1550 19468
rect 1581 19465 1593 19468
rect 1627 19465 1639 19499
rect 1581 19459 1639 19465
rect 2774 19456 2780 19508
rect 2832 19496 2838 19508
rect 3053 19499 3111 19505
rect 3053 19496 3065 19499
rect 2832 19468 3065 19496
rect 2832 19456 2838 19468
rect 3053 19465 3065 19468
rect 3099 19465 3111 19499
rect 3053 19459 3111 19465
rect 4801 19499 4859 19505
rect 4801 19465 4813 19499
rect 4847 19465 4859 19499
rect 4801 19459 4859 19465
rect 4154 19428 4160 19440
rect 1412 19400 4160 19428
rect 1412 19369 1440 19400
rect 4154 19388 4160 19400
rect 4212 19388 4218 19440
rect 4338 19428 4344 19440
rect 4299 19400 4344 19428
rect 4338 19388 4344 19400
rect 4396 19388 4402 19440
rect 4816 19428 4844 19459
rect 4890 19456 4896 19508
rect 4948 19496 4954 19508
rect 6362 19496 6368 19508
rect 4948 19468 4993 19496
rect 6323 19468 6368 19496
rect 4948 19456 4954 19468
rect 6362 19456 6368 19468
rect 6420 19456 6426 19508
rect 6917 19499 6975 19505
rect 6917 19465 6929 19499
rect 6963 19465 6975 19499
rect 6917 19459 6975 19465
rect 5261 19431 5319 19437
rect 5261 19428 5273 19431
rect 4816 19400 5273 19428
rect 5261 19397 5273 19400
rect 5307 19428 5319 19431
rect 6932 19428 6960 19459
rect 8110 19456 8116 19508
rect 8168 19496 8174 19508
rect 8386 19496 8392 19508
rect 8168 19468 8392 19496
rect 8168 19456 8174 19468
rect 8386 19456 8392 19468
rect 8444 19456 8450 19508
rect 9125 19499 9183 19505
rect 9125 19465 9137 19499
rect 9171 19496 9183 19499
rect 9766 19496 9772 19508
rect 9171 19468 9772 19496
rect 9171 19465 9183 19468
rect 9125 19459 9183 19465
rect 9766 19456 9772 19468
rect 9824 19456 9830 19508
rect 10042 19496 10048 19508
rect 10003 19468 10048 19496
rect 10042 19456 10048 19468
rect 10100 19456 10106 19508
rect 10318 19496 10324 19508
rect 10279 19468 10324 19496
rect 10318 19456 10324 19468
rect 10376 19456 10382 19508
rect 11333 19499 11391 19505
rect 11333 19465 11345 19499
rect 11379 19496 11391 19499
rect 11606 19496 11612 19508
rect 11379 19468 11612 19496
rect 11379 19465 11391 19468
rect 11333 19459 11391 19465
rect 11606 19456 11612 19468
rect 11664 19456 11670 19508
rect 11977 19499 12035 19505
rect 11977 19465 11989 19499
rect 12023 19496 12035 19499
rect 14090 19496 14096 19508
rect 12023 19468 14096 19496
rect 12023 19465 12035 19468
rect 11977 19459 12035 19465
rect 14090 19456 14096 19468
rect 14148 19456 14154 19508
rect 14366 19496 14372 19508
rect 14327 19468 14372 19496
rect 14366 19456 14372 19468
rect 14424 19456 14430 19508
rect 15194 19456 15200 19508
rect 15252 19496 15258 19508
rect 16945 19499 17003 19505
rect 15252 19468 16160 19496
rect 15252 19456 15258 19468
rect 7006 19428 7012 19440
rect 5307 19400 6776 19428
rect 6932 19400 7012 19428
rect 5307 19397 5319 19400
rect 5261 19391 5319 19397
rect 1397 19363 1455 19369
rect 1397 19329 1409 19363
rect 1443 19329 1455 19363
rect 1397 19323 1455 19329
rect 1578 19320 1584 19372
rect 1636 19360 1642 19372
rect 1673 19363 1731 19369
rect 1673 19360 1685 19363
rect 1636 19332 1685 19360
rect 1636 19320 1642 19332
rect 1673 19329 1685 19332
rect 1719 19329 1731 19363
rect 1673 19323 1731 19329
rect 1940 19363 1998 19369
rect 1940 19329 1952 19363
rect 1986 19360 1998 19363
rect 3329 19363 3387 19369
rect 3329 19360 3341 19363
rect 1986 19332 3341 19360
rect 1986 19329 1998 19332
rect 1940 19323 1998 19329
rect 3329 19329 3341 19332
rect 3375 19329 3387 19363
rect 3329 19323 3387 19329
rect 3973 19363 4031 19369
rect 3973 19329 3985 19363
rect 4019 19360 4031 19363
rect 4430 19360 4436 19372
rect 4019 19332 4292 19360
rect 4391 19332 4436 19360
rect 4019 19329 4031 19332
rect 3973 19323 4031 19329
rect 4154 19292 4160 19304
rect 4115 19264 4160 19292
rect 4154 19252 4160 19264
rect 4212 19252 4218 19304
rect 4264 19292 4292 19332
rect 4430 19320 4436 19332
rect 4488 19320 4494 19372
rect 5994 19360 6000 19372
rect 5955 19332 6000 19360
rect 5994 19320 6000 19332
rect 6052 19320 6058 19372
rect 6748 19369 6776 19400
rect 7006 19388 7012 19400
rect 7064 19388 7070 19440
rect 7190 19388 7196 19440
rect 7248 19428 7254 19440
rect 7248 19400 7328 19428
rect 7248 19388 7254 19400
rect 7300 19369 7328 19400
rect 8846 19388 8852 19440
rect 8904 19428 8910 19440
rect 10689 19431 10747 19437
rect 8904 19400 9996 19428
rect 8904 19388 8910 19400
rect 6733 19363 6791 19369
rect 6733 19329 6745 19363
rect 6779 19329 6791 19363
rect 6733 19323 6791 19329
rect 7285 19363 7343 19369
rect 7285 19329 7297 19363
rect 7331 19329 7343 19363
rect 7285 19323 7343 19329
rect 7608 19363 7666 19369
rect 7608 19329 7620 19363
rect 7654 19329 7666 19363
rect 9214 19360 9220 19372
rect 9175 19332 9220 19360
rect 7608 19323 7666 19329
rect 4706 19292 4712 19304
rect 4264 19264 4712 19292
rect 4706 19252 4712 19264
rect 4764 19252 4770 19304
rect 4798 19252 4804 19304
rect 4856 19292 4862 19304
rect 5353 19295 5411 19301
rect 5353 19292 5365 19295
rect 4856 19264 5365 19292
rect 4856 19252 4862 19264
rect 5353 19261 5365 19264
rect 5399 19261 5411 19295
rect 5353 19255 5411 19261
rect 5445 19295 5503 19301
rect 5445 19261 5457 19295
rect 5491 19261 5503 19295
rect 5445 19255 5503 19261
rect 3142 19184 3148 19236
rect 3200 19224 3206 19236
rect 3237 19227 3295 19233
rect 3237 19224 3249 19227
rect 3200 19196 3249 19224
rect 3200 19184 3206 19196
rect 3237 19193 3249 19196
rect 3283 19224 3295 19227
rect 3418 19224 3424 19236
rect 3283 19196 3424 19224
rect 3283 19193 3295 19196
rect 3237 19187 3295 19193
rect 3418 19184 3424 19196
rect 3476 19184 3482 19236
rect 4246 19184 4252 19236
rect 4304 19224 4310 19236
rect 5460 19224 5488 19255
rect 7006 19252 7012 19304
rect 7064 19292 7070 19304
rect 7193 19295 7251 19301
rect 7193 19292 7205 19295
rect 7064 19264 7205 19292
rect 7064 19252 7070 19264
rect 7193 19261 7205 19264
rect 7239 19261 7251 19295
rect 7193 19255 7251 19261
rect 7466 19252 7472 19304
rect 7524 19292 7530 19304
rect 7623 19292 7651 19323
rect 9214 19320 9220 19332
rect 9272 19320 9278 19372
rect 9677 19363 9735 19369
rect 9677 19329 9689 19363
rect 9723 19360 9735 19363
rect 9858 19360 9864 19372
rect 9723 19332 9864 19360
rect 9723 19329 9735 19332
rect 9677 19323 9735 19329
rect 9858 19320 9864 19332
rect 9916 19320 9922 19372
rect 9968 19369 9996 19400
rect 10689 19397 10701 19431
rect 10735 19428 10747 19431
rect 11054 19428 11060 19440
rect 10735 19400 11060 19428
rect 10735 19397 10747 19400
rect 10689 19391 10747 19397
rect 11054 19388 11060 19400
rect 11112 19388 11118 19440
rect 16132 19437 16160 19468
rect 16945 19465 16957 19499
rect 16991 19496 17003 19499
rect 18969 19499 19027 19505
rect 16991 19468 18920 19496
rect 16991 19465 17003 19468
rect 16945 19459 17003 19465
rect 13204 19431 13262 19437
rect 13204 19397 13216 19431
rect 13250 19428 13262 19431
rect 15289 19431 15347 19437
rect 15289 19428 15301 19431
rect 13250 19400 15301 19428
rect 13250 19397 13262 19400
rect 13204 19391 13262 19397
rect 15289 19397 15301 19400
rect 15335 19397 15347 19431
rect 15289 19391 15347 19397
rect 16117 19431 16175 19437
rect 16117 19397 16129 19431
rect 16163 19397 16175 19431
rect 18892 19428 18920 19468
rect 18969 19465 18981 19499
rect 19015 19496 19027 19499
rect 19242 19496 19248 19508
rect 19015 19468 19248 19496
rect 19015 19465 19027 19468
rect 18969 19459 19027 19465
rect 19242 19456 19248 19468
rect 19300 19456 19306 19508
rect 21266 19496 21272 19508
rect 19536 19468 21272 19496
rect 19536 19428 19564 19468
rect 21266 19456 21272 19468
rect 21324 19456 21330 19508
rect 21821 19499 21879 19505
rect 21821 19465 21833 19499
rect 21867 19465 21879 19499
rect 22278 19496 22284 19508
rect 22239 19468 22284 19496
rect 21821 19459 21879 19465
rect 18892 19400 19564 19428
rect 16117 19391 16175 19397
rect 20622 19388 20628 19440
rect 20680 19428 20686 19440
rect 21836 19428 21864 19459
rect 22278 19456 22284 19468
rect 22336 19456 22342 19508
rect 23017 19499 23075 19505
rect 23017 19465 23029 19499
rect 23063 19496 23075 19499
rect 23198 19496 23204 19508
rect 23063 19468 23204 19496
rect 23063 19465 23075 19468
rect 23017 19459 23075 19465
rect 23198 19456 23204 19468
rect 23256 19456 23262 19508
rect 23658 19428 23664 19440
rect 20680 19400 21864 19428
rect 22066 19400 23664 19428
rect 20680 19388 20686 19400
rect 9953 19363 10011 19369
rect 9953 19329 9965 19363
rect 9999 19329 10011 19363
rect 10229 19363 10287 19369
rect 10229 19360 10241 19363
rect 9953 19323 10011 19329
rect 10060 19332 10241 19360
rect 7524 19264 7651 19292
rect 7524 19252 7530 19264
rect 7742 19252 7748 19304
rect 7800 19292 7806 19304
rect 7800 19264 7845 19292
rect 7800 19252 7806 19264
rect 7926 19252 7932 19304
rect 7984 19301 7990 19304
rect 7984 19295 8033 19301
rect 7984 19261 7987 19295
rect 8021 19261 8033 19295
rect 7984 19255 8033 19261
rect 7984 19252 7990 19255
rect 8662 19252 8668 19304
rect 8720 19292 8726 19304
rect 10060 19292 10088 19332
rect 10229 19329 10241 19332
rect 10275 19329 10287 19363
rect 11146 19360 11152 19372
rect 11107 19332 11152 19360
rect 10229 19323 10287 19329
rect 11146 19320 11152 19332
rect 11204 19320 11210 19372
rect 11514 19360 11520 19372
rect 11475 19332 11520 19360
rect 11514 19320 11520 19332
rect 11572 19320 11578 19372
rect 11793 19363 11851 19369
rect 11793 19329 11805 19363
rect 11839 19360 11851 19363
rect 12434 19360 12440 19372
rect 11839 19332 12440 19360
rect 11839 19329 11851 19332
rect 11793 19323 11851 19329
rect 12434 19320 12440 19332
rect 12492 19320 12498 19372
rect 13446 19360 13452 19372
rect 13407 19332 13452 19360
rect 13446 19320 13452 19332
rect 13504 19320 13510 19372
rect 13998 19360 14004 19372
rect 13959 19332 14004 19360
rect 13998 19320 14004 19332
rect 14056 19320 14062 19372
rect 14826 19360 14832 19372
rect 14787 19332 14832 19360
rect 14826 19320 14832 19332
rect 14884 19320 14890 19372
rect 14921 19363 14979 19369
rect 14921 19329 14933 19363
rect 14967 19360 14979 19363
rect 15654 19360 15660 19372
rect 14967 19332 15660 19360
rect 14967 19329 14979 19332
rect 14921 19323 14979 19329
rect 15654 19320 15660 19332
rect 15712 19320 15718 19372
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 15764 19332 15945 19360
rect 10778 19292 10784 19304
rect 8720 19264 10088 19292
rect 10739 19264 10784 19292
rect 8720 19252 8726 19264
rect 10778 19252 10784 19264
rect 10836 19252 10842 19304
rect 10873 19295 10931 19301
rect 10873 19261 10885 19295
rect 10919 19261 10931 19295
rect 13725 19295 13783 19301
rect 10873 19255 10931 19261
rect 10980 19264 12480 19292
rect 4304 19196 5488 19224
rect 4304 19184 4310 19196
rect 8846 19184 8852 19236
rect 8904 19224 8910 19236
rect 9493 19227 9551 19233
rect 9493 19224 9505 19227
rect 8904 19196 9505 19224
rect 8904 19184 8910 19196
rect 9493 19193 9505 19196
rect 9539 19193 9551 19227
rect 9493 19187 9551 19193
rect 9858 19184 9864 19236
rect 9916 19224 9922 19236
rect 10888 19224 10916 19255
rect 9916 19196 10916 19224
rect 9916 19184 9922 19196
rect 3510 19116 3516 19168
rect 3568 19156 3574 19168
rect 4522 19156 4528 19168
rect 3568 19128 4528 19156
rect 3568 19116 3574 19128
rect 4522 19116 4528 19128
rect 4580 19116 4586 19168
rect 5810 19156 5816 19168
rect 5771 19128 5816 19156
rect 5810 19116 5816 19128
rect 5868 19116 5874 19168
rect 6178 19156 6184 19168
rect 6139 19128 6184 19156
rect 6178 19116 6184 19128
rect 6236 19116 6242 19168
rect 7006 19116 7012 19168
rect 7064 19156 7070 19168
rect 8386 19156 8392 19168
rect 7064 19128 8392 19156
rect 7064 19116 7070 19128
rect 8386 19116 8392 19128
rect 8444 19116 8450 19168
rect 8662 19116 8668 19168
rect 8720 19156 8726 19168
rect 9030 19156 9036 19168
rect 8720 19128 9036 19156
rect 8720 19116 8726 19128
rect 9030 19116 9036 19128
rect 9088 19116 9094 19168
rect 9122 19116 9128 19168
rect 9180 19156 9186 19168
rect 9401 19159 9459 19165
rect 9401 19156 9413 19159
rect 9180 19128 9413 19156
rect 9180 19116 9186 19128
rect 9401 19125 9413 19128
rect 9447 19125 9459 19159
rect 9401 19119 9459 19125
rect 9769 19159 9827 19165
rect 9769 19125 9781 19159
rect 9815 19156 9827 19159
rect 9950 19156 9956 19168
rect 9815 19128 9956 19156
rect 9815 19125 9827 19128
rect 9769 19119 9827 19125
rect 9950 19116 9956 19128
rect 10008 19116 10014 19168
rect 10502 19116 10508 19168
rect 10560 19156 10566 19168
rect 10980 19156 11008 19264
rect 11790 19184 11796 19236
rect 11848 19224 11854 19236
rect 12452 19224 12480 19264
rect 13725 19261 13737 19295
rect 13771 19261 13783 19295
rect 13725 19255 13783 19261
rect 13740 19224 13768 19255
rect 13814 19252 13820 19304
rect 13872 19292 13878 19304
rect 13909 19295 13967 19301
rect 13909 19292 13921 19295
rect 13872 19264 13921 19292
rect 13872 19252 13878 19264
rect 13909 19261 13921 19264
rect 13955 19261 13967 19295
rect 15010 19292 15016 19304
rect 14971 19264 15016 19292
rect 13909 19255 13967 19261
rect 15010 19252 15016 19264
rect 15068 19252 15074 19304
rect 15764 19292 15792 19332
rect 15933 19329 15945 19332
rect 15979 19329 15991 19363
rect 16761 19363 16819 19369
rect 16761 19360 16773 19363
rect 15933 19323 15991 19329
rect 16408 19332 16773 19360
rect 15120 19264 15792 19292
rect 14274 19224 14280 19236
rect 11848 19196 12204 19224
rect 12452 19196 12572 19224
rect 13740 19196 14280 19224
rect 11848 19184 11854 19196
rect 10560 19128 11008 19156
rect 10560 19116 10566 19128
rect 11238 19116 11244 19168
rect 11296 19156 11302 19168
rect 11514 19156 11520 19168
rect 11296 19128 11520 19156
rect 11296 19116 11302 19128
rect 11514 19116 11520 19128
rect 11572 19116 11578 19168
rect 11698 19156 11704 19168
rect 11659 19128 11704 19156
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 11974 19116 11980 19168
rect 12032 19156 12038 19168
rect 12069 19159 12127 19165
rect 12069 19156 12081 19159
rect 12032 19128 12081 19156
rect 12032 19116 12038 19128
rect 12069 19125 12081 19128
rect 12115 19125 12127 19159
rect 12176 19156 12204 19196
rect 12434 19156 12440 19168
rect 12176 19128 12440 19156
rect 12069 19119 12127 19125
rect 12434 19116 12440 19128
rect 12492 19116 12498 19168
rect 12544 19156 12572 19196
rect 14274 19184 14280 19196
rect 14332 19184 14338 19236
rect 14384 19196 14688 19224
rect 14384 19156 14412 19196
rect 12544 19128 14412 19156
rect 14458 19116 14464 19168
rect 14516 19156 14522 19168
rect 14660 19156 14688 19196
rect 14826 19184 14832 19236
rect 14884 19224 14890 19236
rect 15120 19224 15148 19264
rect 16206 19252 16212 19304
rect 16264 19292 16270 19304
rect 16408 19301 16436 19332
rect 16761 19329 16773 19332
rect 16807 19329 16819 19363
rect 16761 19323 16819 19329
rect 17034 19320 17040 19372
rect 17092 19360 17098 19372
rect 19061 19363 19119 19369
rect 19061 19360 19073 19363
rect 17092 19332 19073 19360
rect 17092 19320 17098 19332
rect 19061 19329 19073 19332
rect 19107 19329 19119 19363
rect 19061 19323 19119 19329
rect 19981 19363 20039 19369
rect 19981 19329 19993 19363
rect 20027 19329 20039 19363
rect 20898 19360 20904 19372
rect 20859 19332 20904 19360
rect 19981 19323 20039 19329
rect 16393 19295 16451 19301
rect 16393 19292 16405 19295
rect 16264 19264 16405 19292
rect 16264 19252 16270 19264
rect 16393 19261 16405 19264
rect 16439 19261 16451 19295
rect 16393 19255 16451 19261
rect 16850 19252 16856 19304
rect 16908 19292 16914 19304
rect 17494 19301 17500 19304
rect 17129 19295 17187 19301
rect 17129 19292 17141 19295
rect 16908 19264 17141 19292
rect 16908 19252 16914 19264
rect 17129 19261 17141 19264
rect 17175 19261 17187 19295
rect 17129 19255 17187 19261
rect 17452 19295 17500 19301
rect 17452 19261 17464 19295
rect 17498 19261 17500 19295
rect 17452 19255 17500 19261
rect 14884 19196 15148 19224
rect 14884 19184 14890 19196
rect 15286 19156 15292 19168
rect 14516 19128 14561 19156
rect 14660 19128 15292 19156
rect 14516 19116 14522 19128
rect 15286 19116 15292 19128
rect 15344 19116 15350 19168
rect 16206 19156 16212 19168
rect 16167 19128 16212 19156
rect 16206 19116 16212 19128
rect 16264 19116 16270 19168
rect 17144 19156 17172 19255
rect 17494 19252 17500 19255
rect 17552 19252 17558 19304
rect 17586 19252 17592 19304
rect 17644 19292 17650 19304
rect 17865 19295 17923 19301
rect 17644 19264 17689 19292
rect 17644 19252 17650 19264
rect 17865 19261 17877 19295
rect 17911 19292 17923 19295
rect 18598 19292 18604 19304
rect 17911 19264 18604 19292
rect 17911 19261 17923 19264
rect 17865 19255 17923 19261
rect 18598 19252 18604 19264
rect 18656 19252 18662 19304
rect 19150 19252 19156 19304
rect 19208 19292 19214 19304
rect 19996 19292 20024 19323
rect 20898 19320 20904 19332
rect 20956 19320 20962 19372
rect 20993 19363 21051 19369
rect 20993 19329 21005 19363
rect 21039 19360 21051 19363
rect 21358 19360 21364 19372
rect 21039 19332 21364 19360
rect 21039 19329 21051 19332
rect 20993 19323 21051 19329
rect 21358 19320 21364 19332
rect 21416 19320 21422 19372
rect 21637 19363 21695 19369
rect 21637 19329 21649 19363
rect 21683 19360 21695 19363
rect 22066 19360 22094 19400
rect 23658 19388 23664 19400
rect 23716 19388 23722 19440
rect 22186 19360 22192 19372
rect 21683 19332 22094 19360
rect 22147 19332 22192 19360
rect 21683 19329 21695 19332
rect 21637 19323 21695 19329
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 22830 19360 22836 19372
rect 22296 19332 22508 19360
rect 22791 19332 22836 19360
rect 19208 19264 20024 19292
rect 19208 19252 19214 19264
rect 19794 19224 19800 19236
rect 19755 19196 19800 19224
rect 19794 19184 19800 19196
rect 19852 19184 19858 19236
rect 19996 19224 20024 19264
rect 21450 19252 21456 19304
rect 21508 19292 21514 19304
rect 22296 19292 22324 19332
rect 21508 19264 22324 19292
rect 22373 19295 22431 19301
rect 21508 19252 21514 19264
rect 22373 19261 22385 19295
rect 22419 19261 22431 19295
rect 22480 19292 22508 19332
rect 22830 19320 22836 19332
rect 22888 19320 22894 19372
rect 22649 19295 22707 19301
rect 22649 19292 22661 19295
rect 22480 19264 22661 19292
rect 22373 19255 22431 19261
rect 22649 19261 22661 19264
rect 22695 19261 22707 19295
rect 22649 19255 22707 19261
rect 19996 19196 21588 19224
rect 19334 19156 19340 19168
rect 17144 19128 19340 19156
rect 19334 19116 19340 19128
rect 19392 19116 19398 19168
rect 19518 19116 19524 19168
rect 19576 19156 19582 19168
rect 19705 19159 19763 19165
rect 19705 19156 19717 19159
rect 19576 19128 19717 19156
rect 19576 19116 19582 19128
rect 19705 19125 19717 19128
rect 19751 19125 19763 19159
rect 20254 19156 20260 19168
rect 20215 19128 20260 19156
rect 19705 19119 19763 19125
rect 20254 19116 20260 19128
rect 20312 19116 20318 19168
rect 21560 19156 21588 19196
rect 21634 19184 21640 19236
rect 21692 19224 21698 19236
rect 22388 19224 22416 19255
rect 21692 19196 22416 19224
rect 21692 19184 21698 19196
rect 22922 19156 22928 19168
rect 21560 19128 22928 19156
rect 22922 19116 22928 19128
rect 22980 19116 22986 19168
rect 1104 19066 23460 19088
rect 1104 19014 3749 19066
rect 3801 19014 3813 19066
rect 3865 19014 3877 19066
rect 3929 19014 3941 19066
rect 3993 19014 4005 19066
rect 4057 19014 9347 19066
rect 9399 19014 9411 19066
rect 9463 19014 9475 19066
rect 9527 19014 9539 19066
rect 9591 19014 9603 19066
rect 9655 19014 14945 19066
rect 14997 19014 15009 19066
rect 15061 19014 15073 19066
rect 15125 19014 15137 19066
rect 15189 19014 15201 19066
rect 15253 19014 20543 19066
rect 20595 19014 20607 19066
rect 20659 19014 20671 19066
rect 20723 19014 20735 19066
rect 20787 19014 20799 19066
rect 20851 19014 23460 19066
rect 1104 18992 23460 19014
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 4430 18952 4436 18964
rect 1728 18924 4436 18952
rect 1728 18912 1734 18924
rect 4430 18912 4436 18924
rect 4488 18912 4494 18964
rect 4798 18952 4804 18964
rect 4759 18924 4804 18952
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 6178 18912 6184 18964
rect 6236 18952 6242 18964
rect 8662 18952 8668 18964
rect 6236 18924 8668 18952
rect 6236 18912 6242 18924
rect 8662 18912 8668 18924
rect 8720 18912 8726 18964
rect 12805 18955 12863 18961
rect 9149 18924 12434 18952
rect 1762 18844 1768 18896
rect 1820 18884 1826 18896
rect 1820 18856 3740 18884
rect 1820 18844 1826 18856
rect 1302 18776 1308 18828
rect 1360 18816 1366 18828
rect 3510 18816 3516 18828
rect 1360 18788 3516 18816
rect 1360 18776 1366 18788
rect 3510 18776 3516 18788
rect 3568 18776 3574 18828
rect 1394 18708 1400 18760
rect 1452 18748 1458 18760
rect 1489 18751 1547 18757
rect 1489 18748 1501 18751
rect 1452 18720 1501 18748
rect 1452 18708 1458 18720
rect 1489 18717 1501 18720
rect 1535 18717 1547 18751
rect 1489 18711 1547 18717
rect 2133 18751 2191 18757
rect 2133 18717 2145 18751
rect 2179 18717 2191 18751
rect 2133 18711 2191 18717
rect 2869 18751 2927 18757
rect 2869 18717 2881 18751
rect 2915 18717 2927 18751
rect 3602 18748 3608 18760
rect 3563 18720 3608 18748
rect 2869 18711 2927 18717
rect 2148 18680 2176 18711
rect 2056 18652 2176 18680
rect 2884 18680 2912 18711
rect 3602 18708 3608 18720
rect 3660 18708 3666 18760
rect 3712 18748 3740 18856
rect 4154 18844 4160 18896
rect 4212 18884 4218 18896
rect 7190 18884 7196 18896
rect 4212 18856 5488 18884
rect 7151 18856 7196 18884
rect 4212 18844 4218 18856
rect 4433 18819 4491 18825
rect 4433 18785 4445 18819
rect 4479 18816 4491 18819
rect 4614 18816 4620 18828
rect 4479 18788 4620 18816
rect 4479 18785 4491 18788
rect 4433 18779 4491 18785
rect 4614 18776 4620 18788
rect 4672 18776 4678 18828
rect 5460 18825 5488 18856
rect 7190 18844 7196 18856
rect 7248 18844 7254 18896
rect 5445 18819 5503 18825
rect 5445 18785 5457 18819
rect 5491 18816 5503 18819
rect 8846 18816 8852 18828
rect 5491 18788 8852 18816
rect 5491 18785 5503 18788
rect 5445 18779 5503 18785
rect 8846 18776 8852 18788
rect 8904 18776 8910 18828
rect 5169 18751 5227 18757
rect 3712 18720 4752 18748
rect 4430 18680 4436 18692
rect 2884 18652 4436 18680
rect 2056 18624 2084 18652
rect 4430 18640 4436 18652
rect 4488 18640 4494 18692
rect 4724 18689 4752 18720
rect 5169 18717 5181 18751
rect 5215 18748 5227 18751
rect 5810 18748 5816 18760
rect 5215 18720 5816 18748
rect 5215 18717 5227 18720
rect 5169 18711 5227 18717
rect 5810 18708 5816 18720
rect 5868 18708 5874 18760
rect 6178 18708 6184 18760
rect 6236 18748 6242 18760
rect 6273 18751 6331 18757
rect 6273 18748 6285 18751
rect 6236 18720 6285 18748
rect 6236 18708 6242 18720
rect 6273 18717 6285 18720
rect 6319 18717 6331 18751
rect 6273 18711 6331 18717
rect 6454 18708 6460 18760
rect 6512 18748 6518 18760
rect 7009 18751 7067 18757
rect 7009 18748 7021 18751
rect 6512 18720 7021 18748
rect 6512 18708 6518 18720
rect 7009 18717 7021 18720
rect 7055 18717 7067 18751
rect 7926 18748 7932 18760
rect 7887 18720 7932 18748
rect 7009 18711 7067 18717
rect 7926 18708 7932 18720
rect 7984 18708 7990 18760
rect 8110 18708 8116 18760
rect 8168 18748 8174 18760
rect 8294 18748 8300 18760
rect 8168 18720 8300 18748
rect 8168 18708 8174 18720
rect 8294 18708 8300 18720
rect 8352 18708 8358 18760
rect 8570 18708 8576 18760
rect 8628 18748 8634 18760
rect 8665 18751 8723 18757
rect 8665 18748 8677 18751
rect 8628 18720 8677 18748
rect 8628 18708 8634 18720
rect 8665 18717 8677 18720
rect 8711 18717 8723 18751
rect 9149 18748 9177 18924
rect 9306 18844 9312 18896
rect 9364 18884 9370 18896
rect 9674 18884 9680 18896
rect 9364 18856 9680 18884
rect 9364 18844 9370 18856
rect 9674 18844 9680 18856
rect 9732 18844 9738 18896
rect 10502 18884 10508 18896
rect 9784 18856 10508 18884
rect 9214 18776 9220 18828
rect 9272 18816 9278 18828
rect 9784 18816 9812 18856
rect 10502 18844 10508 18856
rect 10560 18844 10566 18896
rect 12406 18884 12434 18924
rect 12805 18921 12817 18955
rect 12851 18952 12863 18955
rect 13814 18952 13820 18964
rect 12851 18924 13820 18952
rect 12851 18921 12863 18924
rect 12805 18915 12863 18921
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 13909 18955 13967 18961
rect 13909 18921 13921 18955
rect 13955 18952 13967 18955
rect 13998 18952 14004 18964
rect 13955 18924 14004 18952
rect 13955 18921 13967 18924
rect 13909 18915 13967 18921
rect 13998 18912 14004 18924
rect 14056 18912 14062 18964
rect 14093 18955 14151 18961
rect 14093 18921 14105 18955
rect 14139 18952 14151 18955
rect 14826 18952 14832 18964
rect 14139 18924 14832 18952
rect 14139 18921 14151 18924
rect 14093 18915 14151 18921
rect 14826 18912 14832 18924
rect 14884 18912 14890 18964
rect 15565 18955 15623 18961
rect 15565 18921 15577 18955
rect 15611 18952 15623 18955
rect 15654 18952 15660 18964
rect 15611 18924 15660 18952
rect 15611 18921 15623 18924
rect 15565 18915 15623 18921
rect 15654 18912 15660 18924
rect 15712 18912 15718 18964
rect 15930 18912 15936 18964
rect 15988 18952 15994 18964
rect 17313 18955 17371 18961
rect 15988 18924 16988 18952
rect 15988 18912 15994 18924
rect 14366 18884 14372 18896
rect 12406 18856 14372 18884
rect 14366 18844 14372 18856
rect 14424 18844 14430 18896
rect 9272 18788 9812 18816
rect 10229 18819 10287 18825
rect 10229 18814 10241 18819
rect 9272 18776 9278 18788
rect 10152 18786 10241 18814
rect 8665 18711 8723 18717
rect 8772 18720 9177 18748
rect 9585 18751 9643 18757
rect 4709 18683 4767 18689
rect 4709 18649 4721 18683
rect 4755 18680 4767 18683
rect 8772 18680 8800 18720
rect 9585 18717 9597 18751
rect 9631 18748 9643 18751
rect 9674 18748 9680 18760
rect 9631 18720 9680 18748
rect 9631 18717 9643 18720
rect 9585 18711 9643 18717
rect 9674 18708 9680 18720
rect 9732 18748 9738 18760
rect 10152 18748 10180 18786
rect 10229 18785 10241 18786
rect 10275 18785 10287 18819
rect 10229 18779 10287 18785
rect 11011 18819 11069 18825
rect 11011 18785 11023 18819
rect 11057 18816 11069 18819
rect 11422 18816 11428 18828
rect 11057 18788 11428 18816
rect 11057 18785 11069 18788
rect 11011 18779 11069 18785
rect 11422 18776 11428 18788
rect 11480 18776 11486 18828
rect 11900 18788 13400 18816
rect 10502 18748 10508 18760
rect 9732 18720 10180 18748
rect 10463 18720 10508 18748
rect 9732 18708 9738 18720
rect 10502 18708 10508 18720
rect 10560 18708 10566 18760
rect 10778 18708 10784 18760
rect 10836 18748 10842 18760
rect 11241 18751 11299 18757
rect 11241 18748 11253 18751
rect 10836 18720 11253 18748
rect 10836 18708 10842 18720
rect 11241 18717 11253 18720
rect 11287 18717 11299 18751
rect 11241 18711 11299 18717
rect 4755 18652 8800 18680
rect 8941 18683 8999 18689
rect 4755 18649 4767 18652
rect 4709 18643 4767 18649
rect 8941 18649 8953 18683
rect 8987 18680 8999 18683
rect 10318 18680 10324 18692
rect 8987 18652 10324 18680
rect 8987 18649 8999 18652
rect 8941 18643 8999 18649
rect 10318 18640 10324 18652
rect 10376 18640 10382 18692
rect 2038 18572 2044 18624
rect 2096 18572 2102 18624
rect 2222 18612 2228 18624
rect 2183 18584 2228 18612
rect 2222 18572 2228 18584
rect 2280 18572 2286 18624
rect 2314 18572 2320 18624
rect 2372 18612 2378 18624
rect 2961 18615 3019 18621
rect 2961 18612 2973 18615
rect 2372 18584 2973 18612
rect 2372 18572 2378 18584
rect 2961 18581 2973 18584
rect 3007 18581 3019 18615
rect 2961 18575 3019 18581
rect 3418 18572 3424 18624
rect 3476 18612 3482 18624
rect 3789 18615 3847 18621
rect 3789 18612 3801 18615
rect 3476 18584 3801 18612
rect 3476 18572 3482 18584
rect 3789 18581 3801 18584
rect 3835 18581 3847 18615
rect 4154 18612 4160 18624
rect 4115 18584 4160 18612
rect 3789 18575 3847 18581
rect 4154 18572 4160 18584
rect 4212 18572 4218 18624
rect 4246 18572 4252 18624
rect 4304 18612 4310 18624
rect 5258 18612 5264 18624
rect 4304 18584 4349 18612
rect 5219 18584 5264 18612
rect 4304 18572 4310 18584
rect 5258 18572 5264 18584
rect 5316 18572 5322 18624
rect 5350 18572 5356 18624
rect 5408 18612 5414 18624
rect 5629 18615 5687 18621
rect 5629 18612 5641 18615
rect 5408 18584 5641 18612
rect 5408 18572 5414 18584
rect 5629 18581 5641 18584
rect 5675 18581 5687 18615
rect 5629 18575 5687 18581
rect 5718 18572 5724 18624
rect 5776 18612 5782 18624
rect 6365 18615 6423 18621
rect 6365 18612 6377 18615
rect 5776 18584 6377 18612
rect 5776 18572 5782 18584
rect 6365 18581 6377 18584
rect 6411 18581 6423 18615
rect 6365 18575 6423 18581
rect 7190 18572 7196 18624
rect 7248 18612 7254 18624
rect 7285 18615 7343 18621
rect 7285 18612 7297 18615
rect 7248 18584 7297 18612
rect 7248 18572 7254 18584
rect 7285 18581 7297 18584
rect 7331 18581 7343 18615
rect 7285 18575 7343 18581
rect 8021 18615 8079 18621
rect 8021 18581 8033 18615
rect 8067 18612 8079 18615
rect 8294 18612 8300 18624
rect 8067 18584 8300 18612
rect 8067 18581 8079 18584
rect 8021 18575 8079 18581
rect 8294 18572 8300 18584
rect 8352 18572 8358 18624
rect 9490 18572 9496 18624
rect 9548 18612 9554 18624
rect 9677 18615 9735 18621
rect 9677 18612 9689 18615
rect 9548 18584 9689 18612
rect 9548 18572 9554 18584
rect 9677 18581 9689 18584
rect 9723 18581 9735 18615
rect 10042 18612 10048 18624
rect 10003 18584 10048 18612
rect 9677 18575 9735 18581
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 10137 18615 10195 18621
rect 10137 18581 10149 18615
rect 10183 18612 10195 18615
rect 10870 18612 10876 18624
rect 10183 18584 10876 18612
rect 10183 18581 10195 18584
rect 10137 18575 10195 18581
rect 10870 18572 10876 18584
rect 10928 18572 10934 18624
rect 10962 18572 10968 18624
rect 11020 18621 11026 18624
rect 11020 18612 11029 18621
rect 11900 18612 11928 18788
rect 12618 18748 12624 18760
rect 12579 18720 12624 18748
rect 12618 18708 12624 18720
rect 12676 18708 12682 18760
rect 12894 18748 12900 18760
rect 12855 18720 12900 18748
rect 12894 18708 12900 18720
rect 12952 18708 12958 18760
rect 12434 18680 12440 18692
rect 12360 18652 12440 18680
rect 12360 18621 12388 18652
rect 12434 18640 12440 18652
rect 12492 18680 12498 18692
rect 13262 18680 13268 18692
rect 12492 18652 13268 18680
rect 12492 18640 12498 18652
rect 13262 18640 13268 18652
rect 13320 18640 13326 18692
rect 13372 18680 13400 18788
rect 13446 18776 13452 18828
rect 13504 18816 13510 18828
rect 16960 18816 16988 18924
rect 17313 18921 17325 18955
rect 17359 18952 17371 18955
rect 17586 18952 17592 18964
rect 17359 18924 17592 18952
rect 17359 18921 17371 18924
rect 17313 18915 17371 18921
rect 17586 18912 17592 18924
rect 17644 18912 17650 18964
rect 17770 18912 17776 18964
rect 17828 18952 17834 18964
rect 18230 18952 18236 18964
rect 17828 18924 18236 18952
rect 17828 18912 17834 18924
rect 18230 18912 18236 18924
rect 18288 18912 18294 18964
rect 19886 18912 19892 18964
rect 19944 18952 19950 18964
rect 20438 18952 20444 18964
rect 19944 18924 20444 18952
rect 19944 18912 19950 18924
rect 20438 18912 20444 18924
rect 20496 18952 20502 18964
rect 20533 18955 20591 18961
rect 20533 18952 20545 18955
rect 20496 18924 20545 18952
rect 20496 18912 20502 18924
rect 20533 18921 20545 18924
rect 20579 18921 20591 18955
rect 21910 18952 21916 18964
rect 20533 18915 20591 18921
rect 20640 18924 21916 18952
rect 17221 18887 17279 18893
rect 17221 18853 17233 18887
rect 17267 18884 17279 18887
rect 17402 18884 17408 18896
rect 17267 18856 17408 18884
rect 17267 18853 17279 18856
rect 17221 18847 17279 18853
rect 17402 18844 17408 18856
rect 17460 18844 17466 18896
rect 18877 18887 18935 18893
rect 18877 18884 18889 18887
rect 17512 18856 18889 18884
rect 17512 18816 17540 18856
rect 18877 18853 18889 18856
rect 18923 18853 18935 18887
rect 18877 18847 18935 18853
rect 19334 18844 19340 18896
rect 19392 18884 19398 18896
rect 20346 18884 20352 18896
rect 19392 18856 20352 18884
rect 19392 18844 19398 18856
rect 20346 18844 20352 18856
rect 20404 18844 20410 18896
rect 13504 18788 14504 18816
rect 16960 18788 17540 18816
rect 13504 18776 13510 18788
rect 13725 18751 13783 18757
rect 13725 18717 13737 18751
rect 13771 18748 13783 18751
rect 14090 18748 14096 18760
rect 13771 18720 14096 18748
rect 13771 18717 13783 18720
rect 13725 18711 13783 18717
rect 14090 18708 14096 18720
rect 14148 18708 14154 18760
rect 14476 18748 14504 18788
rect 17586 18776 17592 18828
rect 17644 18816 17650 18828
rect 17865 18819 17923 18825
rect 17865 18816 17877 18819
rect 17644 18788 17877 18816
rect 17644 18776 17650 18788
rect 17865 18785 17877 18788
rect 17911 18785 17923 18819
rect 20640 18816 20668 18924
rect 21910 18912 21916 18924
rect 21968 18912 21974 18964
rect 23017 18955 23075 18961
rect 23017 18921 23029 18955
rect 23063 18952 23075 18955
rect 23106 18952 23112 18964
rect 23063 18924 23112 18952
rect 23063 18921 23075 18924
rect 23017 18915 23075 18921
rect 23106 18912 23112 18924
rect 23164 18912 23170 18964
rect 17865 18779 17923 18785
rect 17972 18788 20668 18816
rect 15470 18748 15476 18760
rect 14476 18720 15476 18748
rect 15470 18708 15476 18720
rect 15528 18748 15534 18760
rect 16945 18751 17003 18757
rect 16945 18748 16957 18751
rect 15528 18720 16957 18748
rect 15528 18708 15534 18720
rect 16945 18717 16957 18720
rect 16991 18717 17003 18751
rect 16945 18711 17003 18717
rect 17037 18751 17095 18757
rect 17037 18717 17049 18751
rect 17083 18748 17095 18751
rect 17126 18748 17132 18760
rect 17083 18720 17132 18748
rect 17083 18717 17095 18720
rect 17037 18711 17095 18717
rect 17126 18708 17132 18720
rect 17184 18708 17190 18760
rect 17770 18748 17776 18760
rect 17731 18720 17776 18748
rect 17770 18708 17776 18720
rect 17828 18708 17834 18760
rect 15228 18683 15286 18689
rect 13372 18652 15148 18680
rect 11020 18584 11928 18612
rect 12345 18615 12403 18621
rect 11020 18575 11029 18584
rect 12345 18581 12357 18615
rect 12391 18581 12403 18615
rect 12526 18612 12532 18624
rect 12487 18584 12532 18612
rect 12345 18575 12403 18581
rect 11020 18572 11026 18575
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 12986 18572 12992 18624
rect 13044 18612 13050 18624
rect 13541 18615 13599 18621
rect 13541 18612 13553 18615
rect 13044 18584 13553 18612
rect 13044 18572 13050 18584
rect 13541 18581 13553 18584
rect 13587 18581 13599 18615
rect 15120 18612 15148 18652
rect 15228 18649 15240 18683
rect 15274 18680 15286 18683
rect 16298 18680 16304 18692
rect 15274 18652 16304 18680
rect 15274 18649 15286 18652
rect 15228 18643 15286 18649
rect 16298 18640 16304 18652
rect 16356 18640 16362 18692
rect 16700 18683 16758 18689
rect 16700 18649 16712 18683
rect 16746 18680 16758 18683
rect 17862 18680 17868 18692
rect 16746 18652 17868 18680
rect 16746 18649 16758 18652
rect 16700 18643 16758 18649
rect 17862 18640 17868 18652
rect 17920 18640 17926 18692
rect 17494 18612 17500 18624
rect 15120 18584 17500 18612
rect 13541 18575 13599 18581
rect 17494 18572 17500 18584
rect 17552 18572 17558 18624
rect 17681 18615 17739 18621
rect 17681 18581 17693 18615
rect 17727 18612 17739 18615
rect 17972 18612 18000 18788
rect 18690 18708 18696 18760
rect 18748 18748 18754 18760
rect 18785 18751 18843 18757
rect 18785 18748 18797 18751
rect 18748 18720 18797 18748
rect 18748 18708 18754 18720
rect 18785 18717 18797 18720
rect 18831 18717 18843 18751
rect 19058 18748 19064 18760
rect 19019 18720 19064 18748
rect 18785 18711 18843 18717
rect 19058 18708 19064 18720
rect 19116 18708 19122 18760
rect 19337 18751 19395 18757
rect 19337 18717 19349 18751
rect 19383 18748 19395 18751
rect 19429 18751 19487 18757
rect 19429 18748 19441 18751
rect 19383 18720 19441 18748
rect 19383 18717 19395 18720
rect 19337 18711 19395 18717
rect 19429 18717 19441 18720
rect 19475 18748 19487 18751
rect 19886 18748 19892 18760
rect 19475 18720 19892 18748
rect 19475 18717 19487 18720
rect 19429 18711 19487 18717
rect 19886 18708 19892 18720
rect 19944 18708 19950 18760
rect 21174 18748 21180 18760
rect 20180 18720 21180 18748
rect 18322 18640 18328 18692
rect 18380 18680 18386 18692
rect 19518 18680 19524 18692
rect 18380 18652 19524 18680
rect 18380 18640 18386 18652
rect 19518 18640 19524 18652
rect 19576 18640 19582 18692
rect 19610 18640 19616 18692
rect 19668 18680 19674 18692
rect 20180 18689 20208 18720
rect 21174 18708 21180 18720
rect 21232 18748 21238 18760
rect 21913 18751 21971 18757
rect 21913 18748 21925 18751
rect 21232 18720 21925 18748
rect 21232 18708 21238 18720
rect 21913 18717 21925 18720
rect 21959 18717 21971 18751
rect 22646 18748 22652 18760
rect 22607 18720 22652 18748
rect 21913 18711 21971 18717
rect 22646 18708 22652 18720
rect 22704 18708 22710 18760
rect 22830 18748 22836 18760
rect 22791 18720 22836 18748
rect 22830 18708 22836 18720
rect 22888 18708 22894 18760
rect 20165 18683 20223 18689
rect 20165 18680 20177 18683
rect 19668 18652 20177 18680
rect 19668 18640 19674 18652
rect 20165 18649 20177 18652
rect 20211 18649 20223 18683
rect 20165 18643 20223 18649
rect 21668 18683 21726 18689
rect 21668 18649 21680 18683
rect 21714 18680 21726 18683
rect 21818 18680 21824 18692
rect 21714 18652 21824 18680
rect 21714 18649 21726 18652
rect 21668 18643 21726 18649
rect 21818 18640 21824 18652
rect 21876 18640 21882 18692
rect 17727 18584 18000 18612
rect 18141 18615 18199 18621
rect 17727 18581 17739 18584
rect 17681 18575 17739 18581
rect 18141 18581 18153 18615
rect 18187 18612 18199 18615
rect 18230 18612 18236 18624
rect 18187 18584 18236 18612
rect 18187 18581 18199 18584
rect 18141 18575 18199 18581
rect 18230 18572 18236 18584
rect 18288 18572 18294 18624
rect 18966 18572 18972 18624
rect 19024 18612 19030 18624
rect 21266 18612 21272 18624
rect 19024 18584 21272 18612
rect 19024 18572 19030 18584
rect 21266 18572 21272 18584
rect 21324 18572 21330 18624
rect 22002 18612 22008 18624
rect 21963 18584 22008 18612
rect 22002 18572 22008 18584
rect 22060 18572 22066 18624
rect 1104 18522 23460 18544
rect 1104 18470 6548 18522
rect 6600 18470 6612 18522
rect 6664 18470 6676 18522
rect 6728 18470 6740 18522
rect 6792 18470 6804 18522
rect 6856 18470 12146 18522
rect 12198 18470 12210 18522
rect 12262 18470 12274 18522
rect 12326 18470 12338 18522
rect 12390 18470 12402 18522
rect 12454 18470 17744 18522
rect 17796 18470 17808 18522
rect 17860 18470 17872 18522
rect 17924 18470 17936 18522
rect 17988 18470 18000 18522
rect 18052 18470 23460 18522
rect 1104 18448 23460 18470
rect 1670 18408 1676 18420
rect 1631 18380 1676 18408
rect 1670 18368 1676 18380
rect 1728 18368 1734 18420
rect 2222 18368 2228 18420
rect 2280 18408 2286 18420
rect 2280 18380 3280 18408
rect 2280 18368 2286 18380
rect 1578 18300 1584 18352
rect 1636 18340 1642 18352
rect 3252 18340 3280 18380
rect 4706 18368 4712 18420
rect 4764 18408 4770 18420
rect 4893 18411 4951 18417
rect 4893 18408 4905 18411
rect 4764 18380 4905 18408
rect 4764 18368 4770 18380
rect 4893 18377 4905 18380
rect 4939 18377 4951 18411
rect 4893 18371 4951 18377
rect 5721 18411 5779 18417
rect 5721 18377 5733 18411
rect 5767 18408 5779 18411
rect 5994 18408 6000 18420
rect 5767 18380 6000 18408
rect 5767 18377 5779 18380
rect 5721 18371 5779 18377
rect 5994 18368 6000 18380
rect 6052 18368 6058 18420
rect 9407 18411 9465 18417
rect 9407 18408 9419 18411
rect 6196 18380 9419 18408
rect 3758 18343 3816 18349
rect 3758 18340 3770 18343
rect 1636 18312 3188 18340
rect 3252 18312 3770 18340
rect 1636 18300 1642 18312
rect 1489 18275 1547 18281
rect 1489 18241 1501 18275
rect 1535 18241 1547 18275
rect 1762 18272 1768 18284
rect 1723 18244 1768 18272
rect 1489 18235 1547 18241
rect 1504 18204 1532 18235
rect 1762 18232 1768 18244
rect 1820 18232 1826 18284
rect 2056 18281 2084 18312
rect 2314 18281 2320 18284
rect 2041 18275 2099 18281
rect 2041 18241 2053 18275
rect 2087 18241 2099 18275
rect 2308 18272 2320 18281
rect 2275 18244 2320 18272
rect 2041 18235 2099 18241
rect 2308 18235 2320 18244
rect 2314 18232 2320 18235
rect 2372 18232 2378 18284
rect 3160 18272 3188 18312
rect 3758 18309 3770 18312
rect 3804 18309 3816 18343
rect 3758 18303 3816 18309
rect 5353 18343 5411 18349
rect 5353 18309 5365 18343
rect 5399 18340 5411 18343
rect 6086 18340 6092 18352
rect 5399 18312 6092 18340
rect 5399 18309 5411 18312
rect 5353 18303 5411 18309
rect 6086 18300 6092 18312
rect 6144 18300 6150 18352
rect 6196 18349 6224 18380
rect 6181 18343 6239 18349
rect 6181 18309 6193 18343
rect 6227 18309 6239 18343
rect 6181 18303 6239 18309
rect 7098 18300 7104 18352
rect 7156 18340 7162 18352
rect 7530 18343 7588 18349
rect 7530 18340 7542 18343
rect 7156 18312 7542 18340
rect 7156 18300 7162 18312
rect 7530 18309 7542 18312
rect 7576 18309 7588 18343
rect 7530 18303 7588 18309
rect 8662 18300 8668 18352
rect 8720 18340 8726 18352
rect 8757 18343 8815 18349
rect 8757 18340 8769 18343
rect 8720 18312 8769 18340
rect 8720 18300 8726 18312
rect 8757 18309 8769 18312
rect 8803 18309 8815 18343
rect 8757 18303 8815 18309
rect 3513 18275 3571 18281
rect 3513 18272 3525 18275
rect 3160 18244 3525 18272
rect 3513 18241 3525 18244
rect 3559 18241 3571 18275
rect 3513 18235 3571 18241
rect 5997 18275 6055 18281
rect 5997 18241 6009 18275
rect 6043 18272 6055 18275
rect 7006 18272 7012 18284
rect 6043 18244 6868 18272
rect 6967 18244 7012 18272
rect 6043 18241 6055 18244
rect 5997 18235 6055 18241
rect 1504 18176 2084 18204
rect 1302 18096 1308 18148
rect 1360 18136 1366 18148
rect 1949 18139 2007 18145
rect 1949 18136 1961 18139
rect 1360 18108 1961 18136
rect 1360 18096 1366 18108
rect 1949 18105 1961 18108
rect 1995 18105 2007 18139
rect 1949 18099 2007 18105
rect 2056 18068 2084 18176
rect 4614 18164 4620 18216
rect 4672 18204 4678 18216
rect 5077 18207 5135 18213
rect 5077 18204 5089 18207
rect 4672 18176 5089 18204
rect 4672 18164 4678 18176
rect 5077 18173 5089 18176
rect 5123 18173 5135 18207
rect 5077 18167 5135 18173
rect 5261 18207 5319 18213
rect 5261 18173 5273 18207
rect 5307 18204 5319 18207
rect 6270 18204 6276 18216
rect 5307 18176 6276 18204
rect 5307 18173 5319 18176
rect 5261 18167 5319 18173
rect 6270 18164 6276 18176
rect 6328 18164 6334 18216
rect 6840 18204 6868 18244
rect 7006 18232 7012 18244
rect 7064 18232 7070 18284
rect 7285 18275 7343 18281
rect 7285 18241 7297 18275
rect 7331 18272 7343 18275
rect 7374 18272 7380 18284
rect 7331 18244 7380 18272
rect 7331 18241 7343 18244
rect 7285 18235 7343 18241
rect 7374 18232 7380 18244
rect 7432 18232 7438 18284
rect 9048 18272 9076 18380
rect 9407 18377 9419 18380
rect 9453 18377 9465 18411
rect 9407 18371 9465 18377
rect 10042 18368 10048 18420
rect 10100 18408 10106 18420
rect 10873 18411 10931 18417
rect 10873 18408 10885 18411
rect 10100 18380 10885 18408
rect 10100 18368 10106 18380
rect 10873 18377 10885 18380
rect 10919 18377 10931 18411
rect 10873 18371 10931 18377
rect 11517 18411 11575 18417
rect 11517 18377 11529 18411
rect 11563 18408 11575 18411
rect 11698 18408 11704 18420
rect 11563 18380 11704 18408
rect 11563 18377 11575 18380
rect 11517 18371 11575 18377
rect 11698 18368 11704 18380
rect 11756 18368 11762 18420
rect 12802 18408 12808 18420
rect 12763 18380 12808 18408
rect 12802 18368 12808 18380
rect 12860 18368 12866 18420
rect 14458 18368 14464 18420
rect 14516 18408 14522 18420
rect 14553 18411 14611 18417
rect 14553 18408 14565 18411
rect 14516 18380 14565 18408
rect 14516 18368 14522 18380
rect 14553 18377 14565 18380
rect 14599 18377 14611 18411
rect 16669 18411 16727 18417
rect 16669 18408 16681 18411
rect 14553 18371 14611 18377
rect 15028 18380 16681 18408
rect 13354 18300 13360 18352
rect 13412 18340 13418 18352
rect 15028 18340 15056 18380
rect 16669 18377 16681 18380
rect 16715 18377 16727 18411
rect 17034 18408 17040 18420
rect 16995 18380 17040 18408
rect 16669 18371 16727 18377
rect 17034 18368 17040 18380
rect 17092 18368 17098 18420
rect 17126 18368 17132 18420
rect 17184 18408 17190 18420
rect 18233 18411 18291 18417
rect 18233 18408 18245 18411
rect 17184 18380 18245 18408
rect 17184 18368 17190 18380
rect 18233 18377 18245 18380
rect 18279 18408 18291 18411
rect 18506 18408 18512 18420
rect 18279 18380 18512 18408
rect 18279 18377 18291 18380
rect 18233 18371 18291 18377
rect 18506 18368 18512 18380
rect 18564 18368 18570 18420
rect 18601 18411 18659 18417
rect 18601 18377 18613 18411
rect 18647 18377 18659 18411
rect 18601 18371 18659 18377
rect 19153 18411 19211 18417
rect 19153 18377 19165 18411
rect 19199 18408 19211 18411
rect 19242 18408 19248 18420
rect 19199 18380 19248 18408
rect 19199 18377 19211 18380
rect 19153 18371 19211 18377
rect 15470 18340 15476 18352
rect 13412 18312 14320 18340
rect 13412 18300 13418 18312
rect 10962 18272 10968 18284
rect 9048 18244 10968 18272
rect 10962 18232 10968 18244
rect 11020 18232 11026 18284
rect 11164 18281 11293 18296
rect 11149 18276 11293 18281
rect 11149 18275 11376 18276
rect 11149 18241 11161 18275
rect 11195 18272 11376 18275
rect 11195 18268 11468 18272
rect 11195 18241 11207 18268
rect 11265 18248 11468 18268
rect 11348 18244 11468 18248
rect 11149 18235 11207 18241
rect 7098 18204 7104 18216
rect 6840 18176 7104 18204
rect 7098 18164 7104 18176
rect 7156 18164 7162 18216
rect 8941 18207 8999 18213
rect 8941 18173 8953 18207
rect 8987 18204 8999 18207
rect 9122 18204 9128 18216
rect 8987 18176 9128 18204
rect 8987 18173 8999 18176
rect 8941 18167 8999 18173
rect 9122 18164 9128 18176
rect 9180 18164 9186 18216
rect 9404 18207 9462 18213
rect 9404 18173 9416 18207
rect 9450 18204 9462 18207
rect 9490 18204 9496 18216
rect 9450 18176 9496 18204
rect 9450 18173 9462 18176
rect 9404 18167 9462 18173
rect 9490 18164 9496 18176
rect 9548 18164 9554 18216
rect 9677 18207 9735 18213
rect 9677 18173 9689 18207
rect 9723 18204 9735 18207
rect 9766 18204 9772 18216
rect 9723 18176 9772 18204
rect 9723 18173 9735 18176
rect 9677 18167 9735 18173
rect 9766 18164 9772 18176
rect 9824 18164 9830 18216
rect 4522 18096 4528 18148
rect 4580 18136 4586 18148
rect 10778 18136 10784 18148
rect 4580 18108 6500 18136
rect 10739 18108 10784 18136
rect 4580 18096 4586 18108
rect 3234 18068 3240 18080
rect 2056 18040 3240 18068
rect 3234 18028 3240 18040
rect 3292 18028 3298 18080
rect 3421 18071 3479 18077
rect 3421 18037 3433 18071
rect 3467 18068 3479 18071
rect 4430 18068 4436 18080
rect 3467 18040 4436 18068
rect 3467 18037 3479 18040
rect 3421 18031 3479 18037
rect 4430 18028 4436 18040
rect 4488 18028 4494 18080
rect 6362 18068 6368 18080
rect 6323 18040 6368 18068
rect 6362 18028 6368 18040
rect 6420 18028 6426 18080
rect 6472 18068 6500 18108
rect 10778 18096 10784 18108
rect 10836 18096 10842 18148
rect 11238 18096 11244 18148
rect 11296 18096 11302 18148
rect 11440 18136 11468 18244
rect 11698 18232 11704 18284
rect 11756 18272 11762 18284
rect 11885 18275 11943 18281
rect 11885 18272 11897 18275
rect 11756 18244 11897 18272
rect 11756 18232 11762 18244
rect 11885 18241 11897 18244
rect 11931 18241 11943 18275
rect 11885 18235 11943 18241
rect 11974 18232 11980 18284
rect 12032 18272 12038 18284
rect 12894 18272 12900 18284
rect 12032 18244 12077 18272
rect 12855 18244 12900 18272
rect 12032 18232 12038 18244
rect 12894 18232 12900 18244
rect 12952 18232 12958 18284
rect 13998 18272 14004 18284
rect 13959 18244 14004 18272
rect 13998 18232 14004 18244
rect 14056 18232 14062 18284
rect 11514 18164 11520 18216
rect 11572 18204 11578 18216
rect 12069 18207 12127 18213
rect 12069 18204 12081 18207
rect 11572 18176 12081 18204
rect 11572 18164 11578 18176
rect 12069 18173 12081 18176
rect 12115 18173 12127 18207
rect 12069 18167 12127 18173
rect 12713 18207 12771 18213
rect 12713 18173 12725 18207
rect 12759 18204 12771 18207
rect 13078 18204 13084 18216
rect 12759 18176 13084 18204
rect 12759 18173 12771 18176
rect 12713 18167 12771 18173
rect 13078 18164 13084 18176
rect 13136 18164 13142 18216
rect 13262 18164 13268 18216
rect 13320 18204 13326 18216
rect 14292 18213 14320 18312
rect 14476 18312 15056 18340
rect 15120 18312 15476 18340
rect 14476 18281 14504 18312
rect 15120 18281 15148 18312
rect 15470 18300 15476 18312
rect 15528 18300 15534 18352
rect 18141 18343 18199 18349
rect 18141 18340 18153 18343
rect 16776 18312 18153 18340
rect 14461 18275 14519 18281
rect 14461 18241 14473 18275
rect 14507 18241 14519 18275
rect 14461 18235 14519 18241
rect 15105 18275 15163 18281
rect 15105 18241 15117 18275
rect 15151 18241 15163 18275
rect 15105 18235 15163 18241
rect 15372 18275 15430 18281
rect 15372 18241 15384 18275
rect 15418 18272 15430 18275
rect 16776 18272 16804 18312
rect 18141 18309 18153 18312
rect 18187 18309 18199 18343
rect 18616 18340 18644 18371
rect 19242 18368 19248 18380
rect 19300 18408 19306 18420
rect 20898 18408 20904 18420
rect 19300 18380 20904 18408
rect 19300 18368 19306 18380
rect 20898 18368 20904 18380
rect 20956 18368 20962 18420
rect 21542 18408 21548 18420
rect 21503 18380 21548 18408
rect 21542 18368 21548 18380
rect 21600 18368 21606 18420
rect 22281 18411 22339 18417
rect 22281 18377 22293 18411
rect 22327 18408 22339 18411
rect 22462 18408 22468 18420
rect 22327 18380 22468 18408
rect 22327 18377 22339 18380
rect 22281 18371 22339 18377
rect 19426 18340 19432 18352
rect 18616 18312 19432 18340
rect 18141 18303 18199 18309
rect 19426 18300 19432 18312
rect 19484 18300 19490 18352
rect 19880 18343 19938 18349
rect 19880 18309 19892 18343
rect 19926 18340 19938 18343
rect 20254 18340 20260 18352
rect 19926 18312 20260 18340
rect 19926 18309 19938 18312
rect 19880 18303 19938 18309
rect 20254 18300 20260 18312
rect 20312 18300 20318 18352
rect 20438 18300 20444 18352
rect 20496 18340 20502 18352
rect 22189 18343 22247 18349
rect 22189 18340 22201 18343
rect 20496 18312 22201 18340
rect 20496 18300 20502 18312
rect 22189 18309 22201 18312
rect 22235 18309 22247 18343
rect 22189 18303 22247 18309
rect 17497 18275 17555 18281
rect 17497 18272 17509 18275
rect 15418 18244 16804 18272
rect 17144 18244 17509 18272
rect 15418 18241 15430 18244
rect 15372 18235 15430 18241
rect 17144 18216 17172 18244
rect 17497 18241 17509 18244
rect 17543 18241 17555 18275
rect 17497 18235 17555 18241
rect 18417 18275 18475 18281
rect 18417 18241 18429 18275
rect 18463 18272 18475 18275
rect 18506 18272 18512 18284
rect 18463 18244 18512 18272
rect 18463 18241 18475 18244
rect 18417 18235 18475 18241
rect 18506 18232 18512 18244
rect 18564 18232 18570 18284
rect 19702 18272 19708 18284
rect 18708 18244 19708 18272
rect 14277 18207 14335 18213
rect 13320 18176 13860 18204
rect 13320 18164 13326 18176
rect 12437 18139 12495 18145
rect 12437 18136 12449 18139
rect 11440 18108 12449 18136
rect 12437 18105 12449 18108
rect 12483 18136 12495 18139
rect 13832 18136 13860 18176
rect 14277 18173 14289 18207
rect 14323 18173 14335 18207
rect 17126 18204 17132 18216
rect 17087 18176 17132 18204
rect 14277 18167 14335 18173
rect 17126 18164 17132 18176
rect 17184 18164 17190 18216
rect 17218 18164 17224 18216
rect 17276 18204 17282 18216
rect 17276 18176 17321 18204
rect 17276 18164 17282 18176
rect 17678 18164 17684 18216
rect 17736 18204 17742 18216
rect 18708 18204 18736 18244
rect 19702 18232 19708 18244
rect 19760 18232 19766 18284
rect 21266 18272 21272 18284
rect 21227 18244 21272 18272
rect 21266 18232 21272 18244
rect 21324 18232 21330 18284
rect 21361 18275 21419 18281
rect 21361 18241 21373 18275
rect 21407 18272 21419 18275
rect 21450 18272 21456 18284
rect 21407 18244 21456 18272
rect 21407 18241 21419 18244
rect 21361 18235 21419 18241
rect 21450 18232 21456 18244
rect 21508 18232 21514 18284
rect 17736 18176 18736 18204
rect 18877 18207 18935 18213
rect 17736 18164 17742 18176
rect 18877 18173 18889 18207
rect 18923 18173 18935 18207
rect 19058 18204 19064 18216
rect 19019 18176 19064 18204
rect 18877 18167 18935 18173
rect 16485 18139 16543 18145
rect 12483 18108 13768 18136
rect 13832 18108 15056 18136
rect 12483 18105 12495 18108
rect 12437 18099 12495 18105
rect 8202 18068 8208 18080
rect 6472 18040 8208 18068
rect 8202 18028 8208 18040
rect 8260 18028 8266 18080
rect 8570 18028 8576 18080
rect 8628 18068 8634 18080
rect 8665 18071 8723 18077
rect 8665 18068 8677 18071
rect 8628 18040 8677 18068
rect 8628 18028 8634 18040
rect 8665 18037 8677 18040
rect 8711 18037 8723 18071
rect 11265 18068 11293 18096
rect 11333 18071 11391 18077
rect 11333 18068 11345 18071
rect 11265 18040 11345 18068
rect 8665 18031 8723 18037
rect 11333 18037 11345 18040
rect 11379 18037 11391 18071
rect 13262 18068 13268 18080
rect 13223 18040 13268 18068
rect 11333 18031 11391 18037
rect 13262 18028 13268 18040
rect 13320 18028 13326 18080
rect 13357 18071 13415 18077
rect 13357 18037 13369 18071
rect 13403 18068 13415 18071
rect 13538 18068 13544 18080
rect 13403 18040 13544 18068
rect 13403 18037 13415 18040
rect 13357 18031 13415 18037
rect 13538 18028 13544 18040
rect 13596 18028 13602 18080
rect 13740 18068 13768 18108
rect 14182 18068 14188 18080
rect 13740 18040 14188 18068
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 14826 18028 14832 18080
rect 14884 18068 14890 18080
rect 14921 18071 14979 18077
rect 14921 18068 14933 18071
rect 14884 18040 14933 18068
rect 14884 18028 14890 18040
rect 14921 18037 14933 18040
rect 14967 18037 14979 18071
rect 15028 18068 15056 18108
rect 16485 18105 16497 18139
rect 16531 18136 16543 18139
rect 17034 18136 17040 18148
rect 16531 18108 17040 18136
rect 16531 18105 16543 18108
rect 16485 18099 16543 18105
rect 17034 18096 17040 18108
rect 17092 18096 17098 18148
rect 18598 18068 18604 18080
rect 15028 18040 18604 18068
rect 14921 18031 14979 18037
rect 18598 18028 18604 18040
rect 18656 18028 18662 18080
rect 18892 18068 18920 18167
rect 19058 18164 19064 18176
rect 19116 18164 19122 18216
rect 19426 18164 19432 18216
rect 19484 18204 19490 18216
rect 19610 18204 19616 18216
rect 19484 18176 19616 18204
rect 19484 18164 19490 18176
rect 19610 18164 19616 18176
rect 19668 18164 19674 18216
rect 20993 18139 21051 18145
rect 20993 18105 21005 18139
rect 21039 18136 21051 18139
rect 22296 18136 22324 18371
rect 22462 18368 22468 18380
rect 22520 18368 22526 18420
rect 22741 18411 22799 18417
rect 22741 18377 22753 18411
rect 22787 18408 22799 18411
rect 22922 18408 22928 18420
rect 22787 18380 22928 18408
rect 22787 18377 22799 18380
rect 22741 18371 22799 18377
rect 22922 18368 22928 18380
rect 22980 18368 22986 18420
rect 22833 18275 22891 18281
rect 22833 18241 22845 18275
rect 22879 18272 22891 18275
rect 22879 18244 22913 18272
rect 22879 18241 22891 18244
rect 22833 18235 22891 18241
rect 22465 18207 22523 18213
rect 22465 18173 22477 18207
rect 22511 18204 22523 18207
rect 22848 18204 22876 18235
rect 22922 18204 22928 18216
rect 22511 18176 22928 18204
rect 22511 18173 22523 18176
rect 22465 18167 22523 18173
rect 22922 18164 22928 18176
rect 22980 18164 22986 18216
rect 21039 18108 22324 18136
rect 21039 18105 21051 18108
rect 20993 18099 21051 18105
rect 19150 18068 19156 18080
rect 18892 18040 19156 18068
rect 19150 18028 19156 18040
rect 19208 18028 19214 18080
rect 19518 18068 19524 18080
rect 19479 18040 19524 18068
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 19610 18028 19616 18080
rect 19668 18068 19674 18080
rect 20346 18068 20352 18080
rect 19668 18040 20352 18068
rect 19668 18028 19674 18040
rect 20346 18028 20352 18040
rect 20404 18068 20410 18080
rect 21085 18071 21143 18077
rect 21085 18068 21097 18071
rect 20404 18040 21097 18068
rect 20404 18028 20410 18040
rect 21085 18037 21097 18040
rect 21131 18037 21143 18071
rect 21085 18031 21143 18037
rect 21266 18028 21272 18080
rect 21324 18068 21330 18080
rect 21821 18071 21879 18077
rect 21821 18068 21833 18071
rect 21324 18040 21833 18068
rect 21324 18028 21330 18040
rect 21821 18037 21833 18040
rect 21867 18037 21879 18071
rect 23014 18068 23020 18080
rect 22975 18040 23020 18068
rect 21821 18031 21879 18037
rect 23014 18028 23020 18040
rect 23072 18028 23078 18080
rect 1104 17978 23460 18000
rect 1104 17926 3749 17978
rect 3801 17926 3813 17978
rect 3865 17926 3877 17978
rect 3929 17926 3941 17978
rect 3993 17926 4005 17978
rect 4057 17926 9347 17978
rect 9399 17926 9411 17978
rect 9463 17926 9475 17978
rect 9527 17926 9539 17978
rect 9591 17926 9603 17978
rect 9655 17926 14945 17978
rect 14997 17926 15009 17978
rect 15061 17926 15073 17978
rect 15125 17926 15137 17978
rect 15189 17926 15201 17978
rect 15253 17926 20543 17978
rect 20595 17926 20607 17978
rect 20659 17926 20671 17978
rect 20723 17926 20735 17978
rect 20787 17926 20799 17978
rect 20851 17926 23460 17978
rect 1104 17904 23460 17926
rect 1673 17867 1731 17873
rect 1673 17833 1685 17867
rect 1719 17864 1731 17867
rect 2498 17864 2504 17876
rect 1719 17836 2504 17864
rect 1719 17833 1731 17836
rect 1673 17827 1731 17833
rect 2498 17824 2504 17836
rect 2556 17824 2562 17876
rect 3145 17867 3203 17873
rect 3145 17833 3157 17867
rect 3191 17864 3203 17867
rect 3602 17864 3608 17876
rect 3191 17836 3608 17864
rect 3191 17833 3203 17836
rect 3145 17827 3203 17833
rect 3602 17824 3608 17836
rect 3660 17824 3666 17876
rect 3973 17867 4031 17873
rect 3973 17833 3985 17867
rect 4019 17864 4031 17867
rect 5258 17864 5264 17876
rect 4019 17836 5264 17864
rect 4019 17833 4031 17836
rect 3973 17827 4031 17833
rect 5258 17824 5264 17836
rect 5316 17824 5322 17876
rect 6454 17864 6460 17876
rect 6415 17836 6460 17864
rect 6454 17824 6460 17836
rect 6512 17824 6518 17876
rect 6733 17867 6791 17873
rect 6733 17833 6745 17867
rect 6779 17864 6791 17867
rect 6914 17864 6920 17876
rect 6779 17836 6920 17864
rect 6779 17833 6791 17836
rect 6733 17827 6791 17833
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 7374 17824 7380 17876
rect 7432 17864 7438 17876
rect 11425 17867 11483 17873
rect 7432 17836 9168 17864
rect 7432 17824 7438 17836
rect 2958 17756 2964 17808
rect 3016 17796 3022 17808
rect 3329 17799 3387 17805
rect 3329 17796 3341 17799
rect 3016 17768 3341 17796
rect 3016 17756 3022 17768
rect 3329 17765 3341 17768
rect 3375 17796 3387 17799
rect 4522 17796 4528 17808
rect 3375 17768 4528 17796
rect 3375 17765 3387 17768
rect 3329 17759 3387 17765
rect 4522 17756 4528 17768
rect 4580 17756 4586 17808
rect 8662 17796 8668 17808
rect 8623 17768 8668 17796
rect 8662 17756 8668 17768
rect 8720 17796 8726 17808
rect 9030 17796 9036 17808
rect 8720 17768 9036 17796
rect 8720 17756 8726 17768
rect 9030 17756 9036 17768
rect 9088 17756 9094 17808
rect 1578 17688 1584 17740
rect 1636 17728 1642 17740
rect 1765 17731 1823 17737
rect 1765 17728 1777 17731
rect 1636 17700 1777 17728
rect 1636 17688 1642 17700
rect 1765 17697 1777 17700
rect 1811 17697 1823 17731
rect 1765 17691 1823 17697
rect 4080 17700 5212 17728
rect 2038 17669 2044 17672
rect 1489 17663 1547 17669
rect 1489 17629 1501 17663
rect 1535 17629 1547 17663
rect 2032 17660 2044 17669
rect 1999 17632 2044 17660
rect 1489 17623 1547 17629
rect 2032 17623 2044 17632
rect 1504 17592 1532 17623
rect 2038 17620 2044 17623
rect 2096 17620 2102 17672
rect 3418 17660 3424 17672
rect 3379 17632 3424 17660
rect 3418 17620 3424 17632
rect 3476 17620 3482 17672
rect 3602 17620 3608 17672
rect 3660 17660 3666 17672
rect 4080 17669 4108 17700
rect 4540 17672 4568 17700
rect 3789 17663 3847 17669
rect 3789 17660 3801 17663
rect 3660 17632 3801 17660
rect 3660 17620 3666 17632
rect 3789 17629 3801 17632
rect 3835 17629 3847 17663
rect 3789 17623 3847 17629
rect 4065 17663 4123 17669
rect 4065 17629 4077 17663
rect 4111 17629 4123 17663
rect 4065 17623 4123 17629
rect 4522 17620 4528 17672
rect 4580 17620 4586 17672
rect 5077 17663 5135 17669
rect 5077 17660 5089 17663
rect 4816 17632 5089 17660
rect 4816 17604 4844 17632
rect 5077 17629 5089 17632
rect 5123 17629 5135 17663
rect 5184 17660 5212 17700
rect 8018 17688 8024 17740
rect 8076 17728 8082 17740
rect 8110 17731 8168 17737
rect 8110 17728 8122 17731
rect 8076 17700 8122 17728
rect 8076 17688 8082 17700
rect 8110 17697 8122 17700
rect 8156 17697 8168 17731
rect 9140 17728 9168 17836
rect 11425 17833 11437 17867
rect 11471 17864 11483 17867
rect 12710 17864 12716 17876
rect 11471 17836 12716 17864
rect 11471 17833 11483 17836
rect 11425 17827 11483 17833
rect 12710 17824 12716 17836
rect 12768 17824 12774 17876
rect 12894 17864 12900 17876
rect 12855 17836 12900 17864
rect 12894 17824 12900 17836
rect 12952 17824 12958 17876
rect 14090 17864 14096 17876
rect 14051 17836 14096 17864
rect 14090 17824 14096 17836
rect 14148 17824 14154 17876
rect 14182 17824 14188 17876
rect 14240 17864 14246 17876
rect 17310 17864 17316 17876
rect 14240 17836 16416 17864
rect 17271 17836 17316 17864
rect 14240 17824 14246 17836
rect 12618 17756 12624 17808
rect 12676 17796 12682 17808
rect 12989 17799 13047 17805
rect 12989 17796 13001 17799
rect 12676 17768 13001 17796
rect 12676 17756 12682 17768
rect 12989 17765 13001 17768
rect 13035 17765 13047 17799
rect 12989 17759 13047 17765
rect 13354 17756 13360 17808
rect 13412 17796 13418 17808
rect 13412 17768 13584 17796
rect 13412 17756 13418 17768
rect 9677 17731 9735 17737
rect 9677 17728 9689 17731
rect 9140 17726 9536 17728
rect 9600 17726 9689 17728
rect 9140 17700 9689 17726
rect 9508 17698 9628 17700
rect 8110 17691 8168 17697
rect 9677 17697 9689 17700
rect 9723 17728 9735 17731
rect 10045 17731 10103 17737
rect 10045 17728 10057 17731
rect 9723 17700 10057 17728
rect 9723 17697 9735 17700
rect 9677 17691 9735 17697
rect 10045 17697 10057 17700
rect 10091 17697 10103 17731
rect 10045 17691 10103 17697
rect 6546 17660 6552 17672
rect 5184 17632 6552 17660
rect 5077 17623 5135 17629
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 7558 17660 7564 17672
rect 6748 17632 7564 17660
rect 3142 17592 3148 17604
rect 1504 17564 3148 17592
rect 3142 17552 3148 17564
rect 3200 17552 3206 17604
rect 4338 17592 4344 17604
rect 3620 17564 4344 17592
rect 3620 17533 3648 17564
rect 4338 17552 4344 17564
rect 4396 17552 4402 17604
rect 4798 17592 4804 17604
rect 4759 17564 4804 17592
rect 4798 17552 4804 17564
rect 4856 17552 4862 17604
rect 5344 17595 5402 17601
rect 5344 17561 5356 17595
rect 5390 17592 5402 17595
rect 6362 17592 6368 17604
rect 5390 17564 6368 17592
rect 5390 17561 5402 17564
rect 5344 17555 5402 17561
rect 6362 17552 6368 17564
rect 6420 17552 6426 17604
rect 3605 17527 3663 17533
rect 3605 17493 3617 17527
rect 3651 17493 3663 17527
rect 3605 17487 3663 17493
rect 4890 17484 4896 17536
rect 4948 17524 4954 17536
rect 6748 17524 6776 17632
rect 7558 17620 7564 17632
rect 7616 17620 7622 17672
rect 7834 17660 7840 17672
rect 7795 17632 7840 17660
rect 7834 17620 7840 17632
rect 7892 17620 7898 17672
rect 8573 17663 8631 17669
rect 8573 17629 8585 17663
rect 8619 17656 8631 17663
rect 9214 17660 9220 17672
rect 8772 17656 9220 17660
rect 8619 17632 9220 17656
rect 8619 17629 8800 17632
rect 8573 17628 8800 17629
rect 8573 17623 8631 17628
rect 9214 17620 9220 17632
rect 9272 17620 9278 17672
rect 10060 17660 10088 17691
rect 13262 17688 13268 17740
rect 13320 17728 13326 17740
rect 13556 17737 13584 17768
rect 14366 17756 14372 17808
rect 14424 17796 14430 17808
rect 14550 17796 14556 17808
rect 14424 17768 14556 17796
rect 14424 17756 14430 17768
rect 14550 17756 14556 17768
rect 14608 17756 14614 17808
rect 16301 17799 16359 17805
rect 16301 17796 16313 17799
rect 14752 17768 16313 17796
rect 13449 17731 13507 17737
rect 13449 17728 13461 17731
rect 13320 17700 13461 17728
rect 13320 17688 13326 17700
rect 13449 17697 13461 17700
rect 13495 17697 13507 17731
rect 13449 17691 13507 17697
rect 13541 17731 13599 17737
rect 13541 17697 13553 17731
rect 13587 17728 13599 17731
rect 14645 17731 14703 17737
rect 14645 17728 14657 17731
rect 13587 17700 14657 17728
rect 13587 17697 13599 17700
rect 13541 17691 13599 17697
rect 14645 17697 14657 17700
rect 14691 17697 14703 17731
rect 14645 17691 14703 17697
rect 11054 17660 11060 17672
rect 10060 17632 11060 17660
rect 11054 17620 11060 17632
rect 11112 17660 11118 17672
rect 11517 17663 11575 17669
rect 11517 17660 11529 17663
rect 11112 17632 11529 17660
rect 11112 17620 11118 17632
rect 11517 17629 11529 17632
rect 11563 17629 11575 17663
rect 11517 17623 11575 17629
rect 11784 17663 11842 17669
rect 11784 17629 11796 17663
rect 11830 17660 11842 17663
rect 12066 17660 12072 17672
rect 11830 17632 12072 17660
rect 11830 17629 11842 17632
rect 11784 17623 11842 17629
rect 12066 17620 12072 17632
rect 12124 17620 12130 17672
rect 14461 17663 14519 17669
rect 14461 17629 14473 17663
rect 14507 17660 14519 17663
rect 14752 17660 14780 17768
rect 16301 17765 16313 17768
rect 16347 17765 16359 17799
rect 16388 17796 16416 17836
rect 17310 17824 17316 17836
rect 17368 17824 17374 17876
rect 19242 17864 19248 17876
rect 17411 17836 18644 17864
rect 19203 17836 19248 17864
rect 17411 17796 17439 17836
rect 16388 17768 17439 17796
rect 17589 17799 17647 17805
rect 16301 17759 16359 17765
rect 17589 17765 17601 17799
rect 17635 17796 17647 17799
rect 17678 17796 17684 17808
rect 17635 17768 17684 17796
rect 17635 17765 17647 17768
rect 17589 17759 17647 17765
rect 17678 17756 17684 17768
rect 17736 17756 17742 17808
rect 18616 17796 18644 17836
rect 19242 17824 19248 17836
rect 19300 17824 19306 17876
rect 21174 17864 21180 17876
rect 19628 17836 21180 17864
rect 19334 17796 19340 17808
rect 18616 17768 19340 17796
rect 19334 17756 19340 17768
rect 19392 17756 19398 17808
rect 14826 17688 14832 17740
rect 14884 17688 14890 17740
rect 15470 17688 15476 17740
rect 15528 17728 15534 17740
rect 16025 17731 16083 17737
rect 16025 17728 16037 17731
rect 15528 17700 16037 17728
rect 15528 17688 15534 17700
rect 16025 17697 16037 17700
rect 16071 17697 16083 17731
rect 16206 17728 16212 17740
rect 16025 17691 16083 17697
rect 16132 17700 16212 17728
rect 14507 17632 14780 17660
rect 14844 17660 14872 17688
rect 15105 17663 15163 17669
rect 15105 17660 15117 17663
rect 14844 17632 15117 17660
rect 14507 17629 14519 17632
rect 14461 17623 14519 17629
rect 15105 17629 15117 17632
rect 15151 17629 15163 17663
rect 15105 17623 15163 17629
rect 15194 17620 15200 17672
rect 15252 17660 15258 17672
rect 16132 17660 16160 17700
rect 16206 17688 16212 17700
rect 16264 17728 16270 17740
rect 16853 17731 16911 17737
rect 16853 17728 16865 17731
rect 16264 17700 16865 17728
rect 16264 17688 16270 17700
rect 16853 17697 16865 17700
rect 16899 17728 16911 17731
rect 17218 17728 17224 17740
rect 16899 17700 17224 17728
rect 16899 17697 16911 17700
rect 16853 17691 16911 17697
rect 17218 17688 17224 17700
rect 17276 17688 17282 17740
rect 18874 17688 18880 17740
rect 18932 17728 18938 17740
rect 19628 17728 19656 17836
rect 21174 17824 21180 17836
rect 21232 17824 21238 17876
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 22833 17867 22891 17873
rect 22833 17864 22845 17867
rect 22152 17836 22845 17864
rect 22152 17824 22158 17836
rect 22833 17833 22845 17836
rect 22879 17833 22891 17867
rect 22833 17827 22891 17833
rect 20622 17756 20628 17808
rect 20680 17796 20686 17808
rect 21361 17799 21419 17805
rect 21361 17796 21373 17799
rect 20680 17768 21373 17796
rect 20680 17756 20686 17768
rect 21361 17765 21373 17768
rect 21407 17765 21419 17799
rect 21361 17759 21419 17765
rect 21450 17728 21456 17740
rect 18932 17700 19656 17728
rect 20640 17700 21456 17728
rect 18932 17688 18938 17700
rect 15252 17632 16160 17660
rect 15252 17620 15258 17632
rect 16482 17620 16488 17672
rect 16540 17660 16546 17672
rect 17129 17663 17187 17669
rect 17129 17660 17141 17663
rect 16540 17632 17141 17660
rect 16540 17620 16546 17632
rect 17129 17629 17141 17632
rect 17175 17629 17187 17663
rect 17129 17623 17187 17629
rect 17405 17663 17463 17669
rect 17405 17629 17417 17663
rect 17451 17629 17463 17663
rect 17405 17623 17463 17629
rect 17681 17663 17739 17669
rect 17681 17629 17693 17663
rect 17727 17660 17739 17663
rect 19426 17660 19432 17672
rect 17727 17632 19432 17660
rect 17727 17629 17739 17632
rect 17681 17623 17739 17629
rect 8941 17595 8999 17601
rect 8941 17561 8953 17595
rect 8987 17592 8999 17595
rect 9030 17592 9036 17604
rect 8987 17564 9036 17592
rect 8987 17561 8999 17564
rect 8941 17555 8999 17561
rect 9030 17552 9036 17564
rect 9088 17552 9094 17604
rect 10318 17601 10324 17604
rect 10312 17592 10324 17601
rect 10279 17564 10324 17592
rect 10312 17555 10324 17564
rect 10318 17552 10324 17555
rect 10376 17552 10382 17604
rect 13909 17595 13967 17601
rect 13909 17561 13921 17595
rect 13955 17592 13967 17595
rect 14826 17592 14832 17604
rect 13955 17564 14832 17592
rect 13955 17561 13967 17564
rect 13909 17555 13967 17561
rect 14826 17552 14832 17564
rect 14884 17592 14890 17604
rect 15289 17595 15347 17601
rect 15289 17592 15301 17595
rect 14884 17564 15301 17592
rect 14884 17552 14890 17564
rect 15289 17561 15301 17564
rect 15335 17561 15347 17595
rect 15289 17555 15347 17561
rect 16574 17552 16580 17604
rect 16632 17592 16638 17604
rect 16761 17595 16819 17601
rect 16761 17592 16773 17595
rect 16632 17564 16773 17592
rect 16632 17552 16638 17564
rect 16761 17561 16773 17564
rect 16807 17561 16819 17595
rect 16761 17555 16819 17561
rect 16942 17552 16948 17604
rect 17000 17592 17006 17604
rect 17420 17592 17448 17623
rect 18156 17604 18184 17632
rect 19426 17620 19432 17632
rect 19484 17660 19490 17672
rect 20640 17669 20668 17700
rect 21450 17688 21456 17700
rect 21508 17688 21514 17740
rect 20625 17663 20683 17669
rect 20625 17660 20637 17663
rect 19484 17632 20637 17660
rect 19484 17620 19490 17632
rect 20625 17629 20637 17632
rect 20671 17629 20683 17663
rect 20625 17623 20683 17629
rect 20714 17620 20720 17672
rect 20772 17660 20778 17672
rect 20772 17632 20817 17660
rect 20772 17620 20778 17632
rect 21542 17620 21548 17672
rect 21600 17660 21606 17672
rect 21709 17663 21767 17669
rect 21709 17660 21721 17663
rect 21600 17632 21721 17660
rect 21600 17620 21606 17632
rect 21709 17629 21721 17632
rect 21755 17629 21767 17663
rect 21709 17623 21767 17629
rect 23109 17663 23167 17669
rect 23109 17629 23121 17663
rect 23155 17660 23167 17663
rect 23290 17660 23296 17672
rect 23155 17632 23296 17660
rect 23155 17629 23167 17632
rect 23109 17623 23167 17629
rect 23290 17620 23296 17632
rect 23348 17620 23354 17672
rect 17000 17564 17448 17592
rect 17948 17595 18006 17601
rect 17000 17552 17006 17564
rect 17948 17561 17960 17595
rect 17994 17592 18006 17595
rect 17994 17564 18092 17592
rect 17994 17561 18006 17564
rect 17948 17555 18006 17561
rect 4948 17496 6776 17524
rect 8106 17527 8164 17533
rect 4948 17484 4954 17496
rect 8106 17493 8118 17527
rect 8152 17524 8164 17527
rect 8202 17524 8208 17536
rect 8152 17496 8208 17524
rect 8152 17493 8164 17496
rect 8106 17487 8164 17493
rect 8202 17484 8208 17496
rect 8260 17484 8266 17536
rect 8662 17484 8668 17536
rect 8720 17524 8726 17536
rect 10594 17524 10600 17536
rect 8720 17496 10600 17524
rect 8720 17484 8726 17496
rect 10594 17484 10600 17496
rect 10652 17484 10658 17536
rect 13354 17524 13360 17536
rect 13315 17496 13360 17524
rect 13354 17484 13360 17496
rect 13412 17484 13418 17536
rect 14550 17484 14556 17536
rect 14608 17524 14614 17536
rect 14608 17496 14653 17524
rect 14608 17484 14614 17496
rect 14734 17484 14740 17536
rect 14792 17524 14798 17536
rect 14921 17527 14979 17533
rect 14921 17524 14933 17527
rect 14792 17496 14933 17524
rect 14792 17484 14798 17496
rect 14921 17493 14933 17496
rect 14967 17493 14979 17527
rect 16666 17524 16672 17536
rect 16627 17496 16672 17524
rect 14921 17487 14979 17493
rect 16666 17484 16672 17496
rect 16724 17484 16730 17536
rect 18064 17524 18092 17564
rect 18138 17552 18144 17604
rect 18196 17552 18202 17604
rect 20380 17595 20438 17601
rect 20380 17561 20392 17595
rect 20426 17592 20438 17595
rect 20530 17592 20536 17604
rect 20426 17564 20536 17592
rect 20426 17561 20438 17564
rect 20380 17555 20438 17561
rect 20530 17552 20536 17564
rect 20588 17552 20594 17604
rect 18230 17524 18236 17536
rect 18064 17496 18236 17524
rect 18230 17484 18236 17496
rect 18288 17484 18294 17536
rect 19058 17524 19064 17536
rect 18971 17496 19064 17524
rect 19058 17484 19064 17496
rect 19116 17524 19122 17536
rect 20714 17524 20720 17536
rect 19116 17496 20720 17524
rect 19116 17484 19122 17496
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 22922 17484 22928 17536
rect 22980 17524 22986 17536
rect 22980 17496 23025 17524
rect 22980 17484 22986 17496
rect 1104 17434 23460 17456
rect 1104 17382 6548 17434
rect 6600 17382 6612 17434
rect 6664 17382 6676 17434
rect 6728 17382 6740 17434
rect 6792 17382 6804 17434
rect 6856 17382 12146 17434
rect 12198 17382 12210 17434
rect 12262 17382 12274 17434
rect 12326 17382 12338 17434
rect 12390 17382 12402 17434
rect 12454 17382 17744 17434
rect 17796 17382 17808 17434
rect 17860 17382 17872 17434
rect 17924 17382 17936 17434
rect 17988 17382 18000 17434
rect 18052 17382 23460 17434
rect 1104 17360 23460 17382
rect 1394 17280 1400 17332
rect 1452 17320 1458 17332
rect 1489 17323 1547 17329
rect 1489 17320 1501 17323
rect 1452 17292 1501 17320
rect 1452 17280 1458 17292
rect 1489 17289 1501 17292
rect 1535 17320 1547 17323
rect 3237 17323 3295 17329
rect 3237 17320 3249 17323
rect 1535 17292 3249 17320
rect 1535 17289 1547 17292
rect 1489 17283 1547 17289
rect 3237 17289 3249 17292
rect 3283 17289 3295 17323
rect 3237 17283 3295 17289
rect 3329 17323 3387 17329
rect 3329 17289 3341 17323
rect 3375 17320 3387 17323
rect 3510 17320 3516 17332
rect 3375 17292 3516 17320
rect 3375 17289 3387 17292
rect 3329 17283 3387 17289
rect 3510 17280 3516 17292
rect 3568 17280 3574 17332
rect 4154 17280 4160 17332
rect 4212 17320 4218 17332
rect 4525 17323 4583 17329
rect 4525 17320 4537 17323
rect 4212 17292 4537 17320
rect 4212 17280 4218 17292
rect 4525 17289 4537 17292
rect 4571 17289 4583 17323
rect 4525 17283 4583 17289
rect 4709 17323 4767 17329
rect 4709 17289 4721 17323
rect 4755 17320 4767 17323
rect 4982 17320 4988 17332
rect 4755 17292 4988 17320
rect 4755 17289 4767 17292
rect 4709 17283 4767 17289
rect 4982 17280 4988 17292
rect 5040 17280 5046 17332
rect 6270 17280 6276 17332
rect 6328 17320 6334 17332
rect 6365 17323 6423 17329
rect 6365 17320 6377 17323
rect 6328 17292 6377 17320
rect 6328 17280 6334 17292
rect 6365 17289 6377 17292
rect 6411 17289 6423 17323
rect 6365 17283 6423 17289
rect 7098 17280 7104 17332
rect 7156 17320 7162 17332
rect 8018 17320 8024 17332
rect 7156 17292 8024 17320
rect 7156 17280 7162 17292
rect 8018 17280 8024 17292
rect 8076 17320 8082 17332
rect 8202 17320 8208 17332
rect 8076 17292 8208 17320
rect 8076 17280 8082 17292
rect 8202 17280 8208 17292
rect 8260 17280 8266 17332
rect 8386 17280 8392 17332
rect 8444 17320 8450 17332
rect 8846 17320 8852 17332
rect 8444 17292 8708 17320
rect 8807 17292 8852 17320
rect 8444 17280 8450 17292
rect 1578 17212 1584 17264
rect 1636 17252 1642 17264
rect 4798 17252 4804 17264
rect 1636 17224 4804 17252
rect 1636 17212 1642 17224
rect 2590 17144 2596 17196
rect 2648 17193 2654 17196
rect 2884 17193 2912 17224
rect 4798 17212 4804 17224
rect 4856 17252 4862 17264
rect 4856 17224 4927 17252
rect 4856 17212 4862 17224
rect 2648 17184 2660 17193
rect 2869 17187 2927 17193
rect 2648 17156 2693 17184
rect 2648 17147 2660 17156
rect 2869 17153 2881 17187
rect 2915 17153 2927 17187
rect 2869 17147 2927 17153
rect 4157 17187 4215 17193
rect 4157 17153 4169 17187
rect 4203 17184 4215 17187
rect 4706 17184 4712 17196
rect 4203 17156 4712 17184
rect 4203 17153 4215 17156
rect 4157 17147 4215 17153
rect 2648 17144 2654 17147
rect 4706 17144 4712 17156
rect 4764 17144 4770 17196
rect 3142 17116 3148 17128
rect 3055 17088 3148 17116
rect 3142 17076 3148 17088
rect 3200 17116 3206 17128
rect 3878 17116 3884 17128
rect 3200 17088 3884 17116
rect 3200 17076 3206 17088
rect 3878 17076 3884 17088
rect 3936 17076 3942 17128
rect 4065 17119 4123 17125
rect 4065 17085 4077 17119
rect 4111 17116 4123 17119
rect 4430 17116 4436 17128
rect 4111 17088 4436 17116
rect 4111 17085 4123 17088
rect 4065 17079 4123 17085
rect 4430 17076 4436 17088
rect 4488 17076 4494 17128
rect 4801 17119 4859 17125
rect 4801 17085 4813 17119
rect 4847 17116 4859 17119
rect 4899 17116 4927 17224
rect 5902 17212 5908 17264
rect 5960 17252 5966 17264
rect 6638 17252 6644 17264
rect 5960 17224 6644 17252
rect 5960 17212 5966 17224
rect 6638 17212 6644 17224
rect 6696 17252 6702 17264
rect 6696 17224 6868 17252
rect 6696 17212 6702 17224
rect 5068 17187 5126 17193
rect 5068 17153 5080 17187
rect 5114 17184 5126 17187
rect 5626 17184 5632 17196
rect 5114 17156 5632 17184
rect 5114 17153 5126 17156
rect 5068 17147 5126 17153
rect 5626 17144 5632 17156
rect 5684 17144 5690 17196
rect 6730 17184 6736 17196
rect 6691 17156 6736 17184
rect 6730 17144 6736 17156
rect 6788 17144 6794 17196
rect 6840 17184 6868 17224
rect 7374 17212 7380 17264
rect 7432 17252 7438 17264
rect 8680 17252 8708 17292
rect 8846 17280 8852 17292
rect 8904 17280 8910 17332
rect 9674 17320 9680 17332
rect 9635 17292 9680 17320
rect 9674 17280 9680 17292
rect 9732 17280 9738 17332
rect 11514 17320 11520 17332
rect 11265 17292 11520 17320
rect 9217 17255 9275 17261
rect 9217 17252 9229 17255
rect 7432 17224 8616 17252
rect 8680 17224 9229 17252
rect 7432 17212 7438 17224
rect 6840 17156 6960 17184
rect 4847 17088 4927 17116
rect 4847 17085 4859 17088
rect 4801 17079 4859 17085
rect 6362 17076 6368 17128
rect 6420 17116 6426 17128
rect 6932 17125 6960 17156
rect 8294 17144 8300 17196
rect 8352 17193 8358 17196
rect 8588 17193 8616 17224
rect 9217 17221 9229 17224
rect 9263 17221 9275 17255
rect 9217 17215 9275 17221
rect 10812 17255 10870 17261
rect 10812 17221 10824 17255
rect 10858 17252 10870 17255
rect 11265 17252 11293 17292
rect 11514 17280 11520 17292
rect 11572 17280 11578 17332
rect 11606 17280 11612 17332
rect 11664 17320 11670 17332
rect 11664 17292 13308 17320
rect 11664 17280 11670 17292
rect 10858 17224 11293 17252
rect 11333 17255 11391 17261
rect 10858 17221 10870 17224
rect 10812 17215 10870 17221
rect 11333 17221 11345 17255
rect 11379 17252 11391 17255
rect 12244 17255 12302 17261
rect 11379 17224 11836 17252
rect 11379 17221 11391 17224
rect 11333 17215 11391 17221
rect 8352 17184 8364 17193
rect 8573 17187 8631 17193
rect 8352 17156 8397 17184
rect 8352 17147 8364 17156
rect 8573 17153 8585 17187
rect 8619 17153 8631 17187
rect 8573 17147 8631 17153
rect 8352 17144 8358 17147
rect 8846 17144 8852 17196
rect 8904 17184 8910 17196
rect 9122 17184 9128 17196
rect 8904 17156 9128 17184
rect 8904 17144 8910 17156
rect 9122 17144 9128 17156
rect 9180 17144 9186 17196
rect 11054 17184 11060 17196
rect 11015 17156 11060 17184
rect 11054 17144 11060 17156
rect 11112 17144 11118 17196
rect 11698 17184 11704 17196
rect 11659 17156 11704 17184
rect 11698 17144 11704 17156
rect 11756 17144 11762 17196
rect 11808 17184 11836 17224
rect 12244 17221 12256 17255
rect 12290 17252 12302 17255
rect 12986 17252 12992 17264
rect 12290 17224 12992 17252
rect 12290 17221 12302 17224
rect 12244 17215 12302 17221
rect 12986 17212 12992 17224
rect 13044 17212 13050 17264
rect 13280 17252 13308 17292
rect 13354 17280 13360 17332
rect 13412 17320 13418 17332
rect 13449 17323 13507 17329
rect 13449 17320 13461 17323
rect 13412 17292 13461 17320
rect 13412 17280 13418 17292
rect 13449 17289 13461 17292
rect 13495 17289 13507 17323
rect 13449 17283 13507 17289
rect 13909 17323 13967 17329
rect 13909 17289 13921 17323
rect 13955 17320 13967 17323
rect 13998 17320 14004 17332
rect 13955 17292 14004 17320
rect 13955 17289 13967 17292
rect 13909 17283 13967 17289
rect 13998 17280 14004 17292
rect 14056 17280 14062 17332
rect 14277 17323 14335 17329
rect 14277 17289 14289 17323
rect 14323 17320 14335 17323
rect 14550 17320 14556 17332
rect 14323 17292 14556 17320
rect 14323 17289 14335 17292
rect 14277 17283 14335 17289
rect 14550 17280 14556 17292
rect 14608 17280 14614 17332
rect 16485 17323 16543 17329
rect 14660 17292 15608 17320
rect 14660 17252 14688 17292
rect 15470 17252 15476 17264
rect 13280 17224 14688 17252
rect 15120 17224 15476 17252
rect 13814 17184 13820 17196
rect 11808 17156 13676 17184
rect 13775 17156 13820 17184
rect 6825 17119 6883 17125
rect 6825 17116 6837 17119
rect 6420 17088 6837 17116
rect 6420 17076 6426 17088
rect 6825 17085 6837 17088
rect 6871 17085 6883 17119
rect 6825 17079 6883 17085
rect 6917 17119 6975 17125
rect 6917 17085 6929 17119
rect 6963 17085 6975 17119
rect 6917 17079 6975 17085
rect 8662 17076 8668 17128
rect 8720 17116 8726 17128
rect 9309 17119 9367 17125
rect 9309 17116 9321 17119
rect 8720 17088 9321 17116
rect 8720 17076 8726 17088
rect 9309 17085 9321 17088
rect 9355 17085 9367 17119
rect 9309 17079 9367 17085
rect 9401 17119 9459 17125
rect 9401 17085 9413 17119
rect 9447 17085 9459 17119
rect 11072 17116 11100 17144
rect 11977 17119 12035 17125
rect 11977 17116 11989 17119
rect 11072 17088 11989 17116
rect 9401 17079 9459 17085
rect 11977 17085 11989 17088
rect 12023 17085 12035 17119
rect 13648 17116 13676 17156
rect 13814 17144 13820 17156
rect 13872 17144 13878 17196
rect 14366 17184 14372 17196
rect 13924 17156 14372 17184
rect 13924 17116 13952 17156
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 14642 17184 14648 17196
rect 14603 17156 14648 17184
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 15120 17193 15148 17224
rect 15470 17212 15476 17224
rect 15528 17212 15534 17264
rect 15580 17252 15608 17292
rect 16485 17289 16497 17323
rect 16531 17320 16543 17323
rect 17126 17320 17132 17332
rect 16531 17292 17132 17320
rect 16531 17289 16543 17292
rect 16485 17283 16543 17289
rect 17126 17280 17132 17292
rect 17184 17280 17190 17332
rect 17405 17323 17463 17329
rect 17405 17289 17417 17323
rect 17451 17320 17463 17323
rect 18690 17320 18696 17332
rect 17451 17292 18696 17320
rect 17451 17289 17463 17292
rect 17405 17283 17463 17289
rect 18690 17280 18696 17292
rect 18748 17320 18754 17332
rect 19245 17323 19303 17329
rect 19245 17320 19257 17323
rect 18748 17292 19257 17320
rect 18748 17280 18754 17292
rect 19245 17289 19257 17292
rect 19291 17289 19303 17323
rect 19245 17283 19303 17289
rect 19518 17280 19524 17332
rect 19576 17320 19582 17332
rect 20073 17323 20131 17329
rect 20073 17320 20085 17323
rect 19576 17292 20085 17320
rect 19576 17280 19582 17292
rect 20073 17289 20085 17292
rect 20119 17289 20131 17323
rect 20073 17283 20131 17289
rect 20809 17323 20867 17329
rect 20809 17289 20821 17323
rect 20855 17289 20867 17323
rect 20809 17283 20867 17289
rect 21177 17323 21235 17329
rect 21177 17289 21189 17323
rect 21223 17320 21235 17323
rect 21821 17323 21879 17329
rect 21821 17320 21833 17323
rect 21223 17292 21833 17320
rect 21223 17289 21235 17292
rect 21177 17283 21235 17289
rect 21821 17289 21833 17292
rect 21867 17289 21879 17323
rect 21821 17283 21879 17289
rect 16758 17252 16764 17264
rect 15580 17224 16764 17252
rect 16758 17212 16764 17224
rect 16816 17212 16822 17264
rect 18138 17212 18144 17264
rect 18196 17252 18202 17264
rect 18196 17224 18828 17252
rect 18196 17212 18202 17224
rect 15105 17187 15163 17193
rect 15105 17153 15117 17187
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 15194 17144 15200 17196
rect 15252 17144 15258 17196
rect 15372 17187 15430 17193
rect 15372 17153 15384 17187
rect 15418 17184 15430 17187
rect 16298 17184 16304 17196
rect 15418 17156 16304 17184
rect 15418 17153 15430 17156
rect 15372 17147 15430 17153
rect 16298 17144 16304 17156
rect 16356 17144 16362 17196
rect 16669 17187 16727 17193
rect 16669 17153 16681 17187
rect 16715 17184 16727 17187
rect 16942 17184 16948 17196
rect 16715 17156 16948 17184
rect 16715 17153 16727 17156
rect 16669 17147 16727 17153
rect 16942 17144 16948 17156
rect 17000 17144 17006 17196
rect 18800 17193 18828 17224
rect 18529 17187 18587 17193
rect 18529 17153 18541 17187
rect 18575 17184 18587 17187
rect 18785 17187 18843 17193
rect 18575 17156 18736 17184
rect 18575 17153 18587 17156
rect 18529 17147 18587 17153
rect 13648 17088 13952 17116
rect 14093 17119 14151 17125
rect 11977 17079 12035 17085
rect 14093 17085 14105 17119
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 3697 17051 3755 17057
rect 3697 17017 3709 17051
rect 3743 17048 3755 17051
rect 4246 17048 4252 17060
rect 3743 17020 4252 17048
rect 3743 17017 3755 17020
rect 3697 17011 3755 17017
rect 4246 17008 4252 17020
rect 4304 17008 4310 17060
rect 6181 17051 6239 17057
rect 4540 17020 4752 17048
rect 2590 16940 2596 16992
rect 2648 16980 2654 16992
rect 4540 16980 4568 17020
rect 2648 16952 4568 16980
rect 4724 16980 4752 17020
rect 6181 17017 6193 17051
rect 6227 17048 6239 17051
rect 7006 17048 7012 17060
rect 6227 17020 7012 17048
rect 6227 17017 6239 17020
rect 6181 17011 6239 17017
rect 7006 17008 7012 17020
rect 7064 17008 7070 17060
rect 9416 17048 9444 17079
rect 14108 17048 14136 17079
rect 14550 17076 14556 17128
rect 14608 17116 14614 17128
rect 14737 17119 14795 17125
rect 14737 17116 14749 17119
rect 14608 17088 14749 17116
rect 14608 17076 14614 17088
rect 14737 17085 14749 17088
rect 14783 17085 14795 17119
rect 14737 17079 14795 17085
rect 14829 17119 14887 17125
rect 14829 17085 14841 17119
rect 14875 17116 14887 17119
rect 15212 17116 15240 17144
rect 14875 17088 15240 17116
rect 18708 17116 18736 17156
rect 18785 17153 18797 17187
rect 18831 17153 18843 17187
rect 19794 17184 19800 17196
rect 18785 17147 18843 17153
rect 19076 17156 19800 17184
rect 18708 17088 18920 17116
rect 14875 17085 14887 17088
rect 14829 17079 14887 17085
rect 14844 17048 14872 17079
rect 8588 17020 9444 17048
rect 13280 17020 14044 17048
rect 14108 17020 14872 17048
rect 5718 16980 5724 16992
rect 4724 16952 5724 16980
rect 2648 16940 2654 16952
rect 5718 16940 5724 16952
rect 5776 16940 5782 16992
rect 7193 16983 7251 16989
rect 7193 16949 7205 16983
rect 7239 16980 7251 16983
rect 7926 16980 7932 16992
rect 7239 16952 7932 16980
rect 7239 16949 7251 16952
rect 7193 16943 7251 16949
rect 7926 16940 7932 16952
rect 7984 16980 7990 16992
rect 8588 16980 8616 17020
rect 7984 16952 8616 16980
rect 8757 16983 8815 16989
rect 7984 16940 7990 16952
rect 8757 16949 8769 16983
rect 8803 16980 8815 16983
rect 9122 16980 9128 16992
rect 8803 16952 9128 16980
rect 8803 16949 8815 16952
rect 8757 16943 8815 16949
rect 9122 16940 9128 16952
rect 9180 16980 9186 16992
rect 11514 16980 11520 16992
rect 9180 16952 11520 16980
rect 9180 16940 9186 16952
rect 11514 16940 11520 16952
rect 11572 16940 11578 16992
rect 11609 16983 11667 16989
rect 11609 16949 11621 16983
rect 11655 16980 11667 16983
rect 11790 16980 11796 16992
rect 11655 16952 11796 16980
rect 11655 16949 11667 16952
rect 11609 16943 11667 16949
rect 11790 16940 11796 16952
rect 11848 16940 11854 16992
rect 11885 16983 11943 16989
rect 11885 16949 11897 16983
rect 11931 16980 11943 16983
rect 13280 16980 13308 17020
rect 11931 16952 13308 16980
rect 13357 16983 13415 16989
rect 11931 16949 11943 16952
rect 11885 16943 11943 16949
rect 13357 16949 13369 16983
rect 13403 16980 13415 16983
rect 13906 16980 13912 16992
rect 13403 16952 13912 16980
rect 13403 16949 13415 16952
rect 13357 16943 13415 16949
rect 13906 16940 13912 16952
rect 13964 16940 13970 16992
rect 14016 16980 14044 17020
rect 16482 17008 16488 17060
rect 16540 17048 16546 17060
rect 16540 17020 17448 17048
rect 16540 17008 16546 17020
rect 16390 16980 16396 16992
rect 14016 16952 16396 16980
rect 16390 16940 16396 16952
rect 16448 16940 16454 16992
rect 17310 16980 17316 16992
rect 17271 16952 17316 16980
rect 17310 16940 17316 16952
rect 17368 16940 17374 16992
rect 17420 16980 17448 17020
rect 18414 16980 18420 16992
rect 17420 16952 18420 16980
rect 18414 16940 18420 16952
rect 18472 16940 18478 16992
rect 18892 16980 18920 17088
rect 18966 17076 18972 17128
rect 19024 17116 19030 17128
rect 19076 17125 19104 17156
rect 19794 17144 19800 17156
rect 19852 17144 19858 17196
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17184 20775 17187
rect 20824 17184 20852 17283
rect 22094 17280 22100 17332
rect 22152 17320 22158 17332
rect 22189 17323 22247 17329
rect 22189 17320 22201 17323
rect 22152 17292 22201 17320
rect 22152 17280 22158 17292
rect 22189 17289 22201 17292
rect 22235 17289 22247 17323
rect 22189 17283 22247 17289
rect 22278 17280 22284 17332
rect 22336 17320 22342 17332
rect 22336 17292 22381 17320
rect 22336 17280 22342 17292
rect 21266 17252 21272 17264
rect 21227 17224 21272 17252
rect 21266 17212 21272 17224
rect 21324 17212 21330 17264
rect 22830 17252 22836 17264
rect 22791 17224 22836 17252
rect 22830 17212 22836 17224
rect 22888 17212 22894 17264
rect 20763 17156 20852 17184
rect 20763 17153 20775 17156
rect 20717 17147 20775 17153
rect 19061 17119 19119 17125
rect 19061 17116 19073 17119
rect 19024 17088 19073 17116
rect 19024 17076 19030 17088
rect 19061 17085 19073 17088
rect 19107 17085 19119 17119
rect 19061 17079 19119 17085
rect 19153 17119 19211 17125
rect 19153 17085 19165 17119
rect 19199 17085 19211 17119
rect 20165 17119 20223 17125
rect 20165 17116 20177 17119
rect 19153 17079 19211 17085
rect 19628 17088 20177 17116
rect 19168 17048 19196 17079
rect 19242 17048 19248 17060
rect 19168 17020 19248 17048
rect 19242 17008 19248 17020
rect 19300 17008 19306 17060
rect 19628 17057 19656 17088
rect 20165 17085 20177 17088
rect 20211 17085 20223 17119
rect 20165 17079 20223 17085
rect 20349 17119 20407 17125
rect 20349 17085 20361 17119
rect 20395 17116 20407 17119
rect 21453 17119 21511 17125
rect 21453 17116 21465 17119
rect 20395 17088 21465 17116
rect 20395 17085 20407 17088
rect 20349 17079 20407 17085
rect 21453 17085 21465 17088
rect 21499 17085 21511 17119
rect 21453 17079 21511 17085
rect 22465 17119 22523 17125
rect 22465 17085 22477 17119
rect 22511 17116 22523 17119
rect 22922 17116 22928 17128
rect 22511 17088 22928 17116
rect 22511 17085 22523 17088
rect 22465 17079 22523 17085
rect 19613 17051 19671 17057
rect 19613 17017 19625 17051
rect 19659 17017 19671 17051
rect 19613 17011 19671 17017
rect 19794 17008 19800 17060
rect 19852 17048 19858 17060
rect 20364 17048 20392 17079
rect 21082 17048 21088 17060
rect 19852 17020 20392 17048
rect 20456 17020 21088 17048
rect 19852 17008 19858 17020
rect 19518 16980 19524 16992
rect 18892 16952 19524 16980
rect 19518 16940 19524 16952
rect 19576 16940 19582 16992
rect 19702 16980 19708 16992
rect 19663 16952 19708 16980
rect 19702 16940 19708 16952
rect 19760 16940 19766 16992
rect 20254 16940 20260 16992
rect 20312 16980 20318 16992
rect 20456 16980 20484 17020
rect 21082 17008 21088 17020
rect 21140 17008 21146 17060
rect 21468 17048 21496 17079
rect 22922 17076 22928 17088
rect 22980 17076 22986 17128
rect 22649 17051 22707 17057
rect 22649 17048 22661 17051
rect 21468 17020 22661 17048
rect 22649 17017 22661 17020
rect 22695 17017 22707 17051
rect 22649 17011 22707 17017
rect 20312 16952 20484 16980
rect 20533 16983 20591 16989
rect 20312 16940 20318 16952
rect 20533 16949 20545 16983
rect 20579 16980 20591 16983
rect 20898 16980 20904 16992
rect 20579 16952 20904 16980
rect 20579 16949 20591 16952
rect 20533 16943 20591 16949
rect 20898 16940 20904 16952
rect 20956 16940 20962 16992
rect 23109 16983 23167 16989
rect 23109 16949 23121 16983
rect 23155 16980 23167 16983
rect 23198 16980 23204 16992
rect 23155 16952 23204 16980
rect 23155 16949 23167 16952
rect 23109 16943 23167 16949
rect 23198 16940 23204 16952
rect 23256 16940 23262 16992
rect 1104 16890 23460 16912
rect 1104 16838 3749 16890
rect 3801 16838 3813 16890
rect 3865 16838 3877 16890
rect 3929 16838 3941 16890
rect 3993 16838 4005 16890
rect 4057 16838 9347 16890
rect 9399 16838 9411 16890
rect 9463 16838 9475 16890
rect 9527 16838 9539 16890
rect 9591 16838 9603 16890
rect 9655 16838 14945 16890
rect 14997 16838 15009 16890
rect 15061 16838 15073 16890
rect 15125 16838 15137 16890
rect 15189 16838 15201 16890
rect 15253 16838 20543 16890
rect 20595 16838 20607 16890
rect 20659 16838 20671 16890
rect 20723 16838 20735 16890
rect 20787 16838 20799 16890
rect 20851 16838 23460 16890
rect 1104 16816 23460 16838
rect 3602 16736 3608 16788
rect 3660 16776 3666 16788
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 3660 16748 3801 16776
rect 3660 16736 3666 16748
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 4798 16776 4804 16788
rect 3789 16739 3847 16745
rect 4632 16748 4804 16776
rect 2685 16643 2743 16649
rect 2685 16609 2697 16643
rect 2731 16640 2743 16643
rect 3142 16640 3148 16652
rect 2731 16612 3148 16640
rect 2731 16609 2743 16612
rect 2685 16603 2743 16609
rect 3142 16600 3148 16612
rect 3200 16600 3206 16652
rect 4433 16643 4491 16649
rect 4433 16609 4445 16643
rect 4479 16640 4491 16643
rect 4522 16640 4528 16652
rect 4479 16612 4528 16640
rect 4479 16609 4491 16612
rect 4433 16603 4491 16609
rect 4522 16600 4528 16612
rect 4580 16600 4586 16652
rect 4632 16649 4660 16748
rect 4798 16736 4804 16748
rect 4856 16736 4862 16788
rect 5997 16779 6055 16785
rect 5997 16745 6009 16779
rect 6043 16776 6055 16779
rect 6178 16776 6184 16788
rect 6043 16748 6184 16776
rect 6043 16745 6055 16748
rect 5997 16739 6055 16745
rect 6178 16736 6184 16748
rect 6236 16776 6242 16788
rect 6730 16776 6736 16788
rect 6236 16748 6736 16776
rect 6236 16736 6242 16748
rect 6730 16736 6736 16748
rect 6788 16736 6794 16788
rect 6914 16736 6920 16788
rect 6972 16776 6978 16788
rect 7282 16776 7288 16788
rect 6972 16748 7288 16776
rect 6972 16736 6978 16748
rect 7282 16736 7288 16748
rect 7340 16736 7346 16788
rect 8113 16779 8171 16785
rect 8113 16745 8125 16779
rect 8159 16776 8171 16779
rect 8662 16776 8668 16788
rect 8159 16748 8668 16776
rect 8159 16745 8171 16748
rect 8113 16739 8171 16745
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 10410 16736 10416 16788
rect 10468 16776 10474 16788
rect 11514 16776 11520 16788
rect 10468 16748 11520 16776
rect 10468 16736 10474 16748
rect 11514 16736 11520 16748
rect 11572 16736 11578 16788
rect 15470 16776 15476 16788
rect 14844 16748 15476 16776
rect 7006 16708 7012 16720
rect 6564 16680 7012 16708
rect 6564 16649 6592 16680
rect 7006 16668 7012 16680
rect 7064 16668 7070 16720
rect 8570 16708 8576 16720
rect 7576 16680 8576 16708
rect 4617 16643 4675 16649
rect 4617 16609 4629 16643
rect 4663 16609 4675 16643
rect 4617 16603 4675 16609
rect 6549 16643 6607 16649
rect 6549 16609 6561 16643
rect 6595 16609 6607 16643
rect 6549 16603 6607 16609
rect 6638 16600 6644 16652
rect 6696 16640 6702 16652
rect 7576 16649 7604 16680
rect 8570 16668 8576 16680
rect 8628 16668 8634 16720
rect 7561 16643 7619 16649
rect 6696 16612 6741 16640
rect 6696 16600 6702 16612
rect 7561 16609 7573 16643
rect 7607 16609 7619 16643
rect 7561 16603 7619 16609
rect 7650 16600 7656 16652
rect 7708 16640 7714 16652
rect 7708 16612 7753 16640
rect 7708 16600 7714 16612
rect 8294 16600 8300 16652
rect 8352 16640 8358 16652
rect 9033 16643 9091 16649
rect 9033 16640 9045 16643
rect 8352 16612 9045 16640
rect 8352 16600 8358 16612
rect 9033 16609 9045 16612
rect 9079 16609 9091 16643
rect 9214 16640 9220 16652
rect 9175 16612 9220 16640
rect 9033 16603 9091 16609
rect 9214 16600 9220 16612
rect 9272 16600 9278 16652
rect 14844 16649 14872 16748
rect 15470 16736 15476 16748
rect 15528 16736 15534 16788
rect 16298 16776 16304 16788
rect 16259 16748 16304 16776
rect 16298 16736 16304 16748
rect 16356 16736 16362 16788
rect 18138 16776 18144 16788
rect 17236 16748 18144 16776
rect 17236 16649 17264 16748
rect 18138 16736 18144 16748
rect 18196 16736 18202 16788
rect 18785 16779 18843 16785
rect 18785 16745 18797 16779
rect 18831 16776 18843 16779
rect 18831 16748 20668 16776
rect 18831 16745 18843 16748
rect 18785 16739 18843 16745
rect 18601 16711 18659 16717
rect 18601 16677 18613 16711
rect 18647 16708 18659 16711
rect 19242 16708 19248 16720
rect 18647 16680 19248 16708
rect 18647 16677 18659 16680
rect 18601 16671 18659 16677
rect 19242 16668 19248 16680
rect 19300 16668 19306 16720
rect 19518 16668 19524 16720
rect 19576 16708 19582 16720
rect 19889 16711 19947 16717
rect 19889 16708 19901 16711
rect 19576 16680 19901 16708
rect 19576 16668 19582 16680
rect 19889 16677 19901 16680
rect 19935 16677 19947 16711
rect 19889 16671 19947 16677
rect 13817 16643 13875 16649
rect 13817 16609 13829 16643
rect 13863 16640 13875 16643
rect 14829 16643 14887 16649
rect 14829 16640 14841 16643
rect 13863 16612 14841 16640
rect 13863 16609 13875 16612
rect 13817 16603 13875 16609
rect 14829 16609 14841 16612
rect 14875 16609 14887 16643
rect 14829 16603 14887 16609
rect 17221 16643 17279 16649
rect 17221 16609 17233 16643
rect 17267 16609 17279 16643
rect 19702 16640 19708 16652
rect 17221 16603 17279 16609
rect 19168 16612 19708 16640
rect 1489 16575 1547 16581
rect 1489 16541 1501 16575
rect 1535 16572 1547 16575
rect 2409 16575 2467 16581
rect 1535 16544 2360 16572
rect 1535 16541 1547 16544
rect 1489 16535 1547 16541
rect 1854 16504 1860 16516
rect 1688 16476 1860 16504
rect 1688 16445 1716 16476
rect 1854 16464 1860 16476
rect 1912 16464 1918 16516
rect 2332 16504 2360 16544
rect 2409 16541 2421 16575
rect 2455 16572 2467 16575
rect 2866 16572 2872 16584
rect 2455 16544 2872 16572
rect 2455 16541 2467 16544
rect 2409 16535 2467 16541
rect 2866 16532 2872 16544
rect 2924 16532 2930 16584
rect 3605 16575 3663 16581
rect 3605 16541 3617 16575
rect 3651 16572 3663 16575
rect 4884 16575 4942 16581
rect 3651 16544 4844 16572
rect 3651 16541 3663 16544
rect 3605 16535 3663 16541
rect 2958 16504 2964 16516
rect 2332 16476 2964 16504
rect 2958 16464 2964 16476
rect 3016 16464 3022 16516
rect 4249 16507 4307 16513
rect 4249 16504 4261 16507
rect 3252 16476 4261 16504
rect 1673 16439 1731 16445
rect 1673 16405 1685 16439
rect 1719 16405 1731 16439
rect 1673 16399 1731 16405
rect 1762 16396 1768 16448
rect 1820 16436 1826 16448
rect 1820 16408 1865 16436
rect 1820 16396 1826 16408
rect 2314 16396 2320 16448
rect 2372 16436 2378 16448
rect 3252 16445 3280 16476
rect 4249 16473 4261 16476
rect 4295 16473 4307 16507
rect 4816 16504 4844 16544
rect 4884 16541 4896 16575
rect 4930 16572 4942 16575
rect 5350 16572 5356 16584
rect 4930 16544 5356 16572
rect 4930 16541 4942 16544
rect 4884 16535 4942 16541
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 6454 16572 6460 16584
rect 6415 16544 6460 16572
rect 6454 16532 6460 16544
rect 6512 16532 6518 16584
rect 7282 16532 7288 16584
rect 7340 16572 7346 16584
rect 7745 16575 7803 16581
rect 7745 16572 7757 16575
rect 7340 16544 7757 16572
rect 7340 16532 7346 16544
rect 7745 16541 7757 16544
rect 7791 16572 7803 16575
rect 7834 16572 7840 16584
rect 7791 16544 7840 16572
rect 7791 16541 7803 16544
rect 7745 16535 7803 16541
rect 7834 16532 7840 16544
rect 7892 16532 7898 16584
rect 8389 16575 8447 16581
rect 8389 16541 8401 16575
rect 8435 16572 8447 16575
rect 8478 16572 8484 16584
rect 8435 16544 8484 16572
rect 8435 16541 8447 16544
rect 8389 16535 8447 16541
rect 8478 16532 8484 16544
rect 8536 16532 8542 16584
rect 11149 16575 11207 16581
rect 11149 16541 11161 16575
rect 11195 16572 11207 16575
rect 11238 16572 11244 16584
rect 11195 16544 11244 16572
rect 11195 16541 11207 16544
rect 11149 16535 11207 16541
rect 11238 16532 11244 16544
rect 11296 16532 11302 16584
rect 12345 16575 12403 16581
rect 12345 16541 12357 16575
rect 12391 16541 12403 16575
rect 12345 16535 12403 16541
rect 8110 16504 8116 16516
rect 4816 16476 8116 16504
rect 4249 16467 4307 16473
rect 8110 16464 8116 16476
rect 8168 16464 8174 16516
rect 10904 16507 10962 16513
rect 10904 16473 10916 16507
rect 10950 16504 10962 16507
rect 12066 16504 12072 16516
rect 10950 16476 12072 16504
rect 10950 16473 10962 16476
rect 10904 16467 10962 16473
rect 12066 16464 12072 16476
rect 12124 16464 12130 16516
rect 2777 16439 2835 16445
rect 2777 16436 2789 16439
rect 2372 16408 2789 16436
rect 2372 16396 2378 16408
rect 2777 16405 2789 16408
rect 2823 16405 2835 16439
rect 2777 16399 2835 16405
rect 3237 16439 3295 16445
rect 3237 16405 3249 16439
rect 3283 16405 3295 16439
rect 3237 16399 3295 16405
rect 3326 16396 3332 16448
rect 3384 16436 3390 16448
rect 3421 16439 3479 16445
rect 3421 16436 3433 16439
rect 3384 16408 3433 16436
rect 3384 16396 3390 16408
rect 3421 16405 3433 16408
rect 3467 16405 3479 16439
rect 3421 16399 3479 16405
rect 3694 16396 3700 16448
rect 3752 16436 3758 16448
rect 4157 16439 4215 16445
rect 4157 16436 4169 16439
rect 3752 16408 4169 16436
rect 3752 16396 3758 16408
rect 4157 16405 4169 16408
rect 4203 16405 4215 16439
rect 4157 16399 4215 16405
rect 6086 16396 6092 16448
rect 6144 16436 6150 16448
rect 7098 16436 7104 16448
rect 6144 16408 6189 16436
rect 7059 16408 7104 16436
rect 6144 16396 6150 16408
rect 7098 16396 7104 16408
rect 7156 16396 7162 16448
rect 8202 16436 8208 16448
rect 8163 16408 8208 16436
rect 8202 16396 8208 16408
rect 8260 16396 8266 16448
rect 9309 16439 9367 16445
rect 9309 16405 9321 16439
rect 9355 16436 9367 16439
rect 9490 16436 9496 16448
rect 9355 16408 9496 16436
rect 9355 16405 9367 16408
rect 9309 16399 9367 16405
rect 9490 16396 9496 16408
rect 9548 16396 9554 16448
rect 9674 16436 9680 16448
rect 9635 16408 9680 16436
rect 9674 16396 9680 16408
rect 9732 16396 9738 16448
rect 9769 16439 9827 16445
rect 9769 16405 9781 16439
rect 9815 16436 9827 16439
rect 9858 16436 9864 16448
rect 9815 16408 9864 16436
rect 9815 16405 9827 16408
rect 9769 16399 9827 16405
rect 9858 16396 9864 16408
rect 9916 16396 9922 16448
rect 10042 16396 10048 16448
rect 10100 16436 10106 16448
rect 11425 16439 11483 16445
rect 11425 16436 11437 16439
rect 10100 16408 11437 16436
rect 10100 16396 10106 16408
rect 11425 16405 11437 16408
rect 11471 16405 11483 16439
rect 11698 16436 11704 16448
rect 11659 16408 11704 16436
rect 11425 16399 11483 16405
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 12360 16436 12388 16535
rect 13538 16532 13544 16584
rect 13596 16581 13602 16584
rect 13596 16572 13608 16581
rect 13596 16544 13641 16572
rect 13596 16535 13608 16544
rect 13596 16532 13602 16535
rect 14550 16532 14556 16584
rect 14608 16572 14614 16584
rect 14737 16575 14795 16581
rect 14737 16572 14749 16575
rect 14608 16544 14749 16572
rect 14608 16532 14614 16544
rect 14737 16541 14749 16544
rect 14783 16541 14795 16575
rect 14737 16535 14795 16541
rect 16666 16532 16672 16584
rect 16724 16572 16730 16584
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 16724 16544 16957 16572
rect 16724 16532 16730 16544
rect 16945 16541 16957 16544
rect 16991 16541 17003 16575
rect 16945 16535 17003 16541
rect 17310 16532 17316 16584
rect 17368 16572 17374 16584
rect 17477 16575 17535 16581
rect 17477 16572 17489 16575
rect 17368 16544 17489 16572
rect 17368 16532 17374 16544
rect 17477 16541 17489 16544
rect 17523 16541 17535 16575
rect 17477 16535 17535 16541
rect 18877 16575 18935 16581
rect 18877 16541 18889 16575
rect 18923 16572 18935 16575
rect 19168 16572 19196 16612
rect 19702 16600 19708 16612
rect 19760 16600 19766 16652
rect 20441 16643 20499 16649
rect 20441 16609 20453 16643
rect 20487 16609 20499 16643
rect 20640 16640 20668 16748
rect 21450 16640 21456 16652
rect 20640 16612 21036 16640
rect 21411 16612 21456 16640
rect 20441 16603 20499 16609
rect 18923 16544 19196 16572
rect 18923 16541 18935 16544
rect 18877 16535 18935 16541
rect 19242 16532 19248 16584
rect 19300 16572 19306 16584
rect 19978 16572 19984 16584
rect 19300 16544 19345 16572
rect 19939 16544 19984 16572
rect 19300 16532 19306 16544
rect 19978 16532 19984 16544
rect 20036 16532 20042 16584
rect 20456 16572 20484 16603
rect 20530 16572 20536 16584
rect 20456 16544 20536 16572
rect 20530 16532 20536 16544
rect 20588 16532 20594 16584
rect 20717 16575 20775 16581
rect 20717 16541 20729 16575
rect 20763 16572 20775 16575
rect 20898 16572 20904 16584
rect 20763 16544 20904 16572
rect 20763 16541 20775 16544
rect 20717 16535 20775 16541
rect 20898 16532 20904 16544
rect 20956 16532 20962 16584
rect 21008 16572 21036 16612
rect 21450 16600 21456 16612
rect 21508 16600 21514 16652
rect 23109 16575 23167 16581
rect 21008 16544 22094 16572
rect 15096 16507 15154 16513
rect 15096 16473 15108 16507
rect 15142 16504 15154 16507
rect 15746 16504 15752 16516
rect 15142 16476 15752 16504
rect 15142 16473 15154 16476
rect 15096 16467 15154 16473
rect 15746 16464 15752 16476
rect 15804 16464 15810 16516
rect 12437 16439 12495 16445
rect 12437 16436 12449 16439
rect 12360 16408 12449 16436
rect 12437 16405 12449 16408
rect 12483 16436 12495 16439
rect 13814 16436 13820 16448
rect 12483 16408 13820 16436
rect 12483 16405 12495 16408
rect 12437 16399 12495 16405
rect 13814 16396 13820 16408
rect 13872 16396 13878 16448
rect 14090 16436 14096 16448
rect 14051 16408 14096 16436
rect 14090 16396 14096 16408
rect 14148 16396 14154 16448
rect 16209 16439 16267 16445
rect 16209 16405 16221 16439
rect 16255 16436 16267 16439
rect 16684 16436 16712 16532
rect 17126 16504 17132 16516
rect 17039 16476 17132 16504
rect 17126 16464 17132 16476
rect 17184 16504 17190 16516
rect 17586 16504 17592 16516
rect 17184 16476 17592 16504
rect 17184 16464 17190 16476
rect 17586 16464 17592 16476
rect 17644 16464 17650 16516
rect 20625 16507 20683 16513
rect 20625 16504 20637 16507
rect 19076 16476 20637 16504
rect 16255 16408 16712 16436
rect 16255 16405 16267 16408
rect 16209 16399 16267 16405
rect 16850 16396 16856 16448
rect 16908 16436 16914 16448
rect 18874 16436 18880 16448
rect 16908 16408 18880 16436
rect 16908 16396 16914 16408
rect 18874 16396 18880 16408
rect 18932 16396 18938 16448
rect 19076 16445 19104 16476
rect 20625 16473 20637 16476
rect 20671 16473 20683 16507
rect 21174 16504 21180 16516
rect 21135 16476 21180 16504
rect 20625 16467 20683 16473
rect 21174 16464 21180 16476
rect 21232 16464 21238 16516
rect 21726 16513 21732 16516
rect 21720 16504 21732 16513
rect 21687 16476 21732 16504
rect 21720 16467 21732 16476
rect 21726 16464 21732 16467
rect 21784 16464 21790 16516
rect 22066 16504 22094 16544
rect 23109 16541 23121 16575
rect 23155 16572 23167 16575
rect 23382 16572 23388 16584
rect 23155 16544 23388 16572
rect 23155 16541 23167 16544
rect 23109 16535 23167 16541
rect 23124 16504 23152 16535
rect 23382 16532 23388 16544
rect 23440 16532 23446 16584
rect 22066 16476 23152 16504
rect 19061 16439 19119 16445
rect 19061 16405 19073 16439
rect 19107 16405 19119 16439
rect 19061 16399 19119 16405
rect 20165 16439 20223 16445
rect 20165 16405 20177 16439
rect 20211 16436 20223 16439
rect 20346 16436 20352 16448
rect 20211 16408 20352 16436
rect 20211 16405 20223 16408
rect 20165 16399 20223 16405
rect 20346 16396 20352 16408
rect 20404 16396 20410 16448
rect 21082 16436 21088 16448
rect 21043 16408 21088 16436
rect 21082 16396 21088 16408
rect 21140 16396 21146 16448
rect 22738 16396 22744 16448
rect 22796 16436 22802 16448
rect 22833 16439 22891 16445
rect 22833 16436 22845 16439
rect 22796 16408 22845 16436
rect 22796 16396 22802 16408
rect 22833 16405 22845 16408
rect 22879 16405 22891 16439
rect 22833 16399 22891 16405
rect 22922 16396 22928 16448
rect 22980 16436 22986 16448
rect 22980 16408 23025 16436
rect 22980 16396 22986 16408
rect 1104 16346 23460 16368
rect 1104 16294 6548 16346
rect 6600 16294 6612 16346
rect 6664 16294 6676 16346
rect 6728 16294 6740 16346
rect 6792 16294 6804 16346
rect 6856 16294 12146 16346
rect 12198 16294 12210 16346
rect 12262 16294 12274 16346
rect 12326 16294 12338 16346
rect 12390 16294 12402 16346
rect 12454 16294 17744 16346
rect 17796 16294 17808 16346
rect 17860 16294 17872 16346
rect 17924 16294 17936 16346
rect 17988 16294 18000 16346
rect 18052 16294 23460 16346
rect 1104 16272 23460 16294
rect 2866 16232 2872 16244
rect 2827 16204 2872 16232
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 3694 16232 3700 16244
rect 3655 16204 3700 16232
rect 3694 16192 3700 16204
rect 3752 16192 3758 16244
rect 5169 16235 5227 16241
rect 5169 16201 5181 16235
rect 5215 16201 5227 16235
rect 5169 16195 5227 16201
rect 5445 16235 5503 16241
rect 5445 16201 5457 16235
rect 5491 16232 5503 16235
rect 5534 16232 5540 16244
rect 5491 16204 5540 16232
rect 5491 16201 5503 16204
rect 5445 16195 5503 16201
rect 3329 16167 3387 16173
rect 3329 16133 3341 16167
rect 3375 16164 3387 16167
rect 4246 16164 4252 16176
rect 3375 16136 4252 16164
rect 3375 16133 3387 16136
rect 3329 16127 3387 16133
rect 4246 16124 4252 16136
rect 4304 16124 4310 16176
rect 5184 16164 5212 16195
rect 5534 16192 5540 16204
rect 5592 16192 5598 16244
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 7208 16204 8033 16232
rect 6362 16164 6368 16176
rect 5184 16136 6368 16164
rect 6362 16124 6368 16136
rect 6420 16124 6426 16176
rect 1756 16099 1814 16105
rect 1756 16065 1768 16099
rect 1802 16096 1814 16099
rect 2038 16096 2044 16108
rect 1802 16068 2044 16096
rect 1802 16065 1814 16068
rect 1756 16059 1814 16065
rect 2038 16056 2044 16068
rect 2096 16056 2102 16108
rect 3142 16096 3148 16108
rect 3068 16068 3148 16096
rect 1486 16028 1492 16040
rect 1447 16000 1492 16028
rect 1486 15988 1492 16000
rect 1544 15988 1550 16040
rect 3068 16037 3096 16068
rect 3142 16056 3148 16068
rect 3200 16056 3206 16108
rect 4056 16099 4114 16105
rect 4056 16065 4068 16099
rect 4102 16096 4114 16099
rect 5166 16096 5172 16108
rect 4102 16068 5172 16096
rect 4102 16065 4114 16068
rect 4056 16059 4114 16065
rect 5166 16056 5172 16068
rect 5224 16056 5230 16108
rect 5261 16099 5319 16105
rect 5261 16065 5273 16099
rect 5307 16096 5319 16099
rect 5537 16099 5595 16105
rect 5307 16068 5396 16096
rect 5307 16065 5319 16068
rect 5261 16059 5319 16065
rect 3053 16031 3111 16037
rect 3053 15997 3065 16031
rect 3099 15997 3111 16031
rect 3234 16028 3240 16040
rect 3195 16000 3240 16028
rect 3053 15991 3111 15997
rect 3234 15988 3240 16000
rect 3292 15988 3298 16040
rect 3789 16031 3847 16037
rect 3789 15997 3801 16031
rect 3835 15997 3847 16031
rect 3789 15991 3847 15997
rect 2866 15920 2872 15972
rect 2924 15960 2930 15972
rect 3804 15960 3832 15991
rect 2924 15932 3832 15960
rect 2924 15920 2930 15932
rect 5368 15892 5396 16068
rect 5537 16065 5549 16099
rect 5583 16096 5595 16099
rect 5626 16096 5632 16108
rect 5583 16068 5632 16096
rect 5583 16065 5595 16068
rect 5537 16059 5595 16065
rect 5626 16056 5632 16068
rect 5684 16056 5690 16108
rect 6178 16096 6184 16108
rect 6139 16068 6184 16096
rect 6178 16056 6184 16068
rect 6236 16056 6242 16108
rect 7208 16105 7236 16204
rect 8021 16201 8033 16204
rect 8067 16232 8079 16235
rect 8294 16232 8300 16244
rect 8067 16204 8300 16232
rect 8067 16201 8079 16204
rect 8021 16195 8079 16201
rect 8294 16192 8300 16204
rect 8352 16192 8358 16244
rect 9490 16232 9496 16244
rect 9451 16204 9496 16232
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 9858 16192 9864 16244
rect 9916 16232 9922 16244
rect 9953 16235 10011 16241
rect 9953 16232 9965 16235
rect 9916 16204 9965 16232
rect 9916 16192 9922 16204
rect 9953 16201 9965 16204
rect 9999 16232 10011 16235
rect 9999 16204 11560 16232
rect 9999 16201 10011 16204
rect 9953 16195 10011 16201
rect 7742 16124 7748 16176
rect 7800 16164 7806 16176
rect 11238 16164 11244 16176
rect 7800 16136 11244 16164
rect 7800 16124 7806 16136
rect 7193 16099 7251 16105
rect 7193 16065 7205 16099
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 7285 16099 7343 16105
rect 7285 16065 7297 16099
rect 7331 16065 7343 16099
rect 9122 16096 9128 16108
rect 9180 16105 9186 16108
rect 9416 16105 9444 16136
rect 11238 16124 11244 16136
rect 11296 16164 11302 16176
rect 11296 16136 11376 16164
rect 11296 16124 11302 16136
rect 9092 16068 9128 16096
rect 7285 16059 7343 16065
rect 5442 15988 5448 16040
rect 5500 16028 5506 16040
rect 6365 16031 6423 16037
rect 6365 16028 6377 16031
rect 5500 16000 6377 16028
rect 5500 15988 5506 16000
rect 6365 15997 6377 16000
rect 6411 15997 6423 16031
rect 6365 15991 6423 15997
rect 6454 15988 6460 16040
rect 6512 16028 6518 16040
rect 7300 16028 7328 16059
rect 9122 16056 9128 16068
rect 9180 16059 9192 16105
rect 9401 16099 9459 16105
rect 9401 16065 9413 16099
rect 9447 16065 9459 16099
rect 11054 16096 11060 16108
rect 11112 16105 11118 16108
rect 11348 16105 11376 16136
rect 11532 16105 11560 16204
rect 12066 16192 12072 16244
rect 12124 16232 12130 16244
rect 12161 16235 12219 16241
rect 12161 16232 12173 16235
rect 12124 16204 12173 16232
rect 12124 16192 12130 16204
rect 12161 16201 12173 16204
rect 12207 16201 12219 16235
rect 12161 16195 12219 16201
rect 13633 16235 13691 16241
rect 13633 16201 13645 16235
rect 13679 16232 13691 16235
rect 14550 16232 14556 16244
rect 13679 16204 14556 16232
rect 13679 16201 13691 16204
rect 13633 16195 13691 16201
rect 14550 16192 14556 16204
rect 14608 16192 14614 16244
rect 14642 16192 14648 16244
rect 14700 16232 14706 16244
rect 15105 16235 15163 16241
rect 15105 16232 15117 16235
rect 14700 16204 15117 16232
rect 14700 16192 14706 16204
rect 15105 16201 15117 16204
rect 15151 16201 15163 16235
rect 15105 16195 15163 16201
rect 16209 16235 16267 16241
rect 16209 16201 16221 16235
rect 16255 16232 16267 16235
rect 21726 16232 21732 16244
rect 16255 16204 21732 16232
rect 16255 16201 16267 16204
rect 16209 16195 16267 16201
rect 13992 16167 14050 16173
rect 12268 16136 13768 16164
rect 12268 16105 12296 16136
rect 13740 16105 13768 16136
rect 13992 16133 14004 16167
rect 14038 16164 14050 16167
rect 14090 16164 14096 16176
rect 14038 16136 14096 16164
rect 14038 16133 14050 16136
rect 13992 16127 14050 16133
rect 14090 16124 14096 16136
rect 14148 16124 14154 16176
rect 11024 16068 11060 16096
rect 9401 16059 9459 16065
rect 9180 16056 9186 16059
rect 11054 16056 11060 16068
rect 11112 16059 11124 16105
rect 11333 16099 11391 16105
rect 11333 16065 11345 16099
rect 11379 16065 11391 16099
rect 11333 16059 11391 16065
rect 11517 16099 11575 16105
rect 11517 16065 11529 16099
rect 11563 16065 11575 16099
rect 11517 16059 11575 16065
rect 12253 16099 12311 16105
rect 12253 16065 12265 16099
rect 12299 16065 12311 16099
rect 12509 16099 12567 16105
rect 12509 16096 12521 16099
rect 12253 16059 12311 16065
rect 12360 16068 12521 16096
rect 11112 16056 11118 16059
rect 6512 16000 7328 16028
rect 6512 15988 6518 16000
rect 11698 15988 11704 16040
rect 11756 16028 11762 16040
rect 12360 16028 12388 16068
rect 12509 16065 12521 16068
rect 12555 16065 12567 16099
rect 12509 16059 12567 16065
rect 13725 16099 13783 16105
rect 13725 16065 13737 16099
rect 13771 16096 13783 16099
rect 13814 16096 13820 16108
rect 13771 16068 13820 16096
rect 13771 16065 13783 16068
rect 13725 16059 13783 16065
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 15120 16096 15148 16195
rect 21726 16192 21732 16204
rect 21784 16192 21790 16244
rect 17126 16164 17132 16176
rect 16040 16136 17132 16164
rect 16040 16105 16068 16136
rect 17126 16124 17132 16136
rect 17184 16124 17190 16176
rect 18080 16167 18138 16173
rect 18080 16133 18092 16167
rect 18126 16164 18138 16167
rect 19889 16167 19947 16173
rect 19889 16164 19901 16167
rect 18126 16136 19901 16164
rect 18126 16133 18138 16136
rect 18080 16127 18138 16133
rect 19889 16133 19901 16136
rect 19935 16133 19947 16167
rect 22738 16164 22744 16176
rect 22699 16136 22744 16164
rect 19889 16127 19947 16133
rect 22738 16124 22744 16136
rect 22796 16124 22802 16176
rect 15197 16099 15255 16105
rect 15197 16096 15209 16099
rect 15120 16068 15209 16096
rect 15197 16065 15209 16068
rect 15243 16065 15255 16099
rect 15197 16059 15255 16065
rect 16025 16099 16083 16105
rect 16025 16065 16037 16099
rect 16071 16065 16083 16099
rect 16025 16059 16083 16065
rect 16301 16099 16359 16105
rect 16301 16065 16313 16099
rect 16347 16096 16359 16099
rect 16390 16096 16396 16108
rect 16347 16068 16396 16096
rect 16347 16065 16359 16068
rect 16301 16059 16359 16065
rect 16390 16056 16396 16068
rect 16448 16056 16454 16108
rect 16669 16099 16727 16105
rect 16669 16065 16681 16099
rect 16715 16096 16727 16099
rect 16758 16096 16764 16108
rect 16715 16068 16764 16096
rect 16715 16065 16727 16068
rect 16669 16059 16727 16065
rect 16758 16056 16764 16068
rect 16816 16056 16822 16108
rect 18230 16056 18236 16108
rect 18288 16096 18294 16108
rect 18325 16099 18383 16105
rect 18325 16096 18337 16099
rect 18288 16068 18337 16096
rect 18288 16056 18294 16068
rect 18325 16065 18337 16068
rect 18371 16065 18383 16099
rect 18782 16096 18788 16108
rect 18743 16068 18788 16096
rect 18325 16059 18383 16065
rect 18782 16056 18788 16068
rect 18840 16056 18846 16108
rect 19242 16096 19248 16108
rect 19203 16068 19248 16096
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 19334 16056 19340 16108
rect 19392 16096 19398 16108
rect 19981 16099 20039 16105
rect 19981 16096 19993 16099
rect 19392 16068 19993 16096
rect 19392 16056 19398 16068
rect 19981 16065 19993 16068
rect 20027 16065 20039 16099
rect 19981 16059 20039 16065
rect 21361 16099 21419 16105
rect 21361 16065 21373 16099
rect 21407 16096 21419 16099
rect 21542 16096 21548 16108
rect 21407 16068 21548 16096
rect 21407 16065 21419 16068
rect 21361 16059 21419 16065
rect 21542 16056 21548 16068
rect 21600 16056 21606 16108
rect 21637 16099 21695 16105
rect 21637 16065 21649 16099
rect 21683 16096 21695 16099
rect 22462 16096 22468 16108
rect 21683 16068 22094 16096
rect 22423 16068 22468 16096
rect 21683 16065 21695 16068
rect 21637 16059 21695 16065
rect 11756 16000 12388 16028
rect 18509 16031 18567 16037
rect 11756 15988 11762 16000
rect 18509 15997 18521 16031
rect 18555 15997 18567 16031
rect 18690 16028 18696 16040
rect 18651 16000 18696 16028
rect 18509 15991 18567 15997
rect 5626 15920 5632 15972
rect 5684 15960 5690 15972
rect 6549 15963 6607 15969
rect 6549 15960 6561 15963
rect 5684 15932 6561 15960
rect 5684 15920 5690 15932
rect 6549 15929 6561 15932
rect 6595 15929 6607 15963
rect 16482 15960 16488 15972
rect 16443 15932 16488 15960
rect 6549 15923 6607 15929
rect 16482 15920 16488 15932
rect 16540 15920 16546 15972
rect 16850 15960 16856 15972
rect 16811 15932 16856 15960
rect 16850 15920 16856 15932
rect 16908 15920 16914 15972
rect 18524 15960 18552 15991
rect 18690 15988 18696 16000
rect 18748 15988 18754 16040
rect 19794 16028 19800 16040
rect 18800 16000 19800 16028
rect 18800 15960 18828 16000
rect 19794 15988 19800 16000
rect 19852 15988 19858 16040
rect 22066 16028 22094 16068
rect 22462 16056 22468 16068
rect 22520 16056 22526 16108
rect 22554 16056 22560 16108
rect 22612 16096 22618 16108
rect 22612 16068 22657 16096
rect 22612 16056 22618 16068
rect 22925 16031 22983 16037
rect 22925 16028 22937 16031
rect 22066 16000 22937 16028
rect 22925 15997 22937 16000
rect 22971 15997 22983 16031
rect 22925 15991 22983 15997
rect 18524 15932 18828 15960
rect 19058 15920 19064 15972
rect 19116 15960 19122 15972
rect 20717 15963 20775 15969
rect 20717 15960 20729 15963
rect 19116 15932 20729 15960
rect 19116 15920 19122 15932
rect 20717 15929 20729 15932
rect 20763 15929 20775 15963
rect 20717 15923 20775 15929
rect 6914 15892 6920 15904
rect 5368 15864 6920 15892
rect 6914 15852 6920 15864
rect 6972 15852 6978 15904
rect 7926 15892 7932 15904
rect 7887 15864 7932 15892
rect 7926 15852 7932 15864
rect 7984 15852 7990 15904
rect 10410 15852 10416 15904
rect 10468 15892 10474 15904
rect 11974 15892 11980 15904
rect 10468 15864 11980 15892
rect 10468 15852 10474 15864
rect 11974 15852 11980 15864
rect 12032 15852 12038 15904
rect 13446 15852 13452 15904
rect 13504 15892 13510 15904
rect 15378 15892 15384 15904
rect 13504 15864 15384 15892
rect 13504 15852 13510 15864
rect 15378 15852 15384 15864
rect 15436 15852 15442 15904
rect 15838 15892 15844 15904
rect 15799 15864 15844 15892
rect 15838 15852 15844 15864
rect 15896 15852 15902 15904
rect 16942 15852 16948 15904
rect 17000 15892 17006 15904
rect 17678 15892 17684 15904
rect 17000 15864 17684 15892
rect 17000 15852 17006 15864
rect 17678 15852 17684 15864
rect 17736 15852 17742 15904
rect 17954 15852 17960 15904
rect 18012 15892 18018 15904
rect 18506 15892 18512 15904
rect 18012 15864 18512 15892
rect 18012 15852 18018 15864
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 18874 15852 18880 15904
rect 18932 15892 18938 15904
rect 19153 15895 19211 15901
rect 19153 15892 19165 15895
rect 18932 15864 19165 15892
rect 18932 15852 18938 15864
rect 19153 15861 19165 15864
rect 19199 15861 19211 15895
rect 19153 15855 19211 15861
rect 20438 15852 20444 15904
rect 20496 15892 20502 15904
rect 20625 15895 20683 15901
rect 20625 15892 20637 15895
rect 20496 15864 20637 15892
rect 20496 15852 20502 15864
rect 20625 15861 20637 15864
rect 20671 15861 20683 15895
rect 21450 15892 21456 15904
rect 21411 15864 21456 15892
rect 20625 15855 20683 15861
rect 21450 15852 21456 15864
rect 21508 15852 21514 15904
rect 21542 15852 21548 15904
rect 21600 15892 21606 15904
rect 21821 15895 21879 15901
rect 21821 15892 21833 15895
rect 21600 15864 21833 15892
rect 21600 15852 21606 15864
rect 21821 15861 21833 15864
rect 21867 15861 21879 15895
rect 23106 15892 23112 15904
rect 23067 15864 23112 15892
rect 21821 15855 21879 15861
rect 23106 15852 23112 15864
rect 23164 15852 23170 15904
rect 1104 15802 23460 15824
rect 1104 15750 3749 15802
rect 3801 15750 3813 15802
rect 3865 15750 3877 15802
rect 3929 15750 3941 15802
rect 3993 15750 4005 15802
rect 4057 15750 9347 15802
rect 9399 15750 9411 15802
rect 9463 15750 9475 15802
rect 9527 15750 9539 15802
rect 9591 15750 9603 15802
rect 9655 15750 14945 15802
rect 14997 15750 15009 15802
rect 15061 15750 15073 15802
rect 15125 15750 15137 15802
rect 15189 15750 15201 15802
rect 15253 15750 20543 15802
rect 20595 15750 20607 15802
rect 20659 15750 20671 15802
rect 20723 15750 20735 15802
rect 20787 15750 20799 15802
rect 20851 15750 23460 15802
rect 1104 15728 23460 15750
rect 2038 15688 2044 15700
rect 1999 15660 2044 15688
rect 2038 15648 2044 15660
rect 2096 15648 2102 15700
rect 2314 15688 2320 15700
rect 2148 15660 2320 15688
rect 2148 15620 2176 15660
rect 2314 15648 2320 15660
rect 2372 15648 2378 15700
rect 3050 15648 3056 15700
rect 3108 15648 3114 15700
rect 3234 15648 3240 15700
rect 3292 15688 3298 15700
rect 3513 15691 3571 15697
rect 3513 15688 3525 15691
rect 3292 15660 3525 15688
rect 3292 15648 3298 15660
rect 3513 15657 3525 15660
rect 3559 15657 3571 15691
rect 3513 15651 3571 15657
rect 4157 15691 4215 15697
rect 4157 15657 4169 15691
rect 4203 15688 4215 15691
rect 4890 15688 4896 15700
rect 4203 15660 4896 15688
rect 4203 15657 4215 15660
rect 4157 15651 4215 15657
rect 1412 15592 2176 15620
rect 3068 15620 3096 15648
rect 3789 15623 3847 15629
rect 3789 15620 3801 15623
rect 3068 15592 3801 15620
rect 1412 15496 1440 15592
rect 3789 15589 3801 15592
rect 3835 15589 3847 15623
rect 3789 15583 3847 15589
rect 1486 15512 1492 15564
rect 1544 15552 1550 15564
rect 2038 15552 2044 15564
rect 1544 15524 2044 15552
rect 1544 15512 1550 15524
rect 2038 15512 2044 15524
rect 2096 15552 2102 15564
rect 2133 15555 2191 15561
rect 2133 15552 2145 15555
rect 2096 15524 2145 15552
rect 2096 15512 2102 15524
rect 2133 15521 2145 15524
rect 2179 15521 2191 15555
rect 4172 15552 4200 15651
rect 4890 15648 4896 15660
rect 4948 15648 4954 15700
rect 5166 15648 5172 15700
rect 5224 15688 5230 15700
rect 5629 15691 5687 15697
rect 5629 15688 5641 15691
rect 5224 15660 5641 15688
rect 5224 15648 5230 15660
rect 5629 15657 5641 15660
rect 5675 15657 5687 15691
rect 5629 15651 5687 15657
rect 8941 15691 8999 15697
rect 8941 15657 8953 15691
rect 8987 15688 8999 15691
rect 10134 15688 10140 15700
rect 8987 15660 10140 15688
rect 8987 15657 8999 15660
rect 8941 15651 8999 15657
rect 10134 15648 10140 15660
rect 10192 15648 10198 15700
rect 10505 15691 10563 15697
rect 10505 15688 10517 15691
rect 10244 15660 10517 15688
rect 6454 15552 6460 15564
rect 2133 15515 2191 15521
rect 3988 15524 4200 15552
rect 6415 15524 6460 15552
rect 1394 15484 1400 15496
rect 1307 15456 1400 15484
rect 1394 15444 1400 15456
rect 1452 15444 1458 15496
rect 3988 15493 4016 15524
rect 6454 15512 6460 15524
rect 6512 15512 6518 15564
rect 6641 15555 6699 15561
rect 6641 15521 6653 15555
rect 6687 15552 6699 15555
rect 7098 15552 7104 15564
rect 6687 15524 7104 15552
rect 6687 15521 6699 15524
rect 6641 15515 6699 15521
rect 7098 15512 7104 15524
rect 7156 15512 7162 15564
rect 9858 15552 9864 15564
rect 9819 15524 9864 15552
rect 9858 15512 9864 15524
rect 9916 15512 9922 15564
rect 9953 15555 10011 15561
rect 9953 15521 9965 15555
rect 9999 15552 10011 15555
rect 10244 15552 10272 15660
rect 10505 15657 10517 15660
rect 10551 15657 10563 15691
rect 10505 15651 10563 15657
rect 11054 15648 11060 15700
rect 11112 15688 11118 15700
rect 12345 15691 12403 15697
rect 12345 15688 12357 15691
rect 11112 15660 12357 15688
rect 11112 15648 11118 15660
rect 12345 15657 12357 15660
rect 12391 15657 12403 15691
rect 13446 15688 13452 15700
rect 13407 15660 13452 15688
rect 12345 15651 12403 15657
rect 13446 15648 13452 15660
rect 13504 15648 13510 15700
rect 13630 15688 13636 15700
rect 13591 15660 13636 15688
rect 13630 15648 13636 15660
rect 13688 15648 13694 15700
rect 13909 15691 13967 15697
rect 13909 15657 13921 15691
rect 13955 15688 13967 15691
rect 15746 15688 15752 15700
rect 13955 15660 15608 15688
rect 15707 15660 15752 15688
rect 13955 15657 13967 15660
rect 13909 15651 13967 15657
rect 10410 15620 10416 15632
rect 10371 15592 10416 15620
rect 10410 15580 10416 15592
rect 10468 15580 10474 15632
rect 11422 15580 11428 15632
rect 11480 15620 11486 15632
rect 11517 15623 11575 15629
rect 11517 15620 11529 15623
rect 11480 15592 11529 15620
rect 11480 15580 11486 15592
rect 11517 15589 11529 15592
rect 11563 15589 11575 15623
rect 15580 15620 15608 15660
rect 15746 15648 15752 15660
rect 15804 15648 15810 15700
rect 17954 15688 17960 15700
rect 16132 15660 17960 15688
rect 16132 15620 16160 15660
rect 17954 15648 17960 15660
rect 18012 15648 18018 15700
rect 18046 15648 18052 15700
rect 18104 15688 18110 15700
rect 18693 15691 18751 15697
rect 18104 15660 18368 15688
rect 18104 15648 18110 15660
rect 18340 15632 18368 15660
rect 18693 15657 18705 15691
rect 18739 15688 18751 15691
rect 18782 15688 18788 15700
rect 18739 15660 18788 15688
rect 18739 15657 18751 15660
rect 18693 15651 18751 15657
rect 18782 15648 18788 15660
rect 18840 15648 18846 15700
rect 19978 15688 19984 15700
rect 19939 15660 19984 15688
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 21085 15691 21143 15697
rect 21085 15657 21097 15691
rect 21131 15688 21143 15691
rect 22094 15688 22100 15700
rect 21131 15660 22100 15688
rect 21131 15657 21143 15660
rect 21085 15651 21143 15657
rect 22094 15648 22100 15660
rect 22152 15648 22158 15700
rect 22646 15648 22652 15700
rect 22704 15688 22710 15700
rect 22833 15691 22891 15697
rect 22833 15688 22845 15691
rect 22704 15660 22845 15688
rect 22704 15648 22710 15660
rect 22833 15657 22845 15660
rect 22879 15657 22891 15691
rect 22833 15651 22891 15657
rect 15580 15592 16160 15620
rect 17865 15623 17923 15629
rect 11517 15583 11575 15589
rect 17865 15589 17877 15623
rect 17911 15620 17923 15623
rect 17911 15592 18276 15620
rect 17911 15589 17923 15592
rect 17865 15583 17923 15589
rect 9999 15524 10272 15552
rect 11149 15555 11207 15561
rect 9999 15521 10011 15524
rect 9953 15515 10011 15521
rect 11149 15521 11161 15555
rect 11195 15552 11207 15555
rect 11606 15552 11612 15564
rect 11195 15524 11612 15552
rect 11195 15521 11207 15524
rect 11149 15515 11207 15521
rect 11606 15512 11612 15524
rect 11664 15552 11670 15564
rect 11664 15524 11744 15552
rect 11664 15512 11670 15524
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 4154 15444 4160 15496
rect 4212 15484 4218 15496
rect 4249 15487 4307 15493
rect 4249 15484 4261 15487
rect 4212 15456 4261 15484
rect 4212 15444 4218 15456
rect 4249 15453 4261 15456
rect 4295 15453 4307 15487
rect 4249 15447 4307 15453
rect 4338 15444 4344 15496
rect 4396 15484 4402 15496
rect 4985 15487 5043 15493
rect 4985 15484 4997 15487
rect 4396 15456 4997 15484
rect 4396 15444 4402 15456
rect 4985 15453 4997 15456
rect 5031 15453 5043 15487
rect 4985 15447 5043 15453
rect 5442 15444 5448 15496
rect 5500 15484 5506 15496
rect 5905 15487 5963 15493
rect 5905 15484 5917 15487
rect 5500 15456 5917 15484
rect 5500 15444 5506 15456
rect 5905 15453 5917 15456
rect 5951 15453 5963 15487
rect 5905 15447 5963 15453
rect 7193 15487 7251 15493
rect 7193 15453 7205 15487
rect 7239 15484 7251 15487
rect 7742 15484 7748 15496
rect 7239 15456 7748 15484
rect 7239 15453 7251 15456
rect 7193 15447 7251 15453
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 9585 15487 9643 15493
rect 9585 15453 9597 15487
rect 9631 15484 9643 15487
rect 9766 15484 9772 15496
rect 9631 15456 9772 15484
rect 9631 15453 9643 15456
rect 9585 15447 9643 15453
rect 9766 15444 9772 15456
rect 9824 15444 9830 15496
rect 10042 15484 10048 15496
rect 10003 15456 10048 15484
rect 10042 15444 10048 15456
rect 10100 15444 10106 15496
rect 10134 15444 10140 15496
rect 10192 15484 10198 15496
rect 10965 15487 11023 15493
rect 10965 15484 10977 15487
rect 10192 15456 10977 15484
rect 10192 15444 10198 15456
rect 10965 15453 10977 15456
rect 11011 15453 11023 15487
rect 11330 15484 11336 15496
rect 11291 15456 11336 15484
rect 10965 15447 11023 15453
rect 11330 15444 11336 15456
rect 11388 15444 11394 15496
rect 11716 15493 11744 15524
rect 13814 15512 13820 15564
rect 13872 15552 13878 15564
rect 14277 15555 14335 15561
rect 14277 15552 14289 15555
rect 13872 15524 14289 15552
rect 13872 15512 13878 15524
rect 14277 15521 14289 15524
rect 14323 15521 14335 15555
rect 18046 15552 18052 15564
rect 18007 15524 18052 15552
rect 14277 15515 14335 15521
rect 18046 15512 18052 15524
rect 18104 15512 18110 15564
rect 18248 15561 18276 15592
rect 18322 15580 18328 15632
rect 18380 15620 18386 15632
rect 18966 15620 18972 15632
rect 18380 15592 18972 15620
rect 18380 15580 18386 15592
rect 18966 15580 18972 15592
rect 19024 15580 19030 15632
rect 20898 15620 20904 15632
rect 20180 15592 20904 15620
rect 18233 15555 18291 15561
rect 18233 15521 18245 15555
rect 18279 15552 18291 15555
rect 19242 15552 19248 15564
rect 18279 15524 19248 15552
rect 18279 15521 18291 15524
rect 18233 15515 18291 15521
rect 19242 15512 19248 15524
rect 19300 15512 19306 15564
rect 19429 15555 19487 15561
rect 19429 15521 19441 15555
rect 19475 15552 19487 15555
rect 19794 15552 19800 15564
rect 19475 15524 19800 15552
rect 19475 15521 19487 15524
rect 19429 15515 19487 15521
rect 19794 15512 19800 15524
rect 19852 15512 19858 15564
rect 20180 15561 20208 15592
rect 20898 15580 20904 15592
rect 20956 15620 20962 15632
rect 21266 15620 21272 15632
rect 20956 15592 21272 15620
rect 20956 15580 20962 15592
rect 21266 15580 21272 15592
rect 21324 15580 21330 15632
rect 20165 15555 20223 15561
rect 20165 15521 20177 15555
rect 20211 15521 20223 15555
rect 20346 15552 20352 15564
rect 20307 15524 20352 15552
rect 20165 15515 20223 15521
rect 20346 15512 20352 15524
rect 20404 15512 20410 15564
rect 20990 15512 20996 15564
rect 21048 15552 21054 15564
rect 21453 15555 21511 15561
rect 21453 15552 21465 15555
rect 21048 15524 21465 15552
rect 21048 15512 21054 15524
rect 21453 15521 21465 15524
rect 21499 15521 21511 15555
rect 21453 15515 21511 15521
rect 11701 15487 11759 15493
rect 11701 15453 11713 15487
rect 11747 15453 11759 15487
rect 11701 15447 11759 15453
rect 13630 15444 13636 15496
rect 13688 15484 13694 15496
rect 13725 15487 13783 15493
rect 13725 15484 13737 15487
rect 13688 15456 13737 15484
rect 13688 15444 13694 15456
rect 13725 15453 13737 15456
rect 13771 15453 13783 15487
rect 13725 15447 13783 15453
rect 14544 15487 14602 15493
rect 14544 15453 14556 15487
rect 14590 15484 14602 15487
rect 15838 15484 15844 15496
rect 14590 15456 15844 15484
rect 14590 15453 14602 15456
rect 14544 15447 14602 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 16393 15487 16451 15493
rect 16393 15453 16405 15487
rect 16439 15453 16451 15487
rect 16393 15447 16451 15453
rect 16485 15487 16543 15493
rect 16485 15453 16497 15487
rect 16531 15484 16543 15487
rect 18138 15484 18144 15496
rect 16531 15456 18144 15484
rect 16531 15453 16543 15456
rect 16485 15447 16543 15453
rect 1762 15376 1768 15428
rect 1820 15416 1826 15428
rect 2378 15419 2436 15425
rect 2378 15416 2390 15419
rect 1820 15388 2390 15416
rect 1820 15376 1826 15388
rect 2378 15385 2390 15388
rect 2424 15385 2436 15419
rect 2378 15379 2436 15385
rect 7460 15419 7518 15425
rect 7460 15385 7472 15419
rect 7506 15416 7518 15419
rect 7926 15416 7932 15428
rect 7506 15388 7932 15416
rect 7506 15385 7518 15388
rect 7460 15379 7518 15385
rect 7926 15376 7932 15388
rect 7984 15376 7990 15428
rect 14185 15419 14243 15425
rect 8036 15388 8708 15416
rect 4890 15348 4896 15360
rect 4851 15320 4896 15348
rect 4890 15308 4896 15320
rect 4948 15308 4954 15360
rect 5721 15351 5779 15357
rect 5721 15317 5733 15351
rect 5767 15348 5779 15351
rect 5902 15348 5908 15360
rect 5767 15320 5908 15348
rect 5767 15317 5779 15320
rect 5721 15311 5779 15317
rect 5902 15308 5908 15320
rect 5960 15308 5966 15360
rect 5994 15308 6000 15360
rect 6052 15348 6058 15360
rect 6052 15320 6097 15348
rect 6052 15308 6058 15320
rect 6362 15308 6368 15360
rect 6420 15348 6426 15360
rect 6549 15351 6607 15357
rect 6549 15348 6561 15351
rect 6420 15320 6561 15348
rect 6420 15308 6426 15320
rect 6549 15317 6561 15320
rect 6595 15317 6607 15351
rect 6549 15311 6607 15317
rect 6914 15308 6920 15360
rect 6972 15348 6978 15360
rect 7027 15351 7085 15357
rect 7027 15348 7039 15351
rect 6972 15320 7039 15348
rect 6972 15308 6978 15320
rect 7027 15317 7039 15320
rect 7073 15348 7085 15351
rect 8036 15348 8064 15388
rect 8570 15348 8576 15360
rect 7073 15320 8064 15348
rect 8531 15320 8576 15348
rect 7073 15317 7085 15320
rect 7027 15311 7085 15317
rect 8570 15308 8576 15320
rect 8628 15308 8634 15360
rect 8680 15348 8708 15388
rect 10704 15388 14136 15416
rect 10704 15348 10732 15388
rect 10870 15348 10876 15360
rect 8680 15320 10732 15348
rect 10831 15320 10876 15348
rect 10870 15308 10876 15320
rect 10928 15308 10934 15360
rect 14108 15348 14136 15388
rect 14185 15385 14197 15419
rect 14231 15416 14243 15419
rect 14458 15416 14464 15428
rect 14231 15388 14464 15416
rect 14231 15385 14243 15388
rect 14185 15379 14243 15385
rect 14458 15376 14464 15388
rect 14516 15376 14522 15428
rect 16408 15416 16436 15447
rect 18138 15444 18144 15456
rect 18196 15444 18202 15496
rect 18874 15484 18880 15496
rect 18835 15456 18880 15484
rect 18874 15444 18880 15456
rect 18932 15444 18938 15496
rect 20898 15484 20904 15496
rect 20859 15456 20904 15484
rect 20898 15444 20904 15456
rect 20956 15444 20962 15496
rect 21169 15487 21227 15493
rect 21169 15484 21181 15487
rect 21100 15456 21181 15484
rect 16574 15416 16580 15428
rect 15672 15388 16580 15416
rect 15562 15348 15568 15360
rect 14108 15320 15568 15348
rect 15562 15308 15568 15320
rect 15620 15308 15626 15360
rect 15672 15357 15700 15388
rect 16574 15376 16580 15388
rect 16632 15376 16638 15428
rect 16752 15419 16810 15425
rect 16752 15385 16764 15419
rect 16798 15416 16810 15419
rect 17586 15416 17592 15428
rect 16798 15388 17592 15416
rect 16798 15385 16810 15388
rect 16752 15379 16810 15385
rect 17586 15376 17592 15388
rect 17644 15376 17650 15428
rect 17678 15376 17684 15428
rect 17736 15416 17742 15428
rect 18325 15419 18383 15425
rect 18325 15416 18337 15419
rect 17736 15388 18337 15416
rect 17736 15376 17742 15388
rect 18325 15385 18337 15388
rect 18371 15385 18383 15419
rect 20441 15419 20499 15425
rect 20441 15416 20453 15419
rect 18325 15379 18383 15385
rect 19076 15388 20453 15416
rect 19076 15357 19104 15388
rect 20441 15385 20453 15388
rect 20487 15385 20499 15419
rect 21100 15416 21128 15456
rect 21169 15453 21181 15456
rect 21215 15453 21227 15487
rect 21169 15447 21227 15453
rect 21266 15444 21272 15496
rect 21324 15484 21330 15496
rect 22738 15484 22744 15496
rect 21324 15456 22744 15484
rect 21324 15444 21330 15456
rect 22738 15444 22744 15456
rect 22796 15444 22802 15496
rect 22830 15444 22836 15496
rect 22888 15484 22894 15496
rect 23109 15487 23167 15493
rect 23109 15484 23121 15487
rect 22888 15456 23121 15484
rect 22888 15444 22894 15456
rect 23109 15453 23121 15456
rect 23155 15453 23167 15487
rect 23109 15447 23167 15453
rect 20441 15379 20499 15385
rect 20824 15388 21128 15416
rect 15657 15351 15715 15357
rect 15657 15317 15669 15351
rect 15703 15317 15715 15351
rect 15657 15311 15715 15317
rect 19061 15351 19119 15357
rect 19061 15317 19073 15351
rect 19107 15317 19119 15351
rect 19518 15348 19524 15360
rect 19479 15320 19524 15348
rect 19061 15311 19119 15317
rect 19518 15308 19524 15320
rect 19576 15308 19582 15360
rect 19610 15308 19616 15360
rect 19668 15348 19674 15360
rect 20824 15357 20852 15388
rect 20809 15351 20867 15357
rect 19668 15320 19713 15348
rect 19668 15308 19674 15320
rect 20809 15317 20821 15351
rect 20855 15317 20867 15351
rect 21100 15348 21128 15388
rect 21720 15419 21778 15425
rect 21720 15385 21732 15419
rect 21766 15416 21778 15419
rect 22370 15416 22376 15428
rect 21766 15388 22376 15416
rect 21766 15385 21778 15388
rect 21720 15379 21778 15385
rect 22370 15376 22376 15388
rect 22428 15376 22434 15428
rect 21266 15348 21272 15360
rect 21100 15320 21272 15348
rect 20809 15311 20867 15317
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 21361 15351 21419 15357
rect 21361 15317 21373 15351
rect 21407 15348 21419 15351
rect 22186 15348 22192 15360
rect 21407 15320 22192 15348
rect 21407 15317 21419 15320
rect 21361 15311 21419 15317
rect 22186 15308 22192 15320
rect 22244 15308 22250 15360
rect 22922 15348 22928 15360
rect 22883 15320 22928 15348
rect 22922 15308 22928 15320
rect 22980 15308 22986 15360
rect 1104 15258 23460 15280
rect 1104 15206 6548 15258
rect 6600 15206 6612 15258
rect 6664 15206 6676 15258
rect 6728 15206 6740 15258
rect 6792 15206 6804 15258
rect 6856 15206 12146 15258
rect 12198 15206 12210 15258
rect 12262 15206 12274 15258
rect 12326 15206 12338 15258
rect 12390 15206 12402 15258
rect 12454 15206 17744 15258
rect 17796 15206 17808 15258
rect 17860 15206 17872 15258
rect 17924 15206 17936 15258
rect 17988 15206 18000 15258
rect 18052 15206 23460 15258
rect 1104 15184 23460 15206
rect 1394 15144 1400 15156
rect 1355 15116 1400 15144
rect 1394 15104 1400 15116
rect 1452 15104 1458 15156
rect 4246 15144 4252 15156
rect 4207 15116 4252 15144
rect 4246 15104 4252 15116
rect 4304 15104 4310 15156
rect 5442 15144 5448 15156
rect 4448 15116 5448 15144
rect 4448 15088 4476 15116
rect 5442 15104 5448 15116
rect 5500 15104 5506 15156
rect 5813 15147 5871 15153
rect 5813 15113 5825 15147
rect 5859 15144 5871 15147
rect 7558 15144 7564 15156
rect 5859 15116 7564 15144
rect 5859 15113 5871 15116
rect 5813 15107 5871 15113
rect 7558 15104 7564 15116
rect 7616 15144 7622 15156
rect 8021 15147 8079 15153
rect 8021 15144 8033 15147
rect 7616 15116 8033 15144
rect 7616 15104 7622 15116
rect 8021 15113 8033 15116
rect 8067 15113 8079 15147
rect 8021 15107 8079 15113
rect 8110 15104 8116 15156
rect 8168 15144 8174 15156
rect 9394 15147 9452 15153
rect 9394 15144 9406 15147
rect 8168 15116 9406 15144
rect 8168 15104 8174 15116
rect 9394 15113 9406 15116
rect 9440 15113 9452 15147
rect 11606 15144 11612 15156
rect 11567 15116 11612 15144
rect 9394 15107 9452 15113
rect 11606 15104 11612 15116
rect 11664 15104 11670 15156
rect 16482 15104 16488 15156
rect 16540 15144 16546 15156
rect 16669 15147 16727 15153
rect 16669 15144 16681 15147
rect 16540 15116 16681 15144
rect 16540 15104 16546 15116
rect 16669 15113 16681 15116
rect 16715 15144 16727 15147
rect 18417 15147 18475 15153
rect 18417 15144 18429 15147
rect 16715 15116 18429 15144
rect 16715 15113 16727 15116
rect 16669 15107 16727 15113
rect 18417 15113 18429 15116
rect 18463 15113 18475 15147
rect 18417 15107 18475 15113
rect 18690 15104 18696 15156
rect 18748 15144 18754 15156
rect 18877 15147 18935 15153
rect 18877 15144 18889 15147
rect 18748 15116 18889 15144
rect 18748 15104 18754 15116
rect 18877 15113 18889 15116
rect 18923 15113 18935 15147
rect 19334 15144 19340 15156
rect 19295 15116 19340 15144
rect 18877 15107 18935 15113
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 19610 15104 19616 15156
rect 19668 15144 19674 15156
rect 19797 15147 19855 15153
rect 19797 15144 19809 15147
rect 19668 15116 19809 15144
rect 19668 15104 19674 15116
rect 19797 15113 19809 15116
rect 19843 15113 19855 15147
rect 20898 15144 20904 15156
rect 20859 15116 20904 15144
rect 19797 15107 19855 15113
rect 20898 15104 20904 15116
rect 20956 15104 20962 15156
rect 21266 15104 21272 15156
rect 21324 15144 21330 15156
rect 21361 15147 21419 15153
rect 21361 15144 21373 15147
rect 21324 15116 21373 15144
rect 21324 15104 21330 15116
rect 21361 15113 21373 15116
rect 21407 15113 21419 15147
rect 22186 15144 22192 15156
rect 22147 15116 22192 15144
rect 21361 15107 21419 15113
rect 22186 15104 22192 15116
rect 22244 15104 22250 15156
rect 22649 15147 22707 15153
rect 22649 15113 22661 15147
rect 22695 15144 22707 15147
rect 23474 15144 23480 15156
rect 22695 15116 23480 15144
rect 22695 15113 22707 15116
rect 22649 15107 22707 15113
rect 23474 15104 23480 15116
rect 23532 15104 23538 15156
rect 2532 15079 2590 15085
rect 2532 15045 2544 15079
rect 2578 15076 2590 15079
rect 4341 15079 4399 15085
rect 2578 15048 4292 15076
rect 2578 15045 2590 15048
rect 2532 15039 2590 15045
rect 2038 14968 2044 15020
rect 2096 15008 2102 15020
rect 2777 15011 2835 15017
rect 2777 15008 2789 15011
rect 2096 14980 2789 15008
rect 2096 14968 2102 14980
rect 2777 14977 2789 14980
rect 2823 15008 2835 15011
rect 2866 15008 2872 15020
rect 2823 14980 2872 15008
rect 2823 14977 2835 14980
rect 2777 14971 2835 14977
rect 2866 14968 2872 14980
rect 2924 14968 2930 15020
rect 2958 14968 2964 15020
rect 3016 15008 3022 15020
rect 3125 15011 3183 15017
rect 3125 15008 3137 15011
rect 3016 14980 3137 15008
rect 3016 14968 3022 14980
rect 3125 14977 3137 14980
rect 3171 14977 3183 15011
rect 4264 15008 4292 15048
rect 4341 15045 4353 15079
rect 4387 15076 4399 15079
rect 4430 15076 4436 15088
rect 4387 15048 4436 15076
rect 4387 15045 4399 15048
rect 4341 15039 4399 15045
rect 4430 15036 4436 15048
rect 4488 15036 4494 15088
rect 4982 15036 4988 15088
rect 5040 15076 5046 15088
rect 5077 15079 5135 15085
rect 5077 15076 5089 15079
rect 5040 15048 5089 15076
rect 5040 15036 5046 15048
rect 5077 15045 5089 15048
rect 5123 15045 5135 15079
rect 5077 15039 5135 15045
rect 5166 15036 5172 15088
rect 5224 15076 5230 15088
rect 7650 15076 7656 15088
rect 5224 15048 7656 15076
rect 5224 15036 5230 15048
rect 7650 15036 7656 15048
rect 7708 15036 7714 15088
rect 10781 15079 10839 15085
rect 10781 15045 10793 15079
rect 10827 15076 10839 15079
rect 11238 15076 11244 15088
rect 10827 15048 11244 15076
rect 10827 15045 10839 15048
rect 10781 15039 10839 15045
rect 11238 15036 11244 15048
rect 11296 15036 11302 15088
rect 14090 15076 14096 15088
rect 14003 15048 14096 15076
rect 14090 15036 14096 15048
rect 14148 15076 14154 15088
rect 14553 15079 14611 15085
rect 14553 15076 14565 15079
rect 14148 15048 14565 15076
rect 14148 15036 14154 15048
rect 14553 15045 14565 15048
rect 14599 15076 14611 15079
rect 14826 15076 14832 15088
rect 14599 15048 14832 15076
rect 14599 15045 14611 15048
rect 14553 15039 14611 15045
rect 14826 15036 14832 15048
rect 14884 15076 14890 15088
rect 22094 15076 22100 15088
rect 14884 15048 19932 15076
rect 22055 15048 22100 15076
rect 14884 15036 14890 15048
rect 19904 15020 19932 15048
rect 22094 15036 22100 15048
rect 22152 15036 22158 15088
rect 5626 15008 5632 15020
rect 4264 14980 5632 15008
rect 3125 14971 3183 14977
rect 5626 14968 5632 14980
rect 5684 14968 5690 15020
rect 5718 14968 5724 15020
rect 5776 15008 5782 15020
rect 6914 15008 6920 15020
rect 5776 14980 5821 15008
rect 5920 14980 6920 15008
rect 5776 14968 5782 14980
rect 5920 14940 5948 14980
rect 6914 14968 6920 14980
rect 6972 14968 6978 15020
rect 7006 14968 7012 15020
rect 7064 15008 7070 15020
rect 7478 15011 7536 15017
rect 7478 15008 7490 15011
rect 7064 14980 7490 15008
rect 7064 14968 7070 14980
rect 7478 14977 7490 14980
rect 7524 14977 7536 15011
rect 7478 14971 7536 14977
rect 9030 14968 9036 15020
rect 9088 15008 9094 15020
rect 9953 15011 10011 15017
rect 9953 15008 9965 15011
rect 9088 14980 9965 15008
rect 9088 14968 9094 14980
rect 9953 14977 9965 14980
rect 9999 15008 10011 15011
rect 11054 15008 11060 15020
rect 9999 14980 11060 15008
rect 9999 14977 10011 14980
rect 9953 14971 10011 14977
rect 11054 14968 11060 14980
rect 11112 14968 11118 15020
rect 11333 15011 11391 15017
rect 11333 14977 11345 15011
rect 11379 15008 11391 15011
rect 11974 15008 11980 15020
rect 11379 14980 11980 15008
rect 11379 14977 11391 14980
rect 11333 14971 11391 14977
rect 11974 14968 11980 14980
rect 12032 14968 12038 15020
rect 12733 15011 12791 15017
rect 12733 14977 12745 15011
rect 12779 15008 12791 15011
rect 12894 15008 12900 15020
rect 12779 14980 12900 15008
rect 12779 14977 12791 14980
rect 12733 14971 12791 14977
rect 12894 14968 12900 14980
rect 12952 14968 12958 15020
rect 12989 15011 13047 15017
rect 12989 14977 13001 15011
rect 13035 15008 13047 15011
rect 13814 15008 13820 15020
rect 13035 14980 13820 15008
rect 13035 14977 13047 14980
rect 12989 14971 13047 14977
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 14369 15011 14427 15017
rect 14369 14977 14381 15011
rect 14415 15008 14427 15011
rect 15378 15008 15384 15020
rect 14415 14980 15384 15008
rect 14415 14977 14427 14980
rect 14369 14971 14427 14977
rect 15378 14968 15384 14980
rect 15436 14968 15442 15020
rect 15749 15011 15807 15017
rect 15749 14977 15761 15011
rect 15795 14977 15807 15011
rect 16482 15008 16488 15020
rect 16443 14980 16488 15008
rect 15749 14971 15807 14977
rect 4172 14912 5948 14940
rect 5997 14943 6055 14949
rect 2406 14764 2412 14816
rect 2464 14804 2470 14816
rect 4172 14804 4200 14912
rect 5997 14909 6009 14943
rect 6043 14909 6055 14943
rect 7742 14940 7748 14952
rect 7703 14912 7748 14940
rect 5997 14903 6055 14909
rect 4246 14832 4252 14884
rect 4304 14872 4310 14884
rect 6012 14872 6040 14903
rect 7742 14900 7748 14912
rect 7800 14900 7806 14952
rect 8754 14900 8760 14952
rect 8812 14940 8818 14952
rect 9125 14943 9183 14949
rect 9125 14940 9137 14943
rect 8812 14912 9137 14940
rect 8812 14900 8818 14912
rect 9125 14909 9137 14912
rect 9171 14909 9183 14943
rect 9398 14940 9404 14952
rect 9359 14912 9404 14940
rect 9125 14903 9183 14909
rect 9398 14900 9404 14912
rect 9456 14900 9462 14952
rect 9674 14900 9680 14952
rect 9732 14940 9738 14952
rect 9861 14943 9919 14949
rect 9861 14940 9873 14943
rect 9732 14912 9873 14940
rect 9732 14900 9738 14912
rect 9861 14909 9873 14912
rect 9907 14909 9919 14943
rect 13832 14940 13860 14968
rect 14826 14940 14832 14952
rect 13832 14912 14832 14940
rect 9861 14903 9919 14909
rect 14826 14900 14832 14912
rect 14884 14940 14890 14952
rect 15289 14943 15347 14949
rect 15289 14940 15301 14943
rect 14884 14912 15301 14940
rect 14884 14900 14890 14912
rect 15289 14909 15301 14912
rect 15335 14909 15347 14943
rect 15764 14940 15792 14971
rect 16482 14968 16488 14980
rect 16540 14968 16546 15020
rect 17793 15011 17851 15017
rect 17793 14977 17805 15011
rect 17839 15008 17851 15011
rect 18049 15011 18107 15017
rect 17839 14980 18000 15008
rect 17839 14977 17851 14980
rect 17793 14971 17851 14977
rect 17034 14940 17040 14952
rect 15764 14912 17040 14940
rect 15289 14903 15347 14909
rect 17034 14900 17040 14912
rect 17092 14900 17098 14952
rect 17972 14940 18000 14980
rect 18049 14977 18061 15011
rect 18095 15008 18107 15011
rect 18138 15008 18144 15020
rect 18095 14980 18144 15008
rect 18095 14977 18107 14980
rect 18049 14971 18107 14977
rect 18138 14968 18144 14980
rect 18196 14968 18202 15020
rect 18506 15008 18512 15020
rect 18467 14980 18512 15008
rect 18506 14968 18512 14980
rect 18564 14968 18570 15020
rect 19426 15008 19432 15020
rect 19387 14980 19432 15008
rect 19426 14968 19432 14980
rect 19484 14968 19490 15020
rect 19886 15008 19892 15020
rect 19847 14980 19892 15008
rect 19886 14968 19892 14980
rect 19944 14968 19950 15020
rect 21174 14968 21180 15020
rect 21232 15008 21238 15020
rect 21269 15011 21327 15017
rect 21269 15008 21281 15011
rect 21232 14980 21281 15008
rect 21232 14968 21238 14980
rect 21269 14977 21281 14980
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 22370 14968 22376 15020
rect 22428 15008 22434 15020
rect 22833 15011 22891 15017
rect 22833 15008 22845 15011
rect 22428 14980 22845 15008
rect 22428 14968 22434 14980
rect 22833 14977 22845 14980
rect 22879 14977 22891 15011
rect 22833 14971 22891 14977
rect 23109 15011 23167 15017
rect 23109 14977 23121 15011
rect 23155 15008 23167 15011
rect 23198 15008 23204 15020
rect 23155 14980 23204 15008
rect 23155 14977 23167 14980
rect 23109 14971 23167 14977
rect 23198 14968 23204 14980
rect 23256 14968 23262 15020
rect 18322 14940 18328 14952
rect 17972 14912 18184 14940
rect 18283 14912 18328 14940
rect 4304 14844 6040 14872
rect 6365 14875 6423 14881
rect 4304 14832 4310 14844
rect 6365 14841 6377 14875
rect 6411 14872 6423 14875
rect 6454 14872 6460 14884
rect 6411 14844 6460 14872
rect 6411 14841 6423 14844
rect 6365 14835 6423 14841
rect 6454 14832 6460 14844
rect 6512 14832 6518 14884
rect 14182 14872 14188 14884
rect 9876 14844 11376 14872
rect 14143 14844 14188 14872
rect 2464 14776 4200 14804
rect 2464 14764 2470 14776
rect 4614 14764 4620 14816
rect 4672 14804 4678 14816
rect 5353 14807 5411 14813
rect 5353 14804 5365 14807
rect 4672 14776 5365 14804
rect 4672 14764 4678 14776
rect 5353 14773 5365 14776
rect 5399 14773 5411 14807
rect 5353 14767 5411 14773
rect 5626 14764 5632 14816
rect 5684 14804 5690 14816
rect 9876 14804 9904 14844
rect 11054 14804 11060 14816
rect 5684 14776 9904 14804
rect 11015 14776 11060 14804
rect 5684 14764 5690 14776
rect 11054 14764 11060 14776
rect 11112 14764 11118 14816
rect 11146 14764 11152 14816
rect 11204 14804 11210 14816
rect 11348 14804 11376 14844
rect 14182 14832 14188 14844
rect 14240 14832 14246 14884
rect 13538 14804 13544 14816
rect 11204 14776 11249 14804
rect 11348 14776 13544 14804
rect 11204 14764 11210 14776
rect 13538 14764 13544 14776
rect 13596 14764 13602 14816
rect 13909 14807 13967 14813
rect 13909 14773 13921 14807
rect 13955 14804 13967 14807
rect 13998 14804 14004 14816
rect 13955 14776 14004 14804
rect 13955 14773 13967 14776
rect 13909 14767 13967 14773
rect 13998 14764 14004 14776
rect 14056 14764 14062 14816
rect 15562 14804 15568 14816
rect 15523 14776 15568 14804
rect 15562 14764 15568 14776
rect 15620 14764 15626 14816
rect 15838 14804 15844 14816
rect 15799 14776 15844 14804
rect 15838 14764 15844 14776
rect 15896 14764 15902 14816
rect 18156 14804 18184 14912
rect 18322 14900 18328 14912
rect 18380 14900 18386 14952
rect 19150 14940 19156 14952
rect 19111 14912 19156 14940
rect 19150 14900 19156 14912
rect 19208 14900 19214 14952
rect 20717 14943 20775 14949
rect 20717 14909 20729 14943
rect 20763 14940 20775 14943
rect 20990 14940 20996 14952
rect 20763 14912 20996 14940
rect 20763 14909 20775 14912
rect 20717 14903 20775 14909
rect 20990 14900 20996 14912
rect 21048 14900 21054 14952
rect 21450 14900 21456 14952
rect 21508 14940 21514 14952
rect 22005 14943 22063 14949
rect 21508 14912 21553 14940
rect 21508 14900 21514 14912
rect 22005 14909 22017 14943
rect 22051 14940 22063 14943
rect 22646 14940 22652 14952
rect 22051 14912 22652 14940
rect 22051 14909 22063 14912
rect 22005 14903 22063 14909
rect 22646 14900 22652 14912
rect 22704 14900 22710 14952
rect 18874 14832 18880 14884
rect 18932 14872 18938 14884
rect 22925 14875 22983 14881
rect 22925 14872 22937 14875
rect 18932 14844 22937 14872
rect 18932 14832 18938 14844
rect 22925 14841 22937 14844
rect 22971 14841 22983 14875
rect 22925 14835 22983 14841
rect 19610 14804 19616 14816
rect 18156 14776 19616 14804
rect 19610 14764 19616 14776
rect 19668 14764 19674 14816
rect 22094 14764 22100 14816
rect 22152 14804 22158 14816
rect 22557 14807 22615 14813
rect 22557 14804 22569 14807
rect 22152 14776 22569 14804
rect 22152 14764 22158 14776
rect 22557 14773 22569 14776
rect 22603 14773 22615 14807
rect 22557 14767 22615 14773
rect 1104 14714 23460 14736
rect 1104 14662 3749 14714
rect 3801 14662 3813 14714
rect 3865 14662 3877 14714
rect 3929 14662 3941 14714
rect 3993 14662 4005 14714
rect 4057 14662 9347 14714
rect 9399 14662 9411 14714
rect 9463 14662 9475 14714
rect 9527 14662 9539 14714
rect 9591 14662 9603 14714
rect 9655 14662 14945 14714
rect 14997 14662 15009 14714
rect 15061 14662 15073 14714
rect 15125 14662 15137 14714
rect 15189 14662 15201 14714
rect 15253 14662 20543 14714
rect 20595 14662 20607 14714
rect 20659 14662 20671 14714
rect 20723 14662 20735 14714
rect 20787 14662 20799 14714
rect 20851 14662 23460 14714
rect 1104 14640 23460 14662
rect 1578 14600 1584 14612
rect 1539 14572 1584 14600
rect 1578 14560 1584 14572
rect 1636 14560 1642 14612
rect 1946 14560 1952 14612
rect 2004 14600 2010 14612
rect 2041 14603 2099 14609
rect 2041 14600 2053 14603
rect 2004 14572 2053 14600
rect 2004 14560 2010 14572
rect 2041 14569 2053 14572
rect 2087 14569 2099 14603
rect 2406 14600 2412 14612
rect 2367 14572 2412 14600
rect 2041 14563 2099 14569
rect 2406 14560 2412 14572
rect 2464 14560 2470 14612
rect 2682 14600 2688 14612
rect 2643 14572 2688 14600
rect 2682 14560 2688 14572
rect 2740 14560 2746 14612
rect 2958 14600 2964 14612
rect 2919 14572 2964 14600
rect 2958 14560 2964 14572
rect 3016 14560 3022 14612
rect 4157 14603 4215 14609
rect 4157 14569 4169 14603
rect 4203 14600 4215 14603
rect 5626 14600 5632 14612
rect 4203 14572 5632 14600
rect 4203 14569 4215 14572
rect 4157 14563 4215 14569
rect 1765 14535 1823 14541
rect 1765 14501 1777 14535
rect 1811 14532 1823 14535
rect 2130 14532 2136 14544
rect 1811 14504 2136 14532
rect 1811 14501 1823 14504
rect 1765 14495 1823 14501
rect 2130 14492 2136 14504
rect 2188 14492 2194 14544
rect 1397 14399 1455 14405
rect 1397 14365 1409 14399
rect 1443 14396 1455 14399
rect 1578 14396 1584 14408
rect 1443 14368 1584 14396
rect 1443 14365 1455 14368
rect 1397 14359 1455 14365
rect 1578 14356 1584 14368
rect 1636 14356 1642 14408
rect 1946 14396 1952 14408
rect 1907 14368 1952 14396
rect 1946 14356 1952 14368
rect 2004 14356 2010 14408
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2424 14396 2452 14560
rect 4172 14532 4200 14563
rect 5626 14560 5632 14572
rect 5684 14560 5690 14612
rect 5718 14560 5724 14612
rect 5776 14600 5782 14612
rect 8941 14603 8999 14609
rect 5776 14572 8340 14600
rect 5776 14560 5782 14572
rect 2884 14504 4200 14532
rect 2884 14405 2912 14504
rect 4614 14464 4620 14476
rect 4575 14436 4620 14464
rect 4614 14424 4620 14436
rect 4672 14424 4678 14476
rect 4801 14467 4859 14473
rect 4801 14433 4813 14467
rect 4847 14433 4859 14467
rect 4982 14464 4988 14476
rect 4943 14436 4988 14464
rect 4801 14427 4859 14433
rect 2271 14368 2452 14396
rect 2593 14399 2651 14405
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2593 14365 2605 14399
rect 2639 14396 2651 14399
rect 2869 14399 2927 14405
rect 2869 14396 2881 14399
rect 2639 14368 2881 14396
rect 2639 14365 2651 14368
rect 2593 14359 2651 14365
rect 2869 14365 2881 14368
rect 2915 14365 2927 14399
rect 2869 14359 2927 14365
rect 3234 14356 3240 14408
rect 3292 14396 3298 14408
rect 3605 14399 3663 14405
rect 3605 14396 3617 14399
rect 3292 14368 3617 14396
rect 3292 14356 3298 14368
rect 3605 14365 3617 14368
rect 3651 14365 3663 14399
rect 3605 14359 3663 14365
rect 3973 14399 4031 14405
rect 3973 14365 3985 14399
rect 4019 14396 4031 14399
rect 4154 14396 4160 14408
rect 4019 14368 4160 14396
rect 4019 14365 4031 14368
rect 3973 14359 4031 14365
rect 4154 14356 4160 14368
rect 4212 14356 4218 14408
rect 4816 14396 4844 14427
rect 4982 14424 4988 14436
rect 5040 14424 5046 14476
rect 7558 14464 7564 14476
rect 7519 14436 7564 14464
rect 7558 14424 7564 14436
rect 7616 14424 7622 14476
rect 7791 14467 7849 14473
rect 7791 14464 7803 14467
rect 7668 14436 7803 14464
rect 5718 14396 5724 14408
rect 4816 14368 5724 14396
rect 5718 14356 5724 14368
rect 5776 14356 5782 14408
rect 6454 14356 6460 14408
rect 6512 14396 6518 14408
rect 7668 14396 7696 14436
rect 7791 14433 7803 14436
rect 7837 14433 7849 14467
rect 8312 14464 8340 14572
rect 8941 14569 8953 14603
rect 8987 14600 8999 14603
rect 9214 14600 9220 14612
rect 8987 14572 9220 14600
rect 8987 14569 8999 14572
rect 8941 14563 8999 14569
rect 9214 14560 9220 14572
rect 9272 14560 9278 14612
rect 10134 14600 10140 14612
rect 10095 14572 10140 14600
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 10413 14603 10471 14609
rect 10413 14569 10425 14603
rect 10459 14600 10471 14603
rect 10870 14600 10876 14612
rect 10459 14572 10876 14600
rect 10459 14569 10471 14572
rect 10413 14563 10471 14569
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 12894 14560 12900 14612
rect 12952 14600 12958 14612
rect 13541 14603 13599 14609
rect 13541 14600 13553 14603
rect 12952 14572 13553 14600
rect 12952 14560 12958 14572
rect 13541 14569 13553 14572
rect 13587 14569 13599 14603
rect 15930 14600 15936 14612
rect 15891 14572 15936 14600
rect 13541 14563 13599 14569
rect 15930 14560 15936 14572
rect 15988 14560 15994 14612
rect 17586 14600 17592 14612
rect 17547 14572 17592 14600
rect 17586 14560 17592 14572
rect 17644 14560 17650 14612
rect 19061 14603 19119 14609
rect 19061 14569 19073 14603
rect 19107 14600 19119 14603
rect 19518 14600 19524 14612
rect 19107 14572 19524 14600
rect 19107 14569 19119 14572
rect 19061 14563 19119 14569
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 19886 14560 19892 14612
rect 19944 14600 19950 14612
rect 20993 14603 21051 14609
rect 20993 14600 21005 14603
rect 19944 14572 21005 14600
rect 19944 14560 19950 14572
rect 20993 14569 21005 14572
rect 21039 14569 21051 14603
rect 20993 14563 21051 14569
rect 22186 14560 22192 14612
rect 22244 14600 22250 14612
rect 22557 14603 22615 14609
rect 22557 14600 22569 14603
rect 22244 14572 22569 14600
rect 22244 14560 22250 14572
rect 22557 14569 22569 14572
rect 22603 14600 22615 14603
rect 23658 14600 23664 14612
rect 22603 14572 23664 14600
rect 22603 14569 22615 14572
rect 22557 14563 22615 14569
rect 23658 14560 23664 14572
rect 23716 14560 23722 14612
rect 10505 14535 10563 14541
rect 10505 14532 10517 14535
rect 9968 14504 10517 14532
rect 7791 14427 7849 14433
rect 8220 14436 8340 14464
rect 6512 14368 7696 14396
rect 6512 14356 6518 14368
rect 5252 14331 5310 14337
rect 5252 14297 5264 14331
rect 5298 14328 5310 14331
rect 5626 14328 5632 14340
rect 5298 14300 5632 14328
rect 5298 14297 5310 14300
rect 5252 14291 5310 14297
rect 5626 14288 5632 14300
rect 5684 14288 5690 14340
rect 4525 14263 4583 14269
rect 4525 14229 4537 14263
rect 4571 14260 4583 14263
rect 5994 14260 6000 14272
rect 4571 14232 6000 14260
rect 4571 14229 4583 14232
rect 4525 14223 4583 14229
rect 5994 14220 6000 14232
rect 6052 14220 6058 14272
rect 6270 14220 6276 14272
rect 6328 14260 6334 14272
rect 6365 14263 6423 14269
rect 6365 14260 6377 14263
rect 6328 14232 6377 14260
rect 6328 14220 6334 14232
rect 6365 14229 6377 14232
rect 6411 14229 6423 14263
rect 6365 14223 6423 14229
rect 6457 14263 6515 14269
rect 6457 14229 6469 14263
rect 6503 14260 6515 14263
rect 7282 14260 7288 14272
rect 6503 14232 7288 14260
rect 6503 14229 6515 14232
rect 6457 14223 6515 14229
rect 7282 14220 7288 14232
rect 7340 14220 7346 14272
rect 7834 14269 7840 14272
rect 7830 14260 7840 14269
rect 7795 14232 7840 14260
rect 7830 14223 7840 14232
rect 7834 14220 7840 14223
rect 7892 14220 7898 14272
rect 8220 14260 8248 14436
rect 8570 14424 8576 14476
rect 8628 14464 8634 14476
rect 9493 14467 9551 14473
rect 9493 14464 9505 14467
rect 8628 14436 9505 14464
rect 8628 14424 8634 14436
rect 9493 14433 9505 14436
rect 9539 14433 9551 14467
rect 9493 14427 9551 14433
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 8846 14396 8852 14408
rect 8343 14368 8852 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 8846 14356 8852 14368
rect 8904 14396 8910 14408
rect 9582 14396 9588 14408
rect 8904 14368 9588 14396
rect 8904 14356 8910 14368
rect 9582 14356 9588 14368
rect 9640 14356 9646 14408
rect 9968 14405 9996 14504
rect 10505 14501 10517 14504
rect 10551 14501 10563 14535
rect 16022 14532 16028 14544
rect 10505 14495 10563 14501
rect 10612 14504 16028 14532
rect 10612 14464 10640 14504
rect 16022 14492 16028 14504
rect 16080 14492 16086 14544
rect 17497 14535 17555 14541
rect 17497 14501 17509 14535
rect 17543 14532 17555 14535
rect 17543 14504 18276 14532
rect 17543 14501 17555 14504
rect 17497 14495 17555 14501
rect 11146 14464 11152 14476
rect 10060 14436 10640 14464
rect 11107 14436 11152 14464
rect 9953 14399 10011 14405
rect 9953 14365 9965 14399
rect 9999 14365 10011 14399
rect 9953 14359 10011 14365
rect 9309 14331 9367 14337
rect 9309 14297 9321 14331
rect 9355 14328 9367 14331
rect 9861 14331 9919 14337
rect 9861 14328 9873 14331
rect 9355 14300 9873 14328
rect 9355 14297 9367 14300
rect 9309 14291 9367 14297
rect 9861 14297 9873 14300
rect 9907 14328 9919 14331
rect 10060 14328 10088 14436
rect 11146 14424 11152 14436
rect 11204 14424 11210 14476
rect 14826 14424 14832 14476
rect 14884 14464 14890 14476
rect 16117 14467 16175 14473
rect 16117 14464 16129 14467
rect 14884 14436 16129 14464
rect 14884 14424 14890 14436
rect 16117 14433 16129 14436
rect 16163 14433 16175 14467
rect 16117 14427 16175 14433
rect 10226 14396 10232 14408
rect 10187 14368 10232 14396
rect 10226 14356 10232 14368
rect 10284 14356 10290 14408
rect 10873 14399 10931 14405
rect 10873 14365 10885 14399
rect 10919 14396 10931 14399
rect 11330 14396 11336 14408
rect 10919 14368 11336 14396
rect 10919 14365 10931 14368
rect 10873 14359 10931 14365
rect 11330 14356 11336 14368
rect 11388 14356 11394 14408
rect 12066 14396 12072 14408
rect 12027 14368 12072 14396
rect 12066 14356 12072 14368
rect 12124 14356 12130 14408
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14396 12219 14399
rect 12618 14396 12624 14408
rect 12207 14368 12624 14396
rect 12207 14365 12219 14368
rect 12161 14359 12219 14365
rect 12618 14356 12624 14368
rect 12676 14356 12682 14408
rect 12894 14396 12900 14408
rect 12855 14368 12900 14396
rect 12894 14356 12900 14368
rect 12952 14356 12958 14408
rect 14734 14396 14740 14408
rect 14695 14368 14740 14396
rect 14734 14356 14740 14368
rect 14792 14356 14798 14408
rect 15470 14396 15476 14408
rect 15431 14368 15476 14396
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 15838 14356 15844 14408
rect 15896 14396 15902 14408
rect 18248 14405 18276 14504
rect 18417 14467 18475 14473
rect 18417 14433 18429 14467
rect 18463 14464 18475 14467
rect 19150 14464 19156 14476
rect 18463 14436 19156 14464
rect 18463 14433 18475 14436
rect 18417 14427 18475 14433
rect 19150 14424 19156 14436
rect 19208 14424 19214 14476
rect 20990 14464 20996 14476
rect 20824 14436 20996 14464
rect 16373 14399 16431 14405
rect 16373 14396 16385 14399
rect 15896 14368 16385 14396
rect 15896 14356 15902 14368
rect 16373 14365 16385 14368
rect 16419 14365 16431 14399
rect 16373 14359 16431 14365
rect 18233 14399 18291 14405
rect 18233 14365 18245 14399
rect 18279 14396 18291 14399
rect 18506 14396 18512 14408
rect 18279 14368 18512 14396
rect 18279 14365 18291 14368
rect 18233 14359 18291 14365
rect 18506 14356 18512 14368
rect 18564 14356 18570 14408
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14396 18751 14399
rect 20070 14396 20076 14408
rect 18739 14368 20076 14396
rect 18739 14365 18751 14368
rect 18693 14359 18751 14365
rect 20070 14356 20076 14368
rect 20128 14356 20134 14408
rect 20346 14356 20352 14408
rect 20404 14405 20410 14408
rect 20404 14396 20416 14405
rect 20625 14399 20683 14405
rect 20404 14368 20449 14396
rect 20404 14359 20416 14368
rect 20625 14365 20637 14399
rect 20671 14396 20683 14399
rect 20714 14396 20720 14408
rect 20671 14368 20720 14396
rect 20671 14365 20683 14368
rect 20625 14359 20683 14365
rect 20404 14356 20410 14359
rect 20714 14356 20720 14368
rect 20772 14396 20778 14408
rect 20824 14396 20852 14436
rect 20990 14424 20996 14436
rect 21048 14464 21054 14476
rect 21177 14467 21235 14473
rect 21177 14464 21189 14467
rect 21048 14436 21189 14464
rect 21048 14424 21054 14436
rect 21177 14433 21189 14436
rect 21223 14433 21235 14467
rect 21177 14427 21235 14433
rect 20772 14368 20852 14396
rect 20772 14356 20778 14368
rect 20898 14356 20904 14408
rect 20956 14396 20962 14408
rect 21444 14399 21502 14405
rect 20956 14368 21001 14396
rect 20956 14356 20962 14368
rect 21444 14365 21456 14399
rect 21490 14396 21502 14399
rect 22002 14396 22008 14408
rect 21490 14368 22008 14396
rect 21490 14365 21502 14368
rect 21444 14359 21502 14365
rect 22002 14356 22008 14368
rect 22060 14356 22066 14408
rect 23106 14396 23112 14408
rect 23067 14368 23112 14396
rect 23106 14356 23112 14368
rect 23164 14356 23170 14408
rect 9907 14300 10088 14328
rect 10244 14328 10272 14356
rect 10965 14331 11023 14337
rect 10965 14328 10977 14331
rect 10244 14300 10977 14328
rect 9907 14297 9919 14300
rect 9861 14291 9919 14297
rect 10965 14297 10977 14300
rect 11011 14297 11023 14331
rect 10965 14291 11023 14297
rect 11790 14288 11796 14340
rect 11848 14328 11854 14340
rect 13906 14328 13912 14340
rect 11848 14300 13912 14328
rect 11848 14288 11854 14300
rect 13906 14288 13912 14300
rect 13964 14288 13970 14340
rect 14458 14288 14464 14340
rect 14516 14328 14522 14340
rect 15565 14331 15623 14337
rect 15565 14328 15577 14331
rect 14516 14300 15577 14328
rect 14516 14288 14522 14300
rect 15565 14297 15577 14300
rect 15611 14297 15623 14331
rect 15565 14291 15623 14297
rect 15749 14331 15807 14337
rect 15749 14297 15761 14331
rect 15795 14328 15807 14331
rect 18874 14328 18880 14340
rect 15795 14300 18880 14328
rect 15795 14297 15807 14300
rect 15749 14291 15807 14297
rect 18874 14288 18880 14300
rect 18932 14288 18938 14340
rect 19150 14288 19156 14340
rect 19208 14328 19214 14340
rect 19208 14300 22968 14328
rect 19208 14288 19214 14300
rect 9401 14263 9459 14269
rect 9401 14260 9413 14263
rect 8220 14232 9413 14260
rect 9401 14229 9413 14232
rect 9447 14229 9459 14263
rect 11422 14260 11428 14272
rect 11383 14232 11428 14260
rect 9401 14223 9459 14229
rect 11422 14220 11428 14232
rect 11480 14220 11486 14272
rect 12802 14260 12808 14272
rect 12763 14232 12808 14260
rect 12802 14220 12808 14232
rect 12860 14220 12866 14272
rect 13722 14220 13728 14272
rect 13780 14260 13786 14272
rect 14093 14263 14151 14269
rect 14093 14260 14105 14263
rect 13780 14232 14105 14260
rect 13780 14220 13786 14232
rect 14093 14229 14105 14232
rect 14139 14229 14151 14263
rect 14093 14223 14151 14229
rect 14829 14263 14887 14269
rect 14829 14229 14841 14263
rect 14875 14260 14887 14263
rect 14918 14260 14924 14272
rect 14875 14232 14924 14260
rect 14875 14229 14887 14232
rect 14829 14223 14887 14229
rect 14918 14220 14924 14232
rect 14976 14220 14982 14272
rect 18598 14260 18604 14272
rect 18559 14232 18604 14260
rect 18598 14220 18604 14232
rect 18656 14220 18662 14272
rect 19245 14263 19303 14269
rect 19245 14229 19257 14263
rect 19291 14260 19303 14263
rect 19426 14260 19432 14272
rect 19291 14232 19432 14260
rect 19291 14229 19303 14232
rect 19245 14223 19303 14229
rect 19426 14220 19432 14232
rect 19484 14260 19490 14272
rect 19978 14260 19984 14272
rect 19484 14232 19984 14260
rect 19484 14220 19490 14232
rect 19978 14220 19984 14232
rect 20036 14220 20042 14272
rect 20162 14220 20168 14272
rect 20220 14260 20226 14272
rect 20717 14263 20775 14269
rect 20717 14260 20729 14263
rect 20220 14232 20729 14260
rect 20220 14220 20226 14232
rect 20717 14229 20729 14232
rect 20763 14229 20775 14263
rect 20717 14223 20775 14229
rect 21726 14220 21732 14272
rect 21784 14260 21790 14272
rect 22278 14260 22284 14272
rect 21784 14232 22284 14260
rect 21784 14220 21790 14232
rect 22278 14220 22284 14232
rect 22336 14220 22342 14272
rect 22646 14220 22652 14272
rect 22704 14260 22710 14272
rect 22940 14269 22968 14300
rect 22925 14263 22983 14269
rect 22704 14232 22749 14260
rect 22704 14220 22710 14232
rect 22925 14229 22937 14263
rect 22971 14229 22983 14263
rect 22925 14223 22983 14229
rect 1104 14170 23460 14192
rect 1104 14118 6548 14170
rect 6600 14118 6612 14170
rect 6664 14118 6676 14170
rect 6728 14118 6740 14170
rect 6792 14118 6804 14170
rect 6856 14118 12146 14170
rect 12198 14118 12210 14170
rect 12262 14118 12274 14170
rect 12326 14118 12338 14170
rect 12390 14118 12402 14170
rect 12454 14118 17744 14170
rect 17796 14118 17808 14170
rect 17860 14118 17872 14170
rect 17924 14118 17936 14170
rect 17988 14118 18000 14170
rect 18052 14118 23460 14170
rect 1104 14096 23460 14118
rect 1946 14016 1952 14068
rect 2004 14056 2010 14068
rect 2777 14059 2835 14065
rect 2777 14056 2789 14059
rect 2004 14028 2789 14056
rect 2004 14016 2010 14028
rect 2777 14025 2789 14028
rect 2823 14056 2835 14059
rect 5166 14056 5172 14068
rect 2823 14028 5172 14056
rect 2823 14025 2835 14028
rect 2777 14019 2835 14025
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 5718 14056 5724 14068
rect 5679 14028 5724 14056
rect 5718 14016 5724 14028
rect 5776 14016 5782 14068
rect 6362 14016 6368 14068
rect 6420 14056 6426 14068
rect 6641 14059 6699 14065
rect 6641 14056 6653 14059
rect 6420 14028 6653 14056
rect 6420 14016 6426 14028
rect 6641 14025 6653 14028
rect 6687 14025 6699 14059
rect 6641 14019 6699 14025
rect 7101 14059 7159 14065
rect 7101 14025 7113 14059
rect 7147 14056 7159 14059
rect 7282 14056 7288 14068
rect 7147 14028 7288 14056
rect 7147 14025 7159 14028
rect 7101 14019 7159 14025
rect 7282 14016 7288 14028
rect 7340 14016 7346 14068
rect 8018 14016 8024 14068
rect 8076 14056 8082 14068
rect 8297 14059 8355 14065
rect 8297 14056 8309 14059
rect 8076 14028 8309 14056
rect 8076 14016 8082 14028
rect 8297 14025 8309 14028
rect 8343 14025 8355 14059
rect 8297 14019 8355 14025
rect 9122 14016 9128 14068
rect 9180 14056 9186 14068
rect 9217 14059 9275 14065
rect 9217 14056 9229 14059
rect 9180 14028 9229 14056
rect 9180 14016 9186 14028
rect 9217 14025 9229 14028
rect 9263 14025 9275 14059
rect 9217 14019 9275 14025
rect 10873 14059 10931 14065
rect 10873 14025 10885 14059
rect 10919 14025 10931 14059
rect 10873 14019 10931 14025
rect 2866 13948 2872 14000
rect 2924 13988 2930 14000
rect 4982 13988 4988 14000
rect 2924 13960 4988 13988
rect 2924 13948 2930 13960
rect 2498 13880 2504 13932
rect 2556 13920 2562 13932
rect 2593 13923 2651 13929
rect 2593 13920 2605 13923
rect 2556 13892 2605 13920
rect 2556 13880 2562 13892
rect 2593 13889 2605 13892
rect 2639 13889 2651 13923
rect 2593 13883 2651 13889
rect 3136 13923 3194 13929
rect 3136 13889 3148 13923
rect 3182 13920 3194 13923
rect 3510 13920 3516 13932
rect 3182 13892 3516 13920
rect 3182 13889 3194 13892
rect 3136 13883 3194 13889
rect 3510 13880 3516 13892
rect 3568 13880 3574 13932
rect 4246 13880 4252 13932
rect 4304 13880 4310 13932
rect 4356 13929 4384 13960
rect 4982 13948 4988 13960
rect 5040 13948 5046 14000
rect 5736 13988 5764 14016
rect 6086 13988 6092 14000
rect 5736 13960 6092 13988
rect 6086 13948 6092 13960
rect 6144 13948 6150 14000
rect 8110 13948 8116 14000
rect 8168 13988 8174 14000
rect 9309 13991 9367 13997
rect 9309 13988 9321 13991
rect 8168 13960 9321 13988
rect 8168 13948 8174 13960
rect 9309 13957 9321 13960
rect 9355 13957 9367 13991
rect 10413 13991 10471 13997
rect 10413 13988 10425 13991
rect 9309 13951 9367 13957
rect 9416 13960 10425 13988
rect 4341 13923 4399 13929
rect 4341 13889 4353 13923
rect 4387 13889 4399 13923
rect 4341 13883 4399 13889
rect 4608 13923 4666 13929
rect 4608 13889 4620 13923
rect 4654 13920 4666 13923
rect 4890 13920 4896 13932
rect 4654 13892 4896 13920
rect 4654 13889 4666 13892
rect 4608 13883 4666 13889
rect 4890 13880 4896 13892
rect 4948 13880 4954 13932
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 5810 13920 5816 13932
rect 5132 13892 5816 13920
rect 5132 13880 5138 13892
rect 5810 13880 5816 13892
rect 5868 13880 5874 13932
rect 5994 13920 6000 13932
rect 5955 13892 6000 13920
rect 5994 13880 6000 13892
rect 6052 13880 6058 13932
rect 6454 13880 6460 13932
rect 6512 13920 6518 13932
rect 7009 13923 7067 13929
rect 7009 13920 7021 13923
rect 6512 13892 7021 13920
rect 6512 13880 6518 13892
rect 7009 13889 7021 13892
rect 7055 13889 7067 13923
rect 7466 13920 7472 13932
rect 7427 13892 7472 13920
rect 7009 13883 7067 13889
rect 7466 13880 7472 13892
rect 7524 13880 7530 13932
rect 7834 13880 7840 13932
rect 7892 13920 7898 13932
rect 8389 13923 8447 13929
rect 8389 13920 8401 13923
rect 7892 13892 8401 13920
rect 7892 13880 7898 13892
rect 8389 13889 8401 13892
rect 8435 13889 8447 13923
rect 8570 13920 8576 13932
rect 8531 13892 8576 13920
rect 8389 13883 8447 13889
rect 8570 13880 8576 13892
rect 8628 13880 8634 13932
rect 9122 13880 9128 13932
rect 9180 13920 9186 13932
rect 9416 13920 9444 13960
rect 10413 13957 10425 13960
rect 10459 13957 10471 13991
rect 10888 13988 10916 14019
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 14090 14056 14096 14068
rect 11112 14028 14096 14056
rect 11112 14016 11118 14028
rect 14090 14016 14096 14028
rect 14148 14016 14154 14068
rect 14553 14059 14611 14065
rect 14553 14025 14565 14059
rect 14599 14056 14611 14059
rect 15470 14056 15476 14068
rect 14599 14028 15476 14056
rect 14599 14025 14611 14028
rect 14553 14019 14611 14025
rect 15470 14016 15476 14028
rect 15528 14016 15534 14068
rect 16117 14059 16175 14065
rect 16117 14025 16129 14059
rect 16163 14056 16175 14059
rect 16666 14056 16672 14068
rect 16163 14028 16672 14056
rect 16163 14025 16175 14028
rect 16117 14019 16175 14025
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 19150 14056 19156 14068
rect 17604 14028 19156 14056
rect 11330 13988 11336 14000
rect 10888 13960 11336 13988
rect 10413 13951 10471 13957
rect 11330 13948 11336 13960
rect 11388 13948 11394 14000
rect 11422 13948 11428 14000
rect 11480 13988 11486 14000
rect 11762 13991 11820 13997
rect 11762 13988 11774 13991
rect 11480 13960 11774 13988
rect 11480 13948 11486 13960
rect 11762 13957 11774 13960
rect 11808 13957 11820 13991
rect 13814 13988 13820 14000
rect 11762 13951 11820 13957
rect 13188 13960 13820 13988
rect 9950 13920 9956 13932
rect 9180 13892 9444 13920
rect 9911 13892 9956 13920
rect 9180 13880 9186 13892
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 10502 13920 10508 13932
rect 10463 13892 10508 13920
rect 10502 13880 10508 13892
rect 10560 13880 10566 13932
rect 11146 13920 11152 13932
rect 11107 13892 11152 13920
rect 11146 13880 11152 13892
rect 11204 13880 11210 13932
rect 11238 13880 11244 13932
rect 11296 13920 11302 13932
rect 13188 13929 13216 13960
rect 13814 13948 13820 13960
rect 13872 13948 13878 14000
rect 16482 13988 16488 14000
rect 16443 13960 16488 13988
rect 16482 13948 16488 13960
rect 16540 13948 16546 14000
rect 11517 13923 11575 13929
rect 11517 13920 11529 13923
rect 11296 13892 11529 13920
rect 11296 13880 11302 13892
rect 11517 13889 11529 13892
rect 11563 13889 11575 13923
rect 11517 13883 11575 13889
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13889 13231 13923
rect 13173 13883 13231 13889
rect 13440 13923 13498 13929
rect 13440 13889 13452 13923
rect 13486 13920 13498 13923
rect 13722 13920 13728 13932
rect 13486 13892 13728 13920
rect 13486 13889 13498 13892
rect 13440 13883 13498 13889
rect 13722 13880 13728 13892
rect 13780 13880 13786 13932
rect 13832 13920 13860 13948
rect 14918 13929 14924 13932
rect 14645 13923 14703 13929
rect 14645 13920 14657 13923
rect 13832 13892 14657 13920
rect 14645 13889 14657 13892
rect 14691 13889 14703 13923
rect 14912 13920 14924 13929
rect 14879 13892 14924 13920
rect 14645 13883 14703 13889
rect 14912 13883 14924 13892
rect 14918 13880 14924 13883
rect 14976 13880 14982 13932
rect 16298 13920 16304 13932
rect 16259 13892 16304 13920
rect 16298 13880 16304 13892
rect 16356 13880 16362 13932
rect 16390 13880 16396 13932
rect 16448 13920 16454 13932
rect 17604 13929 17632 14028
rect 19150 14016 19156 14028
rect 19208 14016 19214 14068
rect 19334 14016 19340 14068
rect 19392 14056 19398 14068
rect 19889 14059 19947 14065
rect 19889 14056 19901 14059
rect 19392 14028 19901 14056
rect 19392 14016 19398 14028
rect 19889 14025 19901 14028
rect 19935 14025 19947 14059
rect 19889 14019 19947 14025
rect 20070 14016 20076 14068
rect 20128 14056 20134 14068
rect 21361 14059 21419 14065
rect 21361 14056 21373 14059
rect 20128 14028 21373 14056
rect 20128 14016 20134 14028
rect 21361 14025 21373 14028
rect 21407 14056 21419 14059
rect 21637 14059 21695 14065
rect 21407 14028 21588 14056
rect 21407 14025 21419 14028
rect 21361 14019 21419 14025
rect 20714 13988 20720 14000
rect 18524 13960 20720 13988
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16448 13892 16681 13920
rect 16448 13880 16454 13892
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 17589 13923 17647 13929
rect 17589 13889 17601 13923
rect 17635 13889 17647 13923
rect 17589 13883 17647 13889
rect 17678 13880 17684 13932
rect 17736 13920 17742 13932
rect 17773 13923 17831 13929
rect 17773 13920 17785 13923
rect 17736 13892 17785 13920
rect 17736 13880 17742 13892
rect 17773 13889 17785 13892
rect 17819 13889 17831 13923
rect 17773 13883 17831 13889
rect 18138 13880 18144 13932
rect 18196 13920 18202 13932
rect 18524 13929 18552 13960
rect 18509 13923 18567 13929
rect 18509 13920 18521 13923
rect 18196 13892 18521 13920
rect 18196 13880 18202 13892
rect 18509 13889 18521 13892
rect 18555 13889 18567 13923
rect 18509 13883 18567 13889
rect 18776 13923 18834 13929
rect 18776 13889 18788 13923
rect 18822 13920 18834 13923
rect 19058 13920 19064 13932
rect 18822 13892 19064 13920
rect 18822 13889 18834 13892
rect 18776 13883 18834 13889
rect 19058 13880 19064 13892
rect 19116 13880 19122 13932
rect 19996 13929 20024 13960
rect 20714 13948 20720 13960
rect 20772 13988 20778 14000
rect 21266 13988 21272 14000
rect 20772 13960 21272 13988
rect 20772 13948 20778 13960
rect 21266 13948 21272 13960
rect 21324 13948 21330 14000
rect 19981 13923 20039 13929
rect 19981 13889 19993 13923
rect 20027 13889 20039 13923
rect 19981 13883 20039 13889
rect 20070 13880 20076 13932
rect 20128 13920 20134 13932
rect 20237 13923 20295 13929
rect 20237 13920 20249 13923
rect 20128 13892 20249 13920
rect 20128 13880 20134 13892
rect 20237 13889 20249 13892
rect 20283 13889 20295 13923
rect 20237 13883 20295 13889
rect 21453 13923 21511 13929
rect 21453 13889 21465 13923
rect 21499 13889 21511 13923
rect 21560 13920 21588 14028
rect 21637 14025 21649 14059
rect 21683 14025 21695 14059
rect 22094 14056 22100 14068
rect 22055 14028 22100 14056
rect 21637 14019 21695 14025
rect 21652 13988 21680 14019
rect 22094 14016 22100 14028
rect 22152 14016 22158 14068
rect 22189 14059 22247 14065
rect 22189 14025 22201 14059
rect 22235 14056 22247 14059
rect 22646 14056 22652 14068
rect 22235 14028 22652 14056
rect 22235 14025 22247 14028
rect 22189 14019 22247 14025
rect 22646 14016 22652 14028
rect 22704 14016 22710 14068
rect 22554 13988 22560 14000
rect 21652 13960 22560 13988
rect 22554 13948 22560 13960
rect 22612 13948 22618 14000
rect 21634 13920 21640 13932
rect 21560 13892 21640 13920
rect 21453 13883 21511 13889
rect 2866 13852 2872 13864
rect 2827 13824 2872 13852
rect 2866 13812 2872 13824
rect 2924 13812 2930 13864
rect 1670 13744 1676 13796
rect 1728 13784 1734 13796
rect 4264 13793 4292 13880
rect 5442 13812 5448 13864
rect 5500 13852 5506 13864
rect 6089 13855 6147 13861
rect 6089 13852 6101 13855
rect 5500 13824 6101 13852
rect 5500 13812 5506 13824
rect 6089 13821 6101 13824
rect 6135 13821 6147 13855
rect 6089 13815 6147 13821
rect 7193 13855 7251 13861
rect 7193 13821 7205 13855
rect 7239 13821 7251 13855
rect 7193 13815 7251 13821
rect 4249 13787 4307 13793
rect 1728 13756 2084 13784
rect 1728 13744 1734 13756
rect 1946 13716 1952 13728
rect 1907 13688 1952 13716
rect 1946 13676 1952 13688
rect 2004 13676 2010 13728
rect 2056 13716 2084 13756
rect 2746 13756 2912 13784
rect 2746 13716 2774 13756
rect 2056 13688 2774 13716
rect 2884 13716 2912 13756
rect 4249 13753 4261 13787
rect 4295 13753 4307 13787
rect 6178 13784 6184 13796
rect 4249 13747 4307 13753
rect 5276 13756 6184 13784
rect 5276 13716 5304 13756
rect 6178 13744 6184 13756
rect 6236 13744 6242 13796
rect 6270 13744 6276 13796
rect 6328 13784 6334 13796
rect 7208 13784 7236 13815
rect 8018 13812 8024 13864
rect 8076 13852 8082 13864
rect 8113 13855 8171 13861
rect 8113 13852 8125 13855
rect 8076 13824 8125 13852
rect 8076 13812 8082 13824
rect 8113 13821 8125 13824
rect 8159 13821 8171 13855
rect 8113 13815 8171 13821
rect 10321 13855 10379 13861
rect 10321 13821 10333 13855
rect 10367 13821 10379 13855
rect 10321 13815 10379 13821
rect 6328 13756 7236 13784
rect 6328 13744 6334 13756
rect 9674 13744 9680 13796
rect 9732 13784 9738 13796
rect 10336 13784 10364 13815
rect 10870 13812 10876 13864
rect 10928 13852 10934 13864
rect 10965 13855 11023 13861
rect 10965 13852 10977 13855
rect 10928 13824 10977 13852
rect 10928 13812 10934 13824
rect 10965 13821 10977 13824
rect 11011 13821 11023 13855
rect 10965 13815 11023 13821
rect 15746 13812 15752 13864
rect 15804 13852 15810 13864
rect 17313 13855 17371 13861
rect 17313 13852 17325 13855
rect 15804 13824 17325 13852
rect 15804 13812 15810 13824
rect 17313 13821 17325 13824
rect 17359 13821 17371 13855
rect 18414 13852 18420 13864
rect 18375 13824 18420 13852
rect 17313 13815 17371 13821
rect 18414 13812 18420 13824
rect 18472 13812 18478 13864
rect 21468 13852 21496 13883
rect 21634 13880 21640 13892
rect 21692 13880 21698 13932
rect 22186 13920 22192 13932
rect 21928 13892 22192 13920
rect 21928 13861 21956 13892
rect 22186 13880 22192 13892
rect 22244 13880 22250 13932
rect 22278 13880 22284 13932
rect 22336 13920 22342 13932
rect 22833 13923 22891 13929
rect 22833 13920 22845 13923
rect 22336 13892 22845 13920
rect 22336 13880 22342 13892
rect 22833 13889 22845 13892
rect 22879 13889 22891 13923
rect 23109 13923 23167 13929
rect 23109 13920 23121 13923
rect 22833 13883 22891 13889
rect 22940 13892 23121 13920
rect 21913 13855 21971 13861
rect 21468 13824 21864 13852
rect 17405 13787 17463 13793
rect 17405 13784 17417 13787
rect 9732 13756 11008 13784
rect 9732 13744 9738 13756
rect 10980 13728 11008 13756
rect 15764 13756 17417 13784
rect 2884 13688 5304 13716
rect 5810 13676 5816 13728
rect 5868 13716 5874 13728
rect 5868 13688 5913 13716
rect 5868 13676 5874 13688
rect 10962 13676 10968 13728
rect 11020 13676 11026 13728
rect 12434 13676 12440 13728
rect 12492 13716 12498 13728
rect 12894 13716 12900 13728
rect 12492 13688 12900 13716
rect 12492 13676 12498 13688
rect 12894 13676 12900 13688
rect 12952 13676 12958 13728
rect 15378 13676 15384 13728
rect 15436 13716 15442 13728
rect 15764 13716 15792 13756
rect 17405 13753 17417 13756
rect 17451 13753 17463 13787
rect 21836 13784 21864 13824
rect 21913 13821 21925 13855
rect 21959 13821 21971 13855
rect 21913 13815 21971 13821
rect 22554 13812 22560 13864
rect 22612 13852 22618 13864
rect 22940 13852 22968 13892
rect 23109 13889 23121 13892
rect 23155 13889 23167 13923
rect 23109 13883 23167 13889
rect 22612 13824 22968 13852
rect 22612 13812 22618 13824
rect 22830 13784 22836 13796
rect 21836 13756 22094 13784
rect 17405 13747 17463 13753
rect 16022 13716 16028 13728
rect 15436 13688 15792 13716
rect 15983 13688 16028 13716
rect 15436 13676 15442 13688
rect 16022 13676 16028 13688
rect 16080 13716 16086 13728
rect 16390 13716 16396 13728
rect 16080 13688 16396 13716
rect 16080 13676 16086 13688
rect 16390 13676 16396 13688
rect 16448 13676 16454 13728
rect 16574 13676 16580 13728
rect 16632 13716 16638 13728
rect 21450 13716 21456 13728
rect 16632 13688 21456 13716
rect 16632 13676 16638 13688
rect 21450 13676 21456 13688
rect 21508 13676 21514 13728
rect 22066 13716 22094 13756
rect 22204 13756 22836 13784
rect 22204 13716 22232 13756
rect 22830 13744 22836 13756
rect 22888 13744 22894 13796
rect 22066 13688 22232 13716
rect 22370 13676 22376 13728
rect 22428 13716 22434 13728
rect 22557 13719 22615 13725
rect 22557 13716 22569 13719
rect 22428 13688 22569 13716
rect 22428 13676 22434 13688
rect 22557 13685 22569 13688
rect 22603 13685 22615 13719
rect 22557 13679 22615 13685
rect 22649 13719 22707 13725
rect 22649 13685 22661 13719
rect 22695 13716 22707 13719
rect 22738 13716 22744 13728
rect 22695 13688 22744 13716
rect 22695 13685 22707 13688
rect 22649 13679 22707 13685
rect 22738 13676 22744 13688
rect 22796 13676 22802 13728
rect 22922 13716 22928 13728
rect 22883 13688 22928 13716
rect 22922 13676 22928 13688
rect 22980 13676 22986 13728
rect 1104 13626 23460 13648
rect 1104 13574 3749 13626
rect 3801 13574 3813 13626
rect 3865 13574 3877 13626
rect 3929 13574 3941 13626
rect 3993 13574 4005 13626
rect 4057 13574 9347 13626
rect 9399 13574 9411 13626
rect 9463 13574 9475 13626
rect 9527 13574 9539 13626
rect 9591 13574 9603 13626
rect 9655 13574 14945 13626
rect 14997 13574 15009 13626
rect 15061 13574 15073 13626
rect 15125 13574 15137 13626
rect 15189 13574 15201 13626
rect 15253 13574 20543 13626
rect 20595 13574 20607 13626
rect 20659 13574 20671 13626
rect 20723 13574 20735 13626
rect 20787 13574 20799 13626
rect 20851 13574 23460 13626
rect 1104 13552 23460 13574
rect 2498 13472 2504 13524
rect 2556 13512 2562 13524
rect 5626 13512 5632 13524
rect 2556 13484 5212 13512
rect 5587 13484 5632 13512
rect 2556 13472 2562 13484
rect 3513 13447 3571 13453
rect 3513 13413 3525 13447
rect 3559 13444 3571 13447
rect 4525 13447 4583 13453
rect 3559 13416 3924 13444
rect 3559 13413 3571 13416
rect 3513 13407 3571 13413
rect 3896 13388 3924 13416
rect 4525 13413 4537 13447
rect 4571 13444 4583 13447
rect 5074 13444 5080 13456
rect 4571 13416 5080 13444
rect 4571 13413 4583 13416
rect 4525 13407 4583 13413
rect 5074 13404 5080 13416
rect 5132 13404 5138 13456
rect 3878 13376 3884 13388
rect 3791 13348 3884 13376
rect 3878 13336 3884 13348
rect 3936 13336 3942 13388
rect 5184 13385 5212 13484
rect 5626 13472 5632 13484
rect 5684 13472 5690 13524
rect 7006 13512 7012 13524
rect 6967 13484 7012 13512
rect 7006 13472 7012 13484
rect 7064 13472 7070 13524
rect 9309 13515 9367 13521
rect 9309 13481 9321 13515
rect 9355 13512 9367 13515
rect 10502 13512 10508 13524
rect 9355 13484 10508 13512
rect 9355 13481 9367 13484
rect 9309 13475 9367 13481
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 11885 13515 11943 13521
rect 11885 13481 11897 13515
rect 11931 13512 11943 13515
rect 12066 13512 12072 13524
rect 11931 13484 12072 13512
rect 11931 13481 11943 13484
rect 11885 13475 11943 13481
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 13909 13515 13967 13521
rect 13909 13481 13921 13515
rect 13955 13512 13967 13515
rect 14366 13512 14372 13524
rect 13955 13484 14372 13512
rect 13955 13481 13967 13484
rect 13909 13475 13967 13481
rect 14366 13472 14372 13484
rect 14424 13512 14430 13524
rect 14734 13512 14740 13524
rect 14424 13484 14740 13512
rect 14424 13472 14430 13484
rect 14734 13472 14740 13484
rect 14792 13472 14798 13524
rect 16117 13515 16175 13521
rect 16117 13481 16129 13515
rect 16163 13512 16175 13515
rect 16298 13512 16304 13524
rect 16163 13484 16304 13512
rect 16163 13481 16175 13484
rect 16117 13475 16175 13481
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 19337 13515 19395 13521
rect 19337 13481 19349 13515
rect 19383 13512 19395 13515
rect 19610 13512 19616 13524
rect 19383 13484 19616 13512
rect 19383 13481 19395 13484
rect 19337 13475 19395 13481
rect 19610 13472 19616 13484
rect 19668 13472 19674 13524
rect 19720 13484 22232 13512
rect 8481 13447 8539 13453
rect 8481 13413 8493 13447
rect 8527 13444 8539 13447
rect 9950 13444 9956 13456
rect 8527 13416 9956 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 9950 13404 9956 13416
rect 10008 13404 10014 13456
rect 10137 13447 10195 13453
rect 10137 13413 10149 13447
rect 10183 13444 10195 13447
rect 10226 13444 10232 13456
rect 10183 13416 10232 13444
rect 10183 13413 10195 13416
rect 10137 13407 10195 13413
rect 10226 13404 10232 13416
rect 10284 13404 10290 13456
rect 11974 13404 11980 13456
rect 12032 13444 12038 13456
rect 12345 13447 12403 13453
rect 12345 13444 12357 13447
rect 12032 13416 12357 13444
rect 12032 13404 12038 13416
rect 12345 13413 12357 13416
rect 12391 13413 12403 13447
rect 12345 13407 12403 13413
rect 5169 13379 5227 13385
rect 5169 13345 5181 13379
rect 5215 13345 5227 13379
rect 9490 13376 9496 13388
rect 9451 13348 9496 13376
rect 5169 13339 5227 13345
rect 9490 13336 9496 13348
rect 9548 13336 9554 13388
rect 9582 13336 9588 13388
rect 9640 13376 9646 13388
rect 18782 13376 18788 13388
rect 9640 13348 10272 13376
rect 18743 13348 18788 13376
rect 9640 13336 9646 13348
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 2038 13268 2044 13320
rect 2096 13308 2102 13320
rect 2133 13311 2191 13317
rect 2133 13308 2145 13311
rect 2096 13280 2145 13308
rect 2096 13268 2102 13280
rect 2133 13277 2145 13280
rect 2179 13308 2191 13311
rect 2866 13308 2872 13320
rect 2179 13280 2872 13308
rect 2179 13277 2191 13280
rect 2133 13271 2191 13277
rect 2866 13268 2872 13280
rect 2924 13268 2930 13320
rect 4154 13308 4160 13320
rect 4115 13280 4160 13308
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 4246 13268 4252 13320
rect 4304 13308 4310 13320
rect 5077 13311 5135 13317
rect 5077 13308 5089 13311
rect 4304 13280 5089 13308
rect 4304 13268 4310 13280
rect 5077 13277 5089 13280
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 6086 13268 6092 13320
rect 6144 13308 6150 13320
rect 6273 13311 6331 13317
rect 6273 13308 6285 13311
rect 6144 13280 6285 13308
rect 6144 13268 6150 13280
rect 6273 13277 6285 13280
rect 6319 13277 6331 13311
rect 6273 13271 6331 13277
rect 6362 13268 6368 13320
rect 6420 13308 6426 13320
rect 7098 13308 7104 13320
rect 6420 13280 6465 13308
rect 7059 13280 7104 13308
rect 6420 13268 6426 13280
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 7190 13268 7196 13320
rect 7248 13308 7254 13320
rect 7357 13311 7415 13317
rect 7357 13308 7369 13311
rect 7248 13280 7369 13308
rect 7248 13268 7254 13280
rect 7357 13277 7369 13280
rect 7403 13277 7415 13311
rect 7357 13271 7415 13277
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13308 8815 13311
rect 8938 13308 8944 13320
rect 8803 13280 8944 13308
rect 8803 13277 8815 13280
rect 8757 13271 8815 13277
rect 8938 13268 8944 13280
rect 8996 13268 9002 13320
rect 9125 13311 9183 13317
rect 9125 13277 9137 13311
rect 9171 13308 9183 13311
rect 10134 13308 10140 13320
rect 9171 13280 10140 13308
rect 9171 13277 9183 13280
rect 9125 13271 9183 13277
rect 10134 13268 10140 13280
rect 10192 13268 10198 13320
rect 10244 13317 10272 13348
rect 18782 13336 18788 13348
rect 18840 13336 18846 13388
rect 19058 13376 19064 13388
rect 19019 13348 19064 13376
rect 19058 13336 19064 13348
rect 19116 13336 19122 13388
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 10505 13311 10563 13317
rect 10505 13277 10517 13311
rect 10551 13277 10563 13311
rect 10505 13271 10563 13277
rect 1946 13200 1952 13252
rect 2004 13240 2010 13252
rect 2378 13243 2436 13249
rect 2378 13240 2390 13243
rect 2004 13212 2390 13240
rect 2004 13200 2010 13212
rect 2378 13209 2390 13212
rect 2424 13209 2436 13243
rect 2378 13203 2436 13209
rect 4065 13243 4123 13249
rect 4065 13209 4077 13243
rect 4111 13240 4123 13243
rect 4111 13212 4660 13240
rect 4111 13209 4123 13212
rect 4065 13203 4123 13209
rect 2041 13175 2099 13181
rect 2041 13141 2053 13175
rect 2087 13172 2099 13175
rect 2130 13172 2136 13184
rect 2087 13144 2136 13172
rect 2087 13141 2099 13144
rect 2041 13135 2099 13141
rect 2130 13132 2136 13144
rect 2188 13132 2194 13184
rect 4632 13181 4660 13212
rect 7742 13200 7748 13252
rect 7800 13240 7806 13252
rect 10520 13240 10548 13271
rect 11882 13268 11888 13320
rect 11940 13308 11946 13320
rect 11977 13311 12035 13317
rect 11977 13308 11989 13311
rect 11940 13280 11989 13308
rect 11940 13268 11946 13280
rect 11977 13277 11989 13280
rect 12023 13277 12035 13311
rect 11977 13271 12035 13277
rect 12161 13311 12219 13317
rect 12161 13277 12173 13311
rect 12207 13308 12219 13311
rect 12434 13308 12440 13320
rect 12207 13280 12440 13308
rect 12207 13277 12219 13280
rect 12161 13271 12219 13277
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 12529 13311 12587 13317
rect 12529 13277 12541 13311
rect 12575 13308 12587 13311
rect 13814 13308 13820 13320
rect 12575 13280 13820 13308
rect 12575 13277 12587 13280
rect 12529 13271 12587 13277
rect 13814 13268 13820 13280
rect 13872 13308 13878 13320
rect 14734 13308 14740 13320
rect 13872 13280 14740 13308
rect 13872 13268 13878 13280
rect 14734 13268 14740 13280
rect 14792 13268 14798 13320
rect 15004 13311 15062 13317
rect 15004 13277 15016 13311
rect 15050 13308 15062 13311
rect 15746 13308 15752 13320
rect 15050 13280 15752 13308
rect 15050 13277 15062 13280
rect 15004 13271 15062 13277
rect 15746 13268 15752 13280
rect 15804 13268 15810 13320
rect 16298 13268 16304 13320
rect 16356 13308 16362 13320
rect 16853 13311 16911 13317
rect 16853 13308 16865 13311
rect 16356 13280 16865 13308
rect 16356 13268 16362 13280
rect 16853 13277 16865 13280
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 16942 13268 16948 13320
rect 17000 13308 17006 13320
rect 17037 13311 17095 13317
rect 17037 13308 17049 13311
rect 17000 13280 17049 13308
rect 17000 13268 17006 13280
rect 17037 13277 17049 13280
rect 17083 13277 17095 13311
rect 17037 13271 17095 13277
rect 17126 13268 17132 13320
rect 17184 13308 17190 13320
rect 17773 13311 17831 13317
rect 17773 13308 17785 13311
rect 17184 13280 17785 13308
rect 17184 13268 17190 13280
rect 17773 13277 17785 13280
rect 17819 13277 17831 13311
rect 17773 13271 17831 13277
rect 7800 13212 10548 13240
rect 7800 13200 7806 13212
rect 10594 13200 10600 13252
rect 10652 13240 10658 13252
rect 12802 13249 12808 13252
rect 10750 13243 10808 13249
rect 10750 13240 10762 13243
rect 10652 13212 10762 13240
rect 10652 13200 10658 13212
rect 10750 13209 10762 13212
rect 10796 13209 10808 13243
rect 12796 13240 12808 13249
rect 10750 13203 10808 13209
rect 12084 13212 12434 13240
rect 12763 13212 12808 13240
rect 4617 13175 4675 13181
rect 4617 13141 4629 13175
rect 4663 13141 4675 13175
rect 4982 13172 4988 13184
rect 4943 13144 4988 13172
rect 4617 13135 4675 13141
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 5810 13132 5816 13184
rect 5868 13172 5874 13184
rect 8202 13172 8208 13184
rect 5868 13144 8208 13172
rect 5868 13132 5874 13144
rect 8202 13132 8208 13144
rect 8260 13132 8266 13184
rect 8570 13172 8576 13184
rect 8531 13144 8576 13172
rect 8570 13132 8576 13144
rect 8628 13132 8634 13184
rect 9674 13172 9680 13184
rect 9635 13144 9680 13172
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 10413 13175 10471 13181
rect 9824 13144 9869 13172
rect 9824 13132 9830 13144
rect 10413 13141 10425 13175
rect 10459 13172 10471 13175
rect 11146 13172 11152 13184
rect 10459 13144 11152 13172
rect 10459 13141 10471 13144
rect 10413 13135 10471 13141
rect 11146 13132 11152 13144
rect 11204 13132 11210 13184
rect 11698 13132 11704 13184
rect 11756 13172 11762 13184
rect 12084 13172 12112 13212
rect 11756 13144 12112 13172
rect 12406 13172 12434 13212
rect 12796 13203 12808 13212
rect 12802 13200 12808 13203
rect 12860 13200 12866 13252
rect 19720 13240 19748 13484
rect 21174 13444 21180 13456
rect 20364 13416 21180 13444
rect 19978 13308 19984 13320
rect 19939 13280 19984 13308
rect 19978 13268 19984 13280
rect 20036 13268 20042 13320
rect 20364 13317 20392 13416
rect 21174 13404 21180 13416
rect 21232 13404 21238 13456
rect 22204 13444 22232 13484
rect 22462 13472 22468 13524
rect 22520 13512 22526 13524
rect 22649 13515 22707 13521
rect 22649 13512 22661 13515
rect 22520 13484 22661 13512
rect 22520 13472 22526 13484
rect 22649 13481 22661 13484
rect 22695 13481 22707 13515
rect 22649 13475 22707 13481
rect 22830 13472 22836 13524
rect 22888 13512 22894 13524
rect 23750 13512 23756 13524
rect 22888 13484 23756 13512
rect 22888 13472 22894 13484
rect 23750 13472 23756 13484
rect 23808 13472 23814 13524
rect 22925 13447 22983 13453
rect 22925 13444 22937 13447
rect 22204 13416 22937 13444
rect 22925 13413 22937 13416
rect 22971 13413 22983 13447
rect 22925 13407 22983 13413
rect 21082 13376 21088 13388
rect 21043 13348 21088 13376
rect 21082 13336 21088 13348
rect 21140 13336 21146 13388
rect 21266 13376 21272 13388
rect 21227 13348 21272 13376
rect 21266 13336 21272 13348
rect 21324 13336 21330 13388
rect 20349 13311 20407 13317
rect 20349 13277 20361 13311
rect 20395 13277 20407 13311
rect 20349 13271 20407 13277
rect 20809 13311 20867 13317
rect 20809 13277 20821 13311
rect 20855 13308 20867 13311
rect 22646 13308 22652 13320
rect 20855 13280 22652 13308
rect 20855 13277 20867 13280
rect 20809 13271 20867 13277
rect 22646 13268 22652 13280
rect 22704 13268 22710 13320
rect 23106 13308 23112 13320
rect 23067 13280 23112 13308
rect 23106 13268 23112 13280
rect 23164 13268 23170 13320
rect 16132 13212 19748 13240
rect 16132 13172 16160 13212
rect 21358 13200 21364 13252
rect 21416 13240 21422 13252
rect 21514 13243 21572 13249
rect 21514 13240 21526 13243
rect 21416 13212 21526 13240
rect 21416 13200 21422 13212
rect 21514 13209 21526 13212
rect 21560 13209 21572 13243
rect 21514 13203 21572 13209
rect 22002 13200 22008 13252
rect 22060 13240 22066 13252
rect 22922 13240 22928 13252
rect 22060 13212 22928 13240
rect 22060 13200 22066 13212
rect 22922 13200 22928 13212
rect 22980 13200 22986 13252
rect 12406 13144 16160 13172
rect 11756 13132 11762 13144
rect 16206 13132 16212 13184
rect 16264 13172 16270 13184
rect 17681 13175 17739 13181
rect 16264 13144 16309 13172
rect 16264 13132 16270 13144
rect 17681 13141 17693 13175
rect 17727 13172 17739 13175
rect 18230 13172 18236 13184
rect 17727 13144 18236 13172
rect 17727 13141 17739 13144
rect 17681 13135 17739 13141
rect 18230 13132 18236 13144
rect 18288 13132 18294 13184
rect 18322 13132 18328 13184
rect 18380 13172 18386 13184
rect 18417 13175 18475 13181
rect 18417 13172 18429 13175
rect 18380 13144 18429 13172
rect 18380 13132 18386 13144
rect 18417 13141 18429 13144
rect 18463 13141 18475 13175
rect 18417 13135 18475 13141
rect 20165 13175 20223 13181
rect 20165 13141 20177 13175
rect 20211 13172 20223 13175
rect 20254 13172 20260 13184
rect 20211 13144 20260 13172
rect 20211 13141 20223 13144
rect 20165 13135 20223 13141
rect 20254 13132 20260 13144
rect 20312 13132 20318 13184
rect 20438 13172 20444 13184
rect 20399 13144 20444 13172
rect 20438 13132 20444 13144
rect 20496 13132 20502 13184
rect 20901 13175 20959 13181
rect 20901 13141 20913 13175
rect 20947 13172 20959 13175
rect 21818 13172 21824 13184
rect 20947 13144 21824 13172
rect 20947 13141 20959 13144
rect 20901 13135 20959 13141
rect 21818 13132 21824 13144
rect 21876 13132 21882 13184
rect 1104 13082 23460 13104
rect 1104 13030 6548 13082
rect 6600 13030 6612 13082
rect 6664 13030 6676 13082
rect 6728 13030 6740 13082
rect 6792 13030 6804 13082
rect 6856 13030 12146 13082
rect 12198 13030 12210 13082
rect 12262 13030 12274 13082
rect 12326 13030 12338 13082
rect 12390 13030 12402 13082
rect 12454 13030 17744 13082
rect 17796 13030 17808 13082
rect 17860 13030 17872 13082
rect 17924 13030 17936 13082
rect 17988 13030 18000 13082
rect 18052 13030 23460 13082
rect 1104 13008 23460 13030
rect 1857 12971 1915 12977
rect 1857 12937 1869 12971
rect 1903 12968 1915 12971
rect 2498 12968 2504 12980
rect 1903 12940 2504 12968
rect 1903 12937 1915 12940
rect 1857 12931 1915 12937
rect 2498 12928 2504 12940
rect 2556 12928 2562 12980
rect 3510 12968 3516 12980
rect 3471 12940 3516 12968
rect 3510 12928 3516 12940
rect 3568 12928 3574 12980
rect 5445 12971 5503 12977
rect 5445 12937 5457 12971
rect 5491 12968 5503 12971
rect 5994 12968 6000 12980
rect 5491 12940 6000 12968
rect 5491 12937 5503 12940
rect 5445 12931 5503 12937
rect 5994 12928 6000 12940
rect 6052 12928 6058 12980
rect 6089 12971 6147 12977
rect 6089 12937 6101 12971
rect 6135 12968 6147 12971
rect 6454 12968 6460 12980
rect 6135 12940 6460 12968
rect 6135 12937 6147 12940
rect 6089 12931 6147 12937
rect 6454 12928 6460 12940
rect 6512 12928 6518 12980
rect 8757 12971 8815 12977
rect 8757 12937 8769 12971
rect 8803 12968 8815 12971
rect 9309 12971 9367 12977
rect 9309 12968 9321 12971
rect 8803 12940 9321 12968
rect 8803 12937 8815 12940
rect 8757 12931 8815 12937
rect 9309 12937 9321 12940
rect 9355 12937 9367 12971
rect 9309 12931 9367 12937
rect 9769 12971 9827 12977
rect 9769 12937 9781 12971
rect 9815 12968 9827 12971
rect 9950 12968 9956 12980
rect 9815 12940 9956 12968
rect 9815 12937 9827 12940
rect 9769 12931 9827 12937
rect 9950 12928 9956 12940
rect 10008 12928 10014 12980
rect 10134 12968 10140 12980
rect 10095 12940 10140 12968
rect 10134 12928 10140 12940
rect 10192 12928 10198 12980
rect 10505 12971 10563 12977
rect 10505 12937 10517 12971
rect 10551 12968 10563 12971
rect 11517 12971 11575 12977
rect 11517 12968 11529 12971
rect 10551 12940 11529 12968
rect 10551 12937 10563 12940
rect 10505 12931 10563 12937
rect 11517 12937 11529 12940
rect 11563 12937 11575 12971
rect 11517 12931 11575 12937
rect 11885 12971 11943 12977
rect 11885 12937 11897 12971
rect 11931 12968 11943 12971
rect 12066 12968 12072 12980
rect 11931 12940 12072 12968
rect 11931 12937 11943 12940
rect 11885 12931 11943 12937
rect 12066 12928 12072 12940
rect 12124 12928 12130 12980
rect 12526 12928 12532 12980
rect 12584 12968 12590 12980
rect 15286 12968 15292 12980
rect 12584 12940 15292 12968
rect 12584 12928 12590 12940
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 18506 12968 18512 12980
rect 16500 12940 18512 12968
rect 2866 12860 2872 12912
rect 2924 12900 2930 12912
rect 2924 12872 3280 12900
rect 2924 12860 2930 12872
rect 2981 12835 3039 12841
rect 2981 12801 2993 12835
rect 3027 12832 3039 12835
rect 3142 12832 3148 12844
rect 3027 12804 3148 12832
rect 3027 12801 3039 12804
rect 2981 12795 3039 12801
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 3252 12841 3280 12872
rect 4614 12860 4620 12912
rect 4672 12900 4678 12912
rect 5810 12909 5816 12912
rect 5629 12903 5687 12909
rect 5629 12900 5641 12903
rect 4672 12872 5641 12900
rect 4672 12860 4678 12872
rect 5629 12869 5641 12872
rect 5675 12869 5687 12903
rect 5629 12863 5687 12869
rect 5794 12903 5816 12909
rect 5794 12869 5806 12903
rect 5794 12863 5816 12869
rect 5810 12860 5816 12863
rect 5868 12860 5874 12912
rect 6178 12860 6184 12912
rect 6236 12900 6242 12912
rect 6236 12872 6868 12900
rect 6236 12860 6242 12872
rect 3237 12835 3295 12841
rect 3237 12801 3249 12835
rect 3283 12801 3295 12835
rect 3237 12795 3295 12801
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 4157 12835 4215 12841
rect 4157 12832 4169 12835
rect 3936 12804 4169 12832
rect 3936 12792 3942 12804
rect 4157 12801 4169 12804
rect 4203 12801 4215 12835
rect 4157 12795 4215 12801
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12832 4859 12835
rect 5350 12832 5356 12844
rect 4847 12804 5356 12832
rect 4847 12801 4859 12804
rect 4801 12795 4859 12801
rect 5350 12792 5356 12804
rect 5408 12832 5414 12844
rect 6840 12841 6868 12872
rect 7098 12860 7104 12912
rect 7156 12900 7162 12912
rect 7742 12900 7748 12912
rect 7156 12872 7748 12900
rect 7156 12860 7162 12872
rect 7742 12860 7748 12872
rect 7800 12900 7806 12912
rect 7800 12872 8432 12900
rect 7800 12860 7806 12872
rect 5905 12835 5963 12841
rect 5905 12832 5917 12835
rect 5408 12804 5917 12832
rect 5408 12792 5414 12804
rect 5905 12801 5917 12804
rect 5951 12801 5963 12835
rect 5905 12795 5963 12801
rect 6365 12835 6423 12841
rect 6365 12801 6377 12835
rect 6411 12801 6423 12835
rect 6365 12795 6423 12801
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 4246 12724 4252 12776
rect 4304 12764 4310 12776
rect 4893 12767 4951 12773
rect 4893 12764 4905 12767
rect 4304 12736 4905 12764
rect 4304 12724 4310 12736
rect 4893 12733 4905 12736
rect 4939 12733 4951 12767
rect 4893 12727 4951 12733
rect 5077 12767 5135 12773
rect 5077 12733 5089 12767
rect 5123 12764 5135 12767
rect 5718 12764 5724 12776
rect 5123 12736 5724 12764
rect 5123 12733 5135 12736
rect 5077 12727 5135 12733
rect 5718 12724 5724 12736
rect 5776 12724 5782 12776
rect 6380 12764 6408 12795
rect 8110 12792 8116 12844
rect 8168 12841 8174 12844
rect 8404 12841 8432 12872
rect 8570 12860 8576 12912
rect 8628 12900 8634 12912
rect 9582 12900 9588 12912
rect 8628 12872 9588 12900
rect 8628 12860 8634 12872
rect 9582 12860 9588 12872
rect 9640 12900 9646 12912
rect 10597 12903 10655 12909
rect 9640 12872 9904 12900
rect 9640 12860 9646 12872
rect 8168 12832 8180 12841
rect 8389 12835 8447 12841
rect 8168 12804 8213 12832
rect 8168 12795 8180 12804
rect 8389 12801 8401 12835
rect 8435 12801 8447 12835
rect 8846 12832 8852 12844
rect 8807 12804 8852 12832
rect 8389 12795 8447 12801
rect 8168 12792 8174 12795
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 9677 12835 9735 12841
rect 9677 12801 9689 12835
rect 9723 12801 9735 12835
rect 9677 12795 9735 12801
rect 5828 12736 6408 12764
rect 8665 12767 8723 12773
rect 4338 12656 4344 12708
rect 4396 12696 4402 12708
rect 5828 12696 5856 12736
rect 8665 12733 8677 12767
rect 8711 12764 8723 12767
rect 8754 12764 8760 12776
rect 8711 12736 8760 12764
rect 8711 12733 8723 12736
rect 8665 12727 8723 12733
rect 8754 12724 8760 12736
rect 8812 12724 8818 12776
rect 9692 12764 9720 12795
rect 9876 12773 9904 12872
rect 10597 12869 10609 12903
rect 10643 12900 10655 12903
rect 11606 12900 11612 12912
rect 10643 12872 11612 12900
rect 10643 12869 10655 12872
rect 10597 12863 10655 12869
rect 11606 12860 11612 12872
rect 11664 12860 11670 12912
rect 13664 12903 13722 12909
rect 13664 12869 13676 12903
rect 13710 12900 13722 12903
rect 14366 12900 14372 12912
rect 13710 12872 14228 12900
rect 14327 12872 14372 12900
rect 13710 12869 13722 12872
rect 13664 12863 13722 12869
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12832 11207 12835
rect 11514 12832 11520 12844
rect 11195 12804 11520 12832
rect 11195 12801 11207 12804
rect 11149 12795 11207 12801
rect 11514 12792 11520 12804
rect 11572 12792 11578 12844
rect 13814 12792 13820 12844
rect 13872 12832 13878 12844
rect 13909 12835 13967 12841
rect 13909 12832 13921 12835
rect 13872 12804 13921 12832
rect 13872 12792 13878 12804
rect 13909 12801 13921 12804
rect 13955 12801 13967 12835
rect 14200 12832 14228 12872
rect 14366 12860 14372 12872
rect 14424 12860 14430 12912
rect 15197 12903 15255 12909
rect 15197 12869 15209 12903
rect 15243 12900 15255 12903
rect 16022 12900 16028 12912
rect 15243 12872 16028 12900
rect 15243 12869 15255 12872
rect 15197 12863 15255 12869
rect 16022 12860 16028 12872
rect 16080 12860 16086 12912
rect 14642 12832 14648 12844
rect 14200 12804 14648 12832
rect 13909 12795 13967 12801
rect 14642 12792 14648 12804
rect 14700 12792 14706 12844
rect 15289 12835 15347 12841
rect 15289 12801 15301 12835
rect 15335 12832 15347 12835
rect 15470 12832 15476 12844
rect 15335 12804 15476 12832
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 15470 12792 15476 12804
rect 15528 12792 15534 12844
rect 16500 12841 16528 12940
rect 18506 12928 18512 12940
rect 18564 12928 18570 12980
rect 18598 12928 18604 12980
rect 18656 12968 18662 12980
rect 18877 12971 18935 12977
rect 18877 12968 18889 12971
rect 18656 12940 18889 12968
rect 18656 12928 18662 12940
rect 18877 12937 18889 12940
rect 18923 12937 18935 12971
rect 18877 12931 18935 12937
rect 19613 12971 19671 12977
rect 19613 12937 19625 12971
rect 19659 12968 19671 12971
rect 20070 12968 20076 12980
rect 19659 12940 20076 12968
rect 19659 12937 19671 12940
rect 19613 12931 19671 12937
rect 18138 12900 18144 12912
rect 17512 12872 18144 12900
rect 16485 12835 16543 12841
rect 16485 12801 16497 12835
rect 16531 12801 16543 12835
rect 16485 12795 16543 12801
rect 16574 12792 16580 12844
rect 16632 12832 16638 12844
rect 17512 12841 17540 12872
rect 18138 12860 18144 12872
rect 18196 12860 18202 12912
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 16632 12804 17049 12832
rect 16632 12792 16638 12804
rect 17037 12801 17049 12804
rect 17083 12801 17095 12835
rect 17037 12795 17095 12801
rect 17497 12835 17555 12841
rect 17497 12801 17509 12835
rect 17543 12801 17555 12835
rect 17497 12795 17555 12801
rect 17764 12835 17822 12841
rect 17764 12801 17776 12835
rect 17810 12832 17822 12835
rect 18892 12832 18920 12931
rect 20070 12928 20076 12940
rect 20128 12928 20134 12980
rect 20257 12971 20315 12977
rect 20257 12937 20269 12971
rect 20303 12968 20315 12971
rect 21082 12968 21088 12980
rect 20303 12940 21088 12968
rect 20303 12937 20315 12940
rect 20257 12931 20315 12937
rect 21082 12928 21088 12940
rect 21140 12928 21146 12980
rect 21818 12968 21824 12980
rect 21779 12940 21824 12968
rect 21818 12928 21824 12940
rect 21876 12928 21882 12980
rect 22646 12968 22652 12980
rect 22607 12940 22652 12968
rect 22646 12928 22652 12940
rect 22704 12928 22710 12980
rect 21266 12860 21272 12912
rect 21324 12900 21330 12912
rect 21324 12872 21680 12900
rect 21324 12860 21330 12872
rect 18969 12835 19027 12841
rect 18969 12832 18981 12835
rect 17810 12804 18828 12832
rect 18892 12804 18981 12832
rect 17810 12801 17822 12804
rect 17764 12795 17822 12801
rect 8864 12736 9720 12764
rect 9861 12767 9919 12773
rect 4396 12668 5856 12696
rect 4396 12656 4402 12668
rect 6362 12656 6368 12708
rect 6420 12696 6426 12708
rect 6641 12699 6699 12705
rect 6641 12696 6653 12699
rect 6420 12668 6653 12696
rect 6420 12656 6426 12668
rect 6641 12665 6653 12668
rect 6687 12665 6699 12699
rect 6641 12659 6699 12665
rect 4430 12628 4436 12640
rect 4391 12600 4436 12628
rect 4430 12588 4436 12600
rect 4488 12588 4494 12640
rect 6454 12588 6460 12640
rect 6512 12628 6518 12640
rect 6549 12631 6607 12637
rect 6549 12628 6561 12631
rect 6512 12600 6561 12628
rect 6512 12588 6518 12600
rect 6549 12597 6561 12600
rect 6595 12597 6607 12631
rect 6549 12591 6607 12597
rect 7009 12631 7067 12637
rect 7009 12597 7021 12631
rect 7055 12628 7067 12631
rect 7466 12628 7472 12640
rect 7055 12600 7472 12628
rect 7055 12597 7067 12600
rect 7009 12591 7067 12597
rect 7466 12588 7472 12600
rect 7524 12628 7530 12640
rect 8864 12628 8892 12736
rect 9861 12733 9873 12767
rect 9907 12733 9919 12767
rect 9861 12727 9919 12733
rect 10781 12767 10839 12773
rect 10781 12733 10793 12767
rect 10827 12764 10839 12767
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 10827 12736 10977 12764
rect 10827 12733 10839 12736
rect 10781 12727 10839 12733
rect 10965 12733 10977 12736
rect 11011 12733 11023 12767
rect 11974 12764 11980 12776
rect 11935 12736 11980 12764
rect 10965 12727 11023 12733
rect 9030 12656 9036 12708
rect 9088 12696 9094 12708
rect 10796 12696 10824 12727
rect 11974 12724 11980 12736
rect 12032 12724 12038 12776
rect 12066 12724 12072 12776
rect 12124 12764 12130 12776
rect 12124 12736 12169 12764
rect 12124 12724 12130 12736
rect 13998 12724 14004 12776
rect 14056 12764 14062 12776
rect 14182 12764 14188 12776
rect 14056 12736 14188 12764
rect 14056 12724 14062 12736
rect 14182 12724 14188 12736
rect 14240 12724 14246 12776
rect 14277 12767 14335 12773
rect 14277 12733 14289 12767
rect 14323 12733 14335 12767
rect 15378 12764 15384 12776
rect 15339 12736 15384 12764
rect 14277 12727 14335 12733
rect 9088 12668 10824 12696
rect 9088 12656 9094 12668
rect 11146 12656 11152 12708
rect 11204 12696 11210 12708
rect 12084 12696 12112 12724
rect 11204 12668 12112 12696
rect 12529 12699 12587 12705
rect 11204 12656 11210 12668
rect 12529 12665 12541 12699
rect 12575 12696 12587 12699
rect 12618 12696 12624 12708
rect 12575 12668 12624 12696
rect 12575 12665 12587 12668
rect 12529 12659 12587 12665
rect 12618 12656 12624 12668
rect 12676 12656 12682 12708
rect 14292 12696 14320 12727
rect 15378 12724 15384 12736
rect 15436 12724 15442 12776
rect 16850 12764 16856 12776
rect 16811 12736 16856 12764
rect 16850 12724 16856 12736
rect 16908 12724 16914 12776
rect 16945 12767 17003 12773
rect 16945 12733 16957 12767
rect 16991 12764 17003 12767
rect 17310 12764 17316 12776
rect 16991 12736 17316 12764
rect 16991 12733 17003 12736
rect 16945 12727 17003 12733
rect 17310 12724 17316 12736
rect 17368 12724 17374 12776
rect 18800 12764 18828 12804
rect 18969 12801 18981 12804
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 19702 12792 19708 12844
rect 19760 12832 19766 12844
rect 19797 12835 19855 12841
rect 19797 12832 19809 12835
rect 19760 12804 19809 12832
rect 19760 12792 19766 12804
rect 19797 12801 19809 12804
rect 19843 12801 19855 12835
rect 19797 12795 19855 12801
rect 21381 12835 21439 12841
rect 21381 12801 21393 12835
rect 21427 12832 21439 12835
rect 21542 12832 21548 12844
rect 21427 12804 21548 12832
rect 21427 12801 21439 12804
rect 21381 12795 21439 12801
rect 21542 12792 21548 12804
rect 21600 12792 21606 12844
rect 21652 12841 21680 12872
rect 21637 12835 21695 12841
rect 21637 12801 21649 12835
rect 21683 12832 21695 12835
rect 21726 12832 21732 12844
rect 21683 12804 21732 12832
rect 21683 12801 21695 12804
rect 21637 12795 21695 12801
rect 21726 12792 21732 12804
rect 21784 12792 21790 12844
rect 22189 12835 22247 12841
rect 22189 12801 22201 12835
rect 22235 12832 22247 12835
rect 22370 12832 22376 12844
rect 22235 12804 22376 12832
rect 22235 12801 22247 12804
rect 22189 12795 22247 12801
rect 22370 12792 22376 12804
rect 22428 12792 22434 12844
rect 22830 12792 22836 12844
rect 22888 12832 22894 12844
rect 23109 12835 23167 12841
rect 23109 12832 23121 12835
rect 22888 12804 23121 12832
rect 22888 12792 22894 12804
rect 23109 12801 23121 12804
rect 23155 12801 23167 12835
rect 23109 12795 23167 12801
rect 19886 12764 19892 12776
rect 18800 12736 19892 12764
rect 19886 12724 19892 12736
rect 19944 12724 19950 12776
rect 21818 12724 21824 12776
rect 21876 12764 21882 12776
rect 22281 12767 22339 12773
rect 22281 12764 22293 12767
rect 21876 12736 22293 12764
rect 21876 12724 21882 12736
rect 22281 12733 22293 12736
rect 22327 12733 22339 12767
rect 22462 12764 22468 12776
rect 22423 12736 22468 12764
rect 22281 12727 22339 12733
rect 22462 12724 22468 12736
rect 22520 12724 22526 12776
rect 14200 12668 14320 12696
rect 17236 12668 17540 12696
rect 7524 12600 8892 12628
rect 7524 12588 7530 12600
rect 8938 12588 8944 12640
rect 8996 12628 9002 12640
rect 9217 12631 9275 12637
rect 9217 12628 9229 12631
rect 8996 12600 9229 12628
rect 8996 12588 9002 12600
rect 9217 12597 9229 12600
rect 9263 12597 9275 12631
rect 12636 12628 12664 12656
rect 14200 12628 14228 12668
rect 12636 12600 14228 12628
rect 9217 12591 9275 12597
rect 14366 12588 14372 12640
rect 14424 12628 14430 12640
rect 14737 12631 14795 12637
rect 14737 12628 14749 12631
rect 14424 12600 14749 12628
rect 14424 12588 14430 12600
rect 14737 12597 14749 12600
rect 14783 12597 14795 12631
rect 14737 12591 14795 12597
rect 14826 12588 14832 12640
rect 14884 12628 14890 12640
rect 15841 12631 15899 12637
rect 14884 12600 14929 12628
rect 14884 12588 14890 12600
rect 15841 12597 15853 12631
rect 15887 12628 15899 12631
rect 17236 12628 17264 12668
rect 17402 12628 17408 12640
rect 15887 12600 17264 12628
rect 17363 12600 17408 12628
rect 15887 12597 15899 12600
rect 15841 12591 15899 12597
rect 17402 12588 17408 12600
rect 17460 12588 17466 12640
rect 17512 12628 17540 12668
rect 19242 12628 19248 12640
rect 17512 12600 19248 12628
rect 19242 12588 19248 12600
rect 19300 12588 19306 12640
rect 19702 12588 19708 12640
rect 19760 12628 19766 12640
rect 19981 12631 20039 12637
rect 19981 12628 19993 12631
rect 19760 12600 19993 12628
rect 19760 12588 19766 12600
rect 19981 12597 19993 12600
rect 20027 12597 20039 12631
rect 19981 12591 20039 12597
rect 20165 12631 20223 12637
rect 20165 12597 20177 12631
rect 20211 12628 20223 12631
rect 22554 12628 22560 12640
rect 20211 12600 22560 12628
rect 20211 12597 20223 12600
rect 20165 12591 20223 12597
rect 22554 12588 22560 12600
rect 22612 12588 22618 12640
rect 22922 12628 22928 12640
rect 22883 12600 22928 12628
rect 22922 12588 22928 12600
rect 22980 12588 22986 12640
rect 1104 12538 23460 12560
rect 1104 12486 3749 12538
rect 3801 12486 3813 12538
rect 3865 12486 3877 12538
rect 3929 12486 3941 12538
rect 3993 12486 4005 12538
rect 4057 12486 9347 12538
rect 9399 12486 9411 12538
rect 9463 12486 9475 12538
rect 9527 12486 9539 12538
rect 9591 12486 9603 12538
rect 9655 12486 14945 12538
rect 14997 12486 15009 12538
rect 15061 12486 15073 12538
rect 15125 12486 15137 12538
rect 15189 12486 15201 12538
rect 15253 12486 20543 12538
rect 20595 12486 20607 12538
rect 20659 12486 20671 12538
rect 20723 12486 20735 12538
rect 20787 12486 20799 12538
rect 20851 12486 23460 12538
rect 1104 12464 23460 12486
rect 3142 12384 3148 12436
rect 3200 12424 3206 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3200 12396 3801 12424
rect 3200 12384 3206 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 3789 12387 3847 12393
rect 9125 12427 9183 12433
rect 9125 12393 9137 12427
rect 9171 12424 9183 12427
rect 9674 12424 9680 12436
rect 9171 12396 9680 12424
rect 9171 12393 9183 12396
rect 9125 12387 9183 12393
rect 9674 12384 9680 12396
rect 9732 12384 9738 12436
rect 10137 12427 10195 12433
rect 10137 12393 10149 12427
rect 10183 12424 10195 12427
rect 11974 12424 11980 12436
rect 10183 12396 11980 12424
rect 10183 12393 10195 12396
rect 10137 12387 10195 12393
rect 3421 12359 3479 12365
rect 3421 12325 3433 12359
rect 3467 12325 3479 12359
rect 3421 12319 3479 12325
rect 8757 12359 8815 12365
rect 8757 12325 8769 12359
rect 8803 12356 8815 12359
rect 9766 12356 9772 12368
rect 8803 12328 9772 12356
rect 8803 12325 8815 12328
rect 8757 12319 8815 12325
rect 2038 12288 2044 12300
rect 1999 12260 2044 12288
rect 2038 12248 2044 12260
rect 2096 12248 2102 12300
rect 3436 12288 3464 12319
rect 9766 12316 9772 12328
rect 9824 12316 9830 12368
rect 4614 12288 4620 12300
rect 3436 12260 4620 12288
rect 2130 12180 2136 12232
rect 2188 12220 2194 12232
rect 4448 12229 4476 12260
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 2297 12223 2355 12229
rect 2297 12220 2309 12223
rect 2188 12192 2309 12220
rect 2188 12180 2194 12192
rect 2297 12189 2309 12192
rect 2343 12189 2355 12223
rect 2297 12183 2355 12189
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12189 4491 12223
rect 4433 12183 4491 12189
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 3694 12112 3700 12164
rect 3752 12152 3758 12164
rect 4540 12152 4568 12183
rect 4890 12180 4896 12232
rect 4948 12220 4954 12232
rect 5445 12223 5503 12229
rect 5445 12220 5457 12223
rect 4948 12192 5457 12220
rect 4948 12180 4954 12192
rect 5445 12189 5457 12192
rect 5491 12189 5503 12223
rect 5445 12183 5503 12189
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 5629 12223 5687 12229
rect 5629 12220 5641 12223
rect 5592 12192 5641 12220
rect 5592 12180 5598 12192
rect 5629 12189 5641 12192
rect 5675 12189 5687 12223
rect 5629 12183 5687 12189
rect 6641 12223 6699 12229
rect 6641 12189 6653 12223
rect 6687 12220 6699 12223
rect 7857 12223 7915 12229
rect 6687 12192 6776 12220
rect 6687 12189 6699 12192
rect 6641 12183 6699 12189
rect 3752 12124 4568 12152
rect 3752 12112 3758 12124
rect 4614 12112 4620 12164
rect 4672 12152 4678 12164
rect 5902 12152 5908 12164
rect 4672 12124 5908 12152
rect 4672 12112 4678 12124
rect 5902 12112 5908 12124
rect 5960 12112 5966 12164
rect 4246 12044 4252 12096
rect 4304 12084 4310 12096
rect 4522 12084 4528 12096
rect 4304 12056 4528 12084
rect 4304 12044 4310 12056
rect 4522 12044 4528 12056
rect 4580 12044 4586 12096
rect 5166 12084 5172 12096
rect 5127 12056 5172 12084
rect 5166 12044 5172 12056
rect 5224 12044 5230 12096
rect 5994 12084 6000 12096
rect 5955 12056 6000 12084
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6748 12093 6776 12192
rect 7857 12189 7869 12223
rect 7903 12220 7915 12223
rect 8018 12220 8024 12232
rect 7903 12192 8024 12220
rect 7903 12189 7915 12192
rect 7857 12183 7915 12189
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 8113 12223 8171 12229
rect 8113 12189 8125 12223
rect 8159 12220 8171 12223
rect 8386 12220 8392 12232
rect 8159 12192 8392 12220
rect 8159 12189 8171 12192
rect 8113 12183 8171 12189
rect 8386 12180 8392 12192
rect 8444 12180 8450 12232
rect 8573 12223 8631 12229
rect 8573 12189 8585 12223
rect 8619 12220 8631 12223
rect 8662 12220 8668 12232
rect 8619 12192 8668 12220
rect 8619 12189 8631 12192
rect 8573 12183 8631 12189
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 8938 12220 8944 12232
rect 8899 12192 8944 12220
rect 8938 12180 8944 12192
rect 8996 12180 9002 12232
rect 10045 12223 10103 12229
rect 10045 12189 10057 12223
rect 10091 12220 10103 12223
rect 10152 12220 10180 12387
rect 11974 12384 11980 12396
rect 12032 12384 12038 12436
rect 14921 12427 14979 12433
rect 14921 12393 14933 12427
rect 14967 12424 14979 12427
rect 14967 12396 16804 12424
rect 14967 12393 14979 12396
rect 14921 12387 14979 12393
rect 16776 12356 16804 12396
rect 16850 12384 16856 12436
rect 16908 12424 16914 12436
rect 17037 12427 17095 12433
rect 17037 12424 17049 12427
rect 16908 12396 17049 12424
rect 16908 12384 16914 12396
rect 17037 12393 17049 12396
rect 17083 12393 17095 12427
rect 17862 12424 17868 12436
rect 17037 12387 17095 12393
rect 17604 12396 17868 12424
rect 17604 12356 17632 12396
rect 17862 12384 17868 12396
rect 17920 12384 17926 12436
rect 18138 12384 18144 12436
rect 18196 12424 18202 12436
rect 19610 12424 19616 12436
rect 18196 12396 18552 12424
rect 19571 12396 19616 12424
rect 18196 12384 18202 12396
rect 16776 12328 17632 12356
rect 13909 12291 13967 12297
rect 13909 12257 13921 12291
rect 13955 12288 13967 12291
rect 14090 12288 14096 12300
rect 13955 12260 14096 12288
rect 13955 12257 13967 12260
rect 13909 12251 13967 12257
rect 14090 12248 14096 12260
rect 14148 12248 14154 12300
rect 14185 12291 14243 12297
rect 14185 12257 14197 12291
rect 14231 12257 14243 12291
rect 14366 12288 14372 12300
rect 14327 12260 14372 12288
rect 14185 12251 14243 12257
rect 11514 12220 11520 12232
rect 10091 12192 10180 12220
rect 11475 12192 11520 12220
rect 10091 12189 10103 12192
rect 10045 12183 10103 12189
rect 11514 12180 11520 12192
rect 11572 12180 11578 12232
rect 9401 12155 9459 12161
rect 9401 12121 9413 12155
rect 9447 12152 9459 12155
rect 10594 12152 10600 12164
rect 9447 12124 10600 12152
rect 9447 12121 9459 12124
rect 9401 12115 9459 12121
rect 10594 12112 10600 12124
rect 10652 12112 10658 12164
rect 11250 12155 11308 12161
rect 11250 12121 11262 12155
rect 11296 12121 11308 12155
rect 11250 12115 11308 12121
rect 6733 12087 6791 12093
rect 6733 12053 6745 12087
rect 6779 12084 6791 12087
rect 8478 12084 8484 12096
rect 6779 12056 8484 12084
rect 6779 12053 6791 12056
rect 6733 12047 6791 12053
rect 8478 12044 8484 12056
rect 8536 12044 8542 12096
rect 11256 12084 11284 12115
rect 11422 12112 11428 12164
rect 11480 12152 11486 12164
rect 12161 12155 12219 12161
rect 12161 12152 12173 12155
rect 11480 12124 12173 12152
rect 11480 12112 11486 12124
rect 12161 12121 12173 12124
rect 12207 12121 12219 12155
rect 14200 12152 14228 12251
rect 14366 12248 14372 12260
rect 14424 12248 14430 12300
rect 14734 12248 14740 12300
rect 14792 12288 14798 12300
rect 18524 12297 18552 12396
rect 19610 12384 19616 12396
rect 19668 12384 19674 12436
rect 19720 12396 21404 12424
rect 18598 12316 18604 12368
rect 18656 12356 18662 12368
rect 19720 12356 19748 12396
rect 18656 12328 19748 12356
rect 21376 12356 21404 12396
rect 21450 12384 21456 12436
rect 21508 12424 21514 12436
rect 21545 12427 21603 12433
rect 21545 12424 21557 12427
rect 21508 12396 21557 12424
rect 21508 12384 21514 12396
rect 21545 12393 21557 12396
rect 21591 12424 21603 12427
rect 22094 12424 22100 12436
rect 21591 12396 22100 12424
rect 21591 12393 21603 12396
rect 21545 12387 21603 12393
rect 22094 12384 22100 12396
rect 22152 12384 22158 12436
rect 21634 12356 21640 12368
rect 21376 12328 21640 12356
rect 18656 12316 18662 12328
rect 21634 12316 21640 12328
rect 21692 12316 21698 12368
rect 20254 12297 20260 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 14792 12260 15669 12288
rect 14792 12248 14798 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 18509 12291 18567 12297
rect 18509 12257 18521 12291
rect 18555 12257 18567 12291
rect 20211 12291 20260 12297
rect 20211 12288 20223 12291
rect 20167 12260 20223 12288
rect 18509 12251 18567 12257
rect 20211 12257 20223 12260
rect 20257 12257 20260 12291
rect 20211 12251 20260 12257
rect 20254 12248 20260 12251
rect 20312 12288 20318 12300
rect 21542 12288 21548 12300
rect 20312 12260 21548 12288
rect 20312 12248 20318 12260
rect 21542 12248 21548 12260
rect 21600 12248 21606 12300
rect 21726 12288 21732 12300
rect 21687 12260 21732 12288
rect 21726 12248 21732 12260
rect 21784 12248 21790 12300
rect 14461 12223 14519 12229
rect 14461 12189 14473 12223
rect 14507 12220 14519 12223
rect 14826 12220 14832 12232
rect 14507 12192 14832 12220
rect 14507 12189 14519 12192
rect 14461 12183 14519 12189
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 15565 12223 15623 12229
rect 15565 12189 15577 12223
rect 15611 12220 15623 12223
rect 15746 12220 15752 12232
rect 15611 12192 15752 12220
rect 15611 12189 15623 12192
rect 15565 12183 15623 12189
rect 15746 12180 15752 12192
rect 15804 12180 15810 12232
rect 15924 12223 15982 12229
rect 15924 12189 15936 12223
rect 15970 12220 15982 12223
rect 16206 12220 16212 12232
rect 15970 12192 16212 12220
rect 15970 12189 15982 12192
rect 15924 12183 15982 12189
rect 16206 12180 16212 12192
rect 16264 12180 16270 12232
rect 18242 12223 18300 12229
rect 18242 12220 18254 12223
rect 18156 12192 18254 12220
rect 18156 12164 18184 12192
rect 18242 12189 18254 12192
rect 18288 12189 18300 12223
rect 19058 12220 19064 12232
rect 19019 12192 19064 12220
rect 18242 12183 18300 12189
rect 19058 12180 19064 12192
rect 19116 12180 19122 12232
rect 19705 12223 19763 12229
rect 19705 12189 19717 12223
rect 19751 12220 19763 12223
rect 19794 12220 19800 12232
rect 19751 12192 19800 12220
rect 19751 12189 19763 12192
rect 19705 12183 19763 12189
rect 19794 12180 19800 12192
rect 19852 12180 19858 12232
rect 20441 12223 20499 12229
rect 20441 12189 20453 12223
rect 20487 12220 20499 12223
rect 21818 12220 21824 12232
rect 20487 12192 21824 12220
rect 20487 12189 20499 12192
rect 20441 12183 20499 12189
rect 21818 12180 21824 12192
rect 21876 12180 21882 12232
rect 22278 12220 22284 12232
rect 21928 12192 22284 12220
rect 14734 12152 14740 12164
rect 14200 12124 14740 12152
rect 12161 12115 12219 12121
rect 14476 12096 14504 12124
rect 14734 12112 14740 12124
rect 14792 12112 14798 12164
rect 18138 12112 18144 12164
rect 18196 12112 18202 12164
rect 18506 12112 18512 12164
rect 18564 12152 18570 12164
rect 18564 12124 19840 12152
rect 18564 12112 18570 12124
rect 11330 12084 11336 12096
rect 11256 12056 11336 12084
rect 11330 12044 11336 12056
rect 11388 12044 11394 12096
rect 14458 12044 14464 12096
rect 14516 12044 14522 12096
rect 14826 12084 14832 12096
rect 14787 12056 14832 12084
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 16942 12044 16948 12096
rect 17000 12084 17006 12096
rect 17126 12084 17132 12096
rect 17000 12056 17132 12084
rect 17000 12044 17006 12056
rect 17126 12044 17132 12056
rect 17184 12044 17190 12096
rect 17218 12044 17224 12096
rect 17276 12084 17282 12096
rect 18601 12087 18659 12093
rect 18601 12084 18613 12087
rect 17276 12056 18613 12084
rect 17276 12044 17282 12056
rect 18601 12053 18613 12056
rect 18647 12053 18659 12087
rect 19426 12084 19432 12096
rect 19387 12056 19432 12084
rect 18601 12047 18659 12053
rect 19426 12044 19432 12056
rect 19484 12044 19490 12096
rect 19812 12084 19840 12124
rect 21726 12112 21732 12164
rect 21784 12152 21790 12164
rect 21928 12152 21956 12192
rect 22278 12180 22284 12192
rect 22336 12180 22342 12232
rect 21784 12124 21956 12152
rect 21996 12155 22054 12161
rect 21784 12112 21790 12124
rect 21996 12121 22008 12155
rect 22042 12152 22054 12155
rect 22462 12152 22468 12164
rect 22042 12124 22468 12152
rect 22042 12121 22054 12124
rect 21996 12115 22054 12121
rect 22462 12112 22468 12124
rect 22520 12112 22526 12164
rect 19978 12084 19984 12096
rect 19812 12056 19984 12084
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 20070 12044 20076 12096
rect 20128 12084 20134 12096
rect 20171 12087 20229 12093
rect 20171 12084 20183 12087
rect 20128 12056 20183 12084
rect 20128 12044 20134 12056
rect 20171 12053 20183 12056
rect 20217 12053 20229 12087
rect 20171 12047 20229 12053
rect 20806 12044 20812 12096
rect 20864 12084 20870 12096
rect 21744 12084 21772 12112
rect 20864 12056 21772 12084
rect 20864 12044 20870 12056
rect 23014 12044 23020 12096
rect 23072 12084 23078 12096
rect 23109 12087 23167 12093
rect 23109 12084 23121 12087
rect 23072 12056 23121 12084
rect 23072 12044 23078 12056
rect 23109 12053 23121 12056
rect 23155 12053 23167 12087
rect 23109 12047 23167 12053
rect 1104 11994 23460 12016
rect 1104 11942 6548 11994
rect 6600 11942 6612 11994
rect 6664 11942 6676 11994
rect 6728 11942 6740 11994
rect 6792 11942 6804 11994
rect 6856 11942 12146 11994
rect 12198 11942 12210 11994
rect 12262 11942 12274 11994
rect 12326 11942 12338 11994
rect 12390 11942 12402 11994
rect 12454 11942 17744 11994
rect 17796 11942 17808 11994
rect 17860 11942 17872 11994
rect 17924 11942 17936 11994
rect 17988 11942 18000 11994
rect 18052 11942 23460 11994
rect 1104 11920 23460 11942
rect 1394 11840 1400 11892
rect 1452 11880 1458 11892
rect 1765 11883 1823 11889
rect 1765 11880 1777 11883
rect 1452 11852 1777 11880
rect 1452 11840 1458 11852
rect 1765 11849 1777 11852
rect 1811 11880 1823 11883
rect 3605 11883 3663 11889
rect 3605 11880 3617 11883
rect 1811 11852 3617 11880
rect 1811 11849 1823 11852
rect 1765 11843 1823 11849
rect 3605 11849 3617 11852
rect 3651 11849 3663 11883
rect 3605 11843 3663 11849
rect 3694 11840 3700 11892
rect 3752 11880 3758 11892
rect 4249 11883 4307 11889
rect 3752 11852 3797 11880
rect 3752 11840 3758 11852
rect 4249 11849 4261 11883
rect 4295 11880 4307 11883
rect 4982 11880 4988 11892
rect 4295 11852 4988 11880
rect 4295 11849 4307 11852
rect 4249 11843 4307 11849
rect 4982 11840 4988 11852
rect 5040 11840 5046 11892
rect 5350 11880 5356 11892
rect 5311 11852 5356 11880
rect 5350 11840 5356 11852
rect 5408 11840 5414 11892
rect 8113 11883 8171 11889
rect 8113 11849 8125 11883
rect 8159 11849 8171 11883
rect 8478 11880 8484 11892
rect 8439 11852 8484 11880
rect 8113 11843 8171 11849
rect 2900 11815 2958 11821
rect 2900 11781 2912 11815
rect 2946 11812 2958 11815
rect 5166 11812 5172 11824
rect 2946 11784 5172 11812
rect 2946 11781 2958 11784
rect 2900 11775 2958 11781
rect 5166 11772 5172 11784
rect 5224 11772 5230 11824
rect 5994 11772 6000 11824
rect 6052 11812 6058 11824
rect 6978 11815 7036 11821
rect 6978 11812 6990 11815
rect 6052 11784 6990 11812
rect 6052 11772 6058 11784
rect 6978 11781 6990 11784
rect 7024 11781 7036 11815
rect 8128 11812 8156 11843
rect 8478 11840 8484 11852
rect 8536 11840 8542 11892
rect 8846 11840 8852 11892
rect 8904 11880 8910 11892
rect 8941 11883 8999 11889
rect 8941 11880 8953 11883
rect 8904 11852 8953 11880
rect 8904 11840 8910 11852
rect 8941 11849 8953 11852
rect 8987 11849 8999 11883
rect 8941 11843 8999 11849
rect 11333 11883 11391 11889
rect 11333 11849 11345 11883
rect 11379 11880 11391 11883
rect 11977 11883 12035 11889
rect 11977 11880 11989 11883
rect 11379 11852 11989 11880
rect 11379 11849 11391 11852
rect 11333 11843 11391 11849
rect 11977 11849 11989 11852
rect 12023 11880 12035 11883
rect 12066 11880 12072 11892
rect 12023 11852 12072 11880
rect 12023 11849 12035 11852
rect 11977 11843 12035 11849
rect 12066 11840 12072 11852
rect 12124 11840 12130 11892
rect 14737 11883 14795 11889
rect 14737 11849 14749 11883
rect 14783 11880 14795 11883
rect 15197 11883 15255 11889
rect 15197 11880 15209 11883
rect 14783 11852 15209 11880
rect 14783 11849 14795 11852
rect 14737 11843 14795 11849
rect 15197 11849 15209 11852
rect 15243 11849 15255 11883
rect 15197 11843 15255 11849
rect 17126 11840 17132 11892
rect 17184 11880 17190 11892
rect 17494 11880 17500 11892
rect 17184 11852 17500 11880
rect 17184 11840 17190 11852
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 17586 11840 17592 11892
rect 17644 11880 17650 11892
rect 18509 11883 18567 11889
rect 18509 11880 18521 11883
rect 17644 11852 18521 11880
rect 17644 11840 17650 11852
rect 18509 11849 18521 11852
rect 18555 11849 18567 11883
rect 18509 11843 18567 11849
rect 18598 11840 18604 11892
rect 18656 11880 18662 11892
rect 18656 11852 19380 11880
rect 18656 11840 18662 11852
rect 8573 11815 8631 11821
rect 8573 11812 8585 11815
rect 8128 11784 8585 11812
rect 6978 11775 7036 11781
rect 8573 11781 8585 11784
rect 8619 11781 8631 11815
rect 11514 11812 11520 11824
rect 8573 11775 8631 11781
rect 9968 11784 11520 11812
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11744 4123 11747
rect 4246 11744 4252 11756
rect 4111 11716 4252 11744
rect 4111 11713 4123 11716
rect 4065 11707 4123 11713
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 4525 11747 4583 11753
rect 4525 11713 4537 11747
rect 4571 11744 4583 11747
rect 4614 11744 4620 11756
rect 4571 11716 4620 11744
rect 4571 11713 4583 11716
rect 4525 11707 4583 11713
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 4982 11744 4988 11756
rect 4943 11716 4988 11744
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 5442 11704 5448 11756
rect 5500 11744 5506 11756
rect 6089 11747 6147 11753
rect 6089 11744 6101 11747
rect 5500 11716 6101 11744
rect 5500 11704 5506 11716
rect 6089 11713 6101 11716
rect 6135 11713 6147 11747
rect 6089 11707 6147 11713
rect 6454 11704 6460 11756
rect 6512 11744 6518 11756
rect 6549 11747 6607 11753
rect 6549 11744 6561 11747
rect 6512 11716 6561 11744
rect 6512 11704 6518 11716
rect 6549 11713 6561 11716
rect 6595 11713 6607 11747
rect 8588 11744 8616 11775
rect 9968 11753 9996 11784
rect 11514 11772 11520 11784
rect 11572 11772 11578 11824
rect 13998 11812 14004 11824
rect 13188 11784 14004 11812
rect 9033 11747 9091 11753
rect 9033 11744 9045 11747
rect 8588 11716 9045 11744
rect 6549 11707 6607 11713
rect 9033 11713 9045 11716
rect 9079 11713 9091 11747
rect 9033 11707 9091 11713
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 10042 11704 10048 11756
rect 10100 11744 10106 11756
rect 10209 11747 10267 11753
rect 10209 11744 10221 11747
rect 10100 11716 10221 11744
rect 10100 11704 10106 11716
rect 10209 11713 10221 11716
rect 10255 11713 10267 11747
rect 10209 11707 10267 11713
rect 11974 11704 11980 11756
rect 12032 11744 12038 11756
rect 12032 11716 12204 11744
rect 12032 11704 12038 11716
rect 3145 11679 3203 11685
rect 3145 11645 3157 11679
rect 3191 11645 3203 11679
rect 3145 11639 3203 11645
rect 3881 11679 3939 11685
rect 3881 11645 3893 11679
rect 3927 11676 3939 11679
rect 4338 11676 4344 11688
rect 3927 11648 4344 11676
rect 3927 11645 3939 11648
rect 3881 11639 3939 11645
rect 3160 11608 3188 11639
rect 4338 11636 4344 11648
rect 4396 11636 4402 11688
rect 4706 11676 4712 11688
rect 4667 11648 4712 11676
rect 4706 11636 4712 11648
rect 4764 11636 4770 11688
rect 4798 11636 4804 11688
rect 4856 11676 4862 11688
rect 4893 11679 4951 11685
rect 4893 11676 4905 11679
rect 4856 11648 4905 11676
rect 4856 11636 4862 11648
rect 4893 11645 4905 11648
rect 4939 11645 4951 11679
rect 4893 11639 4951 11645
rect 6178 11636 6184 11688
rect 6236 11676 6242 11688
rect 6733 11679 6791 11685
rect 6733 11676 6745 11679
rect 6236 11648 6745 11676
rect 6236 11636 6242 11648
rect 6733 11645 6745 11648
rect 6779 11645 6791 11679
rect 6733 11639 6791 11645
rect 8389 11679 8447 11685
rect 8389 11645 8401 11679
rect 8435 11676 8447 11679
rect 8570 11676 8576 11688
rect 8435 11648 8576 11676
rect 8435 11645 8447 11648
rect 8389 11639 8447 11645
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 10962 11636 10968 11688
rect 11020 11676 11026 11688
rect 12176 11685 12204 11716
rect 13188 11685 13216 11784
rect 13998 11772 14004 11784
rect 14056 11772 14062 11824
rect 15562 11812 15568 11824
rect 14568 11784 15568 11812
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11744 13415 11747
rect 13814 11744 13820 11756
rect 13403 11716 13820 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 13814 11704 13820 11716
rect 13872 11704 13878 11756
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11020 11648 12081 11676
rect 11020 11636 11026 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 12161 11679 12219 11685
rect 12161 11645 12173 11679
rect 12207 11645 12219 11679
rect 12161 11639 12219 11645
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 13265 11679 13323 11685
rect 13265 11645 13277 11679
rect 13311 11676 13323 11679
rect 13538 11676 13544 11688
rect 13311 11648 13544 11676
rect 13311 11645 13323 11648
rect 13265 11639 13323 11645
rect 13538 11636 13544 11648
rect 13596 11636 13602 11688
rect 14568 11685 14596 11784
rect 15562 11772 15568 11784
rect 15620 11772 15626 11824
rect 17396 11815 17454 11821
rect 17396 11781 17408 11815
rect 17442 11812 17454 11815
rect 18322 11812 18328 11824
rect 17442 11784 18328 11812
rect 17442 11781 17454 11784
rect 17396 11775 17454 11781
rect 18322 11772 18328 11784
rect 18380 11772 18386 11824
rect 18414 11772 18420 11824
rect 18472 11812 18478 11824
rect 18846 11815 18904 11821
rect 18846 11812 18858 11815
rect 18472 11784 18858 11812
rect 18472 11772 18478 11784
rect 18846 11781 18858 11784
rect 18892 11781 18904 11815
rect 19352 11812 19380 11852
rect 19426 11840 19432 11892
rect 19484 11880 19490 11892
rect 20441 11883 20499 11889
rect 20441 11880 20453 11883
rect 19484 11852 20453 11880
rect 19484 11840 19490 11852
rect 20441 11849 20453 11852
rect 20487 11849 20499 11883
rect 20806 11880 20812 11892
rect 20767 11852 20812 11880
rect 20441 11843 20499 11849
rect 20806 11840 20812 11852
rect 20864 11840 20870 11892
rect 21361 11883 21419 11889
rect 21361 11849 21373 11883
rect 21407 11880 21419 11883
rect 21821 11883 21879 11889
rect 21821 11880 21833 11883
rect 21407 11852 21833 11880
rect 21407 11849 21419 11852
rect 21361 11843 21419 11849
rect 21821 11849 21833 11852
rect 21867 11849 21879 11883
rect 21821 11843 21879 11849
rect 22094 11840 22100 11892
rect 22152 11880 22158 11892
rect 22281 11883 22339 11889
rect 22281 11880 22293 11883
rect 22152 11852 22293 11880
rect 22152 11840 22158 11852
rect 22281 11849 22293 11852
rect 22327 11849 22339 11883
rect 22281 11843 22339 11849
rect 21174 11812 21180 11824
rect 19352 11784 21180 11812
rect 18846 11775 18904 11781
rect 21174 11772 21180 11784
rect 21232 11772 21238 11824
rect 21269 11815 21327 11821
rect 21269 11781 21281 11815
rect 21315 11812 21327 11815
rect 22649 11815 22707 11821
rect 22649 11812 22661 11815
rect 21315 11784 22661 11812
rect 21315 11781 21327 11784
rect 21269 11775 21327 11781
rect 22649 11781 22661 11784
rect 22695 11781 22707 11815
rect 22649 11775 22707 11781
rect 14826 11704 14832 11756
rect 14884 11744 14890 11756
rect 15381 11747 15439 11753
rect 15381 11744 15393 11747
rect 14884 11716 15393 11744
rect 14884 11704 14890 11716
rect 15381 11713 15393 11716
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 15470 11704 15476 11756
rect 15528 11744 15534 11756
rect 15657 11747 15715 11753
rect 15657 11744 15669 11747
rect 15528 11716 15669 11744
rect 15528 11704 15534 11716
rect 15657 11713 15669 11716
rect 15703 11713 15715 11747
rect 16114 11744 16120 11756
rect 16075 11716 16120 11744
rect 15657 11707 15715 11713
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 16666 11704 16672 11756
rect 16724 11744 16730 11756
rect 16853 11747 16911 11753
rect 16853 11744 16865 11747
rect 16724 11716 16865 11744
rect 16724 11704 16730 11716
rect 16853 11713 16865 11716
rect 16899 11713 16911 11747
rect 16853 11707 16911 11713
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 17092 11716 21496 11744
rect 17092 11704 17098 11716
rect 14553 11679 14611 11685
rect 14553 11645 14565 11679
rect 14599 11645 14611 11679
rect 14553 11639 14611 11645
rect 14645 11679 14703 11685
rect 14645 11645 14657 11679
rect 14691 11645 14703 11679
rect 14645 11639 14703 11645
rect 15933 11679 15991 11685
rect 15933 11645 15945 11679
rect 15979 11645 15991 11679
rect 15933 11639 15991 11645
rect 6196 11608 6224 11636
rect 3160 11580 6224 11608
rect 6270 11568 6276 11620
rect 6328 11608 6334 11620
rect 6365 11611 6423 11617
rect 6365 11608 6377 11611
rect 6328 11580 6377 11608
rect 6328 11568 6334 11580
rect 6365 11577 6377 11580
rect 6411 11577 6423 11611
rect 11606 11608 11612 11620
rect 11567 11580 11612 11608
rect 6365 11571 6423 11577
rect 11606 11568 11612 11580
rect 11664 11568 11670 11620
rect 14660 11608 14688 11639
rect 15473 11611 15531 11617
rect 15473 11608 15485 11611
rect 14660 11580 15485 11608
rect 15473 11577 15485 11580
rect 15519 11577 15531 11611
rect 15948 11608 15976 11639
rect 16022 11636 16028 11688
rect 16080 11676 16086 11688
rect 16080 11648 16125 11676
rect 16080 11636 16086 11648
rect 16390 11636 16396 11688
rect 16448 11676 16454 11688
rect 17129 11679 17187 11685
rect 17129 11676 17141 11679
rect 16448 11648 17141 11676
rect 16448 11636 16454 11648
rect 17129 11645 17141 11648
rect 17175 11645 17187 11679
rect 18598 11676 18604 11688
rect 18559 11648 18604 11676
rect 17129 11639 17187 11645
rect 18598 11636 18604 11648
rect 18656 11636 18662 11688
rect 19978 11636 19984 11688
rect 20036 11676 20042 11688
rect 20165 11679 20223 11685
rect 20165 11676 20177 11679
rect 20036 11648 20177 11676
rect 20036 11636 20042 11648
rect 20165 11645 20177 11648
rect 20211 11645 20223 11679
rect 20346 11676 20352 11688
rect 20307 11648 20352 11676
rect 20165 11639 20223 11645
rect 20346 11636 20352 11648
rect 20404 11636 20410 11688
rect 21468 11685 21496 11716
rect 21542 11704 21548 11756
rect 21600 11744 21606 11756
rect 22189 11747 22247 11753
rect 22189 11744 22201 11747
rect 21600 11716 22201 11744
rect 21600 11704 21606 11716
rect 22189 11713 22201 11716
rect 22235 11713 22247 11747
rect 23106 11744 23112 11756
rect 23067 11716 23112 11744
rect 22189 11707 22247 11713
rect 23106 11704 23112 11716
rect 23164 11704 23170 11756
rect 21453 11679 21511 11685
rect 21453 11645 21465 11679
rect 21499 11676 21511 11679
rect 22094 11676 22100 11688
rect 21499 11648 22100 11676
rect 21499 11645 21511 11648
rect 21453 11639 21511 11645
rect 22094 11636 22100 11648
rect 22152 11636 22158 11688
rect 22373 11679 22431 11685
rect 22373 11645 22385 11679
rect 22419 11676 22431 11679
rect 23014 11676 23020 11688
rect 22419 11648 23020 11676
rect 22419 11645 22431 11648
rect 22373 11639 22431 11645
rect 16669 11611 16727 11617
rect 16669 11608 16681 11611
rect 15948 11580 16681 11608
rect 15473 11571 15531 11577
rect 16669 11577 16681 11580
rect 16715 11577 16727 11611
rect 21266 11608 21272 11620
rect 16669 11571 16727 11577
rect 19904 11580 21272 11608
rect 3234 11540 3240 11552
rect 3195 11512 3240 11540
rect 3234 11500 3240 11512
rect 3292 11500 3298 11552
rect 4338 11540 4344 11552
rect 4299 11512 4344 11540
rect 4338 11500 4344 11512
rect 4396 11500 4402 11552
rect 4522 11500 4528 11552
rect 4580 11540 4586 11552
rect 5445 11543 5503 11549
rect 5445 11540 5457 11543
rect 4580 11512 5457 11540
rect 4580 11500 4586 11512
rect 5445 11509 5457 11512
rect 5491 11509 5503 11543
rect 9674 11540 9680 11552
rect 9635 11512 9680 11540
rect 5445 11503 5503 11509
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 13722 11540 13728 11552
rect 13683 11512 13728 11540
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 13909 11543 13967 11549
rect 13909 11509 13921 11543
rect 13955 11540 13967 11543
rect 14550 11540 14556 11552
rect 13955 11512 14556 11540
rect 13955 11509 13967 11512
rect 13909 11503 13967 11509
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 15105 11543 15163 11549
rect 15105 11509 15117 11543
rect 15151 11540 15163 11543
rect 16114 11540 16120 11552
rect 15151 11512 16120 11540
rect 15151 11509 15163 11512
rect 15105 11503 15163 11509
rect 16114 11500 16120 11512
rect 16172 11500 16178 11552
rect 16485 11543 16543 11549
rect 16485 11509 16497 11543
rect 16531 11540 16543 11543
rect 17770 11540 17776 11552
rect 16531 11512 17776 11540
rect 16531 11509 16543 11512
rect 16485 11503 16543 11509
rect 17770 11500 17776 11512
rect 17828 11500 17834 11552
rect 18966 11500 18972 11552
rect 19024 11540 19030 11552
rect 19904 11540 19932 11580
rect 21266 11568 21272 11580
rect 21324 11568 21330 11620
rect 21634 11568 21640 11620
rect 21692 11608 21698 11620
rect 22388 11608 22416 11639
rect 23014 11636 23020 11648
rect 23072 11636 23078 11688
rect 21692 11580 22416 11608
rect 21692 11568 21698 11580
rect 19024 11512 19932 11540
rect 19024 11500 19030 11512
rect 19978 11500 19984 11552
rect 20036 11540 20042 11552
rect 20036 11512 20081 11540
rect 20036 11500 20042 11512
rect 20898 11500 20904 11552
rect 20956 11540 20962 11552
rect 20956 11512 21001 11540
rect 20956 11500 20962 11512
rect 22646 11500 22652 11552
rect 22704 11540 22710 11552
rect 22925 11543 22983 11549
rect 22925 11540 22937 11543
rect 22704 11512 22937 11540
rect 22704 11500 22710 11512
rect 22925 11509 22937 11512
rect 22971 11509 22983 11543
rect 22925 11503 22983 11509
rect 1104 11450 23460 11472
rect 1104 11398 3749 11450
rect 3801 11398 3813 11450
rect 3865 11398 3877 11450
rect 3929 11398 3941 11450
rect 3993 11398 4005 11450
rect 4057 11398 9347 11450
rect 9399 11398 9411 11450
rect 9463 11398 9475 11450
rect 9527 11398 9539 11450
rect 9591 11398 9603 11450
rect 9655 11398 14945 11450
rect 14997 11398 15009 11450
rect 15061 11398 15073 11450
rect 15125 11398 15137 11450
rect 15189 11398 15201 11450
rect 15253 11398 20543 11450
rect 20595 11398 20607 11450
rect 20659 11398 20671 11450
rect 20723 11398 20735 11450
rect 20787 11398 20799 11450
rect 20851 11398 23460 11450
rect 1104 11376 23460 11398
rect 3145 11339 3203 11345
rect 3145 11305 3157 11339
rect 3191 11336 3203 11339
rect 3510 11336 3516 11348
rect 3191 11308 3516 11336
rect 3191 11305 3203 11308
rect 3145 11299 3203 11305
rect 3510 11296 3516 11308
rect 3568 11296 3574 11348
rect 3973 11339 4031 11345
rect 3973 11305 3985 11339
rect 4019 11336 4031 11339
rect 4154 11336 4160 11348
rect 4019 11308 4160 11336
rect 4019 11305 4031 11308
rect 3973 11299 4031 11305
rect 4154 11296 4160 11308
rect 4212 11296 4218 11348
rect 4249 11339 4307 11345
rect 4249 11305 4261 11339
rect 4295 11336 4307 11339
rect 4982 11336 4988 11348
rect 4295 11308 4988 11336
rect 4295 11305 4307 11308
rect 4249 11299 4307 11305
rect 4982 11296 4988 11308
rect 5040 11296 5046 11348
rect 9122 11336 9128 11348
rect 9083 11308 9128 11336
rect 9122 11296 9128 11308
rect 9180 11296 9186 11348
rect 9217 11339 9275 11345
rect 9217 11305 9229 11339
rect 9263 11336 9275 11339
rect 10042 11336 10048 11348
rect 9263 11308 10048 11336
rect 9263 11305 9275 11308
rect 9217 11299 9275 11305
rect 10042 11296 10048 11308
rect 10100 11296 10106 11348
rect 10962 11336 10968 11348
rect 10428 11308 10968 11336
rect 3605 11271 3663 11277
rect 3605 11237 3617 11271
rect 3651 11268 3663 11271
rect 4798 11268 4804 11280
rect 3651 11240 4804 11268
rect 3651 11237 3663 11240
rect 3605 11231 3663 11237
rect 4798 11228 4804 11240
rect 4856 11228 4862 11280
rect 6362 11268 6368 11280
rect 5000 11240 6368 11268
rect 4430 11200 4436 11212
rect 3804 11172 4436 11200
rect 1762 11132 1768 11144
rect 1723 11104 1768 11132
rect 1762 11092 1768 11104
rect 1820 11092 1826 11144
rect 3418 11132 3424 11144
rect 3379 11104 3424 11132
rect 3418 11092 3424 11104
rect 3476 11092 3482 11144
rect 3804 11141 3832 11172
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 4706 11160 4712 11212
rect 4764 11200 4770 11212
rect 5000 11209 5028 11240
rect 6362 11228 6368 11240
rect 6420 11228 6426 11280
rect 9953 11271 10011 11277
rect 9953 11237 9965 11271
rect 9999 11268 10011 11271
rect 10428 11268 10456 11308
rect 10962 11296 10968 11308
rect 11020 11296 11026 11348
rect 11330 11296 11336 11348
rect 11388 11336 11394 11348
rect 11425 11339 11483 11345
rect 11425 11336 11437 11339
rect 11388 11308 11437 11336
rect 11388 11296 11394 11308
rect 11425 11305 11437 11308
rect 11471 11305 11483 11339
rect 11425 11299 11483 11305
rect 13725 11339 13783 11345
rect 13725 11305 13737 11339
rect 13771 11336 13783 11339
rect 13814 11336 13820 11348
rect 13771 11308 13820 11336
rect 13771 11305 13783 11308
rect 13725 11299 13783 11305
rect 13814 11296 13820 11308
rect 13872 11296 13878 11348
rect 13906 11296 13912 11348
rect 13964 11336 13970 11348
rect 14182 11336 14188 11348
rect 13964 11308 14188 11336
rect 13964 11296 13970 11308
rect 14182 11296 14188 11308
rect 14240 11296 14246 11348
rect 14829 11339 14887 11345
rect 14829 11305 14841 11339
rect 14875 11336 14887 11339
rect 15470 11336 15476 11348
rect 14875 11308 15476 11336
rect 14875 11305 14887 11308
rect 14829 11299 14887 11305
rect 15470 11296 15476 11308
rect 15528 11296 15534 11348
rect 15657 11339 15715 11345
rect 15657 11305 15669 11339
rect 15703 11336 15715 11339
rect 16022 11336 16028 11348
rect 15703 11308 16028 11336
rect 15703 11305 15715 11308
rect 15657 11299 15715 11305
rect 9999 11240 10456 11268
rect 9999 11237 10011 11240
rect 9953 11231 10011 11237
rect 4985 11203 5043 11209
rect 4985 11200 4997 11203
rect 4764 11172 4997 11200
rect 4764 11160 4770 11172
rect 4985 11169 4997 11172
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 5813 11163 5871 11169
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11200 6331 11203
rect 6319 11172 7420 11200
rect 6319 11169 6331 11172
rect 6273 11163 6331 11169
rect 3789 11135 3847 11141
rect 3789 11101 3801 11135
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 4065 11135 4123 11141
rect 4065 11101 4077 11135
rect 4111 11101 4123 11135
rect 4614 11132 4620 11144
rect 4065 11095 4123 11101
rect 4356 11104 4620 11132
rect 2032 11067 2090 11073
rect 2032 11033 2044 11067
rect 2078 11064 2090 11067
rect 3142 11064 3148 11076
rect 2078 11036 3148 11064
rect 2078 11033 2090 11036
rect 2032 11027 2090 11033
rect 3142 11024 3148 11036
rect 3200 11024 3206 11076
rect 3510 11024 3516 11076
rect 3568 11064 3574 11076
rect 4080 11064 4108 11095
rect 3568 11036 4108 11064
rect 3568 11024 3574 11036
rect 4356 11005 4384 11104
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 5442 11092 5448 11144
rect 5500 11132 5506 11144
rect 5537 11135 5595 11141
rect 5537 11132 5549 11135
rect 5500 11104 5549 11132
rect 5500 11092 5506 11104
rect 5537 11101 5549 11104
rect 5583 11101 5595 11135
rect 5828 11132 5856 11163
rect 6454 11132 6460 11144
rect 5828 11104 6460 11132
rect 5537 11095 5595 11101
rect 6454 11092 6460 11104
rect 6512 11092 6518 11144
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11132 6975 11135
rect 7392 11132 7420 11172
rect 8386 11132 8392 11144
rect 6963 11104 7052 11132
rect 7392 11104 8064 11132
rect 8299 11104 8392 11132
rect 6963 11101 6975 11104
rect 6917 11095 6975 11101
rect 4706 11064 4712 11076
rect 4667 11036 4712 11064
rect 4706 11024 4712 11036
rect 4764 11024 4770 11076
rect 7024 11008 7052 11104
rect 4341 10999 4399 11005
rect 4341 10965 4353 10999
rect 4387 10965 4399 10999
rect 4341 10959 4399 10965
rect 4522 10956 4528 11008
rect 4580 10996 4586 11008
rect 4801 10999 4859 11005
rect 4801 10996 4813 10999
rect 4580 10968 4813 10996
rect 4580 10956 4586 10968
rect 4801 10965 4813 10968
rect 4847 10965 4859 10999
rect 5166 10996 5172 11008
rect 5127 10968 5172 10996
rect 4801 10959 4859 10965
rect 5166 10956 5172 10968
rect 5224 10956 5230 11008
rect 5629 10999 5687 11005
rect 5629 10965 5641 10999
rect 5675 10996 5687 10999
rect 6086 10996 6092 11008
rect 5675 10968 6092 10996
rect 5675 10965 5687 10968
rect 5629 10959 5687 10965
rect 6086 10956 6092 10968
rect 6144 10956 6150 11008
rect 7006 10996 7012 11008
rect 6967 10968 7012 10996
rect 7006 10956 7012 10968
rect 7064 10956 7070 11008
rect 8036 10996 8064 11104
rect 8386 11092 8392 11104
rect 8444 11132 8450 11144
rect 8570 11132 8576 11144
rect 8444 11104 8576 11132
rect 8444 11092 8450 11104
rect 8570 11092 8576 11104
rect 8628 11092 8634 11144
rect 8938 11132 8944 11144
rect 8899 11104 8944 11132
rect 8938 11092 8944 11104
rect 8996 11092 9002 11144
rect 9861 11135 9919 11141
rect 9861 11101 9873 11135
rect 9907 11132 9919 11135
rect 9968 11132 9996 11231
rect 11333 11203 11391 11209
rect 11333 11169 11345 11203
rect 11379 11200 11391 11203
rect 11514 11200 11520 11212
rect 11379 11172 11520 11200
rect 11379 11169 11391 11172
rect 11333 11163 11391 11169
rect 9907 11104 9996 11132
rect 9907 11101 9919 11104
rect 9861 11095 9919 11101
rect 10502 11092 10508 11144
rect 10560 11132 10566 11144
rect 11348 11132 11376 11163
rect 11514 11160 11520 11172
rect 11572 11160 11578 11212
rect 13906 11200 13912 11212
rect 13648 11172 13912 11200
rect 12066 11132 12072 11144
rect 10560 11104 11376 11132
rect 12027 11104 12072 11132
rect 10560 11092 10566 11104
rect 12066 11092 12072 11104
rect 12124 11092 12130 11144
rect 12345 11135 12403 11141
rect 12345 11101 12357 11135
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 12612 11135 12670 11141
rect 12612 11101 12624 11135
rect 12658 11132 12670 11135
rect 13648 11132 13676 11172
rect 13906 11160 13912 11172
rect 13964 11160 13970 11212
rect 14274 11200 14280 11212
rect 14235 11172 14280 11200
rect 14274 11160 14280 11172
rect 14332 11200 14338 11212
rect 14734 11200 14740 11212
rect 14332 11172 14740 11200
rect 14332 11160 14338 11172
rect 14734 11160 14740 11172
rect 14792 11160 14798 11212
rect 15105 11203 15163 11209
rect 15105 11169 15117 11203
rect 15151 11200 15163 11203
rect 15562 11200 15568 11212
rect 15151 11172 15568 11200
rect 15151 11169 15163 11172
rect 15105 11163 15163 11169
rect 15562 11160 15568 11172
rect 15620 11160 15626 11212
rect 12658 11104 13676 11132
rect 12658 11101 12670 11104
rect 12612 11095 12670 11101
rect 8144 11067 8202 11073
rect 8144 11033 8156 11067
rect 8190 11064 8202 11067
rect 9674 11064 9680 11076
rect 8190 11036 9680 11064
rect 8190 11033 8202 11036
rect 8144 11027 8202 11033
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 10686 11024 10692 11076
rect 10744 11064 10750 11076
rect 11066 11067 11124 11073
rect 11066 11064 11078 11067
rect 10744 11036 11078 11064
rect 10744 11024 10750 11036
rect 11066 11033 11078 11036
rect 11112 11033 11124 11067
rect 11066 11027 11124 11033
rect 8294 10996 8300 11008
rect 8036 10968 8300 10996
rect 8294 10956 8300 10968
rect 8352 10956 8358 11008
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 12360 10996 12388 11095
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 15764 11141 15792 11308
rect 16022 11296 16028 11308
rect 16080 11296 16086 11348
rect 17034 11336 17040 11348
rect 16684 11308 17040 11336
rect 15933 11271 15991 11277
rect 15933 11237 15945 11271
rect 15979 11268 15991 11271
rect 16574 11268 16580 11280
rect 15979 11240 16580 11268
rect 15979 11237 15991 11240
rect 15933 11231 15991 11237
rect 16574 11228 16580 11240
rect 16632 11228 16638 11280
rect 16684 11141 16712 11308
rect 17034 11296 17040 11308
rect 17092 11296 17098 11348
rect 17310 11296 17316 11348
rect 17368 11336 17374 11348
rect 17589 11339 17647 11345
rect 17589 11336 17601 11339
rect 17368 11308 17601 11336
rect 17368 11296 17374 11308
rect 17589 11305 17601 11308
rect 17635 11305 17647 11339
rect 17589 11299 17647 11305
rect 18693 11339 18751 11345
rect 18693 11305 18705 11339
rect 18739 11336 18751 11339
rect 20346 11336 20352 11348
rect 18739 11308 20352 11336
rect 18739 11305 18751 11308
rect 18693 11299 18751 11305
rect 20346 11296 20352 11308
rect 20404 11296 20410 11348
rect 20990 11336 20996 11348
rect 20951 11308 20996 11336
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 23106 11336 23112 11348
rect 21100 11308 23112 11336
rect 17494 11268 17500 11280
rect 17407 11240 17500 11268
rect 17494 11228 17500 11240
rect 17552 11268 17558 11280
rect 18966 11268 18972 11280
rect 17552 11240 18368 11268
rect 18927 11240 18972 11268
rect 17552 11228 17558 11240
rect 16942 11200 16948 11212
rect 16903 11172 16948 11200
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 17037 11203 17095 11209
rect 17037 11169 17049 11203
rect 17083 11200 17095 11203
rect 17402 11200 17408 11212
rect 17083 11172 17408 11200
rect 17083 11169 17095 11172
rect 17037 11163 17095 11169
rect 17402 11160 17408 11172
rect 17460 11160 17466 11212
rect 17586 11160 17592 11212
rect 17644 11200 17650 11212
rect 18049 11203 18107 11209
rect 18049 11200 18061 11203
rect 17644 11172 18061 11200
rect 17644 11160 17650 11172
rect 18049 11169 18061 11172
rect 18095 11169 18107 11203
rect 18049 11163 18107 11169
rect 14461 11135 14519 11141
rect 14461 11132 14473 11135
rect 13780 11104 14473 11132
rect 13780 11092 13786 11104
rect 14461 11101 14473 11104
rect 14507 11101 14519 11135
rect 14461 11095 14519 11101
rect 15749 11135 15807 11141
rect 15749 11101 15761 11135
rect 15795 11101 15807 11135
rect 15749 11095 15807 11101
rect 16669 11135 16727 11141
rect 16669 11101 16681 11135
rect 16715 11101 16727 11135
rect 16669 11095 16727 11101
rect 17129 11135 17187 11141
rect 17129 11101 17141 11135
rect 17175 11132 17187 11135
rect 17218 11132 17224 11144
rect 17175 11104 17224 11132
rect 17175 11101 17187 11104
rect 17129 11095 17187 11101
rect 17218 11092 17224 11104
rect 17276 11092 17282 11144
rect 17770 11132 17776 11144
rect 17731 11104 17776 11132
rect 17770 11092 17776 11104
rect 17828 11092 17834 11144
rect 18340 11141 18368 11240
rect 18966 11228 18972 11240
rect 19024 11228 19030 11280
rect 20438 11228 20444 11280
rect 20496 11268 20502 11280
rect 20625 11271 20683 11277
rect 20625 11268 20637 11271
rect 20496 11240 20637 11268
rect 20496 11228 20502 11240
rect 20625 11237 20637 11240
rect 20671 11237 20683 11271
rect 20625 11231 20683 11237
rect 20809 11271 20867 11277
rect 20809 11237 20821 11271
rect 20855 11268 20867 11271
rect 21100 11268 21128 11308
rect 23106 11296 23112 11308
rect 23164 11296 23170 11348
rect 20855 11240 21128 11268
rect 20855 11237 20867 11240
rect 20809 11231 20867 11237
rect 22094 11228 22100 11280
rect 22152 11268 22158 11280
rect 22465 11271 22523 11277
rect 22465 11268 22477 11271
rect 22152 11240 22477 11268
rect 22152 11228 22158 11240
rect 22465 11237 22477 11240
rect 22511 11237 22523 11271
rect 22465 11231 22523 11237
rect 22741 11271 22799 11277
rect 22741 11237 22753 11271
rect 22787 11237 22799 11271
rect 22741 11231 22799 11237
rect 22925 11271 22983 11277
rect 22925 11237 22937 11271
rect 22971 11268 22983 11271
rect 23198 11268 23204 11280
rect 22971 11240 23204 11268
rect 22971 11237 22983 11240
rect 22925 11231 22983 11237
rect 18598 11160 18604 11212
rect 18656 11200 18662 11212
rect 19245 11203 19303 11209
rect 19245 11200 19257 11203
rect 18656 11172 19257 11200
rect 18656 11160 18662 11172
rect 18984 11144 19012 11172
rect 19245 11169 19257 11172
rect 19291 11169 19303 11203
rect 22756 11200 22784 11231
rect 23198 11228 23204 11240
rect 23256 11228 23262 11280
rect 23566 11200 23572 11212
rect 22756 11172 23572 11200
rect 19245 11163 19303 11169
rect 18325 11135 18383 11141
rect 18325 11101 18337 11135
rect 18371 11101 18383 11135
rect 18325 11095 18383 11101
rect 18966 11092 18972 11144
rect 19024 11092 19030 11144
rect 19260 11132 19288 11163
rect 23566 11160 23572 11172
rect 23624 11160 23630 11212
rect 21085 11135 21143 11141
rect 21085 11132 21097 11135
rect 19260 11104 21097 11132
rect 21085 11101 21097 11104
rect 21131 11101 21143 11135
rect 21085 11095 21143 11101
rect 21174 11092 21180 11144
rect 21232 11132 21238 11144
rect 21341 11135 21399 11141
rect 21341 11132 21353 11135
rect 21232 11104 21353 11132
rect 21232 11092 21238 11104
rect 21341 11101 21353 11104
rect 21387 11101 21399 11135
rect 21341 11095 21399 11101
rect 22186 11092 22192 11144
rect 22244 11132 22250 11144
rect 22557 11135 22615 11141
rect 22557 11132 22569 11135
rect 22244 11104 22569 11132
rect 22244 11092 22250 11104
rect 22557 11101 22569 11104
rect 22603 11101 22615 11135
rect 23106 11132 23112 11144
rect 23067 11104 23112 11132
rect 22557 11095 22615 11101
rect 23106 11092 23112 11104
rect 23164 11092 23170 11144
rect 13630 11024 13636 11076
rect 13688 11064 13694 11076
rect 15197 11067 15255 11073
rect 15197 11064 15209 11067
rect 13688 11036 15209 11064
rect 13688 11024 13694 11036
rect 15197 11033 15209 11036
rect 15243 11033 15255 11067
rect 15197 11027 15255 11033
rect 16025 11067 16083 11073
rect 16025 11033 16037 11067
rect 16071 11064 16083 11067
rect 18233 11067 18291 11073
rect 16071 11036 18184 11064
rect 16071 11033 16083 11036
rect 16025 11027 16083 11033
rect 13354 10996 13360 11008
rect 12124 10968 13360 10996
rect 12124 10956 12130 10968
rect 13354 10956 13360 10968
rect 13412 10956 13418 11008
rect 14366 10996 14372 11008
rect 14327 10968 14372 10996
rect 14366 10956 14372 10968
rect 14424 10956 14430 11008
rect 15289 10999 15347 11005
rect 15289 10965 15301 10999
rect 15335 10996 15347 10999
rect 15378 10996 15384 11008
rect 15335 10968 15384 10996
rect 15335 10965 15347 10968
rect 15289 10959 15347 10965
rect 15378 10956 15384 10968
rect 15436 10956 15442 11008
rect 18156 10996 18184 11036
rect 18233 11033 18245 11067
rect 18279 11064 18291 11067
rect 18690 11064 18696 11076
rect 18279 11036 18696 11064
rect 18279 11033 18291 11036
rect 18233 11027 18291 11033
rect 18690 11024 18696 11036
rect 18748 11024 18754 11076
rect 18877 11067 18935 11073
rect 18877 11033 18889 11067
rect 18923 11064 18935 11067
rect 18923 11036 19196 11064
rect 18923 11033 18935 11036
rect 18877 11027 18935 11033
rect 19058 10996 19064 11008
rect 18156 10968 19064 10996
rect 19058 10956 19064 10968
rect 19116 10956 19122 11008
rect 19168 10996 19196 11036
rect 19242 11024 19248 11076
rect 19300 11064 19306 11076
rect 19490 11067 19548 11073
rect 19490 11064 19502 11067
rect 19300 11036 19502 11064
rect 19300 11024 19306 11036
rect 19490 11033 19502 11036
rect 19536 11033 19548 11067
rect 19490 11027 19548 11033
rect 20548 11036 20852 11064
rect 20548 10996 20576 11036
rect 19168 10968 20576 10996
rect 20824 10996 20852 11036
rect 23014 10996 23020 11008
rect 20824 10968 23020 10996
rect 23014 10956 23020 10968
rect 23072 10956 23078 11008
rect 1104 10906 23460 10928
rect 1104 10854 6548 10906
rect 6600 10854 6612 10906
rect 6664 10854 6676 10906
rect 6728 10854 6740 10906
rect 6792 10854 6804 10906
rect 6856 10854 12146 10906
rect 12198 10854 12210 10906
rect 12262 10854 12274 10906
rect 12326 10854 12338 10906
rect 12390 10854 12402 10906
rect 12454 10854 17744 10906
rect 17796 10854 17808 10906
rect 17860 10854 17872 10906
rect 17924 10854 17936 10906
rect 17988 10854 18000 10906
rect 18052 10854 23460 10906
rect 1104 10832 23460 10854
rect 3418 10752 3424 10804
rect 3476 10792 3482 10804
rect 3973 10795 4031 10801
rect 3973 10792 3985 10795
rect 3476 10764 3985 10792
rect 3476 10752 3482 10764
rect 3973 10761 3985 10764
rect 4019 10761 4031 10795
rect 3973 10755 4031 10761
rect 4341 10795 4399 10801
rect 4341 10761 4353 10795
rect 4387 10792 4399 10795
rect 5166 10792 5172 10804
rect 4387 10764 5172 10792
rect 4387 10761 4399 10764
rect 4341 10755 4399 10761
rect 5166 10752 5172 10764
rect 5224 10752 5230 10804
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 7377 10795 7435 10801
rect 7377 10792 7389 10795
rect 7064 10764 7389 10792
rect 7064 10752 7070 10764
rect 7377 10761 7389 10764
rect 7423 10761 7435 10795
rect 7377 10755 7435 10761
rect 7837 10795 7895 10801
rect 7837 10761 7849 10795
rect 7883 10792 7895 10795
rect 8205 10795 8263 10801
rect 8205 10792 8217 10795
rect 7883 10764 8217 10792
rect 7883 10761 7895 10764
rect 7837 10755 7895 10761
rect 8205 10761 8217 10764
rect 8251 10761 8263 10795
rect 8662 10792 8668 10804
rect 8623 10764 8668 10792
rect 8205 10755 8263 10761
rect 8662 10752 8668 10764
rect 8720 10752 8726 10804
rect 8757 10795 8815 10801
rect 8757 10761 8769 10795
rect 8803 10792 8815 10795
rect 8938 10792 8944 10804
rect 8803 10764 8944 10792
rect 8803 10761 8815 10764
rect 8757 10755 8815 10761
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 9125 10795 9183 10801
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 10597 10795 10655 10801
rect 10597 10792 10609 10795
rect 9171 10764 10609 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 10597 10761 10609 10764
rect 10643 10761 10655 10795
rect 10597 10755 10655 10761
rect 10962 10752 10968 10804
rect 11020 10792 11026 10804
rect 11057 10795 11115 10801
rect 11057 10792 11069 10795
rect 11020 10764 11069 10792
rect 11020 10752 11026 10764
rect 11057 10761 11069 10764
rect 11103 10761 11115 10795
rect 11057 10755 11115 10761
rect 11974 10752 11980 10804
rect 12032 10792 12038 10804
rect 14001 10795 14059 10801
rect 14001 10792 14013 10795
rect 12032 10764 14013 10792
rect 12032 10752 12038 10764
rect 14001 10761 14013 10764
rect 14047 10761 14059 10795
rect 14366 10792 14372 10804
rect 14327 10764 14372 10792
rect 14001 10755 14059 10761
rect 14366 10752 14372 10764
rect 14424 10752 14430 10804
rect 14642 10752 14648 10804
rect 14700 10792 14706 10804
rect 15105 10795 15163 10801
rect 15105 10792 15117 10795
rect 14700 10764 15117 10792
rect 14700 10752 14706 10764
rect 15105 10761 15117 10764
rect 15151 10761 15163 10795
rect 15105 10755 15163 10761
rect 16945 10795 17003 10801
rect 16945 10761 16957 10795
rect 16991 10792 17003 10795
rect 17494 10792 17500 10804
rect 16991 10764 17500 10792
rect 16991 10761 17003 10764
rect 16945 10755 17003 10761
rect 17494 10752 17500 10764
rect 17552 10752 17558 10804
rect 19702 10792 19708 10804
rect 17972 10764 19708 10792
rect 5936 10727 5994 10733
rect 5936 10693 5948 10727
rect 5982 10724 5994 10727
rect 6914 10724 6920 10736
rect 5982 10696 6920 10724
rect 5982 10693 5994 10696
rect 5936 10687 5994 10693
rect 6914 10684 6920 10696
rect 6972 10684 6978 10736
rect 9217 10727 9275 10733
rect 9217 10693 9229 10727
rect 9263 10724 9275 10727
rect 9766 10724 9772 10736
rect 9263 10696 9772 10724
rect 9263 10693 9275 10696
rect 9217 10687 9275 10693
rect 9766 10684 9772 10696
rect 9824 10684 9830 10736
rect 10413 10727 10471 10733
rect 10413 10693 10425 10727
rect 10459 10724 10471 10727
rect 10502 10724 10508 10736
rect 10459 10696 10508 10724
rect 10459 10693 10471 10696
rect 10413 10687 10471 10693
rect 10502 10684 10508 10696
rect 10560 10684 10566 10736
rect 13906 10684 13912 10736
rect 13964 10724 13970 10736
rect 15841 10727 15899 10733
rect 15841 10724 15853 10727
rect 13964 10696 15853 10724
rect 13964 10684 13970 10696
rect 15841 10693 15853 10696
rect 15887 10693 15899 10727
rect 15841 10687 15899 10693
rect 16114 10684 16120 10736
rect 16172 10724 16178 10736
rect 16172 10696 17632 10724
rect 16172 10684 16178 10696
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 2021 10659 2079 10665
rect 2021 10656 2033 10659
rect 1912 10628 2033 10656
rect 1912 10616 1918 10628
rect 2021 10625 2033 10628
rect 2067 10625 2079 10659
rect 2021 10619 2079 10625
rect 3881 10659 3939 10665
rect 3881 10625 3893 10659
rect 3927 10656 3939 10659
rect 4798 10656 4804 10668
rect 3927 10628 4804 10656
rect 3927 10625 3939 10628
rect 3881 10619 3939 10625
rect 4798 10616 4804 10628
rect 4856 10616 4862 10668
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 6178 10656 6184 10668
rect 5408 10628 6184 10656
rect 5408 10616 5414 10628
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 7009 10659 7067 10665
rect 7009 10625 7021 10659
rect 7055 10656 7067 10659
rect 7282 10656 7288 10668
rect 7055 10628 7288 10656
rect 7055 10625 7067 10628
rect 7009 10619 7067 10625
rect 7282 10616 7288 10628
rect 7340 10656 7346 10668
rect 7469 10659 7527 10665
rect 7469 10656 7481 10659
rect 7340 10628 7481 10656
rect 7340 10616 7346 10628
rect 7469 10625 7481 10628
rect 7515 10625 7527 10659
rect 7469 10619 7527 10625
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10656 8355 10659
rect 8938 10656 8944 10668
rect 8343 10628 8944 10656
rect 8343 10625 8355 10628
rect 8297 10619 8355 10625
rect 8938 10616 8944 10628
rect 8996 10616 9002 10668
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10656 9643 10659
rect 10965 10659 11023 10665
rect 9631 10628 9812 10656
rect 9631 10625 9643 10628
rect 9585 10619 9643 10625
rect 1762 10588 1768 10600
rect 1723 10560 1768 10588
rect 1762 10548 1768 10560
rect 1820 10548 1826 10600
rect 4430 10588 4436 10600
rect 4391 10560 4436 10588
rect 4430 10548 4436 10560
rect 4488 10548 4494 10600
rect 4617 10591 4675 10597
rect 4617 10557 4629 10591
rect 4663 10588 4675 10591
rect 4890 10588 4896 10600
rect 4663 10560 4896 10588
rect 4663 10557 4675 10560
rect 4617 10551 4675 10557
rect 4890 10548 4896 10560
rect 4948 10548 4954 10600
rect 7193 10591 7251 10597
rect 7193 10557 7205 10591
rect 7239 10557 7251 10591
rect 7193 10551 7251 10557
rect 8113 10591 8171 10597
rect 8113 10557 8125 10591
rect 8159 10588 8171 10591
rect 8754 10588 8760 10600
rect 8159 10560 8760 10588
rect 8159 10557 8171 10560
rect 8113 10551 8171 10557
rect 3145 10523 3203 10529
rect 3145 10489 3157 10523
rect 3191 10520 3203 10523
rect 4154 10520 4160 10532
rect 3191 10492 4160 10520
rect 3191 10489 3203 10492
rect 3145 10483 3203 10489
rect 4154 10480 4160 10492
rect 4212 10480 4218 10532
rect 7208 10520 7236 10551
rect 8754 10548 8760 10560
rect 8812 10588 8818 10600
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 8812 10560 9321 10588
rect 8812 10548 8818 10560
rect 9309 10557 9321 10560
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 9674 10520 9680 10532
rect 7208 10492 9680 10520
rect 9674 10480 9680 10492
rect 9732 10480 9738 10532
rect 3237 10455 3295 10461
rect 3237 10421 3249 10455
rect 3283 10452 3295 10455
rect 4614 10452 4620 10464
rect 3283 10424 4620 10452
rect 3283 10421 3295 10424
rect 3237 10415 3295 10421
rect 4614 10412 4620 10424
rect 4672 10412 4678 10464
rect 4801 10455 4859 10461
rect 4801 10421 4813 10455
rect 4847 10452 4859 10455
rect 5442 10452 5448 10464
rect 4847 10424 5448 10452
rect 4847 10421 4859 10424
rect 4801 10415 4859 10421
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 6365 10455 6423 10461
rect 6365 10421 6377 10455
rect 6411 10452 6423 10455
rect 7466 10452 7472 10464
rect 6411 10424 7472 10452
rect 6411 10421 6423 10424
rect 6365 10415 6423 10421
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 9784 10452 9812 10628
rect 10965 10625 10977 10659
rect 11011 10656 11023 10659
rect 11330 10656 11336 10668
rect 11011 10628 11336 10656
rect 11011 10625 11023 10628
rect 10965 10619 11023 10625
rect 11330 10616 11336 10628
rect 11388 10616 11394 10668
rect 12066 10616 12072 10668
rect 12124 10656 12130 10668
rect 12161 10659 12219 10665
rect 12161 10656 12173 10659
rect 12124 10628 12173 10656
rect 12124 10616 12130 10628
rect 12161 10625 12173 10628
rect 12207 10625 12219 10659
rect 12161 10619 12219 10625
rect 12428 10659 12486 10665
rect 12428 10625 12440 10659
rect 12474 10656 12486 10659
rect 12710 10656 12716 10668
rect 12474 10628 12716 10656
rect 12474 10625 12486 10628
rect 12428 10619 12486 10625
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 13814 10616 13820 10668
rect 13872 10656 13878 10668
rect 14461 10659 14519 10665
rect 14461 10656 14473 10659
rect 13872 10628 14473 10656
rect 13872 10616 13878 10628
rect 14461 10625 14473 10628
rect 14507 10625 14519 10659
rect 14461 10619 14519 10625
rect 15197 10659 15255 10665
rect 15197 10625 15209 10659
rect 15243 10625 15255 10659
rect 15197 10619 15255 10625
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 17402 10656 17408 10668
rect 17083 10628 17408 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 10870 10548 10876 10600
rect 10928 10588 10934 10600
rect 11149 10591 11207 10597
rect 11149 10588 11161 10591
rect 10928 10560 11161 10588
rect 10928 10548 10934 10560
rect 11149 10557 11161 10560
rect 11195 10557 11207 10591
rect 11149 10551 11207 10557
rect 13725 10591 13783 10597
rect 13725 10557 13737 10591
rect 13771 10557 13783 10591
rect 13906 10588 13912 10600
rect 13867 10560 13912 10588
rect 13725 10551 13783 10557
rect 13538 10520 13544 10532
rect 13499 10492 13544 10520
rect 13538 10480 13544 10492
rect 13596 10480 13602 10532
rect 13740 10520 13768 10551
rect 13906 10548 13912 10560
rect 13964 10548 13970 10600
rect 13998 10520 14004 10532
rect 13740 10492 14004 10520
rect 13998 10480 14004 10492
rect 14056 10480 14062 10532
rect 11514 10452 11520 10464
rect 9784 10424 11520 10452
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 13556 10452 13584 10480
rect 15212 10452 15240 10619
rect 17402 10616 17408 10628
rect 17460 10616 17466 10668
rect 17604 10665 17632 10696
rect 17972 10665 18000 10764
rect 19702 10752 19708 10764
rect 19760 10752 19766 10804
rect 22462 10792 22468 10804
rect 22423 10764 22468 10792
rect 22462 10752 22468 10764
rect 22520 10752 22526 10804
rect 23109 10795 23167 10801
rect 23109 10761 23121 10795
rect 23155 10792 23167 10795
rect 23290 10792 23296 10804
rect 23155 10764 23296 10792
rect 23155 10761 23167 10764
rect 23109 10755 23167 10761
rect 23290 10752 23296 10764
rect 23348 10752 23354 10804
rect 20073 10727 20131 10733
rect 20073 10693 20085 10727
rect 20119 10724 20131 10727
rect 21174 10724 21180 10736
rect 20119 10696 21180 10724
rect 20119 10693 20131 10696
rect 20073 10687 20131 10693
rect 21174 10684 21180 10696
rect 21232 10684 21238 10736
rect 17589 10659 17647 10665
rect 17589 10625 17601 10659
rect 17635 10625 17647 10659
rect 17589 10619 17647 10625
rect 17957 10659 18015 10665
rect 17957 10625 17969 10659
rect 18003 10625 18015 10659
rect 17957 10619 18015 10625
rect 18156 10628 18460 10656
rect 16485 10591 16543 10597
rect 16485 10557 16497 10591
rect 16531 10588 16543 10591
rect 16666 10588 16672 10600
rect 16531 10560 16672 10588
rect 16531 10557 16543 10560
rect 16485 10551 16543 10557
rect 16666 10548 16672 10560
rect 16724 10548 16730 10600
rect 16853 10591 16911 10597
rect 16853 10557 16865 10591
rect 16899 10588 16911 10591
rect 17218 10588 17224 10600
rect 16899 10560 17224 10588
rect 16899 10557 16911 10560
rect 16853 10551 16911 10557
rect 17218 10548 17224 10560
rect 17276 10548 17282 10600
rect 18156 10588 18184 10628
rect 18322 10597 18328 10600
rect 17972 10560 18184 10588
rect 18280 10591 18328 10597
rect 17773 10523 17831 10529
rect 17773 10489 17785 10523
rect 17819 10520 17831 10523
rect 17972 10520 18000 10560
rect 18280 10557 18292 10591
rect 18326 10557 18328 10591
rect 18280 10551 18328 10557
rect 18322 10548 18328 10551
rect 18380 10548 18386 10600
rect 18432 10597 18460 10628
rect 18966 10616 18972 10668
rect 19024 10656 19030 10668
rect 20257 10659 20315 10665
rect 20257 10656 20269 10659
rect 19024 10628 20269 10656
rect 19024 10616 19030 10628
rect 20257 10625 20269 10628
rect 20303 10625 20315 10659
rect 20513 10659 20571 10665
rect 20513 10656 20525 10659
rect 20257 10619 20315 10625
rect 20364 10628 20525 10656
rect 18420 10591 18478 10597
rect 18420 10557 18432 10591
rect 18466 10588 18478 10591
rect 18506 10588 18512 10600
rect 18466 10560 18512 10588
rect 18466 10557 18478 10560
rect 18420 10551 18478 10557
rect 18506 10548 18512 10560
rect 18564 10548 18570 10600
rect 18690 10588 18696 10600
rect 18651 10560 18696 10588
rect 18690 10548 18696 10560
rect 18748 10548 18754 10600
rect 19058 10548 19064 10600
rect 19116 10588 19122 10600
rect 20364 10588 20392 10628
rect 20513 10625 20525 10628
rect 20559 10625 20571 10659
rect 20513 10619 20571 10625
rect 21082 10616 21088 10668
rect 21140 10656 21146 10668
rect 21821 10659 21879 10665
rect 21821 10656 21833 10659
rect 21140 10628 21833 10656
rect 21140 10616 21146 10628
rect 21821 10625 21833 10628
rect 21867 10625 21879 10659
rect 21821 10619 21879 10625
rect 22925 10659 22983 10665
rect 22925 10625 22937 10659
rect 22971 10656 22983 10659
rect 23934 10656 23940 10668
rect 22971 10628 23940 10656
rect 22971 10625 22983 10628
rect 22925 10619 22983 10625
rect 22554 10588 22560 10600
rect 19116 10560 20392 10588
rect 22515 10560 22560 10588
rect 19116 10548 19122 10560
rect 22554 10548 22560 10560
rect 22612 10548 22618 10600
rect 17819 10492 18000 10520
rect 17819 10489 17831 10492
rect 17773 10483 17831 10489
rect 21266 10480 21272 10532
rect 21324 10520 21330 10532
rect 22940 10520 22968 10619
rect 23934 10616 23940 10628
rect 23992 10616 23998 10668
rect 21324 10492 22968 10520
rect 21324 10480 21330 10492
rect 13556 10424 15240 10452
rect 16942 10412 16948 10464
rect 17000 10452 17006 10464
rect 17405 10455 17463 10461
rect 17405 10452 17417 10455
rect 17000 10424 17417 10452
rect 17000 10412 17006 10424
rect 17405 10421 17417 10424
rect 17451 10421 17463 10455
rect 17405 10415 17463 10421
rect 18506 10412 18512 10464
rect 18564 10452 18570 10464
rect 19058 10452 19064 10464
rect 18564 10424 19064 10452
rect 18564 10412 18570 10424
rect 19058 10412 19064 10424
rect 19116 10412 19122 10464
rect 19797 10455 19855 10461
rect 19797 10421 19809 10455
rect 19843 10452 19855 10455
rect 20254 10452 20260 10464
rect 19843 10424 20260 10452
rect 19843 10421 19855 10424
rect 19797 10415 19855 10421
rect 20254 10412 20260 10424
rect 20312 10412 20318 10464
rect 21634 10452 21640 10464
rect 21595 10424 21640 10452
rect 21634 10412 21640 10424
rect 21692 10412 21698 10464
rect 1104 10362 23460 10384
rect 1104 10310 3749 10362
rect 3801 10310 3813 10362
rect 3865 10310 3877 10362
rect 3929 10310 3941 10362
rect 3993 10310 4005 10362
rect 4057 10310 9347 10362
rect 9399 10310 9411 10362
rect 9463 10310 9475 10362
rect 9527 10310 9539 10362
rect 9591 10310 9603 10362
rect 9655 10310 14945 10362
rect 14997 10310 15009 10362
rect 15061 10310 15073 10362
rect 15125 10310 15137 10362
rect 15189 10310 15201 10362
rect 15253 10310 20543 10362
rect 20595 10310 20607 10362
rect 20659 10310 20671 10362
rect 20723 10310 20735 10362
rect 20787 10310 20799 10362
rect 20851 10310 23460 10362
rect 1104 10288 23460 10310
rect 1762 10208 1768 10260
rect 1820 10248 1826 10260
rect 1820 10220 3188 10248
rect 1820 10208 1826 10220
rect 3160 10121 3188 10220
rect 4430 10208 4436 10260
rect 4488 10248 4494 10260
rect 6181 10251 6239 10257
rect 6181 10248 6193 10251
rect 4488 10220 6193 10248
rect 4488 10208 4494 10220
rect 6181 10217 6193 10220
rect 6227 10217 6239 10251
rect 6181 10211 6239 10217
rect 7193 10251 7251 10257
rect 7193 10217 7205 10251
rect 7239 10248 7251 10251
rect 7282 10248 7288 10260
rect 7239 10220 7288 10248
rect 7239 10217 7251 10220
rect 7193 10211 7251 10217
rect 7282 10208 7288 10220
rect 7340 10208 7346 10260
rect 8938 10248 8944 10260
rect 8899 10220 8944 10248
rect 8938 10208 8944 10220
rect 8996 10208 9002 10260
rect 10870 10248 10876 10260
rect 9876 10220 10876 10248
rect 3605 10183 3663 10189
rect 3605 10149 3617 10183
rect 3651 10180 3663 10183
rect 4522 10180 4528 10192
rect 3651 10152 4528 10180
rect 3651 10149 3663 10152
rect 3605 10143 3663 10149
rect 4522 10140 4528 10152
rect 4580 10140 4586 10192
rect 6086 10180 6092 10192
rect 6047 10152 6092 10180
rect 6086 10140 6092 10152
rect 6144 10140 6150 10192
rect 3145 10115 3203 10121
rect 3145 10081 3157 10115
rect 3191 10112 3203 10115
rect 3191 10084 3832 10112
rect 3191 10081 3203 10084
rect 3145 10075 3203 10081
rect 3418 10044 3424 10056
rect 3379 10016 3424 10044
rect 3418 10004 3424 10016
rect 3476 10004 3482 10056
rect 3804 10044 3832 10084
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 4249 10115 4307 10121
rect 4249 10112 4261 10115
rect 3936 10084 4261 10112
rect 3936 10072 3942 10084
rect 4249 10081 4261 10084
rect 4295 10081 4307 10115
rect 4430 10112 4436 10124
rect 4391 10084 4436 10112
rect 4249 10075 4307 10081
rect 4430 10072 4436 10084
rect 4488 10072 4494 10124
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 6733 10115 6791 10121
rect 6733 10112 6745 10115
rect 6512 10084 6745 10112
rect 6512 10072 6518 10084
rect 6733 10081 6745 10084
rect 6779 10081 6791 10115
rect 6733 10075 6791 10081
rect 9493 10115 9551 10121
rect 9493 10081 9505 10115
rect 9539 10112 9551 10115
rect 9674 10112 9680 10124
rect 9539 10084 9680 10112
rect 9539 10081 9551 10084
rect 9493 10075 9551 10081
rect 9674 10072 9680 10084
rect 9732 10112 9738 10124
rect 9876 10112 9904 10220
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 11974 10248 11980 10260
rect 11935 10220 11980 10248
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 13630 10248 13636 10260
rect 13591 10220 13636 10248
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 14277 10251 14335 10257
rect 14277 10217 14289 10251
rect 14323 10248 14335 10251
rect 15378 10248 15384 10260
rect 14323 10220 15384 10248
rect 14323 10217 14335 10220
rect 14277 10211 14335 10217
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 16758 10208 16764 10260
rect 16816 10248 16822 10260
rect 17313 10251 17371 10257
rect 17313 10248 17325 10251
rect 16816 10220 17325 10248
rect 16816 10208 16822 10220
rect 17313 10217 17325 10220
rect 17359 10248 17371 10251
rect 19886 10248 19892 10260
rect 17359 10220 19288 10248
rect 19847 10220 19892 10248
rect 17359 10217 17371 10220
rect 17313 10211 17371 10217
rect 9732 10084 9904 10112
rect 18616 10084 19196 10112
rect 9732 10072 9738 10084
rect 4709 10047 4767 10053
rect 4709 10044 4721 10047
rect 3804 10016 4721 10044
rect 4709 10013 4721 10016
rect 4755 10044 4767 10047
rect 5350 10044 5356 10056
rect 4755 10016 5356 10044
rect 4755 10013 4767 10016
rect 4709 10007 4767 10013
rect 5350 10004 5356 10016
rect 5408 10004 5414 10056
rect 8294 10044 8300 10056
rect 8352 10053 8358 10056
rect 8264 10016 8300 10044
rect 8294 10004 8300 10016
rect 8352 10007 8364 10053
rect 8570 10044 8576 10056
rect 8483 10016 8576 10044
rect 8352 10004 8358 10007
rect 8570 10004 8576 10016
rect 8628 10044 8634 10056
rect 9582 10044 9588 10056
rect 8628 10016 9588 10044
rect 8628 10004 8634 10016
rect 9582 10004 9588 10016
rect 9640 10044 9646 10056
rect 9861 10047 9919 10053
rect 9861 10044 9873 10047
rect 9640 10016 9873 10044
rect 9640 10004 9646 10016
rect 9861 10013 9873 10016
rect 9907 10044 9919 10047
rect 10502 10044 10508 10056
rect 9907 10016 10508 10044
rect 9907 10013 9919 10016
rect 9861 10007 9919 10013
rect 10502 10004 10508 10016
rect 10560 10004 10566 10056
rect 13354 10044 13360 10056
rect 13315 10016 13360 10044
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 13446 10004 13452 10056
rect 13504 10044 13510 10056
rect 13504 10016 13549 10044
rect 13504 10004 13510 10016
rect 13998 10004 14004 10056
rect 14056 10044 14062 10056
rect 14093 10047 14151 10053
rect 14093 10044 14105 10047
rect 14056 10016 14105 10044
rect 14056 10004 14062 10016
rect 14093 10013 14105 10016
rect 14139 10013 14151 10047
rect 14093 10007 14151 10013
rect 15654 10004 15660 10056
rect 15712 10044 15718 10056
rect 15749 10047 15807 10053
rect 15749 10044 15761 10047
rect 15712 10016 15761 10044
rect 15712 10004 15718 10016
rect 15749 10013 15761 10016
rect 15795 10044 15807 10047
rect 15841 10047 15899 10053
rect 15841 10044 15853 10047
rect 15795 10016 15853 10044
rect 15795 10013 15807 10016
rect 15749 10007 15807 10013
rect 15841 10013 15853 10016
rect 15887 10044 15899 10047
rect 16390 10044 16396 10056
rect 15887 10016 16396 10044
rect 15887 10013 15899 10016
rect 15841 10007 15899 10013
rect 16390 10004 16396 10016
rect 16448 10004 16454 10056
rect 16482 10004 16488 10056
rect 16540 10044 16546 10056
rect 18138 10044 18144 10056
rect 16540 10016 18144 10044
rect 16540 10004 16546 10016
rect 18138 10004 18144 10016
rect 18196 10004 18202 10056
rect 18616 10044 18644 10084
rect 18340 10016 18644 10044
rect 18693 10047 18751 10053
rect 2900 9979 2958 9985
rect 2900 9945 2912 9979
rect 2946 9976 2958 9979
rect 4154 9976 4160 9988
rect 2946 9948 4016 9976
rect 4115 9948 4160 9976
rect 2946 9945 2958 9948
rect 2900 9939 2958 9945
rect 1765 9911 1823 9917
rect 1765 9877 1777 9911
rect 1811 9908 1823 9911
rect 2590 9908 2596 9920
rect 1811 9880 2596 9908
rect 1811 9877 1823 9880
rect 1765 9871 1823 9877
rect 2590 9868 2596 9880
rect 2648 9908 2654 9920
rect 3602 9908 3608 9920
rect 2648 9880 3608 9908
rect 2648 9868 2654 9880
rect 3602 9868 3608 9880
rect 3660 9868 3666 9920
rect 3786 9908 3792 9920
rect 3747 9880 3792 9908
rect 3786 9868 3792 9880
rect 3844 9868 3850 9920
rect 3988 9908 4016 9948
rect 4154 9936 4160 9948
rect 4212 9936 4218 9988
rect 4338 9976 4344 9988
rect 4255 9948 4344 9976
rect 4255 9908 4283 9948
rect 4338 9936 4344 9948
rect 4396 9936 4402 9988
rect 4614 9936 4620 9988
rect 4672 9976 4678 9988
rect 4954 9979 5012 9985
rect 4954 9976 4966 9979
rect 4672 9948 4966 9976
rect 4672 9936 4678 9948
rect 4954 9945 4966 9948
rect 5000 9945 5012 9979
rect 4954 9939 5012 9945
rect 9674 9936 9680 9988
rect 9732 9976 9738 9988
rect 10106 9979 10164 9985
rect 10106 9976 10118 9979
rect 9732 9948 10118 9976
rect 9732 9936 9738 9948
rect 10106 9945 10118 9948
rect 10152 9945 10164 9979
rect 10106 9939 10164 9945
rect 13112 9979 13170 9985
rect 13112 9945 13124 9979
rect 13158 9976 13170 9979
rect 15378 9976 15384 9988
rect 13158 9948 15384 9976
rect 13158 9945 13170 9948
rect 13112 9939 13170 9945
rect 15378 9936 15384 9948
rect 15436 9936 15442 9988
rect 15504 9979 15562 9985
rect 15504 9945 15516 9979
rect 15550 9976 15562 9979
rect 16108 9979 16166 9985
rect 15550 9948 16068 9976
rect 15550 9945 15562 9948
rect 15504 9939 15562 9945
rect 3988 9880 4283 9908
rect 4798 9868 4804 9920
rect 4856 9908 4862 9920
rect 6549 9911 6607 9917
rect 6549 9908 6561 9911
rect 4856 9880 6561 9908
rect 4856 9868 4862 9880
rect 6549 9877 6561 9880
rect 6595 9877 6607 9911
rect 6549 9871 6607 9877
rect 6641 9911 6699 9917
rect 6641 9877 6653 9911
rect 6687 9908 6699 9911
rect 6914 9908 6920 9920
rect 6687 9880 6920 9908
rect 6687 9877 6699 9880
rect 6641 9871 6699 9877
rect 6914 9868 6920 9880
rect 6972 9868 6978 9920
rect 8754 9868 8760 9920
rect 8812 9908 8818 9920
rect 9309 9911 9367 9917
rect 9309 9908 9321 9911
rect 8812 9880 9321 9908
rect 8812 9868 8818 9880
rect 9309 9877 9321 9880
rect 9355 9877 9367 9911
rect 9309 9871 9367 9877
rect 9398 9868 9404 9920
rect 9456 9908 9462 9920
rect 11241 9911 11299 9917
rect 9456 9880 9501 9908
rect 9456 9868 9462 9880
rect 11241 9877 11253 9911
rect 11287 9908 11299 9911
rect 11330 9908 11336 9920
rect 11287 9880 11336 9908
rect 11287 9877 11299 9880
rect 11241 9871 11299 9877
rect 11330 9868 11336 9880
rect 11388 9868 11394 9920
rect 13906 9868 13912 9920
rect 13964 9908 13970 9920
rect 14369 9911 14427 9917
rect 14369 9908 14381 9911
rect 13964 9880 14381 9908
rect 13964 9868 13970 9880
rect 14369 9877 14381 9880
rect 14415 9908 14427 9911
rect 15930 9908 15936 9920
rect 14415 9880 15936 9908
rect 14415 9877 14427 9880
rect 14369 9871 14427 9877
rect 15930 9868 15936 9880
rect 15988 9868 15994 9920
rect 16040 9908 16068 9948
rect 16108 9945 16120 9979
rect 16154 9976 16166 9979
rect 18340 9976 18368 10016
rect 18693 10013 18705 10047
rect 18739 10044 18751 10047
rect 18966 10044 18972 10056
rect 18739 10016 18972 10044
rect 18739 10013 18751 10016
rect 18693 10007 18751 10013
rect 18966 10004 18972 10016
rect 19024 10004 19030 10056
rect 19061 10047 19119 10053
rect 19061 10013 19073 10047
rect 19107 10013 19119 10047
rect 19061 10007 19119 10013
rect 16154 9948 18368 9976
rect 16154 9945 16166 9948
rect 16108 9939 16166 9945
rect 18414 9936 18420 9988
rect 18472 9985 18478 9988
rect 18472 9979 18506 9985
rect 18494 9945 18506 9979
rect 18874 9976 18880 9988
rect 18835 9948 18880 9976
rect 18472 9939 18506 9945
rect 18472 9936 18478 9939
rect 18874 9936 18880 9948
rect 18932 9936 18938 9988
rect 17126 9908 17132 9920
rect 16040 9880 17132 9908
rect 17126 9868 17132 9880
rect 17184 9868 17190 9920
rect 17218 9868 17224 9920
rect 17276 9908 17282 9920
rect 18598 9908 18604 9920
rect 17276 9880 18604 9908
rect 17276 9868 17282 9880
rect 18598 9868 18604 9880
rect 18656 9868 18662 9920
rect 19076 9908 19104 10007
rect 19168 9976 19196 10084
rect 19260 10053 19288 10220
rect 19886 10208 19892 10220
rect 19944 10208 19950 10260
rect 20898 10248 20904 10260
rect 19996 10220 20904 10248
rect 19996 10180 20024 10220
rect 20898 10208 20904 10220
rect 20956 10208 20962 10260
rect 21818 10248 21824 10260
rect 21779 10220 21824 10248
rect 21818 10208 21824 10220
rect 21876 10208 21882 10260
rect 21910 10208 21916 10260
rect 21968 10248 21974 10260
rect 22925 10251 22983 10257
rect 22925 10248 22937 10251
rect 21968 10220 22937 10248
rect 21968 10208 21974 10220
rect 22925 10217 22937 10220
rect 22971 10217 22983 10251
rect 22925 10211 22983 10217
rect 19628 10152 20024 10180
rect 19245 10047 19303 10053
rect 19245 10013 19257 10047
rect 19291 10013 19303 10047
rect 19245 10007 19303 10013
rect 19628 9976 19656 10152
rect 21634 10140 21640 10192
rect 21692 10180 21698 10192
rect 22830 10180 22836 10192
rect 21692 10152 22508 10180
rect 22791 10152 22836 10180
rect 21692 10140 21698 10152
rect 20487 10115 20545 10121
rect 20487 10081 20499 10115
rect 20533 10112 20545 10115
rect 21818 10112 21824 10124
rect 20533 10084 21824 10112
rect 20533 10081 20545 10084
rect 20487 10075 20545 10081
rect 21818 10072 21824 10084
rect 21876 10072 21882 10124
rect 22370 10112 22376 10124
rect 22331 10084 22376 10112
rect 22370 10072 22376 10084
rect 22428 10072 22434 10124
rect 22480 10121 22508 10152
rect 22830 10140 22836 10152
rect 22888 10140 22894 10192
rect 22465 10115 22523 10121
rect 22465 10081 22477 10115
rect 22511 10081 22523 10115
rect 22465 10075 22523 10081
rect 19702 10004 19708 10056
rect 19760 10044 19766 10056
rect 19981 10047 20039 10053
rect 19981 10044 19993 10047
rect 19760 10016 19993 10044
rect 19760 10004 19766 10016
rect 19981 10013 19993 10016
rect 20027 10013 20039 10047
rect 19981 10007 20039 10013
rect 20254 10004 20260 10056
rect 20312 10044 20318 10056
rect 20717 10047 20775 10053
rect 20717 10044 20729 10047
rect 20312 10016 20729 10044
rect 20312 10004 20318 10016
rect 20717 10013 20729 10016
rect 20763 10044 20775 10047
rect 20763 10016 22324 10044
rect 20763 10013 20775 10016
rect 20717 10007 20775 10013
rect 22296 9985 22324 10016
rect 23014 10004 23020 10056
rect 23072 10044 23078 10056
rect 23109 10047 23167 10053
rect 23109 10044 23121 10047
rect 23072 10016 23121 10044
rect 23072 10004 23078 10016
rect 23109 10013 23121 10016
rect 23155 10013 23167 10047
rect 23109 10007 23167 10013
rect 19168 9948 19656 9976
rect 22281 9979 22339 9985
rect 22281 9945 22293 9979
rect 22327 9945 22339 9979
rect 22281 9939 22339 9945
rect 19978 9908 19984 9920
rect 19076 9880 19984 9908
rect 19978 9868 19984 9880
rect 20036 9908 20042 9920
rect 20447 9911 20505 9917
rect 20447 9908 20459 9911
rect 20036 9880 20459 9908
rect 20036 9868 20042 9880
rect 20447 9877 20459 9880
rect 20493 9877 20505 9911
rect 20447 9871 20505 9877
rect 21913 9911 21971 9917
rect 21913 9877 21925 9911
rect 21959 9908 21971 9911
rect 22094 9908 22100 9920
rect 21959 9880 22100 9908
rect 21959 9877 21971 9880
rect 21913 9871 21971 9877
rect 22094 9868 22100 9880
rect 22152 9868 22158 9920
rect 1104 9818 23460 9840
rect 1104 9766 6548 9818
rect 6600 9766 6612 9818
rect 6664 9766 6676 9818
rect 6728 9766 6740 9818
rect 6792 9766 6804 9818
rect 6856 9766 12146 9818
rect 12198 9766 12210 9818
rect 12262 9766 12274 9818
rect 12326 9766 12338 9818
rect 12390 9766 12402 9818
rect 12454 9766 17744 9818
rect 17796 9766 17808 9818
rect 17860 9766 17872 9818
rect 17924 9766 17936 9818
rect 17988 9766 18000 9818
rect 18052 9766 23460 9818
rect 1104 9744 23460 9766
rect 2961 9707 3019 9713
rect 2961 9673 2973 9707
rect 3007 9704 3019 9707
rect 3786 9704 3792 9716
rect 3007 9676 3792 9704
rect 3007 9673 3019 9676
rect 2961 9667 3019 9673
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 4798 9704 4804 9716
rect 4759 9676 4804 9704
rect 4798 9664 4804 9676
rect 4856 9664 4862 9716
rect 8757 9707 8815 9713
rect 8757 9704 8769 9707
rect 7300 9676 8769 9704
rect 3053 9639 3111 9645
rect 3053 9605 3065 9639
rect 3099 9636 3111 9639
rect 3234 9636 3240 9648
rect 3099 9608 3240 9636
rect 3099 9605 3111 9608
rect 3053 9599 3111 9605
rect 3234 9596 3240 9608
rect 3292 9596 3298 9648
rect 3973 9639 4031 9645
rect 3973 9605 3985 9639
rect 4019 9636 4031 9639
rect 5350 9636 5356 9648
rect 4019 9608 5356 9636
rect 4019 9605 4031 9608
rect 3973 9599 4031 9605
rect 5350 9596 5356 9608
rect 5408 9636 5414 9648
rect 5408 9608 6224 9636
rect 5408 9596 5414 9608
rect 1394 9568 1400 9580
rect 1355 9540 1400 9568
rect 1394 9528 1400 9540
rect 1452 9568 1458 9580
rect 1673 9571 1731 9577
rect 1673 9568 1685 9571
rect 1452 9540 1685 9568
rect 1452 9528 1458 9540
rect 1673 9537 1685 9540
rect 1719 9537 1731 9571
rect 1673 9531 1731 9537
rect 2593 9571 2651 9577
rect 2593 9537 2605 9571
rect 2639 9568 2651 9571
rect 3326 9568 3332 9580
rect 2639 9540 3332 9568
rect 2639 9537 2651 9540
rect 2593 9531 2651 9537
rect 3326 9528 3332 9540
rect 3384 9528 3390 9580
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9568 3571 9571
rect 4522 9568 4528 9580
rect 3559 9540 4528 9568
rect 3559 9537 3571 9540
rect 3513 9531 3571 9537
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 4709 9571 4767 9577
rect 4709 9537 4721 9571
rect 4755 9568 4767 9571
rect 5534 9568 5540 9580
rect 4755 9540 5540 9568
rect 4755 9537 4767 9540
rect 4709 9531 4767 9537
rect 5534 9528 5540 9540
rect 5592 9528 5598 9580
rect 6196 9577 6224 9608
rect 7300 9577 7328 9676
rect 8757 9673 8769 9676
rect 8803 9704 8815 9707
rect 9398 9704 9404 9716
rect 8803 9676 9404 9704
rect 8803 9673 8815 9676
rect 8757 9667 8815 9673
rect 9398 9664 9404 9676
rect 9456 9664 9462 9716
rect 10962 9704 10968 9716
rect 10923 9676 10968 9704
rect 10962 9664 10968 9676
rect 11020 9664 11026 9716
rect 11514 9664 11520 9716
rect 11572 9704 11578 9716
rect 17135 9707 17193 9713
rect 17135 9704 17147 9707
rect 11572 9676 14136 9704
rect 11572 9664 11578 9676
rect 14108 9648 14136 9676
rect 16592 9676 17147 9704
rect 8570 9636 8576 9648
rect 7392 9608 8576 9636
rect 7392 9577 7420 9608
rect 8570 9596 8576 9608
rect 8628 9596 8634 9648
rect 8849 9639 8907 9645
rect 8849 9605 8861 9639
rect 8895 9636 8907 9639
rect 9674 9636 9680 9648
rect 8895 9608 9680 9636
rect 8895 9605 8907 9608
rect 8849 9599 8907 9605
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 12710 9636 12716 9648
rect 12671 9608 12716 9636
rect 12710 9596 12716 9608
rect 12768 9596 12774 9648
rect 14090 9596 14096 9648
rect 14148 9636 14154 9648
rect 14829 9639 14887 9645
rect 14829 9636 14841 9639
rect 14148 9608 14841 9636
rect 14148 9596 14154 9608
rect 14829 9605 14841 9608
rect 14875 9605 14887 9639
rect 15654 9636 15660 9648
rect 15615 9608 15660 9636
rect 14829 9599 14887 9605
rect 15654 9596 15660 9608
rect 15712 9596 15718 9648
rect 16592 9636 16620 9676
rect 17135 9673 17147 9676
rect 17181 9704 17193 9707
rect 18322 9704 18328 9716
rect 17181 9676 18328 9704
rect 17181 9673 17193 9676
rect 17135 9667 17193 9673
rect 18322 9664 18328 9676
rect 18380 9704 18386 9716
rect 18509 9707 18567 9713
rect 18380 9676 18460 9704
rect 18380 9664 18386 9676
rect 15764 9608 16620 9636
rect 18432 9636 18460 9676
rect 18509 9673 18521 9707
rect 18555 9704 18567 9707
rect 18690 9704 18696 9716
rect 18555 9676 18696 9704
rect 18555 9673 18567 9676
rect 18509 9667 18567 9673
rect 18690 9664 18696 9676
rect 18748 9664 18754 9716
rect 21818 9704 21824 9716
rect 21779 9676 21824 9704
rect 21818 9664 21824 9676
rect 21876 9664 21882 9716
rect 22189 9707 22247 9713
rect 22189 9673 22201 9707
rect 22235 9704 22247 9707
rect 22554 9704 22560 9716
rect 22235 9676 22560 9704
rect 22235 9673 22247 9676
rect 22189 9667 22247 9673
rect 22554 9664 22560 9676
rect 22612 9664 22618 9716
rect 18874 9636 18880 9648
rect 18432 9608 18880 9636
rect 5925 9571 5983 9577
rect 5925 9537 5937 9571
rect 5971 9568 5983 9571
rect 6181 9571 6239 9577
rect 5971 9540 6132 9568
rect 5971 9537 5983 9540
rect 5925 9531 5983 9537
rect 2866 9500 2872 9512
rect 2827 9472 2872 9500
rect 2866 9460 2872 9472
rect 2924 9460 2930 9512
rect 6104 9500 6132 9540
rect 6181 9537 6193 9571
rect 6227 9537 6239 9571
rect 6181 9531 6239 9537
rect 7285 9571 7343 9577
rect 7285 9537 7297 9571
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 7377 9571 7435 9577
rect 7377 9537 7389 9571
rect 7423 9537 7435 9571
rect 7377 9531 7435 9537
rect 7466 9528 7472 9580
rect 7524 9568 7530 9580
rect 7633 9571 7691 9577
rect 7633 9568 7645 9571
rect 7524 9540 7645 9568
rect 7524 9528 7530 9540
rect 7633 9537 7645 9540
rect 7679 9537 7691 9571
rect 7633 9531 7691 9537
rect 9493 9571 9551 9577
rect 9493 9537 9505 9571
rect 9539 9537 9551 9571
rect 9493 9531 9551 9537
rect 7190 9500 7196 9512
rect 6104 9472 7196 9500
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 3421 9435 3479 9441
rect 3421 9401 3433 9435
rect 3467 9432 3479 9435
rect 3510 9432 3516 9444
rect 3467 9404 3516 9432
rect 3467 9401 3479 9404
rect 3421 9395 3479 9401
rect 3510 9392 3516 9404
rect 3568 9392 3574 9444
rect 3697 9435 3755 9441
rect 3697 9401 3709 9435
rect 3743 9432 3755 9435
rect 4706 9432 4712 9444
rect 3743 9404 4712 9432
rect 3743 9401 3755 9404
rect 3697 9395 3755 9401
rect 4706 9392 4712 9404
rect 4764 9392 4770 9444
rect 1486 9324 1492 9376
rect 1544 9364 1550 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 1544 9336 1593 9364
rect 1544 9324 1550 9336
rect 1581 9333 1593 9336
rect 1627 9333 1639 9367
rect 1581 9327 1639 9333
rect 1949 9367 2007 9373
rect 1949 9333 1961 9367
rect 1995 9364 2007 9367
rect 2498 9364 2504 9376
rect 1995 9336 2504 9364
rect 1995 9333 2007 9336
rect 1949 9327 2007 9333
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 6638 9364 6644 9376
rect 6599 9336 6644 9364
rect 6638 9324 6644 9336
rect 6696 9324 6702 9376
rect 9508 9364 9536 9531
rect 9582 9528 9588 9580
rect 9640 9568 9646 9580
rect 9858 9577 9864 9580
rect 9640 9540 9685 9568
rect 9640 9528 9646 9540
rect 9852 9531 9864 9577
rect 9916 9568 9922 9580
rect 9916 9540 9952 9568
rect 9858 9528 9864 9531
rect 9916 9528 9922 9540
rect 11974 9528 11980 9580
rect 12032 9568 12038 9580
rect 12069 9571 12127 9577
rect 12069 9568 12081 9571
rect 12032 9540 12081 9568
rect 12032 9528 12038 9540
rect 12069 9537 12081 9540
rect 12115 9537 12127 9571
rect 13262 9568 13268 9580
rect 13223 9540 13268 9568
rect 12069 9531 12127 9537
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 14366 9568 14372 9580
rect 14327 9540 14372 9568
rect 14366 9528 14372 9540
rect 14424 9528 14430 9580
rect 15764 9568 15792 9608
rect 18874 9596 18880 9608
rect 18932 9596 18938 9648
rect 21174 9636 21180 9648
rect 21135 9608 21180 9636
rect 21174 9596 21180 9608
rect 21232 9596 21238 9648
rect 22094 9596 22100 9648
rect 22152 9636 22158 9648
rect 22281 9639 22339 9645
rect 22281 9636 22293 9639
rect 22152 9608 22293 9636
rect 22152 9596 22158 9608
rect 22281 9605 22293 9608
rect 22327 9605 22339 9639
rect 23106 9636 23112 9648
rect 23067 9608 23112 9636
rect 22281 9599 22339 9605
rect 23106 9596 23112 9608
rect 23164 9596 23170 9648
rect 14844 9540 15792 9568
rect 15841 9571 15899 9577
rect 14844 9512 14872 9540
rect 15841 9537 15853 9571
rect 15887 9568 15899 9571
rect 15930 9568 15936 9580
rect 15887 9540 15936 9568
rect 15887 9537 15899 9540
rect 15841 9531 15899 9537
rect 15930 9528 15936 9540
rect 15988 9528 15994 9580
rect 17402 9568 17408 9580
rect 16592 9540 17408 9568
rect 14458 9500 14464 9512
rect 14419 9472 14464 9500
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 14553 9503 14611 9509
rect 14553 9469 14565 9503
rect 14599 9469 14611 9503
rect 14553 9463 14611 9469
rect 13998 9432 14004 9444
rect 13959 9404 14004 9432
rect 13998 9392 14004 9404
rect 14056 9392 14062 9444
rect 14274 9392 14280 9444
rect 14332 9432 14338 9444
rect 14568 9432 14596 9463
rect 14826 9460 14832 9512
rect 14884 9460 14890 9512
rect 15378 9460 15384 9512
rect 15436 9500 15442 9512
rect 16485 9503 16543 9509
rect 16485 9500 16497 9503
rect 15436 9472 16497 9500
rect 15436 9460 15442 9472
rect 16485 9469 16497 9472
rect 16531 9469 16543 9503
rect 16485 9463 16543 9469
rect 14332 9404 14596 9432
rect 14332 9392 14338 9404
rect 14734 9392 14740 9444
rect 14792 9432 14798 9444
rect 16592 9432 16620 9540
rect 17402 9528 17408 9540
rect 17460 9528 17466 9580
rect 18598 9568 18604 9580
rect 18559 9540 18604 9568
rect 18598 9528 18604 9540
rect 18656 9528 18662 9580
rect 18966 9528 18972 9580
rect 19024 9568 19030 9580
rect 19337 9571 19395 9577
rect 19337 9568 19349 9571
rect 19024 9540 19349 9568
rect 19024 9528 19030 9540
rect 19337 9537 19349 9540
rect 19383 9537 19395 9571
rect 19337 9531 19395 9537
rect 19604 9571 19662 9577
rect 19604 9537 19616 9571
rect 19650 9568 19662 9571
rect 21542 9568 21548 9580
rect 19650 9540 21548 9568
rect 19650 9537 19662 9540
rect 19604 9531 19662 9537
rect 21542 9528 21548 9540
rect 21600 9528 21606 9580
rect 22830 9568 22836 9580
rect 22791 9540 22836 9568
rect 22830 9528 22836 9540
rect 22888 9528 22894 9580
rect 16669 9503 16727 9509
rect 16669 9469 16681 9503
rect 16715 9500 16727 9503
rect 16850 9500 16856 9512
rect 16715 9472 16856 9500
rect 16715 9469 16727 9472
rect 16669 9463 16727 9469
rect 16850 9460 16856 9472
rect 16908 9460 16914 9512
rect 17175 9503 17233 9509
rect 17175 9469 17187 9503
rect 17221 9500 17233 9503
rect 17310 9500 17316 9512
rect 17221 9472 17316 9500
rect 17221 9469 17233 9472
rect 17175 9463 17233 9469
rect 17310 9460 17316 9472
rect 17368 9460 17374 9512
rect 18414 9460 18420 9512
rect 18472 9500 18478 9512
rect 19245 9503 19303 9509
rect 19245 9500 19257 9503
rect 18472 9472 19257 9500
rect 18472 9460 18478 9472
rect 19245 9469 19257 9472
rect 19291 9469 19303 9503
rect 19245 9463 19303 9469
rect 21174 9460 21180 9512
rect 21232 9500 21238 9512
rect 21269 9503 21327 9509
rect 21269 9500 21281 9503
rect 21232 9472 21281 9500
rect 21232 9460 21238 9472
rect 21269 9469 21281 9472
rect 21315 9469 21327 9503
rect 21269 9463 21327 9469
rect 21453 9503 21511 9509
rect 21453 9469 21465 9503
rect 21499 9469 21511 9503
rect 21453 9463 21511 9469
rect 22465 9503 22523 9509
rect 22465 9469 22477 9503
rect 22511 9500 22523 9503
rect 23106 9500 23112 9512
rect 22511 9472 23112 9500
rect 22511 9469 22523 9472
rect 22465 9463 22523 9469
rect 14792 9404 16620 9432
rect 20717 9435 20775 9441
rect 14792 9392 14798 9404
rect 20717 9401 20729 9435
rect 20763 9432 20775 9435
rect 21358 9432 21364 9444
rect 20763 9404 21364 9432
rect 20763 9401 20775 9404
rect 20717 9395 20775 9401
rect 21358 9392 21364 9404
rect 21416 9432 21422 9444
rect 21468 9432 21496 9463
rect 23106 9460 23112 9472
rect 23164 9460 23170 9512
rect 21416 9404 21496 9432
rect 21416 9392 21422 9404
rect 21726 9392 21732 9444
rect 21784 9432 21790 9444
rect 22649 9435 22707 9441
rect 22649 9432 22661 9435
rect 21784 9404 22661 9432
rect 21784 9392 21790 9404
rect 22649 9401 22661 9404
rect 22695 9401 22707 9435
rect 22649 9395 22707 9401
rect 10962 9364 10968 9376
rect 9508 9336 10968 9364
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 13906 9364 13912 9376
rect 13867 9336 13912 9364
rect 13906 9324 13912 9336
rect 13964 9324 13970 9376
rect 16298 9324 16304 9376
rect 16356 9364 16362 9376
rect 17034 9364 17040 9376
rect 16356 9336 17040 9364
rect 16356 9324 16362 9336
rect 17034 9324 17040 9336
rect 17092 9324 17098 9376
rect 20809 9367 20867 9373
rect 20809 9333 20821 9367
rect 20855 9364 20867 9367
rect 20990 9364 20996 9376
rect 20855 9336 20996 9364
rect 20855 9333 20867 9336
rect 20809 9327 20867 9333
rect 20990 9324 20996 9336
rect 21048 9364 21054 9376
rect 21450 9364 21456 9376
rect 21048 9336 21456 9364
rect 21048 9324 21054 9336
rect 21450 9324 21456 9336
rect 21508 9324 21514 9376
rect 1104 9274 23460 9296
rect 1104 9222 3749 9274
rect 3801 9222 3813 9274
rect 3865 9222 3877 9274
rect 3929 9222 3941 9274
rect 3993 9222 4005 9274
rect 4057 9222 9347 9274
rect 9399 9222 9411 9274
rect 9463 9222 9475 9274
rect 9527 9222 9539 9274
rect 9591 9222 9603 9274
rect 9655 9222 14945 9274
rect 14997 9222 15009 9274
rect 15061 9222 15073 9274
rect 15125 9222 15137 9274
rect 15189 9222 15201 9274
rect 15253 9222 20543 9274
rect 20595 9222 20607 9274
rect 20659 9222 20671 9274
rect 20723 9222 20735 9274
rect 20787 9222 20799 9274
rect 20851 9222 23460 9274
rect 1104 9200 23460 9222
rect 1762 9160 1768 9172
rect 1412 9132 1768 9160
rect 1412 9033 1440 9132
rect 1762 9120 1768 9132
rect 1820 9120 1826 9172
rect 3418 9120 3424 9172
rect 3476 9160 3482 9172
rect 3605 9163 3663 9169
rect 3605 9160 3617 9163
rect 3476 9132 3617 9160
rect 3476 9120 3482 9132
rect 3605 9129 3617 9132
rect 3651 9129 3663 9163
rect 4522 9160 4528 9172
rect 4483 9132 4528 9160
rect 3605 9123 3663 9129
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 5445 9163 5503 9169
rect 5445 9129 5457 9163
rect 5491 9160 5503 9163
rect 5534 9160 5540 9172
rect 5491 9132 5540 9160
rect 5491 9129 5503 9132
rect 5445 9123 5503 9129
rect 5534 9120 5540 9132
rect 5592 9120 5598 9172
rect 11422 9160 11428 9172
rect 6886 9132 11428 9160
rect 3142 9052 3148 9104
rect 3200 9092 3206 9104
rect 3789 9095 3847 9101
rect 3789 9092 3801 9095
rect 3200 9064 3801 9092
rect 3200 9052 3206 9064
rect 3789 9061 3801 9064
rect 3835 9061 3847 9095
rect 3789 9055 3847 9061
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 8993 1455 9027
rect 1397 8987 1455 8993
rect 2866 8984 2872 9036
rect 2924 9024 2930 9036
rect 3053 9027 3111 9033
rect 3053 9024 3065 9027
rect 2924 8996 3065 9024
rect 2924 8984 2930 8996
rect 3053 8993 3065 8996
rect 3099 9024 3111 9027
rect 4890 9024 4896 9036
rect 3099 8996 4896 9024
rect 3099 8993 3111 8996
rect 3053 8987 3111 8993
rect 4890 8984 4896 8996
rect 4948 9024 4954 9036
rect 5077 9027 5135 9033
rect 5077 9024 5089 9027
rect 4948 8996 5089 9024
rect 4948 8984 4954 8996
rect 5077 8993 5089 8996
rect 5123 8993 5135 9027
rect 5077 8987 5135 8993
rect 5350 8984 5356 9036
rect 5408 9024 5414 9036
rect 5537 9027 5595 9033
rect 5537 9024 5549 9027
rect 5408 8996 5549 9024
rect 5408 8984 5414 8996
rect 5537 8993 5549 8996
rect 5583 8993 5595 9027
rect 5537 8987 5595 8993
rect 1486 8916 1492 8968
rect 1544 8956 1550 8968
rect 1653 8959 1711 8965
rect 1653 8956 1665 8959
rect 1544 8928 1665 8956
rect 1544 8916 1550 8928
rect 1653 8925 1665 8928
rect 1699 8925 1711 8959
rect 1653 8919 1711 8925
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 4433 8959 4491 8965
rect 4433 8956 4445 8959
rect 4212 8928 4445 8956
rect 4212 8916 4218 8928
rect 4433 8925 4445 8928
rect 4479 8925 4491 8959
rect 6886 8956 6914 9132
rect 11422 9120 11428 9132
rect 11480 9120 11486 9172
rect 13446 9160 13452 9172
rect 13407 9132 13452 9160
rect 13446 9120 13452 9132
rect 13504 9120 13510 9172
rect 14090 9120 14096 9172
rect 14148 9160 14154 9172
rect 14185 9163 14243 9169
rect 14185 9160 14197 9163
rect 14148 9132 14197 9160
rect 14148 9120 14154 9132
rect 14185 9129 14197 9132
rect 14231 9160 14243 9163
rect 18969 9163 19027 9169
rect 18969 9160 18981 9163
rect 14231 9132 18981 9160
rect 14231 9129 14243 9132
rect 14185 9123 14243 9129
rect 18969 9129 18981 9132
rect 19015 9160 19027 9163
rect 19426 9160 19432 9172
rect 19015 9132 19432 9160
rect 19015 9129 19027 9132
rect 18969 9123 19027 9129
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 21542 9160 21548 9172
rect 20364 9132 21036 9160
rect 21503 9132 21548 9160
rect 8386 9052 8392 9104
rect 8444 9092 8450 9104
rect 8754 9092 8760 9104
rect 8444 9064 8760 9092
rect 8444 9052 8450 9064
rect 8754 9052 8760 9064
rect 8812 9052 8818 9104
rect 16850 9052 16856 9104
rect 16908 9092 16914 9104
rect 16908 9064 17071 9092
rect 16908 9052 16914 9064
rect 10502 8984 10508 9036
rect 10560 9024 10566 9036
rect 11241 9027 11299 9033
rect 11241 9024 11253 9027
rect 10560 8996 11253 9024
rect 10560 8984 10566 8996
rect 11241 8993 11253 8996
rect 11287 8993 11299 9027
rect 11241 8987 11299 8993
rect 12897 9027 12955 9033
rect 12897 8993 12909 9027
rect 12943 9024 12955 9027
rect 14274 9024 14280 9036
rect 12943 8996 14280 9024
rect 12943 8993 12955 8996
rect 12897 8987 12955 8993
rect 4433 8919 4491 8925
rect 5644 8928 6914 8956
rect 7377 8959 7435 8965
rect 3145 8891 3203 8897
rect 3145 8857 3157 8891
rect 3191 8888 3203 8891
rect 4338 8888 4344 8900
rect 3191 8860 4344 8888
rect 3191 8857 3203 8860
rect 3145 8851 3203 8857
rect 4338 8848 4344 8860
rect 4396 8848 4402 8900
rect 4706 8848 4712 8900
rect 4764 8888 4770 8900
rect 5644 8888 5672 8928
rect 7377 8925 7389 8959
rect 7423 8956 7435 8959
rect 8386 8956 8392 8968
rect 7423 8928 8392 8956
rect 7423 8925 7435 8928
rect 7377 8919 7435 8925
rect 8386 8916 8392 8928
rect 8444 8956 8450 8968
rect 9125 8959 9183 8965
rect 9125 8956 9137 8959
rect 8444 8928 9137 8956
rect 8444 8916 8450 8928
rect 9125 8925 9137 8928
rect 9171 8956 9183 8959
rect 10520 8956 10548 8984
rect 9171 8928 10548 8956
rect 11256 8956 11284 8987
rect 14274 8984 14280 8996
rect 14332 8984 14338 9036
rect 15378 8984 15384 9036
rect 15436 9024 15442 9036
rect 16758 9024 16764 9036
rect 15436 8996 15884 9024
rect 16719 8996 16764 9024
rect 15436 8984 15442 8996
rect 11974 8956 11980 8968
rect 11256 8928 11980 8956
rect 9171 8925 9183 8928
rect 9125 8919 9183 8925
rect 11974 8916 11980 8928
rect 12032 8916 12038 8968
rect 13446 8916 13452 8968
rect 13504 8956 13510 8968
rect 14369 8959 14427 8965
rect 14369 8956 14381 8959
rect 13504 8928 14381 8956
rect 13504 8916 13510 8928
rect 14369 8925 14381 8928
rect 14415 8956 14427 8959
rect 15654 8956 15660 8968
rect 14415 8928 15660 8956
rect 14415 8925 14427 8928
rect 14369 8919 14427 8925
rect 15654 8916 15660 8928
rect 15712 8916 15718 8968
rect 15856 8965 15884 8996
rect 16758 8984 16764 8996
rect 16816 8984 16822 9036
rect 16942 9024 16948 9036
rect 16903 8996 16948 9024
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 17043 9024 17071 9064
rect 17310 9052 17316 9104
rect 17368 9092 17374 9104
rect 17405 9095 17463 9101
rect 17405 9092 17417 9095
rect 17368 9064 17417 9092
rect 17368 9052 17374 9064
rect 17405 9061 17417 9064
rect 17451 9061 17463 9095
rect 19702 9092 19708 9104
rect 17405 9055 17463 9061
rect 18064 9064 19708 9092
rect 18064 9033 18092 9064
rect 19702 9052 19708 9064
rect 19760 9052 19766 9104
rect 18049 9027 18107 9033
rect 17043 8996 17172 9024
rect 15841 8959 15899 8965
rect 15841 8925 15853 8959
rect 15887 8925 15899 8959
rect 15841 8919 15899 8925
rect 16666 8916 16672 8968
rect 16724 8956 16730 8968
rect 17037 8959 17095 8965
rect 17037 8956 17049 8959
rect 16724 8928 17049 8956
rect 16724 8916 16730 8928
rect 17037 8925 17049 8928
rect 17083 8925 17095 8959
rect 17144 8956 17172 8996
rect 18049 8993 18061 9027
rect 18095 8993 18107 9027
rect 18049 8987 18107 8993
rect 18966 8984 18972 9036
rect 19024 9024 19030 9036
rect 19610 9024 19616 9036
rect 19024 8996 19616 9024
rect 19024 8984 19030 8996
rect 19610 8984 19616 8996
rect 19668 9024 19674 9036
rect 20364 9024 20392 9132
rect 20438 9052 20444 9104
rect 20496 9092 20502 9104
rect 20496 9064 20944 9092
rect 20496 9052 20502 9064
rect 20625 9027 20683 9033
rect 20625 9024 20637 9027
rect 19668 8996 20637 9024
rect 19668 8984 19674 8996
rect 20625 8993 20637 8996
rect 20671 8993 20683 9027
rect 20625 8987 20683 8993
rect 18325 8959 18383 8965
rect 18325 8956 18337 8959
rect 17144 8928 18337 8956
rect 17037 8919 17095 8925
rect 18325 8925 18337 8928
rect 18371 8956 18383 8959
rect 19242 8956 19248 8968
rect 18371 8928 19248 8956
rect 18371 8925 18383 8928
rect 18325 8919 18383 8925
rect 19242 8916 19248 8928
rect 19300 8916 19306 8968
rect 20916 8965 20944 9064
rect 21008 9024 21036 9132
rect 21542 9120 21548 9132
rect 21600 9120 21606 9172
rect 21726 9120 21732 9172
rect 21784 9120 21790 9172
rect 21082 9052 21088 9104
rect 21140 9092 21146 9104
rect 21744 9092 21772 9120
rect 21140 9064 21772 9092
rect 21140 9052 21146 9064
rect 21729 9027 21787 9033
rect 21729 9024 21741 9027
rect 21008 8996 21741 9024
rect 21729 8993 21741 8996
rect 21775 8993 21787 9027
rect 21729 8987 21787 8993
rect 19705 8959 19763 8965
rect 19705 8925 19717 8959
rect 19751 8956 19763 8959
rect 20901 8959 20959 8965
rect 19751 8928 20852 8956
rect 19751 8925 19763 8928
rect 19705 8919 19763 8925
rect 4764 8860 5672 8888
rect 5804 8891 5862 8897
rect 4764 8848 4770 8860
rect 5804 8857 5816 8891
rect 5850 8857 5862 8891
rect 5804 8851 5862 8857
rect 2774 8820 2780 8832
rect 2735 8792 2780 8820
rect 2774 8780 2780 8792
rect 2832 8780 2838 8832
rect 3237 8823 3295 8829
rect 3237 8789 3249 8823
rect 3283 8820 3295 8823
rect 3510 8820 3516 8832
rect 3283 8792 3516 8820
rect 3283 8789 3295 8792
rect 3237 8783 3295 8789
rect 3510 8780 3516 8792
rect 3568 8780 3574 8832
rect 4890 8820 4896 8832
rect 4851 8792 4896 8820
rect 4890 8780 4896 8792
rect 4948 8780 4954 8832
rect 4982 8780 4988 8832
rect 5040 8820 5046 8832
rect 5040 8792 5085 8820
rect 5040 8780 5046 8792
rect 5258 8780 5264 8832
rect 5316 8820 5322 8832
rect 5828 8820 5856 8851
rect 6638 8848 6644 8900
rect 6696 8888 6702 8900
rect 7622 8891 7680 8897
rect 7622 8888 7634 8891
rect 6696 8860 7634 8888
rect 6696 8848 6702 8860
rect 7622 8857 7634 8860
rect 7668 8857 7680 8891
rect 7622 8851 7680 8857
rect 8570 8848 8576 8900
rect 8628 8888 8634 8900
rect 9370 8891 9428 8897
rect 9370 8888 9382 8891
rect 8628 8860 9382 8888
rect 8628 8848 8634 8860
rect 9370 8857 9382 8860
rect 9416 8857 9428 8891
rect 9370 8851 9428 8857
rect 11054 8848 11060 8900
rect 11112 8888 11118 8900
rect 14642 8897 14648 8900
rect 11486 8891 11544 8897
rect 11486 8888 11498 8891
rect 11112 8860 11498 8888
rect 11112 8848 11118 8860
rect 11486 8857 11498 8860
rect 11532 8857 11544 8891
rect 11486 8851 11544 8857
rect 12636 8860 13676 8888
rect 5316 8792 5856 8820
rect 5316 8780 5322 8792
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 10502 8820 10508 8832
rect 6972 8792 7017 8820
rect 10463 8792 10508 8820
rect 6972 8780 6978 8792
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 12636 8829 12664 8860
rect 13648 8832 13676 8860
rect 14636 8851 14648 8897
rect 14700 8888 14706 8900
rect 14700 8860 14736 8888
rect 14642 8848 14648 8851
rect 14700 8848 14706 8860
rect 15286 8848 15292 8900
rect 15344 8888 15350 8900
rect 19429 8891 19487 8897
rect 19429 8888 19441 8891
rect 15344 8860 19441 8888
rect 15344 8848 15350 8860
rect 19429 8857 19441 8860
rect 19475 8857 19487 8891
rect 19429 8851 19487 8857
rect 19518 8848 19524 8900
rect 19576 8888 19582 8900
rect 19889 8891 19947 8897
rect 19889 8888 19901 8891
rect 19576 8860 19901 8888
rect 19576 8848 19582 8860
rect 19889 8857 19901 8860
rect 19935 8857 19947 8891
rect 19889 8851 19947 8857
rect 12621 8823 12679 8829
rect 12621 8789 12633 8823
rect 12667 8789 12679 8823
rect 12986 8820 12992 8832
rect 12947 8792 12992 8820
rect 12621 8783 12679 8789
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 13078 8780 13084 8832
rect 13136 8820 13142 8832
rect 13136 8792 13181 8820
rect 13136 8780 13142 8792
rect 13630 8780 13636 8832
rect 13688 8820 13694 8832
rect 15378 8820 15384 8832
rect 13688 8792 15384 8820
rect 13688 8780 13694 8792
rect 15378 8780 15384 8792
rect 15436 8780 15442 8832
rect 15746 8820 15752 8832
rect 15707 8792 15752 8820
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 15838 8780 15844 8832
rect 15896 8820 15902 8832
rect 16485 8823 16543 8829
rect 16485 8820 16497 8823
rect 15896 8792 16497 8820
rect 15896 8780 15902 8792
rect 16485 8789 16497 8792
rect 16531 8789 16543 8823
rect 20824 8820 20852 8928
rect 20901 8925 20913 8959
rect 20947 8925 20959 8959
rect 20901 8919 20959 8925
rect 21818 8848 21824 8900
rect 21876 8888 21882 8900
rect 21974 8891 22032 8897
rect 21974 8888 21986 8891
rect 21876 8860 21986 8888
rect 21876 8848 21882 8860
rect 21974 8857 21986 8860
rect 22020 8857 22032 8891
rect 21974 8851 22032 8857
rect 22554 8820 22560 8832
rect 20824 8792 22560 8820
rect 16485 8783 16543 8789
rect 22554 8780 22560 8792
rect 22612 8780 22618 8832
rect 23106 8820 23112 8832
rect 23067 8792 23112 8820
rect 23106 8780 23112 8792
rect 23164 8780 23170 8832
rect 1104 8730 23460 8752
rect 1104 8678 6548 8730
rect 6600 8678 6612 8730
rect 6664 8678 6676 8730
rect 6728 8678 6740 8730
rect 6792 8678 6804 8730
rect 6856 8678 12146 8730
rect 12198 8678 12210 8730
rect 12262 8678 12274 8730
rect 12326 8678 12338 8730
rect 12390 8678 12402 8730
rect 12454 8678 17744 8730
rect 17796 8678 17808 8730
rect 17860 8678 17872 8730
rect 17924 8678 17936 8730
rect 17988 8678 18000 8730
rect 18052 8678 23460 8730
rect 1104 8656 23460 8678
rect 3510 8616 3516 8628
rect 3471 8588 3516 8616
rect 3510 8576 3516 8588
rect 3568 8576 3574 8628
rect 3602 8576 3608 8628
rect 3660 8616 3666 8628
rect 3881 8619 3939 8625
rect 3881 8616 3893 8619
rect 3660 8588 3893 8616
rect 3660 8576 3666 8588
rect 3881 8585 3893 8588
rect 3927 8585 3939 8619
rect 4338 8616 4344 8628
rect 4299 8588 4344 8616
rect 3881 8579 3939 8585
rect 4338 8576 4344 8588
rect 4396 8576 4402 8628
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5353 8619 5411 8625
rect 5353 8616 5365 8619
rect 4948 8588 5365 8616
rect 4948 8576 4954 8588
rect 5353 8585 5365 8588
rect 5399 8585 5411 8619
rect 7006 8616 7012 8628
rect 6967 8588 7012 8616
rect 5353 8579 5411 8585
rect 7006 8576 7012 8588
rect 7064 8576 7070 8628
rect 9766 8616 9772 8628
rect 9727 8588 9772 8616
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 10134 8616 10140 8628
rect 10047 8588 10140 8616
rect 10134 8576 10140 8588
rect 10192 8616 10198 8628
rect 10502 8616 10508 8628
rect 10192 8588 10508 8616
rect 10192 8576 10198 8588
rect 10502 8576 10508 8588
rect 10560 8576 10566 8628
rect 10686 8616 10692 8628
rect 10647 8588 10692 8616
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 13262 8576 13268 8628
rect 13320 8616 13326 8628
rect 13357 8619 13415 8625
rect 13357 8616 13369 8619
rect 13320 8588 13369 8616
rect 13320 8576 13326 8588
rect 13357 8585 13369 8588
rect 13403 8616 13415 8619
rect 13403 8588 14320 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 2774 8508 2780 8560
rect 2832 8548 2838 8560
rect 3234 8548 3240 8560
rect 2832 8520 3240 8548
rect 2832 8508 2838 8520
rect 3234 8508 3240 8520
rect 3292 8548 3298 8560
rect 4801 8551 4859 8557
rect 4801 8548 4813 8551
rect 3292 8520 4813 8548
rect 3292 8508 3298 8520
rect 4801 8517 4813 8520
rect 4847 8517 4859 8551
rect 4801 8511 4859 8517
rect 7561 8551 7619 8557
rect 7561 8517 7573 8551
rect 7607 8548 7619 8551
rect 8542 8551 8600 8557
rect 8542 8548 8554 8551
rect 7607 8520 8554 8548
rect 7607 8517 7619 8520
rect 7561 8511 7619 8517
rect 8542 8517 8554 8520
rect 8588 8517 8600 8551
rect 8542 8511 8600 8517
rect 13716 8551 13774 8557
rect 13716 8517 13728 8551
rect 13762 8548 13774 8551
rect 13906 8548 13912 8560
rect 13762 8520 13912 8548
rect 13762 8517 13774 8520
rect 13716 8511 13774 8517
rect 13906 8508 13912 8520
rect 13964 8508 13970 8560
rect 14292 8548 14320 8588
rect 14366 8576 14372 8628
rect 14424 8616 14430 8628
rect 14921 8619 14979 8625
rect 14921 8616 14933 8619
rect 14424 8588 14933 8616
rect 14424 8576 14430 8588
rect 14921 8585 14933 8588
rect 14967 8585 14979 8619
rect 16209 8619 16267 8625
rect 16209 8616 16221 8619
rect 14921 8579 14979 8585
rect 15028 8588 16221 8616
rect 15028 8548 15056 8588
rect 16209 8585 16221 8588
rect 16255 8585 16267 8619
rect 16209 8579 16267 8585
rect 17126 8576 17132 8628
rect 17184 8616 17190 8628
rect 17313 8619 17371 8625
rect 17313 8616 17325 8619
rect 17184 8588 17325 8616
rect 17184 8576 17190 8588
rect 17313 8585 17325 8588
rect 17359 8585 17371 8619
rect 17313 8579 17371 8585
rect 18325 8619 18383 8625
rect 18325 8585 18337 8619
rect 18371 8616 18383 8619
rect 19334 8616 19340 8628
rect 18371 8588 19340 8616
rect 18371 8585 18383 8588
rect 18325 8579 18383 8585
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 20165 8619 20223 8625
rect 20165 8585 20177 8619
rect 20211 8616 20223 8619
rect 20254 8616 20260 8628
rect 20211 8588 20260 8616
rect 20211 8585 20223 8588
rect 20165 8579 20223 8585
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 20625 8619 20683 8625
rect 20625 8585 20637 8619
rect 20671 8616 20683 8619
rect 21174 8616 21180 8628
rect 20671 8588 21180 8616
rect 20671 8585 20683 8588
rect 20625 8579 20683 8585
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 14292 8520 15056 8548
rect 15289 8551 15347 8557
rect 15289 8517 15301 8551
rect 15335 8548 15347 8551
rect 15746 8548 15752 8560
rect 15335 8520 15752 8548
rect 15335 8517 15347 8520
rect 15289 8511 15347 8517
rect 15746 8508 15752 8520
rect 15804 8548 15810 8560
rect 18684 8551 18742 8557
rect 15804 8520 16712 8548
rect 15804 8508 15810 8520
rect 1762 8440 1768 8492
rect 1820 8480 1826 8492
rect 2314 8489 2320 8492
rect 2041 8483 2099 8489
rect 2041 8480 2053 8483
rect 1820 8452 2053 8480
rect 1820 8440 1826 8452
rect 2041 8449 2053 8452
rect 2087 8449 2099 8483
rect 2041 8443 2099 8449
rect 2308 8443 2320 8489
rect 2372 8480 2378 8492
rect 2372 8452 2408 8480
rect 2314 8440 2320 8443
rect 2372 8440 2378 8452
rect 2682 8440 2688 8492
rect 2740 8480 2746 8492
rect 4709 8483 4767 8489
rect 4709 8480 4721 8483
rect 2740 8452 3096 8480
rect 2740 8440 2746 8452
rect 3068 8412 3096 8452
rect 3896 8452 4721 8480
rect 3896 8412 3924 8452
rect 4709 8449 4721 8452
rect 4755 8449 4767 8483
rect 5718 8480 5724 8492
rect 5679 8452 5724 8480
rect 4709 8443 4767 8449
rect 5718 8440 5724 8452
rect 5776 8440 5782 8492
rect 6086 8440 6092 8492
rect 6144 8480 6150 8492
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 6144 8452 6377 8480
rect 6144 8440 6150 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 8202 8480 8208 8492
rect 8163 8452 8208 8480
rect 6365 8443 6423 8449
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 8297 8483 8355 8489
rect 8297 8449 8309 8483
rect 8343 8480 8355 8483
rect 8386 8480 8392 8492
rect 8343 8452 8392 8480
rect 8343 8449 8355 8452
rect 8297 8443 8355 8449
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 11330 8480 11336 8492
rect 11291 8452 11336 8480
rect 11330 8440 11336 8452
rect 11388 8440 11394 8492
rect 11974 8480 11980 8492
rect 11935 8452 11980 8480
rect 11974 8440 11980 8452
rect 12032 8440 12038 8492
rect 12066 8440 12072 8492
rect 12124 8480 12130 8492
rect 12233 8483 12291 8489
rect 12233 8480 12245 8483
rect 12124 8452 12245 8480
rect 12124 8440 12130 8452
rect 12233 8449 12245 8452
rect 12279 8449 12291 8483
rect 13446 8480 13452 8492
rect 13407 8452 13452 8480
rect 12233 8443 12291 8449
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 14550 8440 14556 8492
rect 14608 8480 14614 8492
rect 16114 8480 16120 8492
rect 14608 8452 15516 8480
rect 16075 8452 16120 8480
rect 14608 8440 14614 8452
rect 3068 8384 3924 8412
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8381 4031 8415
rect 3973 8375 4031 8381
rect 4157 8415 4215 8421
rect 4157 8381 4169 8415
rect 4203 8412 4215 8415
rect 4985 8415 5043 8421
rect 4985 8412 4997 8415
rect 4203 8384 4997 8412
rect 4203 8381 4215 8384
rect 4157 8375 4215 8381
rect 4985 8381 4997 8384
rect 5031 8381 5043 8415
rect 5810 8412 5816 8424
rect 5771 8384 5816 8412
rect 4985 8375 5043 8381
rect 3326 8304 3332 8356
rect 3384 8344 3390 8356
rect 3421 8347 3479 8353
rect 3421 8344 3433 8347
rect 3384 8316 3433 8344
rect 3384 8304 3390 8316
rect 3421 8313 3433 8316
rect 3467 8344 3479 8347
rect 3988 8344 4016 8375
rect 3467 8316 4016 8344
rect 5000 8344 5028 8375
rect 5810 8372 5816 8384
rect 5868 8372 5874 8424
rect 5997 8415 6055 8421
rect 5997 8381 6009 8415
rect 6043 8412 6055 8415
rect 6270 8412 6276 8424
rect 6043 8384 6276 8412
rect 6043 8381 6055 8384
rect 5997 8375 6055 8381
rect 5166 8344 5172 8356
rect 5000 8316 5172 8344
rect 3467 8313 3479 8316
rect 3421 8307 3479 8313
rect 5166 8304 5172 8316
rect 5224 8344 5230 8356
rect 6012 8344 6040 8375
rect 6270 8372 6276 8384
rect 6328 8372 6334 8424
rect 10229 8415 10287 8421
rect 10229 8381 10241 8415
rect 10275 8381 10287 8415
rect 10229 8375 10287 8381
rect 10413 8415 10471 8421
rect 10413 8381 10425 8415
rect 10459 8412 10471 8415
rect 10870 8412 10876 8424
rect 10459 8384 10876 8412
rect 10459 8381 10471 8384
rect 10413 8375 10471 8381
rect 9674 8344 9680 8356
rect 5224 8316 6040 8344
rect 9635 8316 9680 8344
rect 5224 8304 5230 8316
rect 9674 8304 9680 8316
rect 9732 8344 9738 8356
rect 10244 8344 10272 8375
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 15378 8412 15384 8424
rect 15339 8384 15384 8412
rect 15378 8372 15384 8384
rect 15436 8372 15442 8424
rect 15488 8421 15516 8452
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16684 8489 16712 8520
rect 18684 8517 18696 8551
rect 18730 8548 18742 8551
rect 22738 8548 22744 8560
rect 18730 8520 22744 8548
rect 18730 8517 18742 8520
rect 18684 8511 18742 8517
rect 22738 8508 22744 8520
rect 22796 8508 22802 8560
rect 16669 8483 16727 8489
rect 16669 8449 16681 8483
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 17405 8483 17463 8489
rect 17405 8449 17417 8483
rect 17451 8480 17463 8483
rect 17494 8480 17500 8492
rect 17451 8452 17500 8480
rect 17451 8449 17463 8452
rect 17405 8443 17463 8449
rect 17494 8440 17500 8452
rect 17552 8440 17558 8492
rect 18417 8483 18475 8489
rect 18417 8449 18429 8483
rect 18463 8480 18475 8483
rect 18966 8480 18972 8492
rect 18463 8452 18972 8480
rect 18463 8449 18475 8452
rect 18417 8443 18475 8449
rect 18966 8440 18972 8452
rect 19024 8440 19030 8492
rect 19058 8440 19064 8492
rect 19116 8480 19122 8492
rect 20257 8483 20315 8489
rect 20257 8480 20269 8483
rect 19116 8452 20269 8480
rect 19116 8440 19122 8452
rect 20257 8449 20269 8452
rect 20303 8449 20315 8483
rect 20257 8443 20315 8449
rect 21358 8440 21364 8492
rect 21416 8480 21422 8492
rect 21416 8452 21461 8480
rect 21416 8440 21422 8452
rect 21726 8440 21732 8492
rect 21784 8480 21790 8492
rect 21821 8483 21879 8489
rect 21821 8480 21833 8483
rect 21784 8452 21833 8480
rect 21784 8440 21790 8452
rect 21821 8449 21833 8452
rect 21867 8449 21879 8483
rect 22554 8480 22560 8492
rect 22515 8452 22560 8480
rect 21821 8443 21879 8449
rect 22554 8440 22560 8452
rect 22612 8440 22618 8492
rect 15473 8415 15531 8421
rect 15473 8381 15485 8415
rect 15519 8412 15531 8415
rect 16301 8415 16359 8421
rect 16301 8412 16313 8415
rect 15519 8384 16313 8412
rect 15519 8381 15531 8384
rect 15473 8375 15531 8381
rect 16301 8381 16313 8384
rect 16347 8381 16359 8415
rect 16301 8375 16359 8381
rect 20073 8415 20131 8421
rect 20073 8381 20085 8415
rect 20119 8412 20131 8415
rect 20438 8412 20444 8424
rect 20119 8384 20444 8412
rect 20119 8381 20131 8384
rect 20073 8375 20131 8381
rect 20438 8372 20444 8384
rect 20496 8372 20502 8424
rect 20717 8415 20775 8421
rect 20717 8381 20729 8415
rect 20763 8412 20775 8415
rect 20806 8412 20812 8424
rect 20763 8384 20812 8412
rect 20763 8381 20775 8384
rect 20717 8375 20775 8381
rect 20806 8372 20812 8384
rect 20864 8372 20870 8424
rect 20898 8372 20904 8424
rect 20956 8412 20962 8424
rect 21453 8415 21511 8421
rect 21453 8412 21465 8415
rect 20956 8384 21465 8412
rect 20956 8372 20962 8384
rect 21453 8381 21465 8384
rect 21499 8381 21511 8415
rect 21453 8375 21511 8381
rect 21542 8372 21548 8424
rect 21600 8412 21606 8424
rect 22465 8415 22523 8421
rect 22465 8412 22477 8415
rect 21600 8384 22477 8412
rect 21600 8372 21606 8384
rect 22465 8381 22477 8384
rect 22511 8381 22523 8415
rect 22465 8375 22523 8381
rect 22741 8415 22799 8421
rect 22741 8381 22753 8415
rect 22787 8381 22799 8415
rect 22741 8375 22799 8381
rect 9732 8316 10272 8344
rect 9732 8304 9738 8316
rect 10686 8304 10692 8356
rect 10744 8344 10750 8356
rect 11698 8344 11704 8356
rect 10744 8316 11704 8344
rect 10744 8304 10750 8316
rect 11698 8304 11704 8316
rect 11756 8304 11762 8356
rect 14458 8304 14464 8356
rect 14516 8344 14522 8356
rect 15749 8347 15807 8353
rect 15749 8344 15761 8347
rect 14516 8316 15761 8344
rect 14516 8304 14522 8316
rect 15749 8313 15761 8316
rect 15795 8313 15807 8347
rect 15749 8307 15807 8313
rect 17586 8304 17592 8356
rect 17644 8344 17650 8356
rect 18049 8347 18107 8353
rect 18049 8344 18061 8347
rect 17644 8316 18061 8344
rect 17644 8304 17650 8316
rect 18049 8313 18061 8316
rect 18095 8313 18107 8347
rect 18049 8307 18107 8313
rect 21174 8304 21180 8356
rect 21232 8344 21238 8356
rect 22756 8344 22784 8375
rect 21232 8316 22784 8344
rect 21232 8304 21238 8316
rect 14829 8279 14887 8285
rect 14829 8245 14841 8279
rect 14875 8276 14887 8279
rect 16114 8276 16120 8288
rect 14875 8248 16120 8276
rect 14875 8245 14887 8248
rect 14829 8239 14887 8245
rect 16114 8236 16120 8248
rect 16172 8236 16178 8288
rect 19797 8279 19855 8285
rect 19797 8245 19809 8279
rect 19843 8276 19855 8279
rect 20254 8276 20260 8288
rect 19843 8248 20260 8276
rect 19843 8245 19855 8248
rect 19797 8239 19855 8245
rect 20254 8236 20260 8248
rect 20312 8276 20318 8288
rect 21726 8276 21732 8288
rect 20312 8248 21732 8276
rect 20312 8236 20318 8248
rect 21726 8236 21732 8248
rect 21784 8236 21790 8288
rect 1104 8186 23460 8208
rect 1104 8134 3749 8186
rect 3801 8134 3813 8186
rect 3865 8134 3877 8186
rect 3929 8134 3941 8186
rect 3993 8134 4005 8186
rect 4057 8134 9347 8186
rect 9399 8134 9411 8186
rect 9463 8134 9475 8186
rect 9527 8134 9539 8186
rect 9591 8134 9603 8186
rect 9655 8134 14945 8186
rect 14997 8134 15009 8186
rect 15061 8134 15073 8186
rect 15125 8134 15137 8186
rect 15189 8134 15201 8186
rect 15253 8134 20543 8186
rect 20595 8134 20607 8186
rect 20659 8134 20671 8186
rect 20723 8134 20735 8186
rect 20787 8134 20799 8186
rect 20851 8134 23460 8186
rect 1104 8112 23460 8134
rect 4617 8075 4675 8081
rect 4617 8041 4629 8075
rect 4663 8072 4675 8075
rect 4982 8072 4988 8084
rect 4663 8044 4988 8072
rect 4663 8041 4675 8044
rect 4617 8035 4675 8041
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5445 8075 5503 8081
rect 5445 8041 5457 8075
rect 5491 8072 5503 8075
rect 5718 8072 5724 8084
rect 5491 8044 5724 8072
rect 5491 8041 5503 8044
rect 5445 8035 5503 8041
rect 3881 8007 3939 8013
rect 3881 7973 3893 8007
rect 3927 8004 3939 8007
rect 5258 8004 5264 8016
rect 3927 7976 5264 8004
rect 3927 7973 3939 7976
rect 3881 7967 3939 7973
rect 5258 7964 5264 7976
rect 5316 7964 5322 8016
rect 1762 7896 1768 7948
rect 1820 7936 1826 7948
rect 2225 7939 2283 7945
rect 2225 7936 2237 7939
rect 1820 7908 2237 7936
rect 1820 7896 1826 7908
rect 2225 7905 2237 7908
rect 2271 7905 2283 7939
rect 5166 7936 5172 7948
rect 5127 7908 5172 7936
rect 2225 7899 2283 7905
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 2130 7868 2136 7880
rect 2091 7840 2136 7868
rect 2130 7828 2136 7840
rect 2188 7828 2194 7880
rect 2498 7877 2504 7880
rect 2492 7868 2504 7877
rect 2459 7840 2504 7868
rect 2492 7831 2504 7840
rect 2498 7828 2504 7831
rect 2556 7828 2562 7880
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 5460 7868 5488 8035
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 7561 8075 7619 8081
rect 7561 8072 7573 8075
rect 7248 8044 7573 8072
rect 7248 8032 7254 8044
rect 7561 8041 7573 8044
rect 7607 8041 7619 8075
rect 7561 8035 7619 8041
rect 8113 8075 8171 8081
rect 8113 8041 8125 8075
rect 8159 8072 8171 8075
rect 8570 8072 8576 8084
rect 8159 8044 8576 8072
rect 8159 8041 8171 8044
rect 8113 8035 8171 8041
rect 8570 8032 8576 8044
rect 8628 8032 8634 8084
rect 9493 8075 9551 8081
rect 9493 8041 9505 8075
rect 9539 8072 9551 8075
rect 9858 8072 9864 8084
rect 9539 8044 9864 8072
rect 9539 8041 9551 8044
rect 9493 8035 9551 8041
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 13078 8032 13084 8084
rect 13136 8072 13142 8084
rect 13173 8075 13231 8081
rect 13173 8072 13185 8075
rect 13136 8044 13185 8072
rect 13136 8032 13142 8044
rect 13173 8041 13185 8044
rect 13219 8041 13231 8075
rect 13173 8035 13231 8041
rect 19150 8032 19156 8084
rect 19208 8072 19214 8084
rect 20898 8072 20904 8084
rect 19208 8044 20904 8072
rect 19208 8032 19214 8044
rect 20898 8032 20904 8044
rect 20956 8032 20962 8084
rect 21358 8072 21364 8084
rect 21319 8044 21364 8072
rect 21358 8032 21364 8044
rect 21416 8032 21422 8084
rect 22830 8032 22836 8084
rect 22888 8072 22894 8084
rect 22925 8075 22983 8081
rect 22925 8072 22937 8075
rect 22888 8044 22937 8072
rect 22888 8032 22894 8044
rect 22925 8041 22937 8044
rect 22971 8041 22983 8075
rect 22925 8035 22983 8041
rect 19061 8007 19119 8013
rect 19061 7973 19073 8007
rect 19107 8004 19119 8007
rect 19107 7976 19288 8004
rect 19107 7973 19119 7976
rect 19061 7967 19119 7973
rect 9950 7896 9956 7948
rect 10008 7936 10014 7948
rect 10229 7939 10287 7945
rect 10229 7936 10241 7939
rect 10008 7908 10241 7936
rect 10008 7896 10014 7908
rect 10229 7905 10241 7908
rect 10275 7905 10287 7939
rect 10229 7899 10287 7905
rect 13081 7939 13139 7945
rect 13081 7905 13093 7939
rect 13127 7936 13139 7939
rect 13446 7936 13452 7948
rect 13127 7908 13452 7936
rect 13127 7905 13139 7908
rect 13081 7899 13139 7905
rect 13446 7896 13452 7908
rect 13504 7896 13510 7948
rect 13630 7936 13636 7948
rect 13591 7908 13636 7936
rect 13630 7896 13636 7908
rect 13688 7896 13694 7948
rect 13725 7939 13783 7945
rect 13725 7905 13737 7939
rect 13771 7936 13783 7939
rect 13814 7936 13820 7948
rect 13771 7908 13820 7936
rect 13771 7905 13783 7908
rect 13725 7899 13783 7905
rect 13814 7896 13820 7908
rect 13872 7936 13878 7948
rect 14458 7936 14464 7948
rect 13872 7908 14464 7936
rect 13872 7896 13878 7908
rect 14458 7896 14464 7908
rect 14516 7896 14522 7948
rect 15473 7939 15531 7945
rect 15473 7905 15485 7939
rect 15519 7936 15531 7939
rect 15654 7936 15660 7948
rect 15519 7908 15660 7936
rect 15519 7905 15531 7908
rect 15473 7899 15531 7905
rect 15654 7896 15660 7908
rect 15712 7896 15718 7948
rect 18509 7939 18567 7945
rect 18509 7905 18521 7939
rect 18555 7936 18567 7939
rect 18598 7936 18604 7948
rect 18555 7908 18604 7936
rect 18555 7905 18567 7908
rect 18509 7899 18567 7905
rect 18598 7896 18604 7908
rect 18656 7896 18662 7948
rect 18966 7936 18972 7948
rect 18708 7908 18972 7936
rect 4571 7840 5488 7868
rect 6825 7871 6883 7877
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 6825 7837 6837 7871
rect 6871 7837 6883 7871
rect 6825 7831 6883 7837
rect 1489 7803 1547 7809
rect 1489 7769 1501 7803
rect 1535 7800 1547 7803
rect 4246 7800 4252 7812
rect 1535 7772 4252 7800
rect 1535 7769 1547 7772
rect 1489 7763 1547 7769
rect 4246 7760 4252 7772
rect 4304 7760 4310 7812
rect 6580 7803 6638 7809
rect 6580 7769 6592 7803
rect 6626 7800 6638 7803
rect 6840 7800 6868 7831
rect 6914 7828 6920 7880
rect 6972 7868 6978 7880
rect 8757 7871 8815 7877
rect 6972 7840 7017 7868
rect 6972 7828 6978 7840
rect 8757 7837 8769 7871
rect 8803 7868 8815 7871
rect 9674 7868 9680 7880
rect 8803 7840 9680 7868
rect 8803 7837 8815 7840
rect 8757 7831 8815 7837
rect 9674 7828 9680 7840
rect 9732 7828 9738 7880
rect 10134 7868 10140 7880
rect 10095 7840 10140 7868
rect 10134 7828 10140 7840
rect 10192 7828 10198 7880
rect 12825 7871 12883 7877
rect 12825 7837 12837 7871
rect 12871 7868 12883 7871
rect 15838 7868 15844 7880
rect 12871 7840 15844 7868
rect 12871 7837 12883 7840
rect 12825 7831 12883 7837
rect 15838 7828 15844 7840
rect 15896 7828 15902 7880
rect 16025 7871 16083 7877
rect 16025 7837 16037 7871
rect 16071 7868 16083 7871
rect 16071 7840 16436 7868
rect 16071 7837 16083 7840
rect 16025 7831 16083 7837
rect 16408 7812 16436 7840
rect 16758 7828 16764 7880
rect 16816 7868 16822 7880
rect 18708 7877 18736 7908
rect 18966 7896 18972 7908
rect 19024 7896 19030 7948
rect 19260 7936 19288 7976
rect 19708 7939 19766 7945
rect 19708 7936 19720 7939
rect 19260 7908 19720 7936
rect 19708 7905 19720 7908
rect 19754 7905 19766 7939
rect 19708 7899 19766 7905
rect 19981 7939 20039 7945
rect 19981 7905 19993 7939
rect 20027 7936 20039 7939
rect 20162 7936 20168 7948
rect 20027 7908 20168 7936
rect 20027 7905 20039 7908
rect 19981 7899 20039 7905
rect 20162 7896 20168 7908
rect 20220 7896 20226 7948
rect 17497 7871 17555 7877
rect 17497 7868 17509 7871
rect 16816 7840 17509 7868
rect 16816 7828 16822 7840
rect 17497 7837 17509 7840
rect 17543 7837 17555 7871
rect 17497 7831 17555 7837
rect 18693 7871 18751 7877
rect 18693 7837 18705 7871
rect 18739 7837 18751 7871
rect 18693 7831 18751 7837
rect 19235 7871 19293 7877
rect 19235 7837 19247 7871
rect 19281 7837 19293 7871
rect 19235 7831 19293 7837
rect 8018 7800 8024 7812
rect 6626 7772 6776 7800
rect 6840 7772 8024 7800
rect 6626 7769 6638 7772
rect 6580 7763 6638 7769
rect 3602 7732 3608 7744
rect 3563 7704 3608 7732
rect 3602 7692 3608 7704
rect 3660 7692 3666 7744
rect 4982 7732 4988 7744
rect 4943 7704 4988 7732
rect 4982 7692 4988 7704
rect 5040 7692 5046 7744
rect 5074 7692 5080 7744
rect 5132 7732 5138 7744
rect 6748 7732 6776 7772
rect 8018 7760 8024 7772
rect 8076 7760 8082 7812
rect 8570 7760 8576 7812
rect 8628 7800 8634 7812
rect 9309 7803 9367 7809
rect 9309 7800 9321 7803
rect 8628 7772 9321 7800
rect 8628 7760 8634 7772
rect 9309 7769 9321 7772
rect 9355 7769 9367 7803
rect 9309 7763 9367 7769
rect 10496 7803 10554 7809
rect 10496 7769 10508 7803
rect 10542 7800 10554 7803
rect 11974 7800 11980 7812
rect 10542 7772 11980 7800
rect 10542 7769 10554 7772
rect 10496 7763 10554 7769
rect 11974 7760 11980 7772
rect 12032 7760 12038 7812
rect 15194 7800 15200 7812
rect 15252 7809 15258 7812
rect 16298 7809 16304 7812
rect 15164 7772 15200 7800
rect 15194 7760 15200 7772
rect 15252 7763 15264 7809
rect 16292 7800 16304 7809
rect 16259 7772 16304 7800
rect 16292 7763 16304 7772
rect 15252 7760 15258 7763
rect 16298 7760 16304 7763
rect 16356 7760 16362 7812
rect 16390 7760 16396 7812
rect 16448 7760 16454 7812
rect 16666 7760 16672 7812
rect 16724 7800 16730 7812
rect 18141 7803 18199 7809
rect 18141 7800 18153 7803
rect 16724 7772 18153 7800
rect 16724 7760 16730 7772
rect 18141 7769 18153 7772
rect 18187 7769 18199 7803
rect 18141 7763 18199 7769
rect 19150 7760 19156 7812
rect 19208 7800 19214 7812
rect 19260 7800 19288 7831
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 21174 7868 21180 7880
rect 19392 7840 21036 7868
rect 21135 7840 21180 7868
rect 19392 7828 19398 7840
rect 19208 7772 19288 7800
rect 21008 7800 21036 7840
rect 21174 7828 21180 7840
rect 21232 7828 21238 7880
rect 21266 7828 21272 7880
rect 21324 7868 21330 7880
rect 21453 7871 21511 7877
rect 21453 7868 21465 7871
rect 21324 7840 21465 7868
rect 21324 7828 21330 7840
rect 21453 7837 21465 7840
rect 21499 7837 21511 7871
rect 21453 7831 21511 7837
rect 23109 7871 23167 7877
rect 23109 7837 23121 7871
rect 23155 7868 23167 7871
rect 23290 7868 23296 7880
rect 23155 7840 23296 7868
rect 23155 7837 23167 7840
rect 23109 7831 23167 7837
rect 23290 7828 23296 7840
rect 23348 7828 23354 7880
rect 21358 7800 21364 7812
rect 21008 7772 21364 7800
rect 19208 7760 19214 7772
rect 21358 7760 21364 7772
rect 21416 7760 21422 7812
rect 21720 7803 21778 7809
rect 21720 7769 21732 7803
rect 21766 7800 21778 7803
rect 22278 7800 22284 7812
rect 21766 7772 22284 7800
rect 21766 7769 21778 7772
rect 21720 7763 21778 7769
rect 22278 7760 22284 7772
rect 22336 7760 22342 7812
rect 7006 7732 7012 7744
rect 5132 7704 5177 7732
rect 6748 7704 7012 7732
rect 5132 7692 5138 7704
rect 7006 7692 7012 7704
rect 7064 7692 7070 7744
rect 9214 7732 9220 7744
rect 9175 7704 9220 7732
rect 9214 7692 9220 7704
rect 9272 7692 9278 7744
rect 11330 7692 11336 7744
rect 11388 7732 11394 7744
rect 11609 7735 11667 7741
rect 11609 7732 11621 7735
rect 11388 7704 11621 7732
rect 11388 7692 11394 7704
rect 11609 7701 11621 7704
rect 11655 7701 11667 7735
rect 11609 7695 11667 7701
rect 11701 7735 11759 7741
rect 11701 7701 11713 7735
rect 11747 7732 11759 7735
rect 12710 7732 12716 7744
rect 11747 7704 12716 7732
rect 11747 7701 11759 7704
rect 11701 7695 11759 7701
rect 12710 7692 12716 7704
rect 12768 7732 12774 7744
rect 13541 7735 13599 7741
rect 13541 7732 13553 7735
rect 12768 7704 13553 7732
rect 12768 7692 12774 7704
rect 13541 7701 13553 7704
rect 13587 7701 13599 7735
rect 13541 7695 13599 7701
rect 14093 7735 14151 7741
rect 14093 7701 14105 7735
rect 14139 7732 14151 7735
rect 15378 7732 15384 7744
rect 14139 7704 15384 7732
rect 14139 7701 14151 7704
rect 14093 7695 14151 7701
rect 15378 7692 15384 7704
rect 15436 7692 15442 7744
rect 17405 7735 17463 7741
rect 17405 7701 17417 7735
rect 17451 7732 17463 7735
rect 17494 7732 17500 7744
rect 17451 7704 17500 7732
rect 17451 7701 17463 7704
rect 17405 7695 17463 7701
rect 17494 7692 17500 7704
rect 17552 7692 17558 7744
rect 18601 7735 18659 7741
rect 18601 7701 18613 7735
rect 18647 7732 18659 7735
rect 18966 7732 18972 7744
rect 18647 7704 18972 7732
rect 18647 7701 18659 7704
rect 18601 7695 18659 7701
rect 18966 7692 18972 7704
rect 19024 7692 19030 7744
rect 19711 7735 19769 7741
rect 19711 7701 19723 7735
rect 19757 7732 19769 7735
rect 19978 7732 19984 7744
rect 19757 7704 19984 7732
rect 19757 7701 19769 7704
rect 19711 7695 19769 7701
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 20806 7692 20812 7744
rect 20864 7732 20870 7744
rect 21085 7735 21143 7741
rect 21085 7732 21097 7735
rect 20864 7704 21097 7732
rect 20864 7692 20870 7704
rect 21085 7701 21097 7704
rect 21131 7701 21143 7735
rect 21085 7695 21143 7701
rect 22738 7692 22744 7744
rect 22796 7732 22802 7744
rect 22833 7735 22891 7741
rect 22833 7732 22845 7735
rect 22796 7704 22845 7732
rect 22796 7692 22802 7704
rect 22833 7701 22845 7704
rect 22879 7701 22891 7735
rect 22833 7695 22891 7701
rect 1104 7642 23460 7664
rect 1104 7590 6548 7642
rect 6600 7590 6612 7642
rect 6664 7590 6676 7642
rect 6728 7590 6740 7642
rect 6792 7590 6804 7642
rect 6856 7590 12146 7642
rect 12198 7590 12210 7642
rect 12262 7590 12274 7642
rect 12326 7590 12338 7642
rect 12390 7590 12402 7642
rect 12454 7590 17744 7642
rect 17796 7590 17808 7642
rect 17860 7590 17872 7642
rect 17924 7590 17936 7642
rect 17988 7590 18000 7642
rect 18052 7590 23460 7642
rect 1104 7568 23460 7590
rect 1397 7531 1455 7537
rect 1397 7497 1409 7531
rect 1443 7528 1455 7531
rect 1578 7528 1584 7540
rect 1443 7500 1584 7528
rect 1443 7497 1455 7500
rect 1397 7491 1455 7497
rect 1578 7488 1584 7500
rect 1636 7488 1642 7540
rect 2130 7488 2136 7540
rect 2188 7528 2194 7540
rect 3237 7531 3295 7537
rect 3237 7528 3249 7531
rect 2188 7500 3249 7528
rect 2188 7488 2194 7500
rect 3237 7497 3249 7500
rect 3283 7528 3295 7531
rect 5074 7528 5080 7540
rect 3283 7500 5080 7528
rect 3283 7497 3295 7500
rect 3237 7491 3295 7497
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 5534 7488 5540 7540
rect 5592 7528 5598 7540
rect 6457 7531 6515 7537
rect 6457 7528 6469 7531
rect 5592 7500 6469 7528
rect 5592 7488 5598 7500
rect 6457 7497 6469 7500
rect 6503 7528 6515 7531
rect 11514 7528 11520 7540
rect 6503 7500 11520 7528
rect 6503 7497 6515 7500
rect 6457 7491 6515 7497
rect 1670 7460 1676 7472
rect 1583 7432 1676 7460
rect 1596 7401 1624 7432
rect 1670 7420 1676 7432
rect 1728 7460 1734 7472
rect 1728 7432 6776 7460
rect 1728 7420 1734 7432
rect 1581 7395 1639 7401
rect 1581 7361 1593 7395
rect 1627 7361 1639 7395
rect 2774 7392 2780 7404
rect 2832 7401 2838 7404
rect 2744 7364 2780 7392
rect 1581 7355 1639 7361
rect 2774 7352 2780 7364
rect 2832 7355 2844 7401
rect 4338 7392 4344 7404
rect 4396 7401 4402 7404
rect 4308 7364 4344 7392
rect 2832 7352 2838 7355
rect 4338 7352 4344 7364
rect 4396 7355 4408 7401
rect 4396 7352 4402 7355
rect 4522 7352 4528 7404
rect 4580 7392 4586 7404
rect 6748 7401 6776 7432
rect 8018 7420 8024 7472
rect 8076 7460 8082 7472
rect 8076 7432 9352 7460
rect 8076 7420 8082 7432
rect 5057 7395 5115 7401
rect 5057 7392 5069 7395
rect 4580 7364 5069 7392
rect 4580 7352 4586 7364
rect 5057 7361 5069 7364
rect 5103 7361 5115 7395
rect 5057 7355 5115 7361
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 9030 7392 9036 7404
rect 9088 7401 9094 7404
rect 9324 7401 9352 7432
rect 9416 7401 9444 7500
rect 11514 7488 11520 7500
rect 11572 7488 11578 7540
rect 11793 7531 11851 7537
rect 11793 7497 11805 7531
rect 11839 7528 11851 7531
rect 11882 7528 11888 7540
rect 11839 7500 11888 7528
rect 11839 7497 11851 7500
rect 11793 7491 11851 7497
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 12621 7531 12679 7537
rect 12621 7497 12633 7531
rect 12667 7528 12679 7531
rect 12986 7528 12992 7540
rect 12667 7500 12992 7528
rect 12667 7497 12679 7500
rect 12621 7491 12679 7497
rect 12986 7488 12992 7500
rect 13044 7488 13050 7540
rect 14553 7531 14611 7537
rect 14553 7497 14565 7531
rect 14599 7528 14611 7531
rect 14642 7528 14648 7540
rect 14599 7500 14648 7528
rect 14599 7497 14611 7500
rect 14553 7491 14611 7497
rect 14642 7488 14648 7500
rect 14700 7488 14706 7540
rect 15194 7488 15200 7540
rect 15252 7528 15258 7540
rect 15289 7531 15347 7537
rect 15289 7528 15301 7531
rect 15252 7500 15301 7528
rect 15252 7488 15258 7500
rect 15289 7497 15301 7500
rect 15335 7497 15347 7531
rect 15289 7491 15347 7497
rect 16117 7531 16175 7537
rect 16117 7497 16129 7531
rect 16163 7528 16175 7531
rect 19334 7528 19340 7540
rect 16163 7500 19340 7528
rect 16163 7497 16175 7500
rect 16117 7491 16175 7497
rect 10689 7463 10747 7469
rect 10689 7429 10701 7463
rect 10735 7460 10747 7463
rect 11054 7460 11060 7472
rect 10735 7432 11060 7460
rect 10735 7429 10747 7432
rect 10689 7423 10747 7429
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 14461 7463 14519 7469
rect 14461 7429 14473 7463
rect 14507 7460 14519 7463
rect 16132 7460 16160 7491
rect 19334 7488 19340 7500
rect 19392 7488 19398 7540
rect 19705 7531 19763 7537
rect 19705 7528 19717 7531
rect 19444 7500 19717 7528
rect 14507 7432 16160 7460
rect 14507 7429 14519 7432
rect 14461 7423 14519 7429
rect 17586 7420 17592 7472
rect 17644 7460 17650 7472
rect 17782 7463 17840 7469
rect 17782 7460 17794 7463
rect 17644 7432 17794 7460
rect 17644 7420 17650 7432
rect 17782 7429 17794 7432
rect 17828 7429 17840 7463
rect 17782 7423 17840 7429
rect 18966 7420 18972 7472
rect 19024 7460 19030 7472
rect 19444 7460 19472 7500
rect 19705 7497 19717 7500
rect 19751 7497 19763 7531
rect 19705 7491 19763 7497
rect 20073 7531 20131 7537
rect 20073 7497 20085 7531
rect 20119 7528 20131 7531
rect 20162 7528 20168 7540
rect 20119 7500 20168 7528
rect 20119 7497 20131 7500
rect 20073 7491 20131 7497
rect 20162 7488 20168 7500
rect 20220 7488 20226 7540
rect 20806 7528 20812 7540
rect 20767 7500 20812 7528
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 21358 7488 21364 7540
rect 21416 7528 21422 7540
rect 21913 7531 21971 7537
rect 21913 7528 21925 7531
rect 21416 7500 21925 7528
rect 21416 7488 21422 7500
rect 21913 7497 21925 7500
rect 21959 7528 21971 7531
rect 22186 7528 22192 7540
rect 21959 7500 22192 7528
rect 21959 7497 21971 7500
rect 21913 7491 21971 7497
rect 22186 7488 22192 7500
rect 22244 7488 22250 7540
rect 21542 7460 21548 7472
rect 19024 7432 19472 7460
rect 19996 7432 21548 7460
rect 19024 7420 19030 7432
rect 6779 7364 6914 7392
rect 9000 7364 9036 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 3050 7324 3056 7336
rect 3011 7296 3056 7324
rect 3050 7284 3056 7296
rect 3108 7284 3114 7336
rect 4614 7324 4620 7336
rect 4575 7296 4620 7324
rect 4614 7284 4620 7296
rect 4672 7324 4678 7336
rect 4801 7327 4859 7333
rect 4801 7324 4813 7327
rect 4672 7296 4813 7324
rect 4672 7284 4678 7296
rect 4801 7293 4813 7296
rect 4847 7293 4859 7327
rect 4801 7287 4859 7293
rect 5810 7216 5816 7268
rect 5868 7256 5874 7268
rect 6181 7259 6239 7265
rect 6181 7256 6193 7259
rect 5868 7228 6193 7256
rect 5868 7216 5874 7228
rect 6181 7225 6193 7228
rect 6227 7256 6239 7259
rect 6362 7256 6368 7268
rect 6227 7228 6368 7256
rect 6227 7225 6239 7228
rect 6181 7219 6239 7225
rect 6362 7216 6368 7228
rect 6420 7216 6426 7268
rect 1673 7191 1731 7197
rect 1673 7157 1685 7191
rect 1719 7188 1731 7191
rect 1762 7188 1768 7200
rect 1719 7160 1768 7188
rect 1719 7157 1731 7160
rect 1673 7151 1731 7157
rect 1762 7148 1768 7160
rect 1820 7188 1826 7200
rect 2682 7188 2688 7200
rect 1820 7160 2688 7188
rect 1820 7148 1826 7160
rect 2682 7148 2688 7160
rect 2740 7148 2746 7200
rect 6886 7188 6914 7364
rect 9030 7352 9036 7364
rect 9088 7355 9100 7401
rect 9309 7395 9367 7401
rect 9309 7361 9321 7395
rect 9355 7361 9367 7395
rect 9309 7355 9367 7361
rect 9401 7395 9459 7401
rect 9401 7361 9413 7395
rect 9447 7361 9459 7395
rect 10594 7392 10600 7404
rect 10555 7364 10600 7392
rect 9401 7355 9459 7361
rect 9088 7352 9094 7355
rect 7285 7327 7343 7333
rect 7285 7293 7297 7327
rect 7331 7324 7343 7327
rect 7374 7324 7380 7336
rect 7331 7296 7380 7324
rect 7331 7293 7343 7296
rect 7285 7287 7343 7293
rect 7374 7284 7380 7296
rect 7432 7324 7438 7336
rect 7834 7324 7840 7336
rect 7432 7296 7840 7324
rect 7432 7284 7438 7296
rect 7834 7284 7840 7296
rect 7892 7284 7898 7336
rect 9324 7324 9352 7355
rect 10594 7352 10600 7364
rect 10652 7352 10658 7404
rect 11330 7392 11336 7404
rect 11291 7364 11336 7392
rect 11330 7352 11336 7364
rect 11388 7392 11394 7404
rect 12253 7395 12311 7401
rect 12253 7392 12265 7395
rect 11388 7364 12265 7392
rect 11388 7352 11394 7364
rect 12253 7361 12265 7364
rect 12299 7361 12311 7395
rect 12253 7355 12311 7361
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7392 15255 7395
rect 15378 7392 15384 7404
rect 15243 7364 15384 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 15378 7352 15384 7364
rect 15436 7352 15442 7404
rect 15933 7395 15991 7401
rect 15933 7361 15945 7395
rect 15979 7392 15991 7395
rect 16114 7392 16120 7404
rect 15979 7364 16120 7392
rect 15979 7361 15991 7364
rect 15933 7355 15991 7361
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 19357 7395 19415 7401
rect 19357 7361 19369 7395
rect 19403 7392 19415 7395
rect 19624 7395 19682 7401
rect 19403 7364 19564 7392
rect 19403 7361 19415 7364
rect 19357 7355 19415 7361
rect 9950 7324 9956 7336
rect 9324 7296 9956 7324
rect 9950 7284 9956 7296
rect 10008 7324 10014 7336
rect 10137 7327 10195 7333
rect 10137 7324 10149 7327
rect 10008 7296 10149 7324
rect 10008 7284 10014 7296
rect 10137 7293 10149 7296
rect 10183 7293 10195 7327
rect 10137 7287 10195 7293
rect 11977 7327 12035 7333
rect 11977 7293 11989 7327
rect 12023 7293 12035 7327
rect 12158 7324 12164 7336
rect 12119 7296 12164 7324
rect 11977 7287 12035 7293
rect 11992 7256 12020 7287
rect 12158 7284 12164 7296
rect 12216 7284 12222 7336
rect 12802 7284 12808 7336
rect 12860 7324 12866 7336
rect 16850 7324 16856 7336
rect 12860 7296 16856 7324
rect 12860 7284 12866 7296
rect 16850 7284 16856 7296
rect 16908 7284 16914 7336
rect 18049 7327 18107 7333
rect 18049 7293 18061 7327
rect 18095 7324 18107 7327
rect 18230 7324 18236 7336
rect 18095 7296 18236 7324
rect 18095 7293 18107 7296
rect 18049 7287 18107 7293
rect 18230 7284 18236 7296
rect 18288 7284 18294 7336
rect 19536 7324 19564 7364
rect 19624 7361 19636 7395
rect 19670 7392 19682 7395
rect 19794 7392 19800 7404
rect 19670 7364 19800 7392
rect 19670 7361 19682 7364
rect 19624 7355 19682 7361
rect 19794 7352 19800 7364
rect 19852 7352 19858 7404
rect 19996 7324 20024 7432
rect 21542 7420 21548 7432
rect 21600 7420 21606 7472
rect 22281 7463 22339 7469
rect 22281 7429 22293 7463
rect 22327 7460 22339 7463
rect 22922 7460 22928 7472
rect 22327 7432 22928 7460
rect 22327 7429 22339 7432
rect 22281 7423 22339 7429
rect 22922 7420 22928 7432
rect 22980 7420 22986 7472
rect 20901 7395 20959 7401
rect 20901 7392 20913 7395
rect 20180 7364 20913 7392
rect 20180 7336 20208 7364
rect 20901 7361 20913 7364
rect 20947 7361 20959 7395
rect 20901 7355 20959 7361
rect 21453 7395 21511 7401
rect 21453 7361 21465 7395
rect 21499 7392 21511 7395
rect 22186 7392 22192 7404
rect 21499 7364 22192 7392
rect 21499 7361 21511 7364
rect 21453 7355 21511 7361
rect 22186 7352 22192 7364
rect 22244 7352 22250 7404
rect 23014 7392 23020 7404
rect 22975 7364 23020 7392
rect 23014 7352 23020 7364
rect 23072 7352 23078 7404
rect 20162 7324 20168 7336
rect 19536 7296 20024 7324
rect 20123 7296 20168 7324
rect 20162 7284 20168 7296
rect 20220 7284 20226 7336
rect 20346 7324 20352 7336
rect 20307 7296 20352 7324
rect 20346 7284 20352 7296
rect 20404 7284 20410 7336
rect 20717 7327 20775 7333
rect 20717 7293 20729 7327
rect 20763 7293 20775 7327
rect 22370 7324 22376 7336
rect 22331 7296 22376 7324
rect 20717 7287 20775 7293
rect 13814 7256 13820 7268
rect 11992 7228 13820 7256
rect 13814 7216 13820 7228
rect 13872 7216 13878 7268
rect 16206 7256 16212 7268
rect 16167 7228 16212 7256
rect 16206 7216 16212 7228
rect 16264 7216 16270 7268
rect 16669 7259 16727 7265
rect 16669 7225 16681 7259
rect 16715 7256 16727 7259
rect 16758 7256 16764 7268
rect 16715 7228 16764 7256
rect 16715 7225 16727 7228
rect 16669 7219 16727 7225
rect 16758 7216 16764 7228
rect 16816 7216 16822 7268
rect 18156 7228 18736 7256
rect 7558 7188 7564 7200
rect 6886 7160 7564 7188
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 7929 7191 7987 7197
rect 7929 7157 7941 7191
rect 7975 7188 7987 7191
rect 8110 7188 8116 7200
rect 7975 7160 8116 7188
rect 7975 7157 7987 7160
rect 7929 7151 7987 7157
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 8570 7148 8576 7200
rect 8628 7188 8634 7200
rect 10413 7191 10471 7197
rect 10413 7188 10425 7191
rect 8628 7160 10425 7188
rect 8628 7148 8634 7160
rect 10413 7157 10425 7160
rect 10459 7157 10471 7191
rect 12986 7188 12992 7200
rect 12947 7160 12992 7188
rect 10413 7151 10471 7157
rect 12986 7148 12992 7160
rect 13044 7148 13050 7200
rect 16485 7191 16543 7197
rect 16485 7157 16497 7191
rect 16531 7188 16543 7191
rect 18156 7188 18184 7228
rect 16531 7160 18184 7188
rect 18233 7191 18291 7197
rect 16531 7157 16543 7160
rect 16485 7151 16543 7157
rect 18233 7157 18245 7191
rect 18279 7188 18291 7191
rect 18598 7188 18604 7200
rect 18279 7160 18604 7188
rect 18279 7157 18291 7160
rect 18233 7151 18291 7157
rect 18598 7148 18604 7160
rect 18656 7148 18662 7200
rect 18708 7188 18736 7228
rect 19610 7216 19616 7268
rect 19668 7256 19674 7268
rect 19794 7256 19800 7268
rect 19668 7228 19800 7256
rect 19668 7216 19674 7228
rect 19794 7216 19800 7228
rect 19852 7216 19858 7268
rect 20254 7216 20260 7268
rect 20312 7256 20318 7268
rect 20732 7256 20760 7287
rect 22370 7284 22376 7296
rect 22428 7284 22434 7336
rect 22557 7327 22615 7333
rect 22557 7293 22569 7327
rect 22603 7324 22615 7327
rect 22738 7324 22744 7336
rect 22603 7296 22744 7324
rect 22603 7293 22615 7296
rect 22557 7287 22615 7293
rect 22738 7284 22744 7296
rect 22796 7284 22802 7336
rect 20312 7228 20760 7256
rect 21637 7259 21695 7265
rect 20312 7216 20318 7228
rect 21637 7225 21649 7259
rect 21683 7256 21695 7259
rect 21683 7228 22048 7256
rect 21683 7225 21695 7228
rect 21637 7219 21695 7225
rect 19334 7188 19340 7200
rect 18708 7160 19340 7188
rect 19334 7148 19340 7160
rect 19392 7148 19398 7200
rect 21269 7191 21327 7197
rect 21269 7157 21281 7191
rect 21315 7188 21327 7191
rect 21726 7188 21732 7200
rect 21315 7160 21732 7188
rect 21315 7157 21327 7160
rect 21269 7151 21327 7157
rect 21726 7148 21732 7160
rect 21784 7148 21790 7200
rect 22020 7188 22048 7228
rect 22094 7216 22100 7268
rect 22152 7256 22158 7268
rect 22833 7259 22891 7265
rect 22833 7256 22845 7259
rect 22152 7228 22845 7256
rect 22152 7216 22158 7228
rect 22833 7225 22845 7228
rect 22879 7225 22891 7259
rect 22833 7219 22891 7225
rect 22738 7188 22744 7200
rect 22020 7160 22744 7188
rect 22738 7148 22744 7160
rect 22796 7148 22802 7200
rect 1104 7098 23460 7120
rect 1104 7046 3749 7098
rect 3801 7046 3813 7098
rect 3865 7046 3877 7098
rect 3929 7046 3941 7098
rect 3993 7046 4005 7098
rect 4057 7046 9347 7098
rect 9399 7046 9411 7098
rect 9463 7046 9475 7098
rect 9527 7046 9539 7098
rect 9591 7046 9603 7098
rect 9655 7046 14945 7098
rect 14997 7046 15009 7098
rect 15061 7046 15073 7098
rect 15125 7046 15137 7098
rect 15189 7046 15201 7098
rect 15253 7046 20543 7098
rect 20595 7046 20607 7098
rect 20659 7046 20671 7098
rect 20723 7046 20735 7098
rect 20787 7046 20799 7098
rect 20851 7046 23460 7098
rect 1104 7024 23460 7046
rect 1670 6984 1676 6996
rect 1631 6956 1676 6984
rect 1670 6944 1676 6956
rect 1728 6944 1734 6996
rect 4614 6984 4620 6996
rect 3988 6956 4620 6984
rect 1854 6848 1860 6860
rect 1815 6820 1860 6848
rect 1854 6808 1860 6820
rect 1912 6808 1918 6860
rect 3050 6808 3056 6860
rect 3108 6848 3114 6860
rect 3988 6857 4016 6956
rect 4614 6944 4620 6956
rect 4672 6984 4678 6996
rect 5442 6984 5448 6996
rect 4672 6956 5448 6984
rect 4672 6944 4678 6956
rect 5442 6944 5448 6956
rect 5500 6984 5506 6996
rect 5500 6956 6224 6984
rect 5500 6944 5506 6956
rect 6196 6860 6224 6956
rect 7558 6944 7564 6996
rect 7616 6984 7622 6996
rect 12158 6984 12164 6996
rect 7616 6956 11744 6984
rect 12119 6956 12164 6984
rect 7616 6944 7622 6956
rect 11716 6916 11744 6956
rect 12158 6944 12164 6956
rect 12216 6944 12222 6996
rect 17957 6987 18015 6993
rect 17957 6984 17969 6987
rect 12268 6956 17969 6984
rect 12268 6916 12296 6956
rect 17957 6953 17969 6956
rect 18003 6953 18015 6987
rect 17957 6947 18015 6953
rect 19061 6987 19119 6993
rect 19061 6953 19073 6987
rect 19107 6984 19119 6987
rect 20162 6984 20168 6996
rect 19107 6956 20168 6984
rect 19107 6953 19119 6956
rect 19061 6947 19119 6953
rect 11716 6888 12296 6916
rect 17972 6916 18000 6947
rect 20162 6944 20168 6956
rect 20220 6944 20226 6996
rect 22094 6984 22100 6996
rect 20824 6956 22100 6984
rect 20824 6928 20852 6956
rect 22094 6944 22100 6956
rect 22152 6944 22158 6996
rect 22186 6944 22192 6996
rect 22244 6984 22250 6996
rect 22557 6987 22615 6993
rect 22557 6984 22569 6987
rect 22244 6956 22569 6984
rect 22244 6944 22250 6956
rect 22557 6953 22569 6956
rect 22603 6953 22615 6987
rect 22557 6947 22615 6953
rect 17972 6888 18552 6916
rect 3973 6851 4031 6857
rect 3973 6848 3985 6851
rect 3108 6820 3985 6848
rect 3108 6808 3114 6820
rect 3973 6817 3985 6820
rect 4019 6817 4031 6851
rect 6178 6848 6184 6860
rect 6091 6820 6184 6848
rect 3973 6811 4031 6817
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 7285 6851 7343 6857
rect 7285 6817 7297 6851
rect 7331 6848 7343 6851
rect 8294 6848 8300 6860
rect 7331 6820 8300 6848
rect 7331 6817 7343 6820
rect 7285 6811 7343 6817
rect 8294 6808 8300 6820
rect 8352 6808 8358 6860
rect 8570 6848 8576 6860
rect 8531 6820 8576 6848
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 12066 6808 12072 6860
rect 12124 6848 12130 6860
rect 12253 6851 12311 6857
rect 12253 6848 12265 6851
rect 12124 6820 12265 6848
rect 12124 6808 12130 6820
rect 12253 6817 12265 6820
rect 12299 6817 12311 6851
rect 14737 6851 14795 6857
rect 14737 6848 14749 6851
rect 12253 6811 12311 6817
rect 12360 6820 13032 6848
rect 2501 6783 2559 6789
rect 2501 6749 2513 6783
rect 2547 6780 2559 6783
rect 2590 6780 2596 6792
rect 2547 6752 2596 6780
rect 2547 6749 2559 6752
rect 2501 6743 2559 6749
rect 2590 6740 2596 6752
rect 2648 6740 2654 6792
rect 4246 6789 4252 6792
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6780 3663 6783
rect 3651 6752 4108 6780
rect 3651 6749 3663 6752
rect 3605 6743 3663 6749
rect 2958 6712 2964 6724
rect 2919 6684 2964 6712
rect 2958 6672 2964 6684
rect 3016 6672 3022 6724
rect 4080 6644 4108 6752
rect 4240 6743 4252 6789
rect 4304 6780 4310 6792
rect 5445 6783 5503 6789
rect 4304 6752 4340 6780
rect 4246 6740 4252 6743
rect 4304 6740 4310 6752
rect 5445 6749 5457 6783
rect 5491 6780 5503 6783
rect 5534 6780 5540 6792
rect 5491 6752 5540 6780
rect 5491 6749 5503 6752
rect 5445 6743 5503 6749
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6749 7251 6783
rect 7193 6743 7251 6749
rect 7929 6783 7987 6789
rect 7929 6749 7941 6783
rect 7975 6780 7987 6783
rect 8662 6780 8668 6792
rect 7975 6752 8668 6780
rect 7975 6749 7987 6752
rect 7929 6743 7987 6749
rect 7208 6712 7236 6743
rect 8662 6740 8668 6752
rect 8720 6780 8726 6792
rect 10321 6783 10379 6789
rect 10321 6780 10333 6783
rect 8720 6752 8984 6780
rect 8720 6740 8726 6752
rect 8110 6712 8116 6724
rect 7208 6684 8116 6712
rect 8110 6672 8116 6684
rect 8168 6712 8174 6724
rect 8481 6715 8539 6721
rect 8481 6712 8493 6715
rect 8168 6684 8493 6712
rect 8168 6672 8174 6684
rect 8481 6681 8493 6684
rect 8527 6681 8539 6715
rect 8481 6675 8539 6681
rect 4982 6644 4988 6656
rect 4080 6616 4988 6644
rect 4982 6604 4988 6616
rect 5040 6644 5046 6656
rect 5353 6647 5411 6653
rect 5353 6644 5365 6647
rect 5040 6616 5365 6644
rect 5040 6604 5046 6616
rect 5353 6613 5365 6616
rect 5399 6613 5411 6647
rect 5353 6607 5411 6613
rect 6549 6647 6607 6653
rect 6549 6613 6561 6647
rect 6595 6644 6607 6647
rect 7190 6644 7196 6656
rect 6595 6616 7196 6644
rect 6595 6613 6607 6616
rect 6549 6607 6607 6613
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 8021 6647 8079 6653
rect 8021 6644 8033 6647
rect 7524 6616 8033 6644
rect 7524 6604 7530 6616
rect 8021 6613 8033 6616
rect 8067 6613 8079 6647
rect 8021 6607 8079 6613
rect 8389 6647 8447 6653
rect 8389 6613 8401 6647
rect 8435 6644 8447 6647
rect 8570 6644 8576 6656
rect 8435 6616 8576 6644
rect 8435 6613 8447 6616
rect 8389 6607 8447 6613
rect 8570 6604 8576 6616
rect 8628 6604 8634 6656
rect 8956 6653 8984 6752
rect 9968 6752 10333 6780
rect 9968 6724 9996 6752
rect 10321 6749 10333 6752
rect 10367 6780 10379 6783
rect 10781 6783 10839 6789
rect 10781 6780 10793 6783
rect 10367 6752 10793 6780
rect 10367 6749 10379 6752
rect 10321 6743 10379 6749
rect 10781 6749 10793 6752
rect 10827 6749 10839 6783
rect 11882 6780 11888 6792
rect 10781 6743 10839 6749
rect 10980 6752 11888 6780
rect 9950 6672 9956 6724
rect 10008 6672 10014 6724
rect 10076 6715 10134 6721
rect 10076 6681 10088 6715
rect 10122 6712 10134 6715
rect 10410 6712 10416 6724
rect 10122 6684 10416 6712
rect 10122 6681 10134 6684
rect 10076 6675 10134 6681
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 10597 6715 10655 6721
rect 10597 6681 10609 6715
rect 10643 6712 10655 6715
rect 10980 6712 11008 6752
rect 11882 6740 11888 6752
rect 11940 6740 11946 6792
rect 12158 6740 12164 6792
rect 12216 6780 12222 6792
rect 12360 6780 12388 6820
rect 12216 6752 12388 6780
rect 12216 6740 12222 6752
rect 12710 6740 12716 6792
rect 12768 6780 12774 6792
rect 13004 6789 13032 6820
rect 13096 6820 14749 6848
rect 12897 6783 12955 6789
rect 12897 6780 12909 6783
rect 12768 6752 12909 6780
rect 12768 6740 12774 6752
rect 12897 6749 12909 6752
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 13000 6783 13058 6789
rect 13000 6749 13012 6783
rect 13046 6749 13058 6783
rect 13000 6743 13058 6749
rect 10643 6684 11008 6712
rect 11048 6715 11106 6721
rect 10643 6681 10655 6684
rect 10597 6675 10655 6681
rect 11048 6681 11060 6715
rect 11094 6712 11106 6715
rect 13096 6712 13124 6820
rect 14737 6817 14749 6820
rect 14783 6817 14795 6851
rect 17494 6848 17500 6860
rect 17455 6820 17500 6848
rect 14737 6811 14795 6817
rect 17494 6808 17500 6820
rect 17552 6808 17558 6860
rect 17589 6851 17647 6857
rect 17589 6817 17601 6851
rect 17635 6817 17647 6851
rect 18414 6848 18420 6860
rect 18375 6820 18420 6848
rect 17589 6811 17647 6817
rect 13630 6740 13636 6792
rect 13688 6780 13694 6792
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13688 6752 14105 6780
rect 13688 6740 13694 6752
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14093 6743 14151 6749
rect 15473 6783 15531 6789
rect 15473 6749 15485 6783
rect 15519 6780 15531 6783
rect 15519 6752 15608 6780
rect 15519 6749 15531 6752
rect 15473 6743 15531 6749
rect 11094 6684 13124 6712
rect 11094 6681 11106 6684
rect 11048 6675 11106 6681
rect 13170 6672 13176 6724
rect 13228 6712 13234 6724
rect 13725 6715 13783 6721
rect 13725 6712 13737 6715
rect 13228 6684 13737 6712
rect 13228 6672 13234 6684
rect 13725 6681 13737 6684
rect 13771 6681 13783 6715
rect 13725 6675 13783 6681
rect 8941 6647 8999 6653
rect 8941 6613 8953 6647
rect 8987 6613 8999 6647
rect 8941 6607 8999 6613
rect 9030 6604 9036 6656
rect 9088 6644 9094 6656
rect 10505 6647 10563 6653
rect 10505 6644 10517 6647
rect 9088 6616 10517 6644
rect 9088 6604 9094 6616
rect 10505 6613 10517 6616
rect 10551 6613 10563 6647
rect 10505 6607 10563 6613
rect 11974 6604 11980 6656
rect 12032 6644 12038 6656
rect 13633 6647 13691 6653
rect 13633 6644 13645 6647
rect 12032 6616 13645 6644
rect 12032 6604 12038 6616
rect 13633 6613 13645 6616
rect 13679 6613 13691 6647
rect 13633 6607 13691 6613
rect 14826 6604 14832 6656
rect 14884 6644 14890 6656
rect 15580 6653 15608 6752
rect 16390 6740 16396 6792
rect 16448 6780 16454 6792
rect 16945 6783 17003 6789
rect 16945 6780 16957 6783
rect 16448 6752 16957 6780
rect 16448 6740 16454 6752
rect 16945 6749 16957 6752
rect 16991 6749 17003 6783
rect 16945 6743 17003 6749
rect 17310 6740 17316 6792
rect 17368 6780 17374 6792
rect 17604 6780 17632 6811
rect 18414 6808 18420 6820
rect 18472 6808 18478 6860
rect 18524 6848 18552 6888
rect 18598 6876 18604 6928
rect 18656 6916 18662 6928
rect 19150 6916 19156 6928
rect 18656 6888 19156 6916
rect 18656 6876 18662 6888
rect 19150 6876 19156 6888
rect 19208 6876 19214 6928
rect 20806 6916 20812 6928
rect 19260 6888 20812 6916
rect 19260 6848 19288 6888
rect 20806 6876 20812 6888
rect 20864 6876 20870 6928
rect 22465 6919 22523 6925
rect 22465 6885 22477 6919
rect 22511 6885 22523 6919
rect 22465 6879 22523 6885
rect 18524 6820 19288 6848
rect 19337 6851 19395 6857
rect 19337 6817 19349 6851
rect 19383 6848 19395 6851
rect 19426 6848 19432 6860
rect 19383 6820 19432 6848
rect 19383 6817 19395 6820
rect 19337 6811 19395 6817
rect 19426 6808 19432 6820
rect 19484 6808 19490 6860
rect 21085 6851 21143 6857
rect 21085 6848 21097 6851
rect 20456 6820 21097 6848
rect 17368 6752 17632 6780
rect 17368 6740 17374 6752
rect 18230 6740 18236 6792
rect 18288 6780 18294 6792
rect 20456 6789 20484 6820
rect 21085 6817 21097 6820
rect 21131 6817 21143 6851
rect 21085 6811 21143 6817
rect 20441 6783 20499 6789
rect 20441 6780 20453 6783
rect 18288 6752 20453 6780
rect 18288 6740 18294 6752
rect 20441 6749 20453 6752
rect 20487 6749 20499 6783
rect 20806 6780 20812 6792
rect 20767 6752 20812 6780
rect 20441 6743 20499 6749
rect 20806 6740 20812 6752
rect 20864 6740 20870 6792
rect 21100 6780 21128 6811
rect 21174 6780 21180 6792
rect 21100 6752 21180 6780
rect 21174 6740 21180 6752
rect 21232 6740 21238 6792
rect 22186 6780 22192 6792
rect 21284 6752 22192 6780
rect 16666 6712 16672 6724
rect 16724 6721 16730 6724
rect 16636 6684 16672 6712
rect 16666 6672 16672 6684
rect 16724 6675 16736 6721
rect 17405 6715 17463 6721
rect 17405 6712 17417 6715
rect 16776 6684 17417 6712
rect 16724 6672 16730 6675
rect 16776 6656 16804 6684
rect 17405 6681 17417 6684
rect 17451 6681 17463 6715
rect 18138 6712 18144 6724
rect 18099 6684 18144 6712
rect 17405 6675 17463 6681
rect 18138 6672 18144 6684
rect 18196 6672 18202 6724
rect 19426 6672 19432 6724
rect 19484 6712 19490 6724
rect 19705 6715 19763 6721
rect 19705 6712 19717 6715
rect 19484 6684 19717 6712
rect 19484 6672 19490 6684
rect 19705 6681 19717 6684
rect 19751 6681 19763 6715
rect 21284 6712 21312 6752
rect 22186 6740 22192 6752
rect 22244 6740 22250 6792
rect 19705 6675 19763 6681
rect 20916 6684 21312 6712
rect 21352 6715 21410 6721
rect 15565 6647 15623 6653
rect 14884 6616 14929 6644
rect 14884 6604 14890 6616
rect 15565 6613 15577 6647
rect 15611 6644 15623 6647
rect 16574 6644 16580 6656
rect 15611 6616 16580 6644
rect 15611 6613 15623 6616
rect 15565 6607 15623 6613
rect 16574 6604 16580 6616
rect 16632 6604 16638 6656
rect 16758 6604 16764 6656
rect 16816 6604 16822 6656
rect 16942 6604 16948 6656
rect 17000 6644 17006 6656
rect 17037 6647 17095 6653
rect 17037 6644 17049 6647
rect 17000 6616 17049 6644
rect 17000 6604 17006 6616
rect 17037 6613 17049 6616
rect 17083 6613 17095 6647
rect 18598 6644 18604 6656
rect 18559 6616 18604 6644
rect 17037 6607 17095 6613
rect 18598 6604 18604 6616
rect 18656 6604 18662 6656
rect 18690 6604 18696 6656
rect 18748 6644 18754 6656
rect 19613 6647 19671 6653
rect 18748 6616 18793 6644
rect 18748 6604 18754 6616
rect 19613 6613 19625 6647
rect 19659 6644 19671 6647
rect 20916 6644 20944 6684
rect 21352 6681 21364 6715
rect 21398 6712 21410 6715
rect 21450 6712 21456 6724
rect 21398 6684 21456 6712
rect 21398 6681 21410 6684
rect 21352 6675 21410 6681
rect 21450 6672 21456 6684
rect 21508 6672 21514 6724
rect 21542 6672 21548 6724
rect 21600 6712 21606 6724
rect 21910 6712 21916 6724
rect 21600 6684 21916 6712
rect 21600 6672 21606 6684
rect 21910 6672 21916 6684
rect 21968 6712 21974 6724
rect 22480 6712 22508 6879
rect 23382 6848 23388 6860
rect 22756 6820 23388 6848
rect 22646 6740 22652 6792
rect 22704 6780 22710 6792
rect 22756 6789 22784 6820
rect 23382 6808 23388 6820
rect 23440 6808 23446 6860
rect 22741 6783 22799 6789
rect 22741 6780 22753 6783
rect 22704 6752 22753 6780
rect 22704 6740 22710 6752
rect 22741 6749 22753 6752
rect 22787 6749 22799 6783
rect 22741 6743 22799 6749
rect 22833 6783 22891 6789
rect 22833 6749 22845 6783
rect 22879 6749 22891 6783
rect 22833 6743 22891 6749
rect 21968 6684 22508 6712
rect 21968 6672 21974 6684
rect 19659 6616 20944 6644
rect 20993 6647 21051 6653
rect 19659 6613 19671 6616
rect 19613 6607 19671 6613
rect 20993 6613 21005 6647
rect 21039 6644 21051 6647
rect 22848 6644 22876 6743
rect 23014 6644 23020 6656
rect 21039 6616 22876 6644
rect 22975 6616 23020 6644
rect 21039 6613 21051 6616
rect 20993 6607 21051 6613
rect 23014 6604 23020 6616
rect 23072 6604 23078 6656
rect 1104 6554 23460 6576
rect 1104 6502 6548 6554
rect 6600 6502 6612 6554
rect 6664 6502 6676 6554
rect 6728 6502 6740 6554
rect 6792 6502 6804 6554
rect 6856 6502 12146 6554
rect 12198 6502 12210 6554
rect 12262 6502 12274 6554
rect 12326 6502 12338 6554
rect 12390 6502 12402 6554
rect 12454 6502 17744 6554
rect 17796 6502 17808 6554
rect 17860 6502 17872 6554
rect 17924 6502 17936 6554
rect 17988 6502 18000 6554
rect 18052 6502 23460 6554
rect 1104 6480 23460 6502
rect 2314 6400 2320 6452
rect 2372 6440 2378 6452
rect 2409 6443 2467 6449
rect 2409 6440 2421 6443
rect 2372 6412 2421 6440
rect 2372 6400 2378 6412
rect 2409 6409 2421 6412
rect 2455 6409 2467 6443
rect 2774 6440 2780 6452
rect 2735 6412 2780 6440
rect 2409 6403 2467 6409
rect 2774 6400 2780 6412
rect 2832 6400 2838 6452
rect 2958 6400 2964 6452
rect 3016 6440 3022 6452
rect 4522 6440 4528 6452
rect 3016 6412 4528 6440
rect 3016 6400 3022 6412
rect 4522 6400 4528 6412
rect 4580 6400 4586 6452
rect 4801 6443 4859 6449
rect 4801 6409 4813 6443
rect 4847 6440 4859 6443
rect 5534 6440 5540 6452
rect 4847 6412 5540 6440
rect 4847 6409 4859 6412
rect 4801 6403 4859 6409
rect 1762 6304 1768 6316
rect 1723 6276 1768 6304
rect 1762 6264 1768 6276
rect 1820 6264 1826 6316
rect 3326 6264 3332 6316
rect 3384 6304 3390 6316
rect 3421 6307 3479 6313
rect 3421 6304 3433 6307
rect 3384 6276 3433 6304
rect 3384 6264 3390 6276
rect 3421 6273 3433 6276
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 4709 6307 4767 6313
rect 4709 6273 4721 6307
rect 4755 6304 4767 6307
rect 4816 6304 4844 6403
rect 5534 6400 5540 6412
rect 5592 6400 5598 6452
rect 7006 6440 7012 6452
rect 6967 6412 7012 6440
rect 7006 6400 7012 6412
rect 7064 6400 7070 6452
rect 7466 6440 7472 6452
rect 7427 6412 7472 6440
rect 7466 6400 7472 6412
rect 7524 6400 7530 6452
rect 7558 6400 7564 6452
rect 7616 6440 7622 6452
rect 11885 6443 11943 6449
rect 7616 6412 11744 6440
rect 7616 6400 7622 6412
rect 5936 6375 5994 6381
rect 5936 6341 5948 6375
rect 5982 6372 5994 6375
rect 5982 6344 6914 6372
rect 5982 6341 5994 6344
rect 5936 6335 5994 6341
rect 6178 6304 6184 6316
rect 4755 6276 4844 6304
rect 6139 6276 6184 6304
rect 4755 6273 4767 6276
rect 4709 6267 4767 6273
rect 6178 6264 6184 6276
rect 6236 6264 6242 6316
rect 6362 6304 6368 6316
rect 6323 6276 6368 6304
rect 6362 6264 6368 6276
rect 6420 6264 6426 6316
rect 6886 6304 6914 6344
rect 7190 6332 7196 6384
rect 7248 6372 7254 6384
rect 8266 6375 8324 6381
rect 8266 6372 8278 6375
rect 7248 6344 8278 6372
rect 7248 6332 7254 6344
rect 8266 6341 8278 6344
rect 8312 6341 8324 6375
rect 9030 6372 9036 6384
rect 8266 6335 8324 6341
rect 8404 6344 9036 6372
rect 7466 6304 7472 6316
rect 6886 6276 7472 6304
rect 7466 6264 7472 6276
rect 7524 6264 7530 6316
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 7834 6304 7840 6316
rect 7607 6276 7840 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 7834 6264 7840 6276
rect 7892 6264 7898 6316
rect 8018 6304 8024 6316
rect 7979 6276 8024 6304
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8404 6304 8432 6344
rect 9030 6332 9036 6344
rect 9088 6332 9094 6384
rect 9214 6332 9220 6384
rect 9272 6372 9278 6384
rect 9585 6375 9643 6381
rect 9585 6372 9597 6375
rect 9272 6344 9597 6372
rect 9272 6332 9278 6344
rect 9585 6341 9597 6344
rect 9631 6341 9643 6375
rect 11716 6372 11744 6412
rect 11885 6409 11897 6443
rect 11931 6440 11943 6443
rect 13078 6440 13084 6452
rect 11931 6412 13084 6440
rect 11931 6409 11943 6412
rect 11885 6403 11943 6409
rect 13078 6400 13084 6412
rect 13136 6400 13142 6452
rect 13170 6400 13176 6452
rect 13228 6440 13234 6452
rect 14734 6440 14740 6452
rect 13228 6412 14740 6440
rect 13228 6400 13234 6412
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 14921 6443 14979 6449
rect 14921 6409 14933 6443
rect 14967 6440 14979 6443
rect 16758 6440 16764 6452
rect 14967 6412 16764 6440
rect 14967 6409 14979 6412
rect 14921 6403 14979 6409
rect 16758 6400 16764 6412
rect 16816 6400 16822 6452
rect 16942 6440 16948 6452
rect 16903 6412 16948 6440
rect 16942 6400 16948 6412
rect 17000 6400 17006 6452
rect 19978 6400 19984 6452
rect 20036 6440 20042 6452
rect 20171 6443 20229 6449
rect 20171 6440 20183 6443
rect 20036 6412 20183 6440
rect 20036 6400 20042 6412
rect 20171 6409 20183 6412
rect 20217 6409 20229 6443
rect 20171 6403 20229 6409
rect 22370 6400 22376 6452
rect 22428 6440 22434 6452
rect 22557 6443 22615 6449
rect 22557 6440 22569 6443
rect 22428 6412 22569 6440
rect 22428 6400 22434 6412
rect 22557 6409 22569 6412
rect 22603 6409 22615 6443
rect 22557 6403 22615 6409
rect 12066 6372 12072 6384
rect 11716 6344 12072 6372
rect 9585 6335 9643 6341
rect 12066 6332 12072 6344
rect 12124 6372 12130 6384
rect 12437 6375 12495 6381
rect 12437 6372 12449 6375
rect 12124 6344 12449 6372
rect 12124 6332 12130 6344
rect 12437 6341 12449 6344
rect 12483 6341 12495 6375
rect 12437 6335 12495 6341
rect 12544 6344 12940 6372
rect 8128 6276 8432 6304
rect 7377 6239 7435 6245
rect 7377 6205 7389 6239
rect 7423 6236 7435 6239
rect 7742 6236 7748 6248
rect 7423 6208 7748 6236
rect 7423 6205 7435 6208
rect 7377 6199 7435 6205
rect 7742 6196 7748 6208
rect 7800 6236 7806 6248
rect 8128 6236 8156 6276
rect 8570 6264 8576 6316
rect 8628 6304 8634 6316
rect 9950 6304 9956 6316
rect 8628 6276 9444 6304
rect 9911 6276 9956 6304
rect 8628 6264 8634 6276
rect 7800 6208 8156 6236
rect 7800 6196 7806 6208
rect 4065 6171 4123 6177
rect 4065 6137 4077 6171
rect 4111 6168 4123 6171
rect 5166 6168 5172 6180
rect 4111 6140 5172 6168
rect 4111 6137 4123 6140
rect 4065 6131 4123 6137
rect 5166 6128 5172 6140
rect 5224 6128 5230 6180
rect 9416 6177 9444 6276
rect 9950 6264 9956 6276
rect 10008 6264 10014 6316
rect 10220 6307 10278 6313
rect 10220 6273 10232 6307
rect 10266 6304 10278 6307
rect 10962 6304 10968 6316
rect 10266 6276 10968 6304
rect 10266 6273 10278 6276
rect 10220 6267 10278 6273
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 11974 6236 11980 6248
rect 11935 6208 11980 6236
rect 11974 6196 11980 6208
rect 12032 6196 12038 6248
rect 12161 6239 12219 6245
rect 12161 6205 12173 6239
rect 12207 6236 12219 6239
rect 12544 6236 12572 6344
rect 12621 6307 12679 6313
rect 12621 6273 12633 6307
rect 12667 6273 12679 6307
rect 12802 6304 12808 6316
rect 12763 6276 12808 6304
rect 12621 6267 12679 6273
rect 12207 6208 12572 6236
rect 12636 6236 12664 6267
rect 12802 6264 12808 6276
rect 12860 6264 12866 6316
rect 12912 6304 12940 6344
rect 14826 6332 14832 6384
rect 14884 6372 14890 6384
rect 15350 6375 15408 6381
rect 15350 6372 15362 6375
rect 14884 6344 15362 6372
rect 14884 6332 14890 6344
rect 15350 6341 15362 6344
rect 15396 6341 15408 6375
rect 18138 6372 18144 6384
rect 18099 6344 18144 6372
rect 15350 6335 15408 6341
rect 18138 6332 18144 6344
rect 18196 6332 18202 6384
rect 22278 6332 22284 6384
rect 22336 6372 22342 6384
rect 22649 6375 22707 6381
rect 22649 6372 22661 6375
rect 22336 6344 22661 6372
rect 22336 6332 22342 6344
rect 22649 6341 22661 6344
rect 22695 6341 22707 6375
rect 22649 6335 22707 6341
rect 13630 6304 13636 6316
rect 12912 6276 13636 6304
rect 13630 6264 13636 6276
rect 13688 6264 13694 6316
rect 15102 6304 15108 6316
rect 15063 6276 15108 6304
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 17034 6304 17040 6316
rect 16995 6276 17040 6304
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 17494 6304 17500 6316
rect 17455 6276 17500 6304
rect 17494 6264 17500 6276
rect 17552 6264 17558 6316
rect 18230 6304 18236 6316
rect 18191 6276 18236 6304
rect 18230 6264 18236 6276
rect 18288 6264 18294 6316
rect 18322 6264 18328 6316
rect 18380 6304 18386 6316
rect 18489 6307 18547 6313
rect 18489 6304 18501 6307
rect 18380 6276 18501 6304
rect 18380 6264 18386 6276
rect 18489 6273 18501 6276
rect 18535 6273 18547 6307
rect 18489 6267 18547 6273
rect 19334 6264 19340 6316
rect 19392 6304 19398 6316
rect 20441 6307 20499 6313
rect 19392 6276 20208 6304
rect 19392 6264 19398 6276
rect 13170 6245 13176 6248
rect 13128 6239 13176 6245
rect 13128 6236 13140 6239
rect 12636 6208 13140 6236
rect 12207 6205 12219 6208
rect 12161 6199 12219 6205
rect 13128 6205 13140 6208
rect 13174 6205 13176 6239
rect 13128 6199 13176 6205
rect 9401 6171 9459 6177
rect 9401 6137 9413 6171
rect 9447 6168 9459 6171
rect 9766 6168 9772 6180
rect 9447 6140 9772 6168
rect 9447 6137 9459 6140
rect 9401 6131 9459 6137
rect 9766 6128 9772 6140
rect 9824 6128 9830 6180
rect 11333 6171 11391 6177
rect 11333 6137 11345 6171
rect 11379 6168 11391 6171
rect 12176 6168 12204 6199
rect 13170 6196 13176 6199
rect 13228 6196 13234 6248
rect 13262 6196 13268 6248
rect 13320 6236 13326 6248
rect 13320 6208 13365 6236
rect 13320 6196 13326 6208
rect 13446 6196 13452 6248
rect 13504 6236 13510 6248
rect 13541 6239 13599 6245
rect 13541 6236 13553 6239
rect 13504 6208 13553 6236
rect 13504 6196 13510 6208
rect 13541 6205 13553 6208
rect 13587 6205 13599 6239
rect 13541 6199 13599 6205
rect 16853 6239 16911 6245
rect 16853 6205 16865 6239
rect 16899 6236 16911 6239
rect 17126 6236 17132 6248
rect 16899 6208 17132 6236
rect 16899 6205 16911 6208
rect 16853 6199 16911 6205
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 19702 6236 19708 6248
rect 19663 6208 19708 6236
rect 19702 6196 19708 6208
rect 19760 6196 19766 6248
rect 20180 6245 20208 6276
rect 20441 6273 20453 6307
rect 20487 6304 20499 6307
rect 20898 6304 20904 6316
rect 20487 6276 20904 6304
rect 20487 6273 20499 6276
rect 20441 6267 20499 6273
rect 20898 6264 20904 6276
rect 20956 6264 20962 6316
rect 22189 6307 22247 6313
rect 22189 6304 22201 6307
rect 21008 6276 22201 6304
rect 20168 6239 20226 6245
rect 20168 6205 20180 6239
rect 20214 6236 20226 6239
rect 21008 6236 21036 6276
rect 22189 6273 22201 6276
rect 22235 6273 22247 6307
rect 22189 6267 22247 6273
rect 22833 6307 22891 6313
rect 22833 6273 22845 6307
rect 22879 6304 22891 6307
rect 23106 6304 23112 6316
rect 22879 6276 23112 6304
rect 22879 6273 22891 6276
rect 22833 6267 22891 6273
rect 23106 6264 23112 6276
rect 23164 6264 23170 6316
rect 21910 6236 21916 6248
rect 20214 6208 21036 6236
rect 21871 6208 21916 6236
rect 20214 6205 20226 6208
rect 20168 6199 20226 6205
rect 21910 6196 21916 6208
rect 21968 6196 21974 6248
rect 22097 6239 22155 6245
rect 22097 6205 22109 6239
rect 22143 6205 22155 6239
rect 22097 6199 22155 6205
rect 11379 6140 12204 6168
rect 14200 6140 14780 6168
rect 11379 6137 11391 6140
rect 11333 6131 11391 6137
rect 7929 6103 7987 6109
rect 7929 6069 7941 6103
rect 7975 6100 7987 6103
rect 8386 6100 8392 6112
rect 7975 6072 8392 6100
rect 7975 6069 7987 6072
rect 7929 6063 7987 6069
rect 8386 6060 8392 6072
rect 8444 6060 8450 6112
rect 9677 6103 9735 6109
rect 9677 6069 9689 6103
rect 9723 6100 9735 6103
rect 9858 6100 9864 6112
rect 9723 6072 9864 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 11517 6103 11575 6109
rect 11517 6069 11529 6103
rect 11563 6100 11575 6103
rect 11882 6100 11888 6112
rect 11563 6072 11888 6100
rect 11563 6069 11575 6072
rect 11517 6063 11575 6069
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 13630 6060 13636 6112
rect 13688 6100 13694 6112
rect 14200 6100 14228 6140
rect 14642 6100 14648 6112
rect 13688 6072 14228 6100
rect 14603 6072 14648 6100
rect 13688 6060 13694 6072
rect 14642 6060 14648 6072
rect 14700 6060 14706 6112
rect 14752 6100 14780 6140
rect 16040 6140 17540 6168
rect 16040 6100 16068 6140
rect 14752 6072 16068 6100
rect 16485 6103 16543 6109
rect 16485 6069 16497 6103
rect 16531 6100 16543 6103
rect 16942 6100 16948 6112
rect 16531 6072 16948 6100
rect 16531 6069 16543 6072
rect 16485 6063 16543 6069
rect 16942 6060 16948 6072
rect 17000 6060 17006 6112
rect 17402 6100 17408 6112
rect 17363 6072 17408 6100
rect 17402 6060 17408 6072
rect 17460 6060 17466 6112
rect 17512 6100 17540 6140
rect 19426 6100 19432 6112
rect 17512 6072 19432 6100
rect 19426 6060 19432 6072
rect 19484 6060 19490 6112
rect 19613 6103 19671 6109
rect 19613 6069 19625 6103
rect 19659 6100 19671 6103
rect 20162 6100 20168 6112
rect 19659 6072 20168 6100
rect 19659 6069 19671 6072
rect 19613 6063 19671 6069
rect 20162 6060 20168 6072
rect 20220 6060 20226 6112
rect 20254 6060 20260 6112
rect 20312 6100 20318 6112
rect 21545 6103 21603 6109
rect 21545 6100 21557 6103
rect 20312 6072 21557 6100
rect 20312 6060 20318 6072
rect 21545 6069 21557 6072
rect 21591 6100 21603 6103
rect 22112 6100 22140 6199
rect 23014 6100 23020 6112
rect 21591 6072 22140 6100
rect 22975 6072 23020 6100
rect 21591 6069 21603 6072
rect 21545 6063 21603 6069
rect 23014 6060 23020 6072
rect 23072 6060 23078 6112
rect 1104 6010 23460 6032
rect 1104 5958 3749 6010
rect 3801 5958 3813 6010
rect 3865 5958 3877 6010
rect 3929 5958 3941 6010
rect 3993 5958 4005 6010
rect 4057 5958 9347 6010
rect 9399 5958 9411 6010
rect 9463 5958 9475 6010
rect 9527 5958 9539 6010
rect 9591 5958 9603 6010
rect 9655 5958 14945 6010
rect 14997 5958 15009 6010
rect 15061 5958 15073 6010
rect 15125 5958 15137 6010
rect 15189 5958 15201 6010
rect 15253 5958 20543 6010
rect 20595 5958 20607 6010
rect 20659 5958 20671 6010
rect 20723 5958 20735 6010
rect 20787 5958 20799 6010
rect 20851 5958 23460 6010
rect 1104 5936 23460 5958
rect 4338 5856 4344 5908
rect 4396 5896 4402 5908
rect 4433 5899 4491 5905
rect 4433 5896 4445 5899
rect 4396 5868 4445 5896
rect 4396 5856 4402 5868
rect 4433 5865 4445 5868
rect 4479 5865 4491 5899
rect 4433 5859 4491 5865
rect 4614 5856 4620 5908
rect 4672 5896 4678 5908
rect 4798 5896 4804 5908
rect 4672 5868 4804 5896
rect 4672 5856 4678 5868
rect 4798 5856 4804 5868
rect 4856 5856 4862 5908
rect 5350 5856 5356 5908
rect 5408 5896 5414 5908
rect 6362 5896 6368 5908
rect 5408 5868 6368 5896
rect 5408 5856 5414 5868
rect 6362 5856 6368 5868
rect 6420 5896 6426 5908
rect 6917 5899 6975 5905
rect 6917 5896 6929 5899
rect 6420 5868 6929 5896
rect 6420 5856 6426 5868
rect 6917 5865 6929 5868
rect 6963 5865 6975 5899
rect 6917 5859 6975 5865
rect 8018 5856 8024 5908
rect 8076 5896 8082 5908
rect 12802 5896 12808 5908
rect 8076 5868 8340 5896
rect 8076 5856 8082 5868
rect 3620 5732 4752 5760
rect 3620 5701 3648 5732
rect 3605 5695 3663 5701
rect 3605 5661 3617 5695
rect 3651 5661 3663 5695
rect 3605 5655 3663 5661
rect 3694 5652 3700 5704
rect 3752 5692 3758 5704
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 3752 5664 3801 5692
rect 3752 5652 3758 5664
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 4724 5692 4752 5732
rect 4798 5720 4804 5772
rect 4856 5760 4862 5772
rect 5442 5760 5448 5772
rect 5500 5769 5506 5772
rect 8312 5769 8340 5868
rect 11440 5868 12808 5896
rect 4856 5732 5448 5760
rect 4856 5720 4862 5732
rect 5442 5720 5448 5732
rect 5500 5760 5510 5769
rect 8297 5763 8355 5769
rect 5500 5732 5545 5760
rect 5500 5723 5510 5732
rect 8297 5729 8309 5763
rect 8343 5760 8355 5763
rect 8478 5760 8484 5772
rect 8343 5732 8484 5760
rect 8343 5729 8355 5732
rect 8297 5723 8355 5729
rect 5500 5720 5506 5723
rect 8478 5720 8484 5732
rect 8536 5760 8542 5772
rect 10318 5760 10324 5772
rect 8536 5732 10324 5760
rect 8536 5720 8542 5732
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 11440 5769 11468 5868
rect 12802 5856 12808 5868
rect 12860 5856 12866 5908
rect 13541 5899 13599 5905
rect 13541 5865 13553 5899
rect 13587 5896 13599 5899
rect 13630 5896 13636 5908
rect 13587 5868 13636 5896
rect 13587 5865 13599 5868
rect 13541 5859 13599 5865
rect 13630 5856 13636 5868
rect 13688 5856 13694 5908
rect 13909 5899 13967 5905
rect 13909 5865 13921 5899
rect 13955 5896 13967 5899
rect 14090 5896 14096 5908
rect 13955 5868 14096 5896
rect 13955 5865 13967 5868
rect 13909 5859 13967 5865
rect 14090 5856 14096 5868
rect 14148 5896 14154 5908
rect 20254 5896 20260 5908
rect 14148 5868 15148 5896
rect 14148 5856 14154 5868
rect 11425 5763 11483 5769
rect 11425 5729 11437 5763
rect 11471 5729 11483 5763
rect 11425 5723 11483 5729
rect 11882 5720 11888 5772
rect 11940 5760 11946 5772
rect 12986 5760 12992 5772
rect 11940 5732 11985 5760
rect 12084 5732 12992 5760
rect 11940 5720 11946 5732
rect 5258 5692 5264 5704
rect 4724 5664 5264 5692
rect 3789 5655 3847 5661
rect 5258 5652 5264 5664
rect 5316 5652 5322 5704
rect 5350 5652 5356 5704
rect 5408 5692 5414 5704
rect 5408 5664 5453 5692
rect 5552 5664 8248 5692
rect 5408 5652 5414 5664
rect 3510 5584 3516 5636
rect 3568 5624 3574 5636
rect 5552 5624 5580 5664
rect 5701 5627 5759 5633
rect 5701 5624 5713 5627
rect 3568 5596 5580 5624
rect 5644 5596 5713 5624
rect 3568 5584 3574 5596
rect 2961 5559 3019 5565
rect 2961 5525 2973 5559
rect 3007 5556 3019 5559
rect 4522 5556 4528 5568
rect 3007 5528 4528 5556
rect 3007 5525 3019 5528
rect 2961 5519 3019 5525
rect 4522 5516 4528 5528
rect 4580 5516 4586 5568
rect 4709 5559 4767 5565
rect 4709 5525 4721 5559
rect 4755 5556 4767 5559
rect 5074 5556 5080 5568
rect 4755 5528 5080 5556
rect 4755 5525 4767 5528
rect 4709 5519 4767 5525
rect 5074 5516 5080 5528
rect 5132 5516 5138 5568
rect 5166 5516 5172 5568
rect 5224 5556 5230 5568
rect 5644 5556 5672 5596
rect 5701 5593 5713 5596
rect 5747 5593 5759 5627
rect 5701 5587 5759 5593
rect 5810 5584 5816 5636
rect 5868 5624 5874 5636
rect 8030 5627 8088 5633
rect 8030 5624 8042 5627
rect 5868 5596 8042 5624
rect 5868 5584 5874 5596
rect 8030 5593 8042 5596
rect 8076 5593 8088 5627
rect 8220 5624 8248 5664
rect 8386 5652 8392 5704
rect 8444 5692 8450 5704
rect 8573 5695 8631 5701
rect 8573 5692 8585 5695
rect 8444 5664 8585 5692
rect 8444 5652 8450 5664
rect 8573 5661 8585 5664
rect 8619 5661 8631 5695
rect 12084 5692 12112 5732
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 15120 5760 15148 5868
rect 15212 5868 20260 5896
rect 15212 5840 15240 5868
rect 20254 5856 20260 5868
rect 20312 5856 20318 5908
rect 21450 5896 21456 5908
rect 20364 5868 21456 5896
rect 15194 5788 15200 5840
rect 15252 5788 15258 5840
rect 16666 5788 16672 5840
rect 16724 5828 16730 5840
rect 19886 5828 19892 5840
rect 16724 5800 16769 5828
rect 19847 5800 19892 5828
rect 16724 5788 16730 5800
rect 19886 5788 19892 5800
rect 19944 5788 19950 5840
rect 20364 5828 20392 5868
rect 21450 5856 21456 5868
rect 21508 5856 21514 5908
rect 20272 5800 20392 5828
rect 15120 5732 16528 5760
rect 8573 5655 8631 5661
rect 11532 5664 12112 5692
rect 12161 5695 12219 5701
rect 9585 5627 9643 5633
rect 9585 5624 9597 5627
rect 8220 5596 9597 5624
rect 8030 5587 8088 5593
rect 9585 5593 9597 5596
rect 9631 5593 9643 5627
rect 9585 5587 9643 5593
rect 11333 5627 11391 5633
rect 11333 5593 11345 5627
rect 11379 5624 11391 5627
rect 11532 5624 11560 5664
rect 12161 5661 12173 5695
rect 12207 5692 12219 5695
rect 12618 5692 12624 5704
rect 12207 5664 12624 5692
rect 12207 5661 12219 5664
rect 12161 5655 12219 5661
rect 12618 5652 12624 5664
rect 12676 5692 12682 5704
rect 14093 5695 14151 5701
rect 12676 5664 14044 5692
rect 12676 5652 12682 5664
rect 13722 5624 13728 5636
rect 11379 5596 11560 5624
rect 13683 5596 13728 5624
rect 11379 5593 11391 5596
rect 11333 5587 11391 5593
rect 13722 5584 13728 5596
rect 13780 5584 13786 5636
rect 5224 5528 5672 5556
rect 5224 5516 5230 5528
rect 6454 5516 6460 5568
rect 6512 5556 6518 5568
rect 6825 5559 6883 5565
rect 6825 5556 6837 5559
rect 6512 5528 6837 5556
rect 6512 5516 6518 5528
rect 6825 5525 6837 5528
rect 6871 5525 6883 5559
rect 6825 5519 6883 5525
rect 8757 5559 8815 5565
rect 8757 5525 8769 5559
rect 8803 5556 8815 5559
rect 10686 5556 10692 5568
rect 8803 5528 10692 5556
rect 8803 5525 8815 5528
rect 8757 5519 8815 5525
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 11891 5559 11949 5565
rect 11891 5525 11903 5559
rect 11937 5556 11949 5559
rect 12066 5556 12072 5568
rect 11937 5528 12072 5556
rect 11937 5525 11949 5528
rect 11891 5519 11949 5525
rect 12066 5516 12072 5528
rect 12124 5516 12130 5568
rect 13265 5559 13323 5565
rect 13265 5525 13277 5559
rect 13311 5556 13323 5559
rect 13354 5556 13360 5568
rect 13311 5528 13360 5556
rect 13311 5525 13323 5528
rect 13265 5519 13323 5525
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 14016 5556 14044 5664
rect 14093 5661 14105 5695
rect 14139 5692 14151 5695
rect 15286 5692 15292 5704
rect 14139 5664 15292 5692
rect 14139 5661 14151 5664
rect 14093 5655 14151 5661
rect 15286 5652 15292 5664
rect 15344 5692 15350 5704
rect 16500 5701 16528 5732
rect 16758 5720 16764 5772
rect 16816 5760 16822 5772
rect 17037 5763 17095 5769
rect 17037 5760 17049 5763
rect 16816 5732 17049 5760
rect 16816 5720 16822 5732
rect 17037 5729 17049 5732
rect 17083 5729 17095 5763
rect 17037 5723 17095 5729
rect 18690 5720 18696 5772
rect 18748 5760 18754 5772
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 18748 5732 19257 5760
rect 18748 5720 18754 5732
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 19426 5720 19432 5772
rect 19484 5760 19490 5772
rect 20272 5760 20300 5800
rect 22922 5760 22928 5772
rect 19484 5732 20300 5760
rect 22883 5732 22928 5760
rect 19484 5720 19490 5732
rect 22922 5720 22928 5732
rect 22980 5720 22986 5772
rect 16485 5695 16543 5701
rect 15344 5664 15792 5692
rect 15344 5652 15350 5664
rect 14360 5627 14418 5633
rect 14360 5593 14372 5627
rect 14406 5624 14418 5627
rect 15378 5624 15384 5636
rect 14406 5596 15384 5624
rect 14406 5593 14418 5596
rect 14360 5587 14418 5593
rect 15378 5584 15384 5596
rect 15436 5584 15442 5636
rect 15764 5633 15792 5664
rect 16485 5661 16497 5695
rect 16531 5661 16543 5695
rect 17402 5692 17408 5704
rect 17363 5664 17408 5692
rect 16485 5655 16543 5661
rect 17402 5652 17408 5664
rect 17460 5652 17466 5704
rect 17681 5695 17739 5701
rect 17681 5661 17693 5695
rect 17727 5692 17739 5695
rect 18230 5692 18236 5704
rect 17727 5664 18236 5692
rect 17727 5661 17739 5664
rect 17681 5655 17739 5661
rect 18230 5652 18236 5664
rect 18288 5652 18294 5704
rect 19521 5695 19579 5701
rect 19521 5661 19533 5695
rect 19567 5692 19579 5695
rect 20714 5692 20720 5704
rect 19567 5664 20720 5692
rect 19567 5661 19579 5664
rect 19521 5655 19579 5661
rect 20714 5652 20720 5664
rect 20772 5652 20778 5704
rect 21174 5652 21180 5704
rect 21232 5692 21238 5704
rect 21269 5695 21327 5701
rect 21269 5692 21281 5695
rect 21232 5664 21281 5692
rect 21232 5652 21238 5664
rect 21269 5661 21281 5664
rect 21315 5692 21327 5695
rect 21453 5695 21511 5701
rect 21453 5692 21465 5695
rect 21315 5664 21465 5692
rect 21315 5661 21327 5664
rect 21269 5655 21327 5661
rect 21453 5661 21465 5664
rect 21499 5661 21511 5695
rect 21453 5655 21511 5661
rect 21542 5652 21548 5704
rect 21600 5692 21606 5704
rect 21709 5695 21767 5701
rect 21709 5692 21721 5695
rect 21600 5664 21721 5692
rect 21600 5652 21606 5664
rect 21709 5661 21721 5664
rect 21755 5661 21767 5695
rect 21709 5655 21767 5661
rect 15749 5627 15807 5633
rect 15749 5593 15761 5627
rect 15795 5624 15807 5627
rect 16390 5624 16396 5636
rect 15795 5596 16396 5624
rect 15795 5593 15807 5596
rect 15749 5587 15807 5593
rect 16390 5584 16396 5596
rect 16448 5584 16454 5636
rect 17218 5624 17224 5636
rect 16684 5596 17224 5624
rect 15194 5556 15200 5568
rect 14016 5528 15200 5556
rect 15194 5516 15200 5528
rect 15252 5516 15258 5568
rect 15473 5559 15531 5565
rect 15473 5525 15485 5559
rect 15519 5556 15531 5559
rect 16684 5556 16712 5596
rect 17218 5584 17224 5596
rect 17276 5584 17282 5636
rect 17948 5627 18006 5633
rect 17948 5593 17960 5627
rect 17994 5624 18006 5627
rect 18138 5624 18144 5636
rect 17994 5596 18144 5624
rect 17994 5593 18006 5596
rect 17948 5587 18006 5593
rect 18138 5584 18144 5596
rect 18196 5584 18202 5636
rect 18874 5584 18880 5636
rect 18932 5624 18938 5636
rect 20254 5624 20260 5636
rect 18932 5596 20260 5624
rect 18932 5584 18938 5596
rect 20254 5584 20260 5596
rect 20312 5584 20318 5636
rect 21024 5627 21082 5633
rect 21024 5593 21036 5627
rect 21070 5624 21082 5627
rect 21070 5596 21588 5624
rect 21070 5593 21082 5596
rect 21024 5587 21082 5593
rect 15519 5528 16712 5556
rect 15519 5525 15531 5528
rect 15473 5519 15531 5525
rect 16758 5516 16764 5568
rect 16816 5556 16822 5568
rect 17129 5559 17187 5565
rect 17129 5556 17141 5559
rect 16816 5528 17141 5556
rect 16816 5516 16822 5528
rect 17129 5525 17141 5528
rect 17175 5525 17187 5559
rect 17586 5556 17592 5568
rect 17547 5528 17592 5556
rect 17129 5519 17187 5525
rect 17586 5516 17592 5528
rect 17644 5516 17650 5568
rect 18414 5516 18420 5568
rect 18472 5556 18478 5568
rect 19061 5559 19119 5565
rect 19061 5556 19073 5559
rect 18472 5528 19073 5556
rect 18472 5516 18478 5528
rect 19061 5525 19073 5528
rect 19107 5525 19119 5559
rect 19702 5556 19708 5568
rect 19663 5528 19708 5556
rect 19061 5519 19119 5525
rect 19702 5516 19708 5528
rect 19760 5516 19766 5568
rect 21560 5556 21588 5596
rect 22094 5584 22100 5636
rect 22152 5624 22158 5636
rect 22152 5596 22876 5624
rect 22152 5584 22158 5596
rect 22370 5556 22376 5568
rect 21560 5528 22376 5556
rect 22370 5516 22376 5528
rect 22428 5516 22434 5568
rect 22848 5565 22876 5596
rect 22833 5559 22891 5565
rect 22833 5525 22845 5559
rect 22879 5525 22891 5559
rect 22833 5519 22891 5525
rect 1104 5466 23460 5488
rect 1104 5414 6548 5466
rect 6600 5414 6612 5466
rect 6664 5414 6676 5466
rect 6728 5414 6740 5466
rect 6792 5414 6804 5466
rect 6856 5414 12146 5466
rect 12198 5414 12210 5466
rect 12262 5414 12274 5466
rect 12326 5414 12338 5466
rect 12390 5414 12402 5466
rect 12454 5414 17744 5466
rect 17796 5414 17808 5466
rect 17860 5414 17872 5466
rect 17924 5414 17936 5466
rect 17988 5414 18000 5466
rect 18052 5414 23460 5466
rect 1104 5392 23460 5414
rect 3237 5355 3295 5361
rect 3237 5321 3249 5355
rect 3283 5352 3295 5355
rect 5166 5352 5172 5364
rect 3283 5324 5172 5352
rect 3283 5321 3295 5324
rect 3237 5315 3295 5321
rect 3344 5225 3372 5324
rect 5166 5312 5172 5324
rect 5224 5312 5230 5364
rect 5258 5312 5264 5364
rect 5316 5352 5322 5364
rect 6178 5352 6184 5364
rect 5316 5324 6184 5352
rect 5316 5312 5322 5324
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 6454 5312 6460 5364
rect 6512 5352 6518 5364
rect 6733 5355 6791 5361
rect 6733 5352 6745 5355
rect 6512 5324 6745 5352
rect 6512 5312 6518 5324
rect 6733 5321 6745 5324
rect 6779 5321 6791 5355
rect 6733 5315 6791 5321
rect 7101 5355 7159 5361
rect 7101 5321 7113 5355
rect 7147 5352 7159 5355
rect 7653 5355 7711 5361
rect 7653 5352 7665 5355
rect 7147 5324 7665 5352
rect 7147 5321 7159 5324
rect 7101 5315 7159 5321
rect 7653 5321 7665 5324
rect 7699 5321 7711 5355
rect 7653 5315 7711 5321
rect 7834 5312 7840 5364
rect 7892 5352 7898 5364
rect 8113 5355 8171 5361
rect 8113 5352 8125 5355
rect 7892 5324 8125 5352
rect 7892 5312 7898 5324
rect 8113 5321 8125 5324
rect 8159 5321 8171 5355
rect 8113 5315 8171 5321
rect 8481 5355 8539 5361
rect 8481 5321 8493 5355
rect 8527 5352 8539 5355
rect 8846 5352 8852 5364
rect 8527 5324 8852 5352
rect 8527 5321 8539 5324
rect 8481 5315 8539 5321
rect 8846 5312 8852 5324
rect 8904 5352 8910 5364
rect 8941 5355 8999 5361
rect 8941 5352 8953 5355
rect 8904 5324 8953 5352
rect 8904 5312 8910 5324
rect 8941 5321 8953 5324
rect 8987 5321 8999 5355
rect 10686 5352 10692 5364
rect 10647 5324 10692 5352
rect 8941 5315 8999 5321
rect 10686 5312 10692 5324
rect 10744 5312 10750 5364
rect 11974 5312 11980 5364
rect 12032 5352 12038 5364
rect 12069 5355 12127 5361
rect 12069 5352 12081 5355
rect 12032 5324 12081 5352
rect 12032 5312 12038 5324
rect 12069 5321 12081 5324
rect 12115 5321 12127 5355
rect 12069 5315 12127 5321
rect 12437 5355 12495 5361
rect 12437 5321 12449 5355
rect 12483 5352 12495 5355
rect 12618 5352 12624 5364
rect 12483 5324 12624 5352
rect 12483 5321 12495 5324
rect 12437 5315 12495 5321
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 16482 5352 16488 5364
rect 16408 5324 16488 5352
rect 5074 5293 5080 5296
rect 3973 5287 4031 5293
rect 3973 5253 3985 5287
rect 4019 5284 4031 5287
rect 5068 5284 5080 5293
rect 4019 5256 4936 5284
rect 5035 5256 5080 5284
rect 4019 5253 4031 5256
rect 3973 5247 4031 5253
rect 3329 5219 3387 5225
rect 3329 5185 3341 5219
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5216 4123 5219
rect 4614 5216 4620 5228
rect 4111 5188 4620 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 4798 5216 4804 5228
rect 4759 5188 4804 5216
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 4908 5216 4936 5256
rect 5068 5247 5080 5256
rect 5074 5244 5080 5247
rect 5132 5244 5138 5296
rect 5534 5244 5540 5296
rect 5592 5284 5598 5296
rect 6641 5287 6699 5293
rect 6641 5284 6653 5287
rect 5592 5256 6653 5284
rect 5592 5244 5598 5256
rect 6641 5253 6653 5256
rect 6687 5253 6699 5287
rect 6641 5247 6699 5253
rect 7374 5244 7380 5296
rect 7432 5284 7438 5296
rect 8573 5287 8631 5293
rect 7432 5256 8248 5284
rect 7432 5244 7438 5256
rect 4908 5188 6776 5216
rect 6362 5108 6368 5160
rect 6420 5148 6426 5160
rect 6457 5151 6515 5157
rect 6457 5148 6469 5151
rect 6420 5120 6469 5148
rect 6420 5108 6426 5120
rect 6457 5117 6469 5120
rect 6503 5117 6515 5151
rect 6748 5148 6776 5188
rect 6914 5176 6920 5228
rect 6972 5216 6978 5228
rect 7561 5219 7619 5225
rect 7561 5216 7573 5219
rect 6972 5188 7573 5216
rect 6972 5176 6978 5188
rect 7561 5185 7573 5188
rect 7607 5185 7619 5219
rect 7561 5179 7619 5185
rect 7742 5148 7748 5160
rect 6748 5120 7604 5148
rect 7703 5120 7748 5148
rect 6457 5111 6515 5117
rect 6472 5080 6500 5111
rect 7374 5080 7380 5092
rect 6472 5052 7380 5080
rect 7374 5040 7380 5052
rect 7432 5040 7438 5092
rect 4709 5015 4767 5021
rect 4709 4981 4721 5015
rect 4755 5012 4767 5015
rect 5442 5012 5448 5024
rect 4755 4984 5448 5012
rect 4755 4981 4767 4984
rect 4709 4975 4767 4981
rect 5442 4972 5448 4984
rect 5500 4972 5506 5024
rect 7098 4972 7104 5024
rect 7156 5012 7162 5024
rect 7193 5015 7251 5021
rect 7193 5012 7205 5015
rect 7156 4984 7205 5012
rect 7156 4972 7162 4984
rect 7193 4981 7205 4984
rect 7239 4981 7251 5015
rect 7576 5012 7604 5120
rect 7742 5108 7748 5120
rect 7800 5108 7806 5160
rect 8220 5148 8248 5256
rect 8573 5253 8585 5287
rect 8619 5284 8631 5287
rect 8662 5284 8668 5296
rect 8619 5256 8668 5284
rect 8619 5253 8631 5256
rect 8573 5247 8631 5253
rect 8662 5244 8668 5256
rect 8720 5244 8726 5296
rect 9674 5244 9680 5296
rect 9732 5284 9738 5296
rect 10781 5287 10839 5293
rect 10781 5284 10793 5287
rect 9732 5256 10793 5284
rect 9732 5244 9738 5256
rect 10781 5253 10793 5256
rect 10827 5253 10839 5287
rect 10781 5247 10839 5253
rect 12529 5287 12587 5293
rect 12529 5253 12541 5287
rect 12575 5284 12587 5287
rect 12802 5284 12808 5296
rect 12575 5256 12808 5284
rect 12575 5253 12587 5256
rect 12529 5247 12587 5253
rect 12802 5244 12808 5256
rect 12860 5244 12866 5296
rect 12986 5284 12992 5296
rect 12947 5256 12992 5284
rect 12986 5244 12992 5256
rect 13044 5244 13050 5296
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 10054 5219 10112 5225
rect 10054 5216 10066 5219
rect 8352 5188 10066 5216
rect 8352 5176 8358 5188
rect 10054 5185 10066 5188
rect 10100 5185 10112 5219
rect 10318 5216 10324 5228
rect 10279 5188 10324 5216
rect 10054 5179 10112 5185
rect 10318 5176 10324 5188
rect 10376 5176 10382 5228
rect 11330 5176 11336 5228
rect 11388 5216 11394 5228
rect 11517 5219 11575 5225
rect 11517 5216 11529 5219
rect 11388 5188 11529 5216
rect 11388 5176 11394 5188
rect 11517 5185 11529 5188
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 15953 5219 16011 5225
rect 15953 5185 15965 5219
rect 15999 5216 16011 5219
rect 16114 5216 16120 5228
rect 15999 5188 16120 5216
rect 15999 5185 16011 5188
rect 15953 5179 16011 5185
rect 16114 5176 16120 5188
rect 16172 5176 16178 5228
rect 16301 5220 16359 5225
rect 16408 5220 16436 5324
rect 16482 5312 16488 5324
rect 16540 5312 16546 5364
rect 16574 5312 16580 5364
rect 16632 5352 16638 5364
rect 16945 5355 17003 5361
rect 16945 5352 16957 5355
rect 16632 5324 16957 5352
rect 16632 5312 16638 5324
rect 16945 5321 16957 5324
rect 16991 5321 17003 5355
rect 16945 5315 17003 5321
rect 17034 5312 17040 5364
rect 17092 5352 17098 5364
rect 17405 5355 17463 5361
rect 17405 5352 17417 5355
rect 17092 5324 17417 5352
rect 17092 5312 17098 5324
rect 17405 5321 17417 5324
rect 17451 5321 17463 5355
rect 17405 5315 17463 5321
rect 17586 5312 17592 5364
rect 17644 5352 17650 5364
rect 17773 5355 17831 5361
rect 17773 5352 17785 5355
rect 17644 5324 17785 5352
rect 17644 5312 17650 5324
rect 17773 5321 17785 5324
rect 17819 5321 17831 5355
rect 18598 5352 18604 5364
rect 18559 5324 18604 5352
rect 17773 5315 17831 5321
rect 18598 5312 18604 5324
rect 18656 5312 18662 5364
rect 18874 5312 18880 5364
rect 18932 5352 18938 5364
rect 19334 5352 19340 5364
rect 18932 5324 19340 5352
rect 18932 5312 18938 5324
rect 19334 5312 19340 5324
rect 19392 5312 19398 5364
rect 19429 5355 19487 5361
rect 19429 5321 19441 5355
rect 19475 5321 19487 5355
rect 20254 5352 20260 5364
rect 20215 5324 20260 5352
rect 19429 5315 19487 5321
rect 19444 5284 19472 5315
rect 20254 5312 20260 5324
rect 20312 5312 20318 5364
rect 20993 5355 21051 5361
rect 20993 5321 21005 5355
rect 21039 5352 21051 5355
rect 21818 5352 21824 5364
rect 21039 5324 21824 5352
rect 21039 5321 21051 5324
rect 20993 5315 21051 5321
rect 21818 5312 21824 5324
rect 21876 5312 21882 5364
rect 22186 5352 22192 5364
rect 22147 5324 22192 5352
rect 22186 5312 22192 5324
rect 22244 5312 22250 5364
rect 18340 5256 19472 5284
rect 16301 5219 16436 5220
rect 16301 5185 16313 5219
rect 16347 5192 16436 5219
rect 16347 5185 16359 5192
rect 16301 5179 16359 5185
rect 16942 5176 16948 5228
rect 17000 5216 17006 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 17000 5188 17049 5216
rect 17000 5176 17006 5188
rect 17037 5185 17049 5188
rect 17083 5185 17095 5219
rect 17037 5179 17095 5185
rect 17678 5176 17684 5228
rect 17736 5216 17742 5228
rect 18340 5225 18368 5256
rect 19518 5244 19524 5296
rect 19576 5284 19582 5296
rect 19576 5256 20944 5284
rect 19576 5244 19582 5256
rect 17865 5219 17923 5225
rect 17865 5216 17877 5219
rect 17736 5188 17877 5216
rect 17736 5176 17742 5188
rect 17865 5185 17877 5188
rect 17911 5185 17923 5219
rect 17865 5179 17923 5185
rect 18325 5219 18383 5225
rect 18325 5185 18337 5219
rect 18371 5185 18383 5219
rect 18966 5216 18972 5228
rect 18927 5188 18972 5216
rect 18325 5179 18383 5185
rect 18966 5176 18972 5188
rect 19024 5176 19030 5228
rect 19426 5176 19432 5228
rect 19484 5216 19490 5228
rect 20916 5225 20944 5256
rect 21726 5244 21732 5296
rect 21784 5284 21790 5296
rect 22281 5287 22339 5293
rect 22281 5284 22293 5287
rect 21784 5256 22293 5284
rect 21784 5244 21790 5256
rect 22281 5253 22293 5256
rect 22327 5253 22339 5287
rect 22281 5247 22339 5253
rect 22649 5287 22707 5293
rect 22649 5253 22661 5287
rect 22695 5284 22707 5287
rect 23198 5284 23204 5296
rect 22695 5256 23204 5284
rect 22695 5253 22707 5256
rect 22649 5247 22707 5253
rect 23198 5244 23204 5256
rect 23256 5244 23262 5296
rect 19797 5219 19855 5225
rect 19797 5216 19809 5219
rect 19484 5188 19809 5216
rect 19484 5176 19490 5188
rect 19797 5185 19809 5188
rect 19843 5185 19855 5219
rect 19797 5179 19855 5185
rect 20901 5219 20959 5225
rect 20901 5185 20913 5219
rect 20947 5185 20959 5219
rect 21634 5216 21640 5228
rect 21595 5188 21640 5216
rect 20901 5179 20959 5185
rect 21634 5176 21640 5188
rect 21692 5176 21698 5228
rect 22830 5216 22836 5228
rect 22791 5188 22836 5216
rect 22830 5176 22836 5188
rect 22888 5176 22894 5228
rect 8665 5151 8723 5157
rect 8665 5148 8677 5151
rect 8220 5120 8677 5148
rect 8665 5117 8677 5120
rect 8711 5148 8723 5151
rect 9214 5148 9220 5160
rect 8711 5120 9220 5148
rect 8711 5117 8723 5120
rect 8665 5111 8723 5117
rect 9214 5108 9220 5120
rect 9272 5108 9278 5160
rect 10502 5148 10508 5160
rect 10463 5120 10508 5148
rect 10502 5108 10508 5120
rect 10560 5108 10566 5160
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5148 12035 5151
rect 12618 5148 12624 5160
rect 12023 5120 12624 5148
rect 12023 5117 12035 5120
rect 11977 5111 12035 5117
rect 12618 5108 12624 5120
rect 12676 5108 12682 5160
rect 12713 5151 12771 5157
rect 12713 5117 12725 5151
rect 12759 5148 12771 5151
rect 14734 5148 14740 5160
rect 12759 5120 14596 5148
rect 14695 5120 14740 5148
rect 12759 5117 12771 5120
rect 12713 5111 12771 5117
rect 14458 5080 14464 5092
rect 11072 5052 14464 5080
rect 11072 5012 11100 5052
rect 14458 5040 14464 5052
rect 14516 5040 14522 5092
rect 14568 5080 14596 5120
rect 14734 5108 14740 5120
rect 14792 5108 14798 5160
rect 16209 5151 16267 5157
rect 16209 5117 16221 5151
rect 16255 5148 16267 5151
rect 16390 5148 16396 5160
rect 16255 5120 16396 5148
rect 16255 5117 16267 5120
rect 16209 5111 16267 5117
rect 16390 5108 16396 5120
rect 16448 5108 16454 5160
rect 16853 5151 16911 5157
rect 16853 5117 16865 5151
rect 16899 5148 16911 5151
rect 17310 5148 17316 5160
rect 16899 5120 17316 5148
rect 16899 5117 16911 5120
rect 16853 5111 16911 5117
rect 17310 5108 17316 5120
rect 17368 5108 17374 5160
rect 17586 5148 17592 5160
rect 17547 5120 17592 5148
rect 17586 5108 17592 5120
rect 17644 5108 17650 5160
rect 19061 5151 19119 5157
rect 19061 5148 19073 5151
rect 18524 5120 19073 5148
rect 16485 5083 16543 5089
rect 14568 5052 14872 5080
rect 7576 4984 11100 5012
rect 11149 5015 11207 5021
rect 7193 4975 7251 4981
rect 11149 4981 11161 5015
rect 11195 5012 11207 5015
rect 11422 5012 11428 5024
rect 11195 4984 11428 5012
rect 11195 4981 11207 4984
rect 11149 4975 11207 4981
rect 11422 4972 11428 4984
rect 11480 4972 11486 5024
rect 11701 5015 11759 5021
rect 11701 4981 11713 5015
rect 11747 5012 11759 5015
rect 13262 5012 13268 5024
rect 11747 4984 13268 5012
rect 11747 4981 11759 4984
rect 11701 4975 11759 4981
rect 13262 4972 13268 4984
rect 13320 5012 13326 5024
rect 13446 5012 13452 5024
rect 13320 4984 13452 5012
rect 13320 4972 13326 4984
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 14844 5021 14872 5052
rect 16485 5049 16497 5083
rect 16531 5080 16543 5083
rect 17604 5080 17632 5108
rect 18524 5089 18552 5120
rect 19061 5117 19073 5120
rect 19107 5117 19119 5151
rect 19061 5111 19119 5117
rect 19153 5151 19211 5157
rect 19153 5117 19165 5151
rect 19199 5117 19211 5151
rect 19153 5111 19211 5117
rect 19889 5151 19947 5157
rect 19889 5117 19901 5151
rect 19935 5117 19947 5151
rect 19889 5111 19947 5117
rect 20073 5151 20131 5157
rect 20073 5117 20085 5151
rect 20119 5148 20131 5151
rect 21818 5148 21824 5160
rect 20119 5120 21824 5148
rect 20119 5117 20131 5120
rect 20073 5111 20131 5117
rect 16531 5052 17632 5080
rect 18509 5083 18567 5089
rect 16531 5049 16543 5052
rect 16485 5043 16543 5049
rect 18509 5049 18521 5083
rect 18555 5049 18567 5083
rect 18509 5043 18567 5049
rect 18782 5040 18788 5092
rect 18840 5080 18846 5092
rect 19168 5080 19196 5111
rect 19242 5080 19248 5092
rect 18840 5052 19248 5080
rect 18840 5040 18846 5052
rect 19242 5040 19248 5052
rect 19300 5080 19306 5092
rect 19794 5080 19800 5092
rect 19300 5052 19800 5080
rect 19300 5040 19306 5052
rect 19794 5040 19800 5052
rect 19852 5040 19858 5092
rect 19904 5024 19932 5111
rect 21818 5108 21824 5120
rect 21876 5108 21882 5160
rect 22278 5108 22284 5160
rect 22336 5148 22342 5160
rect 22373 5151 22431 5157
rect 22373 5148 22385 5151
rect 22336 5120 22385 5148
rect 22336 5108 22342 5120
rect 22373 5117 22385 5120
rect 22419 5117 22431 5151
rect 22373 5111 22431 5117
rect 19978 5040 19984 5092
rect 20036 5080 20042 5092
rect 21726 5080 21732 5092
rect 20036 5052 21732 5080
rect 20036 5040 20042 5052
rect 21726 5040 21732 5052
rect 21784 5040 21790 5092
rect 14829 5015 14887 5021
rect 14829 4981 14841 5015
rect 14875 5012 14887 5015
rect 17494 5012 17500 5024
rect 14875 4984 17500 5012
rect 14875 4981 14887 4984
rect 14829 4975 14887 4981
rect 17494 4972 17500 4984
rect 17552 4972 17558 5024
rect 18233 5015 18291 5021
rect 18233 4981 18245 5015
rect 18279 5012 18291 5015
rect 19886 5012 19892 5024
rect 18279 4984 19892 5012
rect 18279 4981 18291 4984
rect 18233 4975 18291 4981
rect 19886 4972 19892 4984
rect 19944 4972 19950 5024
rect 21634 4972 21640 5024
rect 21692 5012 21698 5024
rect 21821 5015 21879 5021
rect 21821 5012 21833 5015
rect 21692 4984 21833 5012
rect 21692 4972 21698 4984
rect 21821 4981 21833 4984
rect 21867 4981 21879 5015
rect 21821 4975 21879 4981
rect 23017 5015 23075 5021
rect 23017 4981 23029 5015
rect 23063 5012 23075 5015
rect 23106 5012 23112 5024
rect 23063 4984 23112 5012
rect 23063 4981 23075 4984
rect 23017 4975 23075 4981
rect 23106 4972 23112 4984
rect 23164 4972 23170 5024
rect 1104 4922 23460 4944
rect 1104 4870 3749 4922
rect 3801 4870 3813 4922
rect 3865 4870 3877 4922
rect 3929 4870 3941 4922
rect 3993 4870 4005 4922
rect 4057 4870 9347 4922
rect 9399 4870 9411 4922
rect 9463 4870 9475 4922
rect 9527 4870 9539 4922
rect 9591 4870 9603 4922
rect 9655 4870 14945 4922
rect 14997 4870 15009 4922
rect 15061 4870 15073 4922
rect 15125 4870 15137 4922
rect 15189 4870 15201 4922
rect 15253 4870 20543 4922
rect 20595 4870 20607 4922
rect 20659 4870 20671 4922
rect 20723 4870 20735 4922
rect 20787 4870 20799 4922
rect 20851 4870 23460 4922
rect 1104 4848 23460 4870
rect 3881 4811 3939 4817
rect 3881 4777 3893 4811
rect 3927 4808 3939 4811
rect 4154 4808 4160 4820
rect 3927 4780 4160 4808
rect 3927 4777 3939 4780
rect 3881 4771 3939 4777
rect 2866 4604 2872 4616
rect 2827 4576 2872 4604
rect 2866 4564 2872 4576
rect 2924 4564 2930 4616
rect 3605 4607 3663 4613
rect 3605 4573 3617 4607
rect 3651 4604 3663 4607
rect 3896 4604 3924 4771
rect 4154 4768 4160 4780
rect 4212 4768 4218 4820
rect 5445 4811 5503 4817
rect 5445 4777 5457 4811
rect 5491 4808 5503 4811
rect 5810 4808 5816 4820
rect 5491 4780 5816 4808
rect 5491 4777 5503 4780
rect 5445 4771 5503 4777
rect 5810 4768 5816 4780
rect 5868 4768 5874 4820
rect 6178 4768 6184 4820
rect 6236 4808 6242 4820
rect 6546 4808 6552 4820
rect 6236 4780 6552 4808
rect 6236 4768 6242 4780
rect 6546 4768 6552 4780
rect 6604 4768 6610 4820
rect 6914 4768 6920 4820
rect 6972 4808 6978 4820
rect 6972 4780 7017 4808
rect 6972 4768 6978 4780
rect 7466 4768 7472 4820
rect 7524 4808 7530 4820
rect 8113 4811 8171 4817
rect 8113 4808 8125 4811
rect 7524 4780 8125 4808
rect 7524 4768 7530 4780
rect 8113 4777 8125 4780
rect 8159 4777 8171 4811
rect 9858 4808 9864 4820
rect 8113 4771 8171 4777
rect 8404 4780 9864 4808
rect 4709 4743 4767 4749
rect 4709 4709 4721 4743
rect 4755 4740 4767 4743
rect 4755 4712 7604 4740
rect 4755 4709 4767 4712
rect 4709 4703 4767 4709
rect 6362 4672 6368 4684
rect 6323 4644 6368 4672
rect 6362 4632 6368 4644
rect 6420 4632 6426 4684
rect 3651 4576 3924 4604
rect 4617 4607 4675 4613
rect 3651 4573 3663 4576
rect 3605 4567 3663 4573
rect 4617 4573 4629 4607
rect 4663 4573 4675 4607
rect 5350 4604 5356 4616
rect 5311 4576 5356 4604
rect 4617 4567 4675 4573
rect 2958 4536 2964 4548
rect 2919 4508 2964 4536
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 4632 4536 4660 4567
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 6089 4607 6147 4613
rect 6089 4573 6101 4607
rect 6135 4604 6147 4607
rect 6454 4604 6460 4616
rect 6135 4576 6460 4604
rect 6135 4573 6147 4576
rect 6089 4567 6147 4573
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 6604 4576 6649 4604
rect 6604 4564 6610 4576
rect 6178 4536 6184 4548
rect 4632 4508 6184 4536
rect 6178 4496 6184 4508
rect 6236 4496 6242 4548
rect 7190 4496 7196 4548
rect 7248 4536 7254 4548
rect 7469 4539 7527 4545
rect 7469 4536 7481 4539
rect 7248 4508 7481 4536
rect 7248 4496 7254 4508
rect 7469 4505 7481 4508
rect 7515 4505 7527 4539
rect 7576 4536 7604 4712
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4672 7711 4675
rect 8404 4672 8432 4780
rect 9858 4768 9864 4780
rect 9916 4768 9922 4820
rect 10410 4808 10416 4820
rect 10371 4780 10416 4808
rect 10410 4768 10416 4780
rect 10468 4768 10474 4820
rect 10594 4808 10600 4820
rect 10555 4780 10600 4808
rect 10594 4768 10600 4780
rect 10652 4768 10658 4820
rect 10965 4811 11023 4817
rect 10965 4808 10977 4811
rect 10796 4780 10977 4808
rect 10226 4740 10232 4752
rect 8772 4712 10232 4740
rect 8772 4672 8800 4712
rect 10226 4700 10232 4712
rect 10284 4700 10290 4752
rect 7699 4644 8432 4672
rect 8680 4644 8800 4672
rect 9125 4675 9183 4681
rect 7699 4641 7711 4644
rect 7653 4635 7711 4641
rect 7834 4604 7840 4616
rect 7795 4576 7840 4604
rect 7834 4564 7840 4576
rect 7892 4564 7898 4616
rect 8680 4604 8708 4644
rect 9125 4641 9137 4675
rect 9171 4672 9183 4675
rect 10502 4672 10508 4684
rect 9171 4644 10508 4672
rect 9171 4641 9183 4644
rect 9125 4635 9183 4641
rect 10502 4632 10508 4644
rect 10560 4632 10566 4684
rect 10796 4672 10824 4780
rect 10965 4777 10977 4780
rect 11011 4777 11023 4811
rect 10965 4771 11023 4777
rect 11790 4768 11796 4820
rect 11848 4808 11854 4820
rect 12253 4811 12311 4817
rect 12253 4808 12265 4811
rect 11848 4780 12265 4808
rect 11848 4768 11854 4780
rect 10873 4743 10931 4749
rect 10873 4709 10885 4743
rect 10919 4740 10931 4743
rect 10919 4712 11560 4740
rect 10919 4709 10931 4712
rect 10873 4703 10931 4709
rect 11532 4681 11560 4712
rect 10612 4644 10824 4672
rect 11517 4675 11575 4681
rect 7944 4576 8708 4604
rect 8757 4607 8815 4613
rect 7944 4536 7972 4576
rect 8757 4573 8769 4607
rect 8803 4604 8815 4607
rect 8846 4604 8852 4616
rect 8803 4576 8852 4604
rect 8803 4573 8815 4576
rect 8757 4567 8815 4573
rect 8846 4564 8852 4576
rect 8904 4564 8910 4616
rect 9214 4564 9220 4616
rect 9272 4604 9278 4616
rect 9766 4604 9772 4616
rect 9272 4576 9444 4604
rect 9727 4576 9772 4604
rect 9272 4564 9278 4576
rect 9309 4539 9367 4545
rect 9309 4536 9321 4539
rect 7576 4508 7972 4536
rect 8036 4508 9321 4536
rect 7469 4499 7527 4505
rect 2222 4468 2228 4480
rect 2183 4440 2228 4468
rect 2222 4428 2228 4440
rect 2280 4428 2286 4480
rect 3973 4471 4031 4477
rect 3973 4437 3985 4471
rect 4019 4468 4031 4471
rect 5074 4468 5080 4480
rect 4019 4440 5080 4468
rect 4019 4437 4031 4440
rect 3973 4431 4031 4437
rect 5074 4428 5080 4440
rect 5132 4428 5138 4480
rect 6270 4428 6276 4480
rect 6328 4468 6334 4480
rect 6457 4471 6515 4477
rect 6457 4468 6469 4471
rect 6328 4440 6469 4468
rect 6328 4428 6334 4440
rect 6457 4437 6469 4440
rect 6503 4437 6515 4471
rect 6457 4431 6515 4437
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 7374 4468 7380 4480
rect 7064 4440 7109 4468
rect 7335 4440 7380 4468
rect 7064 4428 7070 4440
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 8036 4477 8064 4508
rect 9309 4505 9321 4508
rect 9355 4505 9367 4539
rect 9416 4536 9444 4576
rect 9766 4564 9772 4576
rect 9824 4564 9830 4616
rect 10612 4536 10640 4644
rect 11517 4641 11529 4675
rect 11563 4641 11575 4675
rect 11517 4635 11575 4641
rect 12176 4613 12204 4780
rect 12253 4777 12265 4780
rect 12299 4777 12311 4811
rect 12253 4771 12311 4777
rect 14829 4811 14887 4817
rect 14829 4777 14841 4811
rect 14875 4808 14887 4811
rect 16482 4808 16488 4820
rect 14875 4780 16488 4808
rect 14875 4777 14887 4780
rect 14829 4771 14887 4777
rect 16482 4768 16488 4780
rect 16540 4768 16546 4820
rect 18046 4808 18052 4820
rect 18007 4780 18052 4808
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 18874 4768 18880 4820
rect 18932 4808 18938 4820
rect 19061 4811 19119 4817
rect 19061 4808 19073 4811
rect 18932 4780 19073 4808
rect 18932 4768 18938 4780
rect 19061 4777 19073 4780
rect 19107 4777 19119 4811
rect 19242 4808 19248 4820
rect 19203 4780 19248 4808
rect 19061 4771 19119 4777
rect 19242 4768 19248 4780
rect 19300 4768 19306 4820
rect 19426 4808 19432 4820
rect 19387 4780 19432 4808
rect 19426 4768 19432 4780
rect 19484 4768 19490 4820
rect 19518 4768 19524 4820
rect 19576 4808 19582 4820
rect 21542 4808 21548 4820
rect 19576 4780 20760 4808
rect 21503 4780 21548 4808
rect 19576 4768 19582 4780
rect 15010 4740 15016 4752
rect 14971 4712 15016 4740
rect 15010 4700 15016 4712
rect 15068 4700 15074 4752
rect 17126 4740 17132 4752
rect 16776 4712 17132 4740
rect 14277 4675 14335 4681
rect 14277 4641 14289 4675
rect 14323 4672 14335 4675
rect 15470 4672 15476 4684
rect 14323 4644 15476 4672
rect 14323 4641 14335 4644
rect 14277 4635 14335 4641
rect 15470 4632 15476 4644
rect 15528 4632 15534 4684
rect 16776 4681 16804 4712
rect 17126 4700 17132 4712
rect 17184 4740 17190 4752
rect 18230 4740 18236 4752
rect 17184 4712 18236 4740
rect 17184 4700 17190 4712
rect 18230 4700 18236 4712
rect 18288 4700 18294 4752
rect 18966 4700 18972 4752
rect 19024 4740 19030 4752
rect 20257 4743 20315 4749
rect 20257 4740 20269 4743
rect 19024 4712 20269 4740
rect 19024 4700 19030 4712
rect 20257 4709 20269 4712
rect 20303 4709 20315 4743
rect 20257 4703 20315 4709
rect 16761 4675 16819 4681
rect 16761 4641 16773 4675
rect 16807 4641 16819 4675
rect 16761 4635 16819 4641
rect 16942 4632 16948 4684
rect 17000 4672 17006 4684
rect 17000 4644 17540 4672
rect 17000 4632 17006 4644
rect 10689 4607 10747 4613
rect 10689 4573 10701 4607
rect 10735 4604 10747 4607
rect 11793 4607 11851 4613
rect 11793 4604 11805 4607
rect 10735 4576 11805 4604
rect 10735 4573 10747 4576
rect 10689 4567 10747 4573
rect 11793 4573 11805 4576
rect 11839 4573 11851 4607
rect 11793 4567 11851 4573
rect 12161 4607 12219 4613
rect 12161 4573 12173 4607
rect 12207 4573 12219 4607
rect 12161 4567 12219 4573
rect 12526 4564 12532 4616
rect 12584 4604 12590 4616
rect 13081 4607 13139 4613
rect 13081 4604 13093 4607
rect 12584 4576 13093 4604
rect 12584 4564 12590 4576
rect 13081 4573 13093 4576
rect 13127 4573 13139 4607
rect 13081 4567 13139 4573
rect 13909 4607 13967 4613
rect 13909 4573 13921 4607
rect 13955 4604 13967 4607
rect 13955 4576 15148 4604
rect 13955 4573 13967 4576
rect 13909 4567 13967 4573
rect 9416 4508 10640 4536
rect 9309 4499 9367 4505
rect 11054 4496 11060 4548
rect 11112 4536 11118 4548
rect 11977 4539 12035 4545
rect 11977 4536 11989 4539
rect 11112 4508 11989 4536
rect 11112 4496 11118 4508
rect 11977 4505 11989 4508
rect 12023 4505 12035 4539
rect 11977 4499 12035 4505
rect 13446 4496 13452 4548
rect 13504 4536 13510 4548
rect 14461 4539 14519 4545
rect 14461 4536 14473 4539
rect 13504 4508 14473 4536
rect 13504 4496 13510 4508
rect 14461 4505 14473 4508
rect 14507 4505 14519 4539
rect 14461 4499 14519 4505
rect 8021 4471 8079 4477
rect 8021 4437 8033 4471
rect 8067 4437 8079 4471
rect 8021 4431 8079 4437
rect 8386 4428 8392 4480
rect 8444 4468 8450 4480
rect 9217 4471 9275 4477
rect 9217 4468 9229 4471
rect 8444 4440 9229 4468
rect 8444 4428 8450 4440
rect 9217 4437 9229 4440
rect 9263 4437 9275 4471
rect 9217 4431 9275 4437
rect 9677 4471 9735 4477
rect 9677 4437 9689 4471
rect 9723 4468 9735 4471
rect 11330 4468 11336 4480
rect 9723 4440 11336 4468
rect 9723 4437 9735 4440
rect 9677 4431 9735 4437
rect 11330 4428 11336 4440
rect 11388 4428 11394 4480
rect 11422 4428 11428 4480
rect 11480 4468 11486 4480
rect 12437 4471 12495 4477
rect 11480 4440 11525 4468
rect 11480 4428 11486 4440
rect 12437 4437 12449 4471
rect 12483 4468 12495 4471
rect 12618 4468 12624 4480
rect 12483 4440 12624 4468
rect 12483 4437 12495 4440
rect 12437 4431 12495 4437
rect 12618 4428 12624 4440
rect 12676 4428 12682 4480
rect 13265 4471 13323 4477
rect 13265 4437 13277 4471
rect 13311 4468 13323 4471
rect 14274 4468 14280 4480
rect 13311 4440 14280 4468
rect 13311 4437 13323 4440
rect 13265 4431 13323 4437
rect 14274 4428 14280 4440
rect 14332 4428 14338 4480
rect 14369 4471 14427 4477
rect 14369 4437 14381 4471
rect 14415 4468 14427 4471
rect 14642 4468 14648 4480
rect 14415 4440 14648 4468
rect 14415 4437 14427 4440
rect 14369 4431 14427 4437
rect 14642 4428 14648 4440
rect 14700 4428 14706 4480
rect 15120 4477 15148 4576
rect 16390 4564 16396 4616
rect 16448 4604 16454 4616
rect 16485 4607 16543 4613
rect 16485 4604 16497 4607
rect 16448 4576 16497 4604
rect 16448 4564 16454 4576
rect 16485 4573 16497 4576
rect 16531 4573 16543 4607
rect 16485 4567 16543 4573
rect 17218 4564 17224 4616
rect 17276 4604 17282 4616
rect 17405 4607 17463 4613
rect 17405 4604 17417 4607
rect 17276 4576 17417 4604
rect 17276 4564 17282 4576
rect 17405 4573 17417 4576
rect 17451 4573 17463 4607
rect 17512 4604 17540 4644
rect 17586 4632 17592 4684
rect 17644 4672 17650 4684
rect 20732 4681 20760 4780
rect 21542 4768 21548 4780
rect 21600 4768 21606 4820
rect 19981 4675 20039 4681
rect 19981 4672 19993 4675
rect 17644 4644 19993 4672
rect 17644 4632 17650 4644
rect 19981 4641 19993 4644
rect 20027 4641 20039 4675
rect 19981 4635 20039 4641
rect 20717 4675 20775 4681
rect 20717 4641 20729 4675
rect 20763 4672 20775 4675
rect 21082 4672 21088 4684
rect 20763 4644 21088 4672
rect 20763 4641 20775 4644
rect 20717 4635 20775 4641
rect 21082 4632 21088 4644
rect 21140 4632 21146 4684
rect 21174 4632 21180 4684
rect 21232 4672 21238 4684
rect 21729 4675 21787 4681
rect 21729 4672 21741 4675
rect 21232 4644 21741 4672
rect 21232 4632 21238 4644
rect 21729 4641 21741 4644
rect 21775 4641 21787 4675
rect 21729 4635 21787 4641
rect 18141 4607 18199 4613
rect 18141 4604 18153 4607
rect 17512 4576 18153 4604
rect 17405 4567 17463 4573
rect 18141 4573 18153 4576
rect 18187 4573 18199 4607
rect 18141 4567 18199 4573
rect 18877 4607 18935 4613
rect 18877 4573 18889 4607
rect 18923 4604 18935 4607
rect 19426 4604 19432 4616
rect 18923 4576 19432 4604
rect 18923 4573 18935 4576
rect 18877 4567 18935 4573
rect 19426 4564 19432 4576
rect 19484 4564 19490 4616
rect 19886 4564 19892 4616
rect 19944 4604 19950 4616
rect 20441 4607 20499 4613
rect 20441 4604 20453 4607
rect 19944 4576 20453 4604
rect 19944 4564 19950 4576
rect 20441 4573 20453 4576
rect 20487 4573 20499 4607
rect 20441 4567 20499 4573
rect 20809 4607 20867 4613
rect 20809 4573 20821 4607
rect 20855 4604 20867 4607
rect 20898 4604 20904 4616
rect 20855 4576 20904 4604
rect 20855 4573 20867 4576
rect 20809 4567 20867 4573
rect 20898 4564 20904 4576
rect 20956 4564 20962 4616
rect 21266 4564 21272 4616
rect 21324 4604 21330 4616
rect 21361 4607 21419 4613
rect 21361 4604 21373 4607
rect 21324 4576 21373 4604
rect 21324 4564 21330 4576
rect 21361 4573 21373 4576
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 21450 4564 21456 4616
rect 21508 4604 21514 4616
rect 21985 4607 22043 4613
rect 21985 4604 21997 4607
rect 21508 4576 21997 4604
rect 21508 4564 21514 4576
rect 21985 4573 21997 4576
rect 22031 4573 22043 4607
rect 21985 4567 22043 4573
rect 16240 4539 16298 4545
rect 16240 4505 16252 4539
rect 16286 4536 16298 4539
rect 18785 4539 18843 4545
rect 18785 4536 18797 4539
rect 16286 4508 18797 4536
rect 16286 4505 16298 4508
rect 16240 4499 16298 4505
rect 18785 4505 18797 4508
rect 18831 4505 18843 4539
rect 21082 4536 21088 4548
rect 18785 4499 18843 4505
rect 19904 4508 21088 4536
rect 15105 4471 15163 4477
rect 15105 4437 15117 4471
rect 15151 4468 15163 4471
rect 16574 4468 16580 4480
rect 15151 4440 16580 4468
rect 15151 4437 15163 4440
rect 15105 4431 15163 4437
rect 16574 4428 16580 4440
rect 16632 4428 16638 4480
rect 16850 4468 16856 4480
rect 16811 4440 16856 4468
rect 16850 4428 16856 4440
rect 16908 4428 16914 4480
rect 16942 4428 16948 4480
rect 17000 4468 17006 4480
rect 17313 4471 17371 4477
rect 17000 4440 17045 4468
rect 17000 4428 17006 4440
rect 17313 4437 17325 4471
rect 17359 4468 17371 4471
rect 17494 4468 17500 4480
rect 17359 4440 17500 4468
rect 17359 4437 17371 4440
rect 17313 4431 17371 4437
rect 17494 4428 17500 4440
rect 17552 4428 17558 4480
rect 18230 4428 18236 4480
rect 18288 4468 18294 4480
rect 19518 4468 19524 4480
rect 18288 4440 19524 4468
rect 18288 4428 18294 4440
rect 19518 4428 19524 4440
rect 19576 4428 19582 4480
rect 19794 4468 19800 4480
rect 19755 4440 19800 4468
rect 19794 4428 19800 4440
rect 19852 4428 19858 4480
rect 19904 4477 19932 4508
rect 21082 4496 21088 4508
rect 21140 4496 21146 4548
rect 21284 4508 21680 4536
rect 19889 4471 19947 4477
rect 19889 4437 19901 4471
rect 19935 4437 19947 4471
rect 19889 4431 19947 4437
rect 20901 4471 20959 4477
rect 20901 4437 20913 4471
rect 20947 4468 20959 4471
rect 20990 4468 20996 4480
rect 20947 4440 20996 4468
rect 20947 4437 20959 4440
rect 20901 4431 20959 4437
rect 20990 4428 20996 4440
rect 21048 4428 21054 4480
rect 21284 4477 21312 4508
rect 21269 4471 21327 4477
rect 21269 4437 21281 4471
rect 21315 4437 21327 4471
rect 21652 4468 21680 4508
rect 21726 4496 21732 4548
rect 21784 4536 21790 4548
rect 21784 4508 23152 4536
rect 21784 4496 21790 4508
rect 23014 4468 23020 4480
rect 21652 4440 23020 4468
rect 21269 4431 21327 4437
rect 23014 4428 23020 4440
rect 23072 4428 23078 4480
rect 23124 4477 23152 4508
rect 23109 4471 23167 4477
rect 23109 4437 23121 4471
rect 23155 4437 23167 4471
rect 23109 4431 23167 4437
rect 1104 4378 23460 4400
rect 1104 4326 6548 4378
rect 6600 4326 6612 4378
rect 6664 4326 6676 4378
rect 6728 4326 6740 4378
rect 6792 4326 6804 4378
rect 6856 4326 12146 4378
rect 12198 4326 12210 4378
rect 12262 4326 12274 4378
rect 12326 4326 12338 4378
rect 12390 4326 12402 4378
rect 12454 4326 17744 4378
rect 17796 4326 17808 4378
rect 17860 4326 17872 4378
rect 17924 4326 17936 4378
rect 17988 4326 18000 4378
rect 18052 4326 23460 4378
rect 1104 4304 23460 4326
rect 2866 4224 2872 4276
rect 2924 4264 2930 4276
rect 2961 4267 3019 4273
rect 2961 4264 2973 4267
rect 2924 4236 2973 4264
rect 2924 4224 2930 4236
rect 2961 4233 2973 4236
rect 3007 4233 3019 4267
rect 2961 4227 3019 4233
rect 5166 4224 5172 4276
rect 5224 4264 5230 4276
rect 6917 4267 6975 4273
rect 5224 4236 5304 4264
rect 5224 4224 5230 4236
rect 5046 4199 5104 4205
rect 5046 4196 5058 4199
rect 4632 4168 5058 4196
rect 3329 4131 3387 4137
rect 3329 4097 3341 4131
rect 3375 4097 3387 4131
rect 3329 4091 3387 4097
rect 3237 3927 3295 3933
rect 3237 3893 3249 3927
rect 3283 3924 3295 3927
rect 3344 3924 3372 4091
rect 4522 4088 4528 4140
rect 4580 4128 4586 4140
rect 4632 4128 4660 4168
rect 5046 4165 5058 4168
rect 5092 4165 5104 4199
rect 5276 4196 5304 4236
rect 6917 4233 6929 4267
rect 6963 4264 6975 4267
rect 7006 4264 7012 4276
rect 6963 4236 7012 4264
rect 6963 4233 6975 4236
rect 6917 4227 6975 4233
rect 7006 4224 7012 4236
rect 7064 4224 7070 4276
rect 7282 4264 7288 4276
rect 7243 4236 7288 4264
rect 7282 4224 7288 4236
rect 7340 4224 7346 4276
rect 7745 4267 7803 4273
rect 7745 4233 7757 4267
rect 7791 4264 7803 4267
rect 7834 4264 7840 4276
rect 7791 4236 7840 4264
rect 7791 4233 7803 4236
rect 7745 4227 7803 4233
rect 7834 4224 7840 4236
rect 7892 4224 7898 4276
rect 8938 4264 8944 4276
rect 8036 4236 8944 4264
rect 8036 4196 8064 4236
rect 8938 4224 8944 4236
rect 8996 4224 9002 4276
rect 10229 4267 10287 4273
rect 10229 4233 10241 4267
rect 10275 4264 10287 4267
rect 10965 4267 11023 4273
rect 10965 4264 10977 4267
rect 10275 4236 10977 4264
rect 10275 4233 10287 4236
rect 10229 4227 10287 4233
rect 10965 4233 10977 4236
rect 11011 4233 11023 4267
rect 10965 4227 11023 4233
rect 12802 4224 12808 4276
rect 12860 4264 12866 4276
rect 13446 4264 13452 4276
rect 12860 4236 13452 4264
rect 12860 4224 12866 4236
rect 13446 4224 13452 4236
rect 13504 4224 13510 4276
rect 16669 4267 16727 4273
rect 16669 4233 16681 4267
rect 16715 4264 16727 4267
rect 16850 4264 16856 4276
rect 16715 4236 16856 4264
rect 16715 4233 16727 4236
rect 16669 4227 16727 4233
rect 16850 4224 16856 4236
rect 16908 4224 16914 4276
rect 17037 4267 17095 4273
rect 17037 4233 17049 4267
rect 17083 4264 17095 4267
rect 17083 4236 17540 4264
rect 17083 4233 17095 4236
rect 17037 4227 17095 4233
rect 5276 4168 8064 4196
rect 8113 4199 8171 4205
rect 5046 4159 5104 4165
rect 8113 4165 8125 4199
rect 8159 4196 8171 4199
rect 9030 4196 9036 4208
rect 8159 4168 9036 4196
rect 8159 4165 8171 4168
rect 8113 4159 8171 4165
rect 9030 4156 9036 4168
rect 9088 4156 9094 4208
rect 11422 4196 11428 4208
rect 10428 4168 11428 4196
rect 4580 4100 4660 4128
rect 4709 4131 4767 4137
rect 4580 4088 4586 4100
rect 4709 4097 4721 4131
rect 4755 4128 4767 4131
rect 7190 4128 7196 4140
rect 4755 4100 7196 4128
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 7190 4088 7196 4100
rect 7248 4088 7254 4140
rect 7282 4088 7288 4140
rect 7340 4128 7346 4140
rect 7469 4131 7527 4137
rect 7469 4128 7481 4131
rect 7340 4100 7481 4128
rect 7340 4088 7346 4100
rect 7469 4097 7481 4100
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 7742 4088 7748 4140
rect 7800 4128 7806 4140
rect 7800 4100 8340 4128
rect 7800 4088 7806 4100
rect 4798 4060 4804 4072
rect 4759 4032 4804 4060
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 6733 4063 6791 4069
rect 6733 4029 6745 4063
rect 6779 4029 6791 4063
rect 6733 4023 6791 4029
rect 6825 4063 6883 4069
rect 6825 4029 6837 4063
rect 6871 4060 6883 4063
rect 7006 4060 7012 4072
rect 6871 4032 7012 4060
rect 6871 4029 6883 4032
rect 6825 4023 6883 4029
rect 3970 3992 3976 4004
rect 3931 3964 3976 3992
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 5810 3952 5816 4004
rect 5868 3992 5874 4004
rect 6178 3992 6184 4004
rect 5868 3964 6184 3992
rect 5868 3952 5874 3964
rect 6178 3952 6184 3964
rect 6236 3952 6242 4004
rect 6748 3992 6776 4023
rect 7006 4020 7012 4032
rect 7064 4020 7070 4072
rect 7760 4060 7788 4088
rect 8202 4060 8208 4072
rect 7208 4032 7788 4060
rect 8163 4032 8208 4060
rect 7208 3992 7236 4032
rect 8202 4020 8208 4032
rect 8260 4020 8266 4072
rect 8312 4069 8340 4100
rect 8478 4088 8484 4140
rect 8536 4128 8542 4140
rect 8573 4131 8631 4137
rect 8573 4128 8585 4131
rect 8536 4100 8585 4128
rect 8536 4088 8542 4100
rect 8573 4097 8585 4100
rect 8619 4097 8631 4131
rect 8829 4131 8887 4137
rect 8829 4128 8841 4131
rect 8573 4091 8631 4097
rect 8680 4100 8841 4128
rect 8297 4063 8355 4069
rect 8297 4029 8309 4063
rect 8343 4029 8355 4063
rect 8680 4060 8708 4100
rect 8829 4097 8841 4100
rect 8875 4097 8887 4131
rect 8829 4091 8887 4097
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4128 10103 4131
rect 10428 4128 10456 4168
rect 11422 4156 11428 4168
rect 11480 4156 11486 4208
rect 16574 4156 16580 4208
rect 16632 4196 16638 4208
rect 17129 4199 17187 4205
rect 17129 4196 17141 4199
rect 16632 4168 17141 4196
rect 16632 4156 16638 4168
rect 17129 4165 17141 4168
rect 17175 4165 17187 4199
rect 17129 4159 17187 4165
rect 10091 4100 10456 4128
rect 10505 4131 10563 4137
rect 10091 4097 10103 4100
rect 10045 4091 10103 4097
rect 10505 4097 10517 4131
rect 10551 4128 10563 4131
rect 10594 4128 10600 4140
rect 10551 4100 10600 4128
rect 10551 4097 10563 4100
rect 10505 4091 10563 4097
rect 10594 4088 10600 4100
rect 10652 4088 10658 4140
rect 11330 4088 11336 4140
rect 11388 4128 11394 4140
rect 12630 4131 12688 4137
rect 12630 4128 12642 4131
rect 11388 4100 12642 4128
rect 11388 4088 11394 4100
rect 12630 4097 12642 4100
rect 12676 4097 12688 4131
rect 13354 4128 13360 4140
rect 13315 4100 13360 4128
rect 12630 4091 12688 4097
rect 13354 4088 13360 4100
rect 13412 4088 13418 4140
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 13909 4131 13967 4137
rect 13909 4128 13921 4131
rect 13872 4100 13921 4128
rect 13872 4088 13878 4100
rect 13909 4097 13921 4100
rect 13955 4097 13967 4131
rect 13909 4091 13967 4097
rect 14274 4088 14280 4140
rect 14332 4128 14338 4140
rect 15361 4131 15419 4137
rect 15361 4128 15373 4131
rect 14332 4100 15373 4128
rect 14332 4088 14338 4100
rect 15361 4097 15373 4100
rect 15407 4097 15419 4131
rect 17236 4128 17264 4236
rect 17512 4196 17540 4236
rect 17586 4224 17592 4276
rect 17644 4264 17650 4276
rect 17681 4267 17739 4273
rect 17681 4264 17693 4267
rect 17644 4236 17693 4264
rect 17644 4224 17650 4236
rect 17681 4233 17693 4236
rect 17727 4233 17739 4267
rect 19150 4264 19156 4276
rect 17681 4227 17739 4233
rect 18708 4236 19156 4264
rect 17862 4196 17868 4208
rect 17512 4168 17868 4196
rect 17862 4156 17868 4168
rect 17920 4156 17926 4208
rect 17494 4128 17500 4140
rect 15361 4091 15419 4097
rect 17144 4100 17264 4128
rect 17455 4100 17500 4128
rect 8297 4023 8355 4029
rect 8496 4032 8708 4060
rect 10689 4063 10747 4069
rect 6748 3964 7236 3992
rect 7653 3995 7711 4001
rect 7653 3961 7665 3995
rect 7699 3992 7711 3995
rect 8386 3992 8392 4004
rect 7699 3964 8392 3992
rect 7699 3961 7711 3964
rect 7653 3955 7711 3961
rect 8386 3952 8392 3964
rect 8444 3952 8450 4004
rect 3418 3924 3424 3936
rect 3283 3896 3424 3924
rect 3283 3893 3295 3896
rect 3237 3887 3295 3893
rect 3418 3884 3424 3896
rect 3476 3884 3482 3936
rect 4065 3927 4123 3933
rect 4065 3893 4077 3927
rect 4111 3924 4123 3927
rect 6086 3924 6092 3936
rect 4111 3896 6092 3924
rect 4111 3893 4123 3896
rect 4065 3887 4123 3893
rect 6086 3884 6092 3896
rect 6144 3884 6150 3936
rect 6914 3884 6920 3936
rect 6972 3924 6978 3936
rect 8496 3924 8524 4032
rect 10689 4029 10701 4063
rect 10735 4029 10747 4063
rect 10870 4060 10876 4072
rect 10831 4032 10876 4060
rect 10689 4023 10747 4029
rect 10321 3995 10379 4001
rect 10321 3961 10333 3995
rect 10367 3992 10379 3995
rect 10502 3992 10508 4004
rect 10367 3964 10508 3992
rect 10367 3961 10379 3964
rect 10321 3955 10379 3961
rect 10502 3952 10508 3964
rect 10560 3952 10566 4004
rect 10704 3992 10732 4023
rect 10870 4020 10876 4032
rect 10928 4020 10934 4072
rect 12897 4063 12955 4069
rect 12897 4029 12909 4063
rect 12943 4029 12955 4063
rect 12897 4023 12955 4029
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 13998 4060 14004 4072
rect 13311 4032 14004 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 12912 3992 12940 4023
rect 13998 4020 14004 4032
rect 14056 4020 14062 4072
rect 14090 4020 14096 4072
rect 14148 4060 14154 4072
rect 14645 4063 14703 4069
rect 14645 4060 14657 4063
rect 14148 4032 14657 4060
rect 14148 4020 14154 4032
rect 14645 4029 14657 4032
rect 14691 4029 14703 4063
rect 14645 4023 14703 4029
rect 15105 4063 15163 4069
rect 15105 4029 15117 4063
rect 15151 4029 15163 4063
rect 15105 4023 15163 4029
rect 15120 3992 15148 4023
rect 10704 3964 11560 3992
rect 11532 3936 11560 3964
rect 12912 3964 15148 3992
rect 16485 3995 16543 4001
rect 6972 3896 8524 3924
rect 6972 3884 6978 3896
rect 9858 3884 9864 3936
rect 9916 3924 9922 3936
rect 9953 3927 10011 3933
rect 9953 3924 9965 3927
rect 9916 3896 9965 3924
rect 9916 3884 9922 3896
rect 9953 3893 9965 3896
rect 9999 3893 10011 3927
rect 9953 3887 10011 3893
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 11333 3927 11391 3933
rect 11333 3924 11345 3927
rect 11296 3896 11345 3924
rect 11296 3884 11302 3896
rect 11333 3893 11345 3896
rect 11379 3893 11391 3927
rect 11514 3924 11520 3936
rect 11475 3896 11520 3924
rect 11333 3887 11391 3893
rect 11514 3884 11520 3896
rect 11572 3884 11578 3936
rect 12526 3884 12532 3936
rect 12584 3924 12590 3936
rect 12912 3924 12940 3964
rect 16485 3961 16497 3995
rect 16531 3992 16543 3995
rect 17144 3992 17172 4100
rect 17494 4088 17500 4100
rect 17552 4088 17558 4140
rect 17773 4131 17831 4137
rect 17773 4097 17785 4131
rect 17819 4128 17831 4131
rect 18322 4128 18328 4140
rect 17819 4100 18328 4128
rect 17819 4097 17831 4100
rect 17773 4091 17831 4097
rect 18322 4088 18328 4100
rect 18380 4088 18386 4140
rect 18414 4088 18420 4140
rect 18472 4128 18478 4140
rect 18708 4128 18736 4236
rect 19150 4224 19156 4236
rect 19208 4224 19214 4276
rect 19610 4224 19616 4276
rect 19668 4264 19674 4276
rect 19705 4267 19763 4273
rect 19705 4264 19717 4267
rect 19668 4236 19717 4264
rect 19668 4224 19674 4236
rect 19705 4233 19717 4236
rect 19751 4233 19763 4267
rect 19705 4227 19763 4233
rect 19794 4224 19800 4276
rect 19852 4264 19858 4276
rect 22925 4267 22983 4273
rect 22925 4264 22937 4267
rect 19852 4236 22937 4264
rect 19852 4224 19858 4236
rect 22925 4233 22937 4236
rect 22971 4233 22983 4267
rect 22925 4227 22983 4233
rect 19996 4168 20300 4196
rect 18472 4100 18517 4128
rect 18616 4100 18736 4128
rect 18785 4131 18843 4137
rect 18472 4088 18478 4100
rect 17310 4060 17316 4072
rect 17223 4032 17316 4060
rect 17310 4020 17316 4032
rect 17368 4060 17374 4072
rect 17678 4060 17684 4072
rect 17368 4032 17684 4060
rect 17368 4020 17374 4032
rect 17678 4020 17684 4032
rect 17736 4020 17742 4072
rect 18616 4060 18644 4100
rect 18785 4097 18797 4131
rect 18831 4128 18843 4131
rect 18966 4128 18972 4140
rect 18831 4100 18972 4128
rect 18831 4097 18843 4100
rect 18785 4091 18843 4097
rect 18966 4088 18972 4100
rect 19024 4088 19030 4140
rect 19242 4088 19248 4140
rect 19300 4128 19306 4140
rect 19300 4100 19345 4128
rect 19300 4088 19306 4100
rect 19058 4060 19064 4072
rect 17779 4032 18644 4060
rect 19019 4032 19064 4060
rect 16531 3964 17172 3992
rect 16531 3961 16543 3964
rect 16485 3955 16543 3961
rect 12584 3896 12940 3924
rect 13817 3927 13875 3933
rect 12584 3884 12590 3896
rect 13817 3893 13829 3927
rect 13863 3924 13875 3927
rect 13906 3924 13912 3936
rect 13863 3896 13912 3924
rect 13863 3893 13875 3896
rect 13817 3887 13875 3893
rect 13906 3884 13912 3896
rect 13964 3884 13970 3936
rect 14550 3924 14556 3936
rect 14511 3896 14556 3924
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 14826 3884 14832 3936
rect 14884 3924 14890 3936
rect 14921 3927 14979 3933
rect 14921 3924 14933 3927
rect 14884 3896 14933 3924
rect 14884 3884 14890 3896
rect 14921 3893 14933 3896
rect 14967 3893 14979 3927
rect 14921 3887 14979 3893
rect 15286 3884 15292 3936
rect 15344 3924 15350 3936
rect 17779 3924 17807 4032
rect 19058 4020 19064 4032
rect 19116 4020 19122 4072
rect 19996 4060 20024 4168
rect 20070 4088 20076 4140
rect 20128 4128 20134 4140
rect 20165 4131 20223 4137
rect 20165 4128 20177 4131
rect 20128 4100 20177 4128
rect 20128 4088 20134 4100
rect 20165 4097 20177 4100
rect 20211 4097 20223 4131
rect 20272 4128 20300 4168
rect 20346 4156 20352 4208
rect 20404 4196 20410 4208
rect 20502 4199 20560 4205
rect 20502 4196 20514 4199
rect 20404 4168 20514 4196
rect 20404 4156 20410 4168
rect 20502 4165 20514 4168
rect 20548 4165 20560 4199
rect 20502 4159 20560 4165
rect 20990 4156 20996 4208
rect 21048 4196 21054 4208
rect 21358 4196 21364 4208
rect 21048 4168 21364 4196
rect 21048 4156 21054 4168
rect 21358 4156 21364 4168
rect 21416 4156 21422 4208
rect 21450 4156 21456 4208
rect 21508 4196 21514 4208
rect 21634 4196 21640 4208
rect 21508 4168 21640 4196
rect 21508 4156 21514 4168
rect 21634 4156 21640 4168
rect 21692 4156 21698 4208
rect 22462 4156 22468 4208
rect 22520 4196 22526 4208
rect 22738 4196 22744 4208
rect 22520 4168 22744 4196
rect 22520 4156 22526 4168
rect 22738 4156 22744 4168
rect 22796 4156 22802 4208
rect 21821 4131 21879 4137
rect 21821 4128 21833 4131
rect 20272 4100 21833 4128
rect 20165 4091 20223 4097
rect 21821 4097 21833 4100
rect 21867 4097 21879 4131
rect 21821 4091 21879 4097
rect 23014 4088 23020 4140
rect 23072 4128 23078 4140
rect 23109 4131 23167 4137
rect 23109 4128 23121 4131
rect 23072 4100 23121 4128
rect 23072 4088 23078 4100
rect 23109 4097 23121 4100
rect 23155 4097 23167 4131
rect 23109 4091 23167 4097
rect 20254 4060 20260 4072
rect 19168 4032 20024 4060
rect 20215 4032 20260 4060
rect 17862 3952 17868 4004
rect 17920 3992 17926 4004
rect 19168 3992 19196 4032
rect 20254 4020 20260 4032
rect 20312 4020 20318 4072
rect 21266 4020 21272 4072
rect 21324 4060 21330 4072
rect 21324 4032 22048 4060
rect 21324 4020 21330 4032
rect 22020 4004 22048 4032
rect 19978 3992 19984 4004
rect 17920 3964 19196 3992
rect 19939 3964 19984 3992
rect 17920 3952 17926 3964
rect 19978 3952 19984 3964
rect 20036 3952 20042 4004
rect 21560 3964 21864 3992
rect 15344 3896 17807 3924
rect 18601 3927 18659 3933
rect 15344 3884 15350 3896
rect 18601 3893 18613 3927
rect 18647 3924 18659 3927
rect 19058 3924 19064 3936
rect 18647 3896 19064 3924
rect 18647 3893 18659 3896
rect 18601 3887 18659 3893
rect 19058 3884 19064 3896
rect 19116 3884 19122 3936
rect 19610 3924 19616 3936
rect 19571 3896 19616 3924
rect 19610 3884 19616 3896
rect 19668 3884 19674 3936
rect 19794 3884 19800 3936
rect 19852 3924 19858 3936
rect 21560 3924 21588 3964
rect 19852 3896 21588 3924
rect 21637 3927 21695 3933
rect 19852 3884 19858 3896
rect 21637 3893 21649 3927
rect 21683 3924 21695 3927
rect 21726 3924 21732 3936
rect 21683 3896 21732 3924
rect 21683 3893 21695 3896
rect 21637 3887 21695 3893
rect 21726 3884 21732 3896
rect 21784 3884 21790 3936
rect 21836 3924 21864 3964
rect 22002 3952 22008 4004
rect 22060 3992 22066 4004
rect 22557 3995 22615 4001
rect 22557 3992 22569 3995
rect 22060 3964 22569 3992
rect 22060 3952 22066 3964
rect 22557 3961 22569 3964
rect 22603 3961 22615 3995
rect 22557 3955 22615 3961
rect 22465 3927 22523 3933
rect 22465 3924 22477 3927
rect 21836 3896 22477 3924
rect 22465 3893 22477 3896
rect 22511 3893 22523 3927
rect 22465 3887 22523 3893
rect 1104 3834 23460 3856
rect 1104 3782 3749 3834
rect 3801 3782 3813 3834
rect 3865 3782 3877 3834
rect 3929 3782 3941 3834
rect 3993 3782 4005 3834
rect 4057 3782 9347 3834
rect 9399 3782 9411 3834
rect 9463 3782 9475 3834
rect 9527 3782 9539 3834
rect 9591 3782 9603 3834
rect 9655 3782 14945 3834
rect 14997 3782 15009 3834
rect 15061 3782 15073 3834
rect 15125 3782 15137 3834
rect 15189 3782 15201 3834
rect 15253 3782 20543 3834
rect 20595 3782 20607 3834
rect 20659 3782 20671 3834
rect 20723 3782 20735 3834
rect 20787 3782 20799 3834
rect 20851 3782 23460 3834
rect 1104 3760 23460 3782
rect 3436 3692 13768 3720
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3584 2283 3587
rect 2271 3556 3372 3584
rect 2271 3553 2283 3556
rect 2225 3547 2283 3553
rect 1581 3519 1639 3525
rect 1581 3485 1593 3519
rect 1627 3516 1639 3519
rect 2038 3516 2044 3528
rect 1627 3488 2044 3516
rect 1627 3485 1639 3488
rect 1581 3479 1639 3485
rect 2038 3476 2044 3488
rect 2096 3476 2102 3528
rect 2869 3519 2927 3525
rect 2869 3485 2881 3519
rect 2915 3516 2927 3519
rect 2915 3488 3188 3516
rect 2915 3485 2927 3488
rect 2869 3479 2927 3485
rect 1394 3380 1400 3392
rect 1355 3352 1400 3380
rect 1394 3340 1400 3352
rect 1452 3340 1458 3392
rect 2958 3380 2964 3392
rect 2919 3352 2964 3380
rect 2958 3340 2964 3352
rect 3016 3340 3022 3392
rect 3160 3380 3188 3488
rect 3344 3448 3372 3556
rect 3436 3516 3464 3692
rect 6917 3655 6975 3661
rect 6917 3621 6929 3655
rect 6963 3652 6975 3655
rect 7190 3652 7196 3664
rect 6963 3624 7196 3652
rect 6963 3621 6975 3624
rect 6917 3615 6975 3621
rect 7190 3612 7196 3624
rect 7248 3612 7254 3664
rect 10965 3655 11023 3661
rect 10965 3621 10977 3655
rect 11011 3652 11023 3655
rect 11054 3652 11060 3664
rect 11011 3624 11060 3652
rect 11011 3621 11023 3624
rect 10965 3615 11023 3621
rect 11054 3612 11060 3624
rect 11112 3612 11118 3664
rect 12066 3612 12072 3664
rect 12124 3652 12130 3664
rect 12434 3652 12440 3664
rect 12124 3624 12440 3652
rect 12124 3612 12130 3624
rect 12434 3612 12440 3624
rect 12492 3612 12498 3664
rect 13740 3652 13768 3692
rect 13814 3680 13820 3732
rect 13872 3720 13878 3732
rect 13909 3723 13967 3729
rect 13909 3720 13921 3723
rect 13872 3692 13921 3720
rect 13872 3680 13878 3692
rect 13909 3689 13921 3692
rect 13955 3689 13967 3723
rect 15286 3720 15292 3732
rect 13909 3683 13967 3689
rect 14108 3692 15292 3720
rect 14108 3652 14136 3692
rect 15286 3680 15292 3692
rect 15344 3680 15350 3732
rect 15470 3720 15476 3732
rect 15431 3692 15476 3720
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 16942 3680 16948 3732
rect 17000 3720 17006 3732
rect 17037 3723 17095 3729
rect 17037 3720 17049 3723
rect 17000 3692 17049 3720
rect 17000 3680 17006 3692
rect 17037 3689 17049 3692
rect 17083 3689 17095 3723
rect 19794 3720 19800 3732
rect 17037 3683 17095 3689
rect 18524 3692 19800 3720
rect 18524 3652 18552 3692
rect 19794 3680 19800 3692
rect 19852 3680 19858 3732
rect 20165 3723 20223 3729
rect 20165 3689 20177 3723
rect 20211 3720 20223 3723
rect 22646 3720 22652 3732
rect 20211 3692 22652 3720
rect 20211 3689 20223 3692
rect 20165 3683 20223 3689
rect 22646 3680 22652 3692
rect 22704 3680 22710 3732
rect 22830 3680 22836 3732
rect 22888 3720 22894 3732
rect 23109 3723 23167 3729
rect 23109 3720 23121 3723
rect 22888 3692 23121 3720
rect 22888 3680 22894 3692
rect 23109 3689 23121 3692
rect 23155 3689 23167 3723
rect 23109 3683 23167 3689
rect 13740 3624 14136 3652
rect 16868 3624 18552 3652
rect 18601 3655 18659 3661
rect 3510 3544 3516 3596
rect 3568 3584 3574 3596
rect 4617 3587 4675 3593
rect 3568 3556 3832 3584
rect 3568 3544 3574 3556
rect 3804 3525 3832 3556
rect 4617 3553 4629 3587
rect 4663 3584 4675 3587
rect 4706 3584 4712 3596
rect 4663 3556 4712 3584
rect 4663 3553 4675 3556
rect 4617 3547 4675 3553
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 4798 3544 4804 3596
rect 4856 3584 4862 3596
rect 5537 3587 5595 3593
rect 5537 3584 5549 3587
rect 4856 3556 5549 3584
rect 4856 3544 4862 3556
rect 5537 3553 5549 3556
rect 5583 3553 5595 3587
rect 9585 3587 9643 3593
rect 9585 3584 9597 3587
rect 5537 3547 5595 3553
rect 8496 3556 9597 3584
rect 8496 3528 8524 3556
rect 9585 3553 9597 3556
rect 9631 3553 9643 3587
rect 9585 3547 9643 3553
rect 3605 3519 3663 3525
rect 3605 3516 3617 3519
rect 3436 3488 3617 3516
rect 3605 3485 3617 3488
rect 3651 3485 3663 3519
rect 3605 3479 3663 3485
rect 3789 3519 3847 3525
rect 3789 3485 3801 3519
rect 3835 3485 3847 3519
rect 7098 3516 7104 3528
rect 7059 3488 7104 3516
rect 3789 3479 3847 3485
rect 7098 3476 7104 3488
rect 7156 3476 7162 3528
rect 7377 3519 7435 3525
rect 7377 3485 7389 3519
rect 7423 3516 7435 3519
rect 8478 3516 8484 3528
rect 7423 3488 8484 3516
rect 7423 3485 7435 3488
rect 7377 3479 7435 3485
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 9214 3476 9220 3528
rect 9272 3516 9278 3528
rect 9309 3519 9367 3525
rect 9309 3516 9321 3519
rect 9272 3488 9321 3516
rect 9272 3476 9278 3488
rect 9309 3485 9321 3488
rect 9355 3485 9367 3519
rect 9600 3516 9628 3547
rect 10594 3516 10600 3528
rect 9600 3488 10600 3516
rect 9309 3479 9367 3485
rect 10594 3476 10600 3488
rect 10652 3516 10658 3528
rect 11057 3519 11115 3525
rect 11057 3516 11069 3519
rect 10652 3488 11069 3516
rect 10652 3476 10658 3488
rect 11057 3485 11069 3488
rect 11103 3485 11115 3519
rect 12526 3516 12532 3528
rect 12487 3488 12532 3516
rect 11057 3479 11115 3485
rect 12526 3476 12532 3488
rect 12584 3516 12590 3528
rect 14093 3519 14151 3525
rect 14093 3516 14105 3519
rect 12584 3488 14105 3516
rect 12584 3476 12590 3488
rect 14093 3485 14105 3488
rect 14139 3516 14151 3519
rect 15565 3519 15623 3525
rect 15565 3516 15577 3519
rect 14139 3488 15577 3516
rect 14139 3485 14151 3488
rect 14093 3479 14151 3485
rect 15565 3485 15577 3488
rect 15611 3516 15623 3519
rect 16390 3516 16396 3528
rect 15611 3488 16396 3516
rect 15611 3485 15623 3488
rect 15565 3479 15623 3485
rect 16390 3476 16396 3488
rect 16448 3476 16454 3528
rect 5782 3451 5840 3457
rect 5782 3448 5794 3451
rect 3344 3420 5794 3448
rect 5782 3417 5794 3420
rect 5828 3417 5840 3451
rect 5782 3411 5840 3417
rect 5902 3408 5908 3460
rect 5960 3448 5966 3460
rect 7622 3451 7680 3457
rect 7622 3448 7634 3451
rect 5960 3420 7634 3448
rect 5960 3408 5966 3420
rect 7622 3417 7634 3420
rect 7668 3417 7680 3451
rect 9674 3448 9680 3460
rect 7622 3411 7680 3417
rect 8312 3420 9680 3448
rect 6178 3380 6184 3392
rect 3160 3352 6184 3380
rect 6178 3340 6184 3352
rect 6236 3340 6242 3392
rect 6454 3340 6460 3392
rect 6512 3380 6518 3392
rect 6914 3380 6920 3392
rect 6512 3352 6920 3380
rect 6512 3340 6518 3352
rect 6914 3340 6920 3352
rect 6972 3340 6978 3392
rect 7285 3383 7343 3389
rect 7285 3349 7297 3383
rect 7331 3380 7343 3383
rect 8312 3380 8340 3420
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 9852 3451 9910 3457
rect 9852 3417 9864 3451
rect 9898 3448 9910 3451
rect 11146 3448 11152 3460
rect 9898 3420 11152 3448
rect 9898 3417 9910 3420
rect 9852 3411 9910 3417
rect 11146 3408 11152 3420
rect 11204 3408 11210 3460
rect 11324 3451 11382 3457
rect 11324 3417 11336 3451
rect 11370 3448 11382 3451
rect 12066 3448 12072 3460
rect 11370 3420 12072 3448
rect 11370 3417 11382 3420
rect 11324 3411 11382 3417
rect 12066 3408 12072 3420
rect 12124 3408 12130 3460
rect 12796 3451 12854 3457
rect 12796 3417 12808 3451
rect 12842 3448 12854 3451
rect 14182 3448 14188 3460
rect 12842 3420 14188 3448
rect 12842 3417 12854 3420
rect 12796 3411 12854 3417
rect 14182 3408 14188 3420
rect 14240 3408 14246 3460
rect 14360 3451 14418 3457
rect 14360 3417 14372 3451
rect 14406 3448 14418 3451
rect 14550 3448 14556 3460
rect 14406 3420 14556 3448
rect 14406 3417 14418 3420
rect 14360 3411 14418 3417
rect 14550 3408 14556 3420
rect 14608 3408 14614 3460
rect 15832 3451 15890 3457
rect 15832 3417 15844 3451
rect 15878 3448 15890 3451
rect 16868 3448 16896 3624
rect 18601 3621 18613 3655
rect 18647 3652 18659 3655
rect 18647 3624 19564 3652
rect 18647 3621 18659 3624
rect 18601 3615 18659 3621
rect 17678 3584 17684 3596
rect 17639 3556 17684 3584
rect 17678 3544 17684 3556
rect 17736 3544 17742 3596
rect 18049 3587 18107 3593
rect 18049 3553 18061 3587
rect 18095 3584 18107 3587
rect 19426 3584 19432 3596
rect 18095 3556 18920 3584
rect 19387 3556 19432 3584
rect 18095 3553 18107 3556
rect 18049 3547 18107 3553
rect 17497 3519 17555 3525
rect 17497 3485 17509 3519
rect 17543 3516 17555 3519
rect 18230 3516 18236 3528
rect 17543 3488 18236 3516
rect 17543 3485 17555 3488
rect 17497 3479 17555 3485
rect 17512 3448 17540 3479
rect 18230 3476 18236 3488
rect 18288 3476 18294 3528
rect 18892 3525 18920 3556
rect 19426 3544 19432 3556
rect 19484 3544 19490 3596
rect 19536 3593 19564 3624
rect 19521 3587 19579 3593
rect 19521 3553 19533 3587
rect 19567 3553 19579 3587
rect 20254 3584 20260 3596
rect 20167 3556 20260 3584
rect 19521 3547 19579 3553
rect 20254 3544 20260 3556
rect 20312 3544 20318 3596
rect 18877 3519 18935 3525
rect 18877 3485 18889 3519
rect 18923 3516 18935 3519
rect 18966 3516 18972 3528
rect 18923 3488 18972 3516
rect 18923 3485 18935 3488
rect 18877 3479 18935 3485
rect 18966 3476 18972 3488
rect 19024 3476 19030 3528
rect 19610 3516 19616 3528
rect 19571 3488 19616 3516
rect 19610 3476 19616 3488
rect 19668 3476 19674 3528
rect 20272 3516 20300 3544
rect 21266 3516 21272 3528
rect 20272 3488 21272 3516
rect 21266 3476 21272 3488
rect 21324 3516 21330 3528
rect 21729 3519 21787 3525
rect 21729 3516 21741 3519
rect 21324 3488 21741 3516
rect 21324 3476 21330 3488
rect 21729 3485 21741 3488
rect 21775 3485 21787 3519
rect 21729 3479 21787 3485
rect 15878 3420 16896 3448
rect 16960 3420 17540 3448
rect 15878 3417 15890 3420
rect 15832 3411 15890 3417
rect 7331 3352 8340 3380
rect 7331 3349 7343 3352
rect 7285 3343 7343 3349
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 8757 3383 8815 3389
rect 8757 3380 8769 3383
rect 8444 3352 8769 3380
rect 8444 3340 8450 3352
rect 8757 3349 8769 3352
rect 8803 3349 8815 3383
rect 8757 3343 8815 3349
rect 9493 3383 9551 3389
rect 9493 3349 9505 3383
rect 9539 3380 9551 3383
rect 10870 3380 10876 3392
rect 9539 3352 10876 3380
rect 9539 3349 9551 3352
rect 9493 3343 9551 3349
rect 10870 3340 10876 3352
rect 10928 3340 10934 3392
rect 10962 3340 10968 3392
rect 11020 3380 11026 3392
rect 13630 3380 13636 3392
rect 11020 3352 13636 3380
rect 11020 3340 11026 3352
rect 13630 3340 13636 3352
rect 13688 3340 13694 3392
rect 13722 3340 13728 3392
rect 13780 3380 13786 3392
rect 16758 3380 16764 3392
rect 13780 3352 16764 3380
rect 13780 3340 13786 3352
rect 16758 3340 16764 3352
rect 16816 3340 16822 3392
rect 16960 3389 16988 3420
rect 17678 3408 17684 3460
rect 17736 3448 17742 3460
rect 20530 3457 20536 3460
rect 18693 3451 18751 3457
rect 18693 3448 18705 3451
rect 17736 3420 18705 3448
rect 17736 3408 17742 3420
rect 18693 3417 18705 3420
rect 18739 3417 18751 3451
rect 18693 3411 18751 3417
rect 19996 3420 20484 3448
rect 16945 3383 17003 3389
rect 16945 3349 16957 3383
rect 16991 3349 17003 3383
rect 17402 3380 17408 3392
rect 17363 3352 17408 3380
rect 16945 3343 17003 3349
rect 17402 3340 17408 3352
rect 17460 3340 17466 3392
rect 18138 3380 18144 3392
rect 18099 3352 18144 3380
rect 18138 3340 18144 3352
rect 18196 3340 18202 3392
rect 18233 3383 18291 3389
rect 18233 3349 18245 3383
rect 18279 3380 18291 3383
rect 18322 3380 18328 3392
rect 18279 3352 18328 3380
rect 18279 3349 18291 3352
rect 18233 3343 18291 3349
rect 18322 3340 18328 3352
rect 18380 3340 18386 3392
rect 19996 3389 20024 3420
rect 19981 3383 20039 3389
rect 19981 3349 19993 3383
rect 20027 3349 20039 3383
rect 20456 3380 20484 3420
rect 20524 3411 20536 3457
rect 20588 3448 20594 3460
rect 20588 3420 20624 3448
rect 20530 3408 20536 3411
rect 20588 3408 20594 3420
rect 20714 3408 20720 3460
rect 20772 3448 20778 3460
rect 21974 3451 22032 3457
rect 21974 3448 21986 3451
rect 20772 3420 21986 3448
rect 20772 3408 20778 3420
rect 21974 3417 21986 3420
rect 22020 3417 22032 3451
rect 21974 3411 22032 3417
rect 21266 3380 21272 3392
rect 20456 3352 21272 3380
rect 19981 3343 20039 3349
rect 21266 3340 21272 3352
rect 21324 3340 21330 3392
rect 21634 3380 21640 3392
rect 21595 3352 21640 3380
rect 21634 3340 21640 3352
rect 21692 3340 21698 3392
rect 1104 3290 23460 3312
rect 1104 3238 6548 3290
rect 6600 3238 6612 3290
rect 6664 3238 6676 3290
rect 6728 3238 6740 3290
rect 6792 3238 6804 3290
rect 6856 3238 12146 3290
rect 12198 3238 12210 3290
rect 12262 3238 12274 3290
rect 12326 3238 12338 3290
rect 12390 3238 12402 3290
rect 12454 3238 17744 3290
rect 17796 3238 17808 3290
rect 17860 3238 17872 3290
rect 17924 3238 17936 3290
rect 17988 3238 18000 3290
rect 18052 3238 23460 3290
rect 1104 3216 23460 3238
rect 2498 3176 2504 3188
rect 2459 3148 2504 3176
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 3234 3176 3240 3188
rect 3195 3148 3240 3176
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 4065 3179 4123 3185
rect 4065 3145 4077 3179
rect 4111 3176 4123 3179
rect 5902 3176 5908 3188
rect 4111 3148 5908 3176
rect 4111 3145 4123 3148
rect 4065 3139 4123 3145
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 5994 3136 6000 3188
rect 6052 3176 6058 3188
rect 6178 3176 6184 3188
rect 6052 3148 6184 3176
rect 6052 3136 6058 3148
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 6365 3179 6423 3185
rect 6365 3145 6377 3179
rect 6411 3176 6423 3179
rect 6454 3176 6460 3188
rect 6411 3148 6460 3176
rect 6411 3145 6423 3148
rect 6365 3139 6423 3145
rect 6454 3136 6460 3148
rect 6512 3136 6518 3188
rect 10962 3176 10968 3188
rect 6932 3148 10968 3176
rect 2038 3108 2044 3120
rect 1999 3080 2044 3108
rect 2038 3068 2044 3080
rect 2096 3068 2102 3120
rect 3510 3108 3516 3120
rect 2332 3080 3516 3108
rect 1489 3043 1547 3049
rect 1489 3009 1501 3043
rect 1535 3040 1547 3043
rect 1578 3040 1584 3052
rect 1535 3012 1584 3040
rect 1535 3009 1547 3012
rect 1489 3003 1547 3009
rect 1578 3000 1584 3012
rect 1636 3000 1642 3052
rect 2332 3049 2360 3080
rect 3510 3068 3516 3080
rect 3568 3068 3574 3120
rect 6932 3108 6960 3148
rect 10962 3136 10968 3148
rect 11020 3136 11026 3188
rect 11330 3176 11336 3188
rect 11291 3148 11336 3176
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 12066 3136 12072 3188
rect 12124 3176 12130 3188
rect 12161 3179 12219 3185
rect 12161 3176 12173 3179
rect 12124 3148 12173 3176
rect 12124 3136 12130 3148
rect 12161 3145 12173 3148
rect 12207 3145 12219 3179
rect 12526 3176 12532 3188
rect 12161 3139 12219 3145
rect 12268 3148 12532 3176
rect 3988 3080 6960 3108
rect 2317 3043 2375 3049
rect 2317 3009 2329 3043
rect 2363 3009 2375 3043
rect 2317 3003 2375 3009
rect 2498 3000 2504 3052
rect 2556 3040 2562 3052
rect 3988 3049 4016 3080
rect 7190 3068 7196 3120
rect 7248 3108 7254 3120
rect 7346 3111 7404 3117
rect 7346 3108 7358 3111
rect 7248 3080 7358 3108
rect 7248 3068 7254 3080
rect 7346 3077 7358 3080
rect 7392 3077 7404 3111
rect 8938 3108 8944 3120
rect 8851 3080 8944 3108
rect 7346 3071 7404 3077
rect 8938 3068 8944 3080
rect 8996 3108 9002 3120
rect 8996 3080 11192 3108
rect 8996 3068 9002 3080
rect 2593 3043 2651 3049
rect 2593 3040 2605 3043
rect 2556 3012 2605 3040
rect 2556 3000 2562 3012
rect 2593 3009 2605 3012
rect 2639 3009 2651 3043
rect 2593 3003 2651 3009
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3009 4031 3043
rect 3973 3003 4031 3009
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3009 4767 3043
rect 4709 3003 4767 3009
rect 1765 2839 1823 2845
rect 1765 2805 1777 2839
rect 1811 2836 1823 2839
rect 1854 2836 1860 2848
rect 1811 2808 1860 2836
rect 1811 2805 1823 2808
rect 1765 2799 1823 2805
rect 1854 2796 1860 2808
rect 1912 2796 1918 2848
rect 3326 2796 3332 2848
rect 3384 2836 3390 2848
rect 4724 2836 4752 3003
rect 4798 3000 4804 3052
rect 4856 3040 4862 3052
rect 5074 3049 5080 3052
rect 5068 3040 5080 3049
rect 4856 3012 4901 3040
rect 5035 3012 5080 3040
rect 4856 3000 4862 3012
rect 5068 3003 5080 3012
rect 5074 3000 5080 3003
rect 5132 3000 5138 3052
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3040 7067 3043
rect 8386 3040 8392 3052
rect 7055 3012 8392 3040
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 8386 3000 8392 3012
rect 8444 3000 8450 3052
rect 10318 3040 10324 3052
rect 10376 3049 10382 3052
rect 10288 3012 10324 3040
rect 10318 3000 10324 3012
rect 10376 3003 10388 3049
rect 10594 3040 10600 3052
rect 10555 3012 10600 3040
rect 10376 3000 10382 3003
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3040 10747 3043
rect 11054 3040 11060 3052
rect 10735 3012 11060 3040
rect 10735 3009 10747 3012
rect 10689 3003 10747 3009
rect 11054 3000 11060 3012
rect 11112 3000 11118 3052
rect 6362 2932 6368 2984
rect 6420 2972 6426 2984
rect 7101 2975 7159 2981
rect 7101 2972 7113 2975
rect 6420 2944 7113 2972
rect 6420 2932 6426 2944
rect 7101 2941 7113 2944
rect 7147 2941 7159 2975
rect 9122 2972 9128 2984
rect 9083 2944 9128 2972
rect 7101 2935 7159 2941
rect 9122 2932 9128 2944
rect 9180 2932 9186 2984
rect 6822 2904 6828 2916
rect 6104 2876 6828 2904
rect 6104 2836 6132 2876
rect 6822 2864 6828 2876
rect 6880 2864 6886 2916
rect 8573 2907 8631 2913
rect 8573 2904 8585 2907
rect 8036 2876 8585 2904
rect 3384 2808 3429 2836
rect 4724 2808 6132 2836
rect 3384 2796 3390 2808
rect 6270 2796 6276 2848
rect 6328 2836 6334 2848
rect 8036 2836 8064 2876
rect 8573 2873 8585 2876
rect 8619 2873 8631 2907
rect 8573 2867 8631 2873
rect 6328 2808 8064 2836
rect 6328 2796 6334 2808
rect 8294 2796 8300 2848
rect 8352 2836 8358 2848
rect 8481 2839 8539 2845
rect 8481 2836 8493 2839
rect 8352 2808 8493 2836
rect 8352 2796 8358 2808
rect 8481 2805 8493 2808
rect 8527 2805 8539 2839
rect 8481 2799 8539 2805
rect 9217 2839 9275 2845
rect 9217 2805 9229 2839
rect 9263 2836 9275 2839
rect 9674 2836 9680 2848
rect 9263 2808 9680 2836
rect 9263 2805 9275 2808
rect 9217 2799 9275 2805
rect 9674 2796 9680 2808
rect 9732 2796 9738 2848
rect 11164 2836 11192 3080
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 12268 3049 12296 3148
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 13906 3176 13912 3188
rect 13867 3148 13912 3176
rect 13906 3136 13912 3148
rect 13964 3136 13970 3188
rect 14550 3176 14556 3188
rect 14511 3148 14556 3176
rect 14550 3136 14556 3148
rect 14608 3136 14614 3188
rect 14734 3136 14740 3188
rect 14792 3176 14798 3188
rect 20806 3176 20812 3188
rect 14792 3148 20812 3176
rect 14792 3136 14798 3148
rect 20806 3136 20812 3148
rect 20864 3136 20870 3188
rect 21358 3136 21364 3188
rect 21416 3176 21422 3188
rect 21821 3179 21879 3185
rect 21821 3176 21833 3179
rect 21416 3148 21833 3176
rect 21416 3136 21422 3148
rect 21821 3145 21833 3148
rect 21867 3145 21879 3179
rect 21821 3139 21879 3145
rect 12618 3068 12624 3120
rect 12676 3068 12682 3120
rect 13814 3108 13820 3120
rect 13775 3080 13820 3108
rect 13814 3068 13820 3080
rect 13872 3068 13878 3120
rect 14090 3108 14096 3120
rect 14051 3080 14096 3108
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 16914 3111 16972 3117
rect 16914 3108 16926 3111
rect 14384 3080 16926 3108
rect 12253 3043 12311 3049
rect 12253 3009 12265 3043
rect 12299 3009 12311 3043
rect 12253 3003 12311 3009
rect 12520 3043 12578 3049
rect 12520 3009 12532 3043
rect 12566 3040 12578 3043
rect 12636 3040 12664 3068
rect 12566 3012 12664 3040
rect 12566 3009 12578 3012
rect 12520 3003 12578 3009
rect 14090 2932 14096 2984
rect 14148 2972 14154 2984
rect 14384 2972 14412 3080
rect 16914 3077 16926 3080
rect 16960 3077 16972 3111
rect 19334 3108 19340 3120
rect 16914 3071 16972 3077
rect 18156 3080 19340 3108
rect 14642 3000 14648 3052
rect 14700 3040 14706 3052
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 14700 3012 14841 3040
rect 14700 3000 14706 3012
rect 14829 3009 14841 3012
rect 14875 3040 14887 3043
rect 15654 3040 15660 3052
rect 14875 3012 15660 3040
rect 14875 3009 14887 3012
rect 14829 3003 14887 3009
rect 15654 3000 15660 3012
rect 15712 3000 15718 3052
rect 16206 3040 16212 3052
rect 16264 3049 16270 3052
rect 16176 3012 16212 3040
rect 16206 3000 16212 3012
rect 16264 3003 16276 3049
rect 16264 3000 16270 3003
rect 16390 3000 16396 3052
rect 16448 3040 16454 3052
rect 16485 3043 16543 3049
rect 16485 3040 16497 3043
rect 16448 3012 16497 3040
rect 16448 3000 16454 3012
rect 16485 3009 16497 3012
rect 16531 3040 16543 3043
rect 16574 3040 16580 3052
rect 16531 3012 16580 3040
rect 16531 3009 16543 3012
rect 16485 3003 16543 3009
rect 16574 3000 16580 3012
rect 16632 3040 16638 3052
rect 16669 3043 16727 3049
rect 16669 3040 16681 3043
rect 16632 3012 16681 3040
rect 16632 3000 16638 3012
rect 16669 3009 16681 3012
rect 16715 3009 16727 3043
rect 16669 3003 16727 3009
rect 16758 3000 16764 3052
rect 16816 3040 16822 3052
rect 18156 3049 18184 3080
rect 19334 3068 19340 3080
rect 19392 3108 19398 3120
rect 21174 3108 21180 3120
rect 19392 3080 21180 3108
rect 19392 3068 19398 3080
rect 18414 3049 18420 3052
rect 18141 3043 18199 3049
rect 16816 3012 17724 3040
rect 16816 3000 16822 3012
rect 14148 2944 14412 2972
rect 14148 2932 14154 2944
rect 14458 2932 14464 2984
rect 14516 2972 14522 2984
rect 14921 2975 14979 2981
rect 14921 2972 14933 2975
rect 14516 2944 14933 2972
rect 14516 2932 14522 2944
rect 14921 2941 14933 2944
rect 14967 2941 14979 2975
rect 14921 2935 14979 2941
rect 13633 2907 13691 2913
rect 13633 2873 13645 2907
rect 13679 2904 13691 2907
rect 13998 2904 14004 2916
rect 13679 2876 14004 2904
rect 13679 2873 13691 2876
rect 13633 2867 13691 2873
rect 13998 2864 14004 2876
rect 14056 2864 14062 2916
rect 14274 2864 14280 2916
rect 14332 2904 14338 2916
rect 14332 2876 15148 2904
rect 14332 2864 14338 2876
rect 13722 2836 13728 2848
rect 11164 2808 13728 2836
rect 13722 2796 13728 2808
rect 13780 2796 13786 2848
rect 14366 2836 14372 2848
rect 14327 2808 14372 2836
rect 14366 2796 14372 2808
rect 14424 2796 14430 2848
rect 15120 2845 15148 2876
rect 15105 2839 15163 2845
rect 15105 2805 15117 2839
rect 15151 2836 15163 2839
rect 17402 2836 17408 2848
rect 15151 2808 17408 2836
rect 15151 2805 15163 2808
rect 15105 2799 15163 2805
rect 17402 2796 17408 2808
rect 17460 2796 17466 2848
rect 17696 2836 17724 3012
rect 18141 3009 18153 3043
rect 18187 3009 18199 3043
rect 18141 3003 18199 3009
rect 18408 3003 18420 3049
rect 18472 3040 18478 3052
rect 18472 3012 18508 3040
rect 18414 3000 18420 3003
rect 18472 3000 18478 3012
rect 20438 3000 20444 3052
rect 20496 3040 20502 3052
rect 21008 3049 21036 3080
rect 21174 3068 21180 3080
rect 21232 3068 21238 3120
rect 21542 3068 21548 3120
rect 21600 3108 21606 3120
rect 22281 3111 22339 3117
rect 22281 3108 22293 3111
rect 21600 3080 22293 3108
rect 21600 3068 21606 3080
rect 22281 3077 22293 3080
rect 22327 3077 22339 3111
rect 22281 3071 22339 3077
rect 20726 3043 20784 3049
rect 20726 3040 20738 3043
rect 20496 3012 20738 3040
rect 20496 3000 20502 3012
rect 20726 3009 20738 3012
rect 20772 3009 20784 3043
rect 20726 3003 20784 3009
rect 20993 3043 21051 3049
rect 20993 3009 21005 3043
rect 21039 3009 21051 3043
rect 21266 3040 21272 3052
rect 21227 3012 21272 3040
rect 20993 3003 21051 3009
rect 21266 3000 21272 3012
rect 21324 3000 21330 3052
rect 21358 3000 21364 3052
rect 21416 3040 21422 3052
rect 22189 3043 22247 3049
rect 21416 3012 21461 3040
rect 21416 3000 21422 3012
rect 22189 3009 22201 3043
rect 22235 3009 22247 3043
rect 22646 3040 22652 3052
rect 22607 3012 22652 3040
rect 22189 3003 22247 3009
rect 22094 2972 22100 2984
rect 19168 2944 19748 2972
rect 18049 2907 18107 2913
rect 18049 2873 18061 2907
rect 18095 2904 18107 2907
rect 18138 2904 18144 2916
rect 18095 2876 18144 2904
rect 18095 2873 18107 2876
rect 18049 2867 18107 2873
rect 18138 2864 18144 2876
rect 18196 2864 18202 2916
rect 19168 2904 19196 2944
rect 19076 2876 19196 2904
rect 19076 2836 19104 2876
rect 19242 2864 19248 2916
rect 19300 2904 19306 2916
rect 19300 2876 19656 2904
rect 19300 2864 19306 2876
rect 17696 2808 19104 2836
rect 19150 2796 19156 2848
rect 19208 2836 19214 2848
rect 19628 2845 19656 2876
rect 19521 2839 19579 2845
rect 19521 2836 19533 2839
rect 19208 2808 19533 2836
rect 19208 2796 19214 2808
rect 19521 2805 19533 2808
rect 19567 2805 19579 2839
rect 19521 2799 19579 2805
rect 19613 2839 19671 2845
rect 19613 2805 19625 2839
rect 19659 2805 19671 2839
rect 19720 2836 19748 2944
rect 21008 2944 22100 2972
rect 21008 2836 21036 2944
rect 22094 2932 22100 2944
rect 22152 2972 22158 2984
rect 22204 2972 22232 3003
rect 22646 3000 22652 3012
rect 22704 3000 22710 3052
rect 22462 2972 22468 2984
rect 22152 2944 22232 2972
rect 22423 2944 22468 2972
rect 22152 2932 22158 2944
rect 22462 2932 22468 2944
rect 22520 2932 22526 2984
rect 22830 2972 22836 2984
rect 22791 2944 22836 2972
rect 22830 2932 22836 2944
rect 22888 2932 22894 2984
rect 19720 2808 21036 2836
rect 19613 2799 19671 2805
rect 21082 2796 21088 2848
rect 21140 2836 21146 2848
rect 21542 2836 21548 2848
rect 21140 2808 21185 2836
rect 21503 2808 21548 2836
rect 21140 2796 21146 2808
rect 21542 2796 21548 2808
rect 21600 2796 21606 2848
rect 1104 2746 23460 2768
rect 1104 2694 3749 2746
rect 3801 2694 3813 2746
rect 3865 2694 3877 2746
rect 3929 2694 3941 2746
rect 3993 2694 4005 2746
rect 4057 2694 9347 2746
rect 9399 2694 9411 2746
rect 9463 2694 9475 2746
rect 9527 2694 9539 2746
rect 9591 2694 9603 2746
rect 9655 2694 14945 2746
rect 14997 2694 15009 2746
rect 15061 2694 15073 2746
rect 15125 2694 15137 2746
rect 15189 2694 15201 2746
rect 15253 2694 20543 2746
rect 20595 2694 20607 2746
rect 20659 2694 20671 2746
rect 20723 2694 20735 2746
rect 20787 2694 20799 2746
rect 20851 2694 23460 2746
rect 1104 2672 23460 2694
rect 4798 2592 4804 2644
rect 4856 2632 4862 2644
rect 7006 2632 7012 2644
rect 4856 2604 6040 2632
rect 4856 2592 4862 2604
rect 5902 2564 5908 2576
rect 5644 2536 5908 2564
rect 5644 2505 5672 2536
rect 5902 2524 5908 2536
rect 5960 2524 5966 2576
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2465 5687 2499
rect 5629 2459 5687 2465
rect 5721 2499 5779 2505
rect 5721 2465 5733 2499
rect 5767 2496 5779 2499
rect 5810 2496 5816 2508
rect 5767 2468 5816 2496
rect 5767 2465 5779 2468
rect 5721 2459 5779 2465
rect 5810 2456 5816 2468
rect 5868 2456 5874 2508
rect 6012 2496 6040 2604
rect 6380 2604 7012 2632
rect 6181 2567 6239 2573
rect 6181 2533 6193 2567
rect 6227 2564 6239 2567
rect 6380 2564 6408 2604
rect 7006 2592 7012 2604
rect 7064 2592 7070 2644
rect 7098 2592 7104 2644
rect 7156 2632 7162 2644
rect 7156 2604 7328 2632
rect 7156 2592 7162 2604
rect 6227 2536 6408 2564
rect 7300 2564 7328 2604
rect 7374 2592 7380 2644
rect 7432 2632 7438 2644
rect 7745 2635 7803 2641
rect 7745 2632 7757 2635
rect 7432 2604 7757 2632
rect 7432 2592 7438 2604
rect 7745 2601 7757 2604
rect 7791 2601 7803 2635
rect 7745 2595 7803 2601
rect 8021 2635 8079 2641
rect 8021 2601 8033 2635
rect 8067 2632 8079 2635
rect 8202 2632 8208 2644
rect 8067 2604 8208 2632
rect 8067 2601 8079 2604
rect 8021 2595 8079 2601
rect 8202 2592 8208 2604
rect 8260 2592 8266 2644
rect 9030 2592 9036 2644
rect 9088 2632 9094 2644
rect 9401 2635 9459 2641
rect 9401 2632 9413 2635
rect 9088 2604 9413 2632
rect 9088 2592 9094 2604
rect 9401 2601 9413 2604
rect 9447 2601 9459 2635
rect 9950 2632 9956 2644
rect 9401 2595 9459 2601
rect 9508 2604 9956 2632
rect 9508 2564 9536 2604
rect 9950 2592 9956 2604
rect 10008 2592 10014 2644
rect 10318 2592 10324 2644
rect 10376 2632 10382 2644
rect 10873 2635 10931 2641
rect 10873 2632 10885 2635
rect 10376 2604 10885 2632
rect 10376 2592 10382 2604
rect 10873 2601 10885 2604
rect 10919 2601 10931 2635
rect 10873 2595 10931 2601
rect 11146 2592 11152 2644
rect 11204 2632 11210 2644
rect 12161 2635 12219 2641
rect 12161 2632 12173 2635
rect 11204 2604 12173 2632
rect 11204 2592 11210 2604
rect 12161 2601 12173 2604
rect 12207 2601 12219 2635
rect 12161 2595 12219 2601
rect 12989 2635 13047 2641
rect 12989 2601 13001 2635
rect 13035 2632 13047 2635
rect 13446 2632 13452 2644
rect 13035 2604 13452 2632
rect 13035 2601 13047 2604
rect 12989 2595 13047 2601
rect 13446 2592 13452 2604
rect 13504 2592 13510 2644
rect 14182 2592 14188 2644
rect 14240 2632 14246 2644
rect 14737 2635 14795 2641
rect 14737 2632 14749 2635
rect 14240 2604 14749 2632
rect 14240 2592 14246 2604
rect 14737 2601 14749 2604
rect 14783 2601 14795 2635
rect 14737 2595 14795 2601
rect 15013 2635 15071 2641
rect 15013 2601 15025 2635
rect 15059 2632 15071 2635
rect 17494 2632 17500 2644
rect 15059 2604 17500 2632
rect 15059 2601 15071 2604
rect 15013 2595 15071 2601
rect 17494 2592 17500 2604
rect 17552 2592 17558 2644
rect 22830 2632 22836 2644
rect 17880 2604 22836 2632
rect 7300 2536 9536 2564
rect 9692 2536 10180 2564
rect 6227 2533 6239 2536
rect 6181 2527 6239 2533
rect 6362 2496 6368 2508
rect 6012 2468 6368 2496
rect 6362 2456 6368 2468
rect 6420 2456 6426 2508
rect 8294 2456 8300 2508
rect 8352 2496 8358 2508
rect 8680 2505 8708 2536
rect 8481 2499 8539 2505
rect 8481 2496 8493 2499
rect 8352 2468 8493 2496
rect 8352 2456 8358 2468
rect 8481 2465 8493 2468
rect 8527 2465 8539 2499
rect 8481 2459 8539 2465
rect 8665 2499 8723 2505
rect 8665 2465 8677 2499
rect 8711 2465 8723 2499
rect 9692 2496 9720 2536
rect 9858 2496 9864 2508
rect 8665 2459 8723 2465
rect 9048 2468 9720 2496
rect 9819 2468 9864 2496
rect 1854 2428 1860 2440
rect 1815 2400 1860 2428
rect 1854 2388 1860 2400
rect 1912 2388 1918 2440
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2397 2927 2431
rect 3602 2428 3608 2440
rect 3563 2400 3608 2428
rect 2869 2391 2927 2397
rect 2038 2292 2044 2304
rect 1999 2264 2044 2292
rect 2038 2252 2044 2264
rect 2096 2252 2102 2304
rect 2222 2292 2228 2304
rect 2183 2264 2228 2292
rect 2222 2252 2228 2264
rect 2280 2252 2286 2304
rect 2884 2292 2912 2391
rect 3602 2388 3608 2400
rect 3660 2388 3666 2440
rect 4614 2428 4620 2440
rect 4575 2400 4620 2428
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 5350 2428 5356 2440
rect 5311 2400 5356 2428
rect 5350 2388 5356 2400
rect 5408 2388 5414 2440
rect 8202 2428 8208 2440
rect 5736 2400 8208 2428
rect 2961 2363 3019 2369
rect 2961 2329 2973 2363
rect 3007 2360 3019 2363
rect 4709 2363 4767 2369
rect 3007 2332 4660 2360
rect 3007 2329 3019 2332
rect 2961 2323 3019 2329
rect 3786 2292 3792 2304
rect 2884 2264 3792 2292
rect 3786 2252 3792 2264
rect 3844 2252 3850 2304
rect 3970 2292 3976 2304
rect 3931 2264 3976 2292
rect 3970 2252 3976 2264
rect 4028 2252 4034 2304
rect 4632 2292 4660 2332
rect 4709 2329 4721 2363
rect 4755 2360 4767 2363
rect 5736 2360 5764 2400
rect 8202 2388 8208 2400
rect 8260 2388 8266 2440
rect 8386 2428 8392 2440
rect 8347 2400 8392 2428
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 4755 2332 5764 2360
rect 4755 2329 4767 2332
rect 4709 2323 4767 2329
rect 5810 2320 5816 2372
rect 5868 2360 5874 2372
rect 5868 2332 5913 2360
rect 5868 2320 5874 2332
rect 6086 2320 6092 2372
rect 6144 2360 6150 2372
rect 6610 2363 6668 2369
rect 6610 2360 6622 2363
rect 6144 2332 6622 2360
rect 6144 2320 6150 2332
rect 6610 2329 6622 2332
rect 6656 2329 6668 2363
rect 6610 2323 6668 2329
rect 6822 2320 6828 2372
rect 6880 2320 6886 2372
rect 8110 2320 8116 2372
rect 8168 2360 8174 2372
rect 9048 2360 9076 2468
rect 9858 2456 9864 2468
rect 9916 2456 9922 2508
rect 9950 2456 9956 2508
rect 10008 2496 10014 2508
rect 10152 2496 10180 2536
rect 10226 2524 10232 2576
rect 10284 2564 10290 2576
rect 11057 2567 11115 2573
rect 11057 2564 11069 2567
rect 10284 2536 11069 2564
rect 10284 2524 10290 2536
rect 11057 2533 11069 2536
rect 11103 2533 11115 2567
rect 11057 2527 11115 2533
rect 11238 2524 11244 2576
rect 11296 2564 11302 2576
rect 13265 2567 13323 2573
rect 11296 2536 12572 2564
rect 11296 2524 11302 2536
rect 10008 2468 10053 2496
rect 10152 2468 11652 2496
rect 10008 2456 10014 2468
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9876 2428 9904 2456
rect 11256 2437 11284 2468
rect 10229 2431 10287 2437
rect 10229 2428 10241 2431
rect 9876 2400 10241 2428
rect 9769 2391 9827 2397
rect 10229 2397 10241 2400
rect 10275 2397 10287 2431
rect 10229 2391 10287 2397
rect 11241 2431 11299 2437
rect 11241 2397 11253 2431
rect 11287 2397 11299 2431
rect 11241 2391 11299 2397
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 11624 2428 11652 2468
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 11756 2468 12020 2496
rect 11756 2456 11762 2468
rect 11624 2400 11928 2428
rect 11517 2391 11575 2397
rect 8168 2332 9076 2360
rect 8168 2320 8174 2332
rect 9122 2320 9128 2372
rect 9180 2360 9186 2372
rect 9784 2360 9812 2391
rect 11532 2360 11560 2391
rect 11698 2360 11704 2372
rect 9180 2332 9720 2360
rect 9784 2332 11560 2360
rect 11624 2332 11704 2360
rect 9180 2320 9186 2332
rect 6840 2292 6868 2320
rect 9306 2292 9312 2304
rect 4632 2264 6868 2292
rect 9267 2264 9312 2292
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 9692 2292 9720 2332
rect 11624 2292 11652 2332
rect 11698 2320 11704 2332
rect 11756 2320 11762 2372
rect 9692 2264 11652 2292
rect 11900 2292 11928 2400
rect 11992 2360 12020 2468
rect 12066 2456 12072 2508
rect 12124 2496 12130 2508
rect 12544 2505 12572 2536
rect 13265 2533 13277 2567
rect 13311 2564 13323 2567
rect 14090 2564 14096 2576
rect 13311 2536 14096 2564
rect 13311 2533 13323 2536
rect 13265 2527 13323 2533
rect 14090 2524 14096 2536
rect 14148 2524 14154 2576
rect 15286 2564 15292 2576
rect 15247 2536 15292 2564
rect 15286 2524 15292 2536
rect 15344 2524 15350 2576
rect 15378 2524 15384 2576
rect 15436 2564 15442 2576
rect 16117 2567 16175 2573
rect 16117 2564 16129 2567
rect 15436 2536 16129 2564
rect 15436 2524 15442 2536
rect 16117 2533 16129 2536
rect 16163 2533 16175 2567
rect 16390 2564 16396 2576
rect 16351 2536 16396 2564
rect 16117 2527 16175 2533
rect 16390 2524 16396 2536
rect 16448 2524 16454 2576
rect 12345 2499 12403 2505
rect 12345 2496 12357 2499
rect 12124 2468 12357 2496
rect 12124 2456 12130 2468
rect 12345 2465 12357 2468
rect 12391 2465 12403 2499
rect 12345 2459 12403 2465
rect 12529 2499 12587 2505
rect 12529 2465 12541 2499
rect 12575 2465 12587 2499
rect 14274 2496 14280 2508
rect 12529 2459 12587 2465
rect 13924 2468 14280 2496
rect 12621 2431 12679 2437
rect 12621 2397 12633 2431
rect 12667 2428 12679 2431
rect 12710 2428 12716 2440
rect 12667 2400 12716 2428
rect 12667 2397 12679 2400
rect 12621 2391 12679 2397
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 13924 2437 13952 2468
rect 14274 2456 14280 2468
rect 14332 2456 14338 2508
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 14424 2468 15148 2496
rect 14424 2456 14430 2468
rect 13909 2431 13967 2437
rect 13909 2397 13921 2431
rect 13955 2397 13967 2431
rect 13909 2391 13967 2397
rect 13998 2388 14004 2440
rect 14056 2428 14062 2440
rect 15120 2437 15148 2468
rect 16574 2456 16580 2508
rect 16632 2496 16638 2508
rect 16761 2499 16819 2505
rect 16761 2496 16773 2499
rect 16632 2468 16773 2496
rect 16632 2456 16638 2468
rect 16761 2465 16773 2468
rect 16807 2465 16819 2499
rect 16761 2459 16819 2465
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 14056 2400 14105 2428
rect 14056 2388 14062 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 15105 2431 15163 2437
rect 15105 2397 15117 2431
rect 15151 2397 15163 2431
rect 15470 2428 15476 2440
rect 15431 2400 15476 2428
rect 15105 2391 15163 2397
rect 14844 2360 14872 2391
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 16206 2428 16212 2440
rect 16167 2400 16212 2428
rect 16206 2388 16212 2400
rect 16264 2388 16270 2440
rect 17880 2428 17908 2604
rect 22830 2592 22836 2604
rect 22888 2592 22894 2644
rect 20714 2564 20720 2576
rect 20675 2536 20720 2564
rect 20714 2524 20720 2536
rect 20772 2524 20778 2576
rect 20809 2567 20867 2573
rect 20809 2533 20821 2567
rect 20855 2564 20867 2567
rect 20898 2564 20904 2576
rect 20855 2536 20904 2564
rect 20855 2533 20867 2536
rect 20809 2527 20867 2533
rect 20898 2524 20904 2536
rect 20956 2524 20962 2576
rect 22370 2524 22376 2576
rect 22428 2564 22434 2576
rect 22465 2567 22523 2573
rect 22465 2564 22477 2567
rect 22428 2536 22477 2564
rect 22428 2524 22434 2536
rect 22465 2533 22477 2536
rect 22511 2533 22523 2567
rect 22738 2564 22744 2576
rect 22699 2536 22744 2564
rect 22465 2527 22523 2533
rect 22738 2524 22744 2536
rect 22796 2524 22802 2576
rect 19334 2496 19340 2508
rect 19295 2468 19340 2496
rect 19334 2456 19340 2468
rect 19392 2456 19398 2508
rect 20346 2456 20352 2508
rect 20404 2496 20410 2508
rect 21453 2499 21511 2505
rect 20404 2468 21312 2496
rect 20404 2456 20410 2468
rect 18230 2428 18236 2440
rect 16776 2400 17908 2428
rect 18191 2400 18236 2428
rect 16776 2360 16804 2400
rect 18230 2388 18236 2400
rect 18288 2388 18294 2440
rect 18966 2388 18972 2440
rect 19024 2428 19030 2440
rect 20438 2428 20444 2440
rect 19024 2400 20444 2428
rect 19024 2388 19030 2400
rect 20438 2388 20444 2400
rect 20496 2388 20502 2440
rect 21284 2428 21312 2468
rect 21453 2465 21465 2499
rect 21499 2496 21511 2499
rect 22002 2496 22008 2508
rect 21499 2468 22008 2496
rect 21499 2465 21511 2468
rect 21453 2459 21511 2465
rect 22002 2456 22008 2468
rect 22060 2456 22066 2508
rect 21821 2431 21879 2437
rect 21821 2428 21833 2431
rect 21284 2400 21833 2428
rect 21821 2397 21833 2400
rect 21867 2397 21879 2431
rect 21821 2391 21879 2397
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 22557 2431 22615 2437
rect 22557 2428 22569 2431
rect 21968 2400 22569 2428
rect 21968 2388 21974 2400
rect 22557 2397 22569 2400
rect 22603 2397 22615 2431
rect 23106 2428 23112 2440
rect 23067 2400 23112 2428
rect 22557 2391 22615 2397
rect 23106 2388 23112 2400
rect 23164 2388 23170 2440
rect 17034 2369 17040 2372
rect 11992 2332 13216 2360
rect 14844 2332 16804 2360
rect 12894 2292 12900 2304
rect 11900 2264 12900 2292
rect 12894 2252 12900 2264
rect 12952 2292 12958 2304
rect 13081 2295 13139 2301
rect 13081 2292 13093 2295
rect 12952 2264 13093 2292
rect 12952 2252 12958 2264
rect 13081 2261 13093 2264
rect 13127 2261 13139 2295
rect 13188 2292 13216 2332
rect 17028 2323 17040 2369
rect 17092 2360 17098 2372
rect 17092 2332 17128 2360
rect 18064 2332 19288 2360
rect 17034 2320 17040 2323
rect 17092 2320 17098 2332
rect 18064 2292 18092 2332
rect 13188 2264 18092 2292
rect 18141 2295 18199 2301
rect 13081 2255 13139 2261
rect 18141 2261 18153 2295
rect 18187 2292 18199 2295
rect 18230 2292 18236 2304
rect 18187 2264 18236 2292
rect 18187 2261 18199 2264
rect 18141 2255 18199 2261
rect 18230 2252 18236 2264
rect 18288 2252 18294 2304
rect 18874 2292 18880 2304
rect 18835 2264 18880 2292
rect 18874 2252 18880 2264
rect 18932 2252 18938 2304
rect 18966 2252 18972 2304
rect 19024 2292 19030 2304
rect 19260 2292 19288 2332
rect 19334 2320 19340 2372
rect 19392 2360 19398 2372
rect 19582 2363 19640 2369
rect 19582 2360 19594 2363
rect 19392 2332 19594 2360
rect 19392 2320 19398 2332
rect 19582 2329 19594 2332
rect 19628 2329 19640 2363
rect 19582 2323 19640 2329
rect 20806 2320 20812 2372
rect 20864 2360 20870 2372
rect 21269 2363 21327 2369
rect 21269 2360 21281 2363
rect 20864 2332 21281 2360
rect 20864 2320 20870 2332
rect 21269 2329 21281 2332
rect 21315 2329 21327 2363
rect 21269 2323 21327 2329
rect 21177 2295 21235 2301
rect 21177 2292 21189 2295
rect 19024 2264 19069 2292
rect 19260 2264 21189 2292
rect 19024 2252 19030 2264
rect 21177 2261 21189 2264
rect 21223 2292 21235 2295
rect 21634 2292 21640 2304
rect 21223 2264 21640 2292
rect 21223 2261 21235 2264
rect 21177 2255 21235 2261
rect 21634 2252 21640 2264
rect 21692 2252 21698 2304
rect 21818 2252 21824 2304
rect 21876 2292 21882 2304
rect 22925 2295 22983 2301
rect 22925 2292 22937 2295
rect 21876 2264 22937 2292
rect 21876 2252 21882 2264
rect 22925 2261 22937 2264
rect 22971 2261 22983 2295
rect 22925 2255 22983 2261
rect 1104 2202 23460 2224
rect 1104 2150 6548 2202
rect 6600 2150 6612 2202
rect 6664 2150 6676 2202
rect 6728 2150 6740 2202
rect 6792 2150 6804 2202
rect 6856 2150 12146 2202
rect 12198 2150 12210 2202
rect 12262 2150 12274 2202
rect 12326 2150 12338 2202
rect 12390 2150 12402 2202
rect 12454 2150 17744 2202
rect 17796 2150 17808 2202
rect 17860 2150 17872 2202
rect 17924 2150 17936 2202
rect 17988 2150 18000 2202
rect 18052 2150 23460 2202
rect 1104 2128 23460 2150
rect 3786 2048 3792 2100
rect 3844 2088 3850 2100
rect 9306 2088 9312 2100
rect 3844 2060 9312 2088
rect 3844 2048 3850 2060
rect 9306 2048 9312 2060
rect 9364 2088 9370 2100
rect 9364 2060 17448 2088
rect 9364 2048 9370 2060
rect 2222 1980 2228 2032
rect 2280 2020 2286 2032
rect 2280 1992 8156 2020
rect 2280 1980 2286 1992
rect 4614 1912 4620 1964
rect 4672 1952 4678 1964
rect 7926 1952 7932 1964
rect 4672 1924 7932 1952
rect 4672 1912 4678 1924
rect 7926 1912 7932 1924
rect 7984 1912 7990 1964
rect 8128 1952 8156 1992
rect 8202 1980 8208 2032
rect 8260 2020 8266 2032
rect 17034 2020 17040 2032
rect 8260 1992 17040 2020
rect 8260 1980 8266 1992
rect 17034 1980 17040 1992
rect 17092 1980 17098 2032
rect 17420 2020 17448 2060
rect 17494 2048 17500 2100
rect 17552 2088 17558 2100
rect 22462 2088 22468 2100
rect 17552 2060 22468 2088
rect 17552 2048 17558 2060
rect 22462 2048 22468 2060
rect 22520 2048 22526 2100
rect 20714 2020 20720 2032
rect 17420 1992 20720 2020
rect 20714 1980 20720 1992
rect 20772 1980 20778 2032
rect 14826 1952 14832 1964
rect 8128 1924 14832 1952
rect 14826 1912 14832 1924
rect 14884 1912 14890 1964
rect 16390 1912 16396 1964
rect 16448 1952 16454 1964
rect 20254 1952 20260 1964
rect 16448 1924 20260 1952
rect 16448 1912 16454 1924
rect 20254 1912 20260 1924
rect 20312 1912 20318 1964
rect 3602 1844 3608 1896
rect 3660 1884 3666 1896
rect 7374 1884 7380 1896
rect 3660 1856 7380 1884
rect 3660 1844 3666 1856
rect 7374 1844 7380 1856
rect 7432 1844 7438 1896
rect 16298 1844 16304 1896
rect 16356 1884 16362 1896
rect 18874 1884 18880 1896
rect 16356 1856 18880 1884
rect 16356 1844 16362 1856
rect 18874 1844 18880 1856
rect 18932 1844 18938 1896
rect 3418 1776 3424 1828
rect 3476 1816 3482 1828
rect 9122 1816 9128 1828
rect 3476 1788 9128 1816
rect 3476 1776 3482 1788
rect 9122 1776 9128 1788
rect 9180 1776 9186 1828
rect 15286 1776 15292 1828
rect 15344 1816 15350 1828
rect 20162 1816 20168 1828
rect 15344 1788 20168 1816
rect 15344 1776 15350 1788
rect 20162 1776 20168 1788
rect 20220 1776 20226 1828
rect 18230 1748 18236 1760
rect 16546 1720 18236 1748
rect 7926 1572 7932 1624
rect 7984 1612 7990 1624
rect 16546 1612 16574 1720
rect 18230 1708 18236 1720
rect 18288 1708 18294 1760
rect 7984 1584 16574 1612
rect 7984 1572 7990 1584
<< via1 >>
rect 6000 22924 6052 22976
rect 6736 22924 6788 22976
rect 20260 22380 20312 22432
rect 21916 22380 21968 22432
rect 3749 22278 3801 22330
rect 3813 22278 3865 22330
rect 3877 22278 3929 22330
rect 3941 22278 3993 22330
rect 4005 22278 4057 22330
rect 9347 22278 9399 22330
rect 9411 22278 9463 22330
rect 9475 22278 9527 22330
rect 9539 22278 9591 22330
rect 9603 22278 9655 22330
rect 14945 22278 14997 22330
rect 15009 22278 15061 22330
rect 15073 22278 15125 22330
rect 15137 22278 15189 22330
rect 15201 22278 15253 22330
rect 20543 22278 20595 22330
rect 20607 22278 20659 22330
rect 20671 22278 20723 22330
rect 20735 22278 20787 22330
rect 20799 22278 20851 22330
rect 8484 22176 8536 22228
rect 1952 22040 2004 22092
rect 1860 21972 1912 22024
rect 4988 22040 5040 22092
rect 3056 21972 3108 22024
rect 3332 22015 3384 22024
rect 3332 21981 3341 22015
rect 3341 21981 3375 22015
rect 3375 21981 3384 22015
rect 4068 22015 4120 22024
rect 3332 21972 3384 21981
rect 4068 21981 4077 22015
rect 4077 21981 4111 22015
rect 4111 21981 4120 22015
rect 4068 21972 4120 21981
rect 4528 21972 4580 22024
rect 5172 21972 5224 22024
rect 6460 21972 6512 22024
rect 2044 21904 2096 21956
rect 6368 21904 6420 21956
rect 6736 21904 6788 21956
rect 296 21836 348 21888
rect 1584 21836 1636 21888
rect 2228 21836 2280 21888
rect 2872 21879 2924 21888
rect 2872 21845 2881 21879
rect 2881 21845 2915 21879
rect 2915 21845 2924 21879
rect 2872 21836 2924 21845
rect 2964 21836 3016 21888
rect 3516 21879 3568 21888
rect 3516 21845 3525 21879
rect 3525 21845 3559 21879
rect 3559 21845 3568 21879
rect 3516 21836 3568 21845
rect 4160 21836 4212 21888
rect 4712 21836 4764 21888
rect 4804 21879 4856 21888
rect 4804 21845 4813 21879
rect 4813 21845 4847 21879
rect 4847 21845 4856 21879
rect 5540 21879 5592 21888
rect 4804 21836 4856 21845
rect 5540 21845 5549 21879
rect 5549 21845 5583 21879
rect 5583 21845 5592 21879
rect 5540 21836 5592 21845
rect 5632 21836 5684 21888
rect 7380 21972 7432 22024
rect 8484 21972 8536 22024
rect 8668 21972 8720 22024
rect 9128 21972 9180 22024
rect 10324 22015 10376 22024
rect 10324 21981 10333 22015
rect 10333 21981 10367 22015
rect 10367 21981 10376 22015
rect 12532 22176 12584 22228
rect 17684 22176 17736 22228
rect 13084 22108 13136 22160
rect 10324 21972 10376 21981
rect 12164 22015 12216 22024
rect 12164 21981 12173 22015
rect 12173 21981 12207 22015
rect 12207 21981 12216 22015
rect 12164 21972 12216 21981
rect 13360 21972 13412 22024
rect 13912 22015 13964 22024
rect 13912 21981 13921 22015
rect 13921 21981 13955 22015
rect 13955 21981 13964 22015
rect 13912 21972 13964 21981
rect 8116 21904 8168 21956
rect 8392 21904 8444 21956
rect 11520 21904 11572 21956
rect 8484 21879 8536 21888
rect 8484 21845 8493 21879
rect 8493 21845 8527 21879
rect 8527 21845 8536 21879
rect 8484 21836 8536 21845
rect 8760 21879 8812 21888
rect 8760 21845 8769 21879
rect 8769 21845 8803 21879
rect 8803 21845 8812 21879
rect 8760 21836 8812 21845
rect 9956 21836 10008 21888
rect 10508 21836 10560 21888
rect 11060 21836 11112 21888
rect 11796 21879 11848 21888
rect 11796 21845 11805 21879
rect 11805 21845 11839 21879
rect 11839 21845 11848 21879
rect 11796 21836 11848 21845
rect 12072 21879 12124 21888
rect 12072 21845 12081 21879
rect 12081 21845 12115 21879
rect 12115 21845 12124 21879
rect 12072 21836 12124 21845
rect 12440 21904 12492 21956
rect 12992 21947 13044 21956
rect 12992 21913 13001 21947
rect 13001 21913 13035 21947
rect 13035 21913 13044 21947
rect 12992 21904 13044 21913
rect 13636 21904 13688 21956
rect 15660 21972 15712 22024
rect 16304 22015 16356 22024
rect 16304 21981 16313 22015
rect 16313 21981 16347 22015
rect 16347 21981 16356 22015
rect 16304 21972 16356 21981
rect 13728 21836 13780 21888
rect 13820 21836 13872 21888
rect 16580 21904 16632 21956
rect 17224 21972 17276 22024
rect 17684 22015 17736 22024
rect 17684 21981 17693 22015
rect 17693 21981 17727 22015
rect 17727 21981 17736 22015
rect 17684 21972 17736 21981
rect 18144 21972 18196 22024
rect 18512 21972 18564 22024
rect 19248 21972 19300 22024
rect 19432 22015 19484 22024
rect 19432 21981 19441 22015
rect 19441 21981 19475 22015
rect 19475 21981 19484 22015
rect 22560 22176 22612 22228
rect 21916 22108 21968 22160
rect 19984 22040 20036 22092
rect 19432 21972 19484 21981
rect 19708 21904 19760 21956
rect 14740 21879 14792 21888
rect 14740 21845 14749 21879
rect 14749 21845 14783 21879
rect 14783 21845 14792 21879
rect 14740 21836 14792 21845
rect 14832 21836 14884 21888
rect 15844 21836 15896 21888
rect 16396 21879 16448 21888
rect 16396 21845 16405 21879
rect 16405 21845 16439 21879
rect 16439 21845 16448 21879
rect 16396 21836 16448 21845
rect 16672 21879 16724 21888
rect 16672 21845 16681 21879
rect 16681 21845 16715 21879
rect 16715 21845 16724 21879
rect 16672 21836 16724 21845
rect 16948 21879 17000 21888
rect 16948 21845 16957 21879
rect 16957 21845 16991 21879
rect 16991 21845 17000 21879
rect 16948 21836 17000 21845
rect 18696 21879 18748 21888
rect 18696 21845 18705 21879
rect 18705 21845 18739 21879
rect 18739 21845 18748 21879
rect 18696 21836 18748 21845
rect 19064 21836 19116 21888
rect 19248 21836 19300 21888
rect 19892 21879 19944 21888
rect 19892 21845 19901 21879
rect 19901 21845 19935 21879
rect 19935 21845 19944 21879
rect 19892 21836 19944 21845
rect 20444 21879 20496 21888
rect 20444 21845 20453 21879
rect 20453 21845 20487 21879
rect 20487 21845 20496 21879
rect 20444 21836 20496 21845
rect 20628 22015 20680 22024
rect 20628 21981 20637 22015
rect 20637 21981 20671 22015
rect 20671 21981 20680 22015
rect 20904 22015 20956 22024
rect 20628 21972 20680 21981
rect 20904 21981 20913 22015
rect 20913 21981 20947 22015
rect 20947 21981 20956 22015
rect 20904 21972 20956 21981
rect 22192 22040 22244 22092
rect 21824 22015 21876 22024
rect 21824 21981 21833 22015
rect 21833 21981 21867 22015
rect 21867 21981 21876 22015
rect 21824 21972 21876 21981
rect 22100 21972 22152 22024
rect 22744 21972 22796 22024
rect 21732 21836 21784 21888
rect 22928 21904 22980 21956
rect 22376 21836 22428 21888
rect 6548 21734 6600 21786
rect 6612 21734 6664 21786
rect 6676 21734 6728 21786
rect 6740 21734 6792 21786
rect 6804 21734 6856 21786
rect 12146 21734 12198 21786
rect 12210 21734 12262 21786
rect 12274 21734 12326 21786
rect 12338 21734 12390 21786
rect 12402 21734 12454 21786
rect 17744 21734 17796 21786
rect 17808 21734 17860 21786
rect 17872 21734 17924 21786
rect 17936 21734 17988 21786
rect 18000 21734 18052 21786
rect 940 21632 992 21684
rect 2872 21632 2924 21684
rect 4252 21632 4304 21684
rect 2504 21564 2556 21616
rect 4068 21564 4120 21616
rect 4988 21607 5040 21616
rect 4988 21573 4997 21607
rect 4997 21573 5031 21607
rect 5031 21573 5040 21607
rect 4988 21564 5040 21573
rect 5172 21607 5224 21616
rect 5172 21573 5181 21607
rect 5181 21573 5215 21607
rect 5215 21573 5224 21607
rect 5172 21564 5224 21573
rect 1768 21539 1820 21548
rect 1768 21505 1777 21539
rect 1777 21505 1811 21539
rect 1811 21505 1820 21539
rect 1768 21496 1820 21505
rect 2964 21496 3016 21548
rect 4712 21496 4764 21548
rect 2596 21471 2648 21480
rect 2596 21437 2605 21471
rect 2605 21437 2639 21471
rect 2639 21437 2648 21471
rect 2596 21428 2648 21437
rect 2780 21471 2832 21480
rect 2780 21437 2789 21471
rect 2789 21437 2823 21471
rect 2823 21437 2832 21471
rect 3424 21471 3476 21480
rect 2780 21428 2832 21437
rect 3424 21437 3433 21471
rect 3433 21437 3467 21471
rect 3467 21437 3476 21471
rect 3424 21428 3476 21437
rect 4436 21428 4488 21480
rect 5632 21632 5684 21684
rect 6368 21632 6420 21684
rect 6920 21632 6972 21684
rect 5540 21564 5592 21616
rect 2688 21360 2740 21412
rect 5724 21496 5776 21548
rect 7380 21496 7432 21548
rect 8944 21632 8996 21684
rect 8116 21564 8168 21616
rect 9220 21564 9272 21616
rect 6460 21428 6512 21480
rect 7196 21428 7248 21480
rect 9036 21496 9088 21548
rect 9128 21496 9180 21548
rect 9864 21632 9916 21684
rect 10324 21632 10376 21684
rect 12992 21632 13044 21684
rect 14188 21632 14240 21684
rect 10232 21564 10284 21616
rect 10600 21564 10652 21616
rect 12532 21564 12584 21616
rect 9680 21539 9732 21548
rect 9680 21505 9689 21539
rect 9689 21505 9723 21539
rect 9723 21505 9732 21539
rect 9680 21496 9732 21505
rect 11244 21496 11296 21548
rect 12164 21539 12216 21548
rect 12164 21505 12173 21539
rect 12173 21505 12207 21539
rect 12207 21505 12216 21539
rect 12164 21496 12216 21505
rect 10048 21428 10100 21480
rect 11336 21471 11388 21480
rect 11336 21437 11345 21471
rect 11345 21437 11379 21471
rect 11379 21437 11388 21471
rect 11336 21428 11388 21437
rect 2320 21292 2372 21344
rect 3240 21335 3292 21344
rect 3240 21301 3249 21335
rect 3249 21301 3283 21335
rect 3283 21301 3292 21335
rect 3240 21292 3292 21301
rect 5080 21292 5132 21344
rect 7104 21292 7156 21344
rect 8668 21335 8720 21344
rect 8668 21301 8677 21335
rect 8677 21301 8711 21335
rect 8711 21301 8720 21335
rect 8668 21292 8720 21301
rect 9772 21360 9824 21412
rect 12072 21360 12124 21412
rect 12900 21360 12952 21412
rect 13268 21496 13320 21548
rect 14096 21496 14148 21548
rect 13360 21471 13412 21480
rect 13360 21437 13369 21471
rect 13369 21437 13403 21471
rect 13403 21437 13412 21471
rect 13360 21428 13412 21437
rect 13544 21471 13596 21480
rect 13544 21437 13553 21471
rect 13553 21437 13587 21471
rect 13587 21437 13596 21471
rect 13544 21428 13596 21437
rect 13728 21428 13780 21480
rect 13176 21360 13228 21412
rect 10416 21292 10468 21344
rect 13728 21292 13780 21344
rect 13820 21292 13872 21344
rect 16580 21632 16632 21684
rect 16948 21607 17000 21616
rect 16948 21573 16982 21607
rect 16982 21573 17000 21607
rect 16948 21564 17000 21573
rect 18144 21632 18196 21684
rect 19432 21632 19484 21684
rect 19616 21632 19668 21684
rect 22008 21632 22060 21684
rect 18696 21564 18748 21616
rect 19064 21564 19116 21616
rect 24124 21564 24176 21616
rect 15936 21496 15988 21548
rect 20352 21496 20404 21548
rect 20904 21496 20956 21548
rect 21088 21539 21140 21548
rect 21088 21505 21097 21539
rect 21097 21505 21131 21539
rect 21131 21505 21140 21539
rect 21088 21496 21140 21505
rect 21640 21539 21692 21548
rect 21640 21505 21649 21539
rect 21649 21505 21683 21539
rect 21683 21505 21692 21539
rect 21640 21496 21692 21505
rect 22468 21539 22520 21548
rect 22468 21505 22477 21539
rect 22477 21505 22511 21539
rect 22511 21505 22520 21539
rect 22468 21496 22520 21505
rect 15568 21428 15620 21480
rect 18144 21471 18196 21480
rect 18144 21437 18153 21471
rect 18153 21437 18187 21471
rect 18187 21437 18196 21471
rect 18144 21428 18196 21437
rect 20996 21471 21048 21480
rect 20996 21437 21005 21471
rect 21005 21437 21039 21471
rect 21039 21437 21048 21471
rect 20996 21428 21048 21437
rect 21364 21428 21416 21480
rect 21824 21428 21876 21480
rect 22652 21496 22704 21548
rect 23480 21428 23532 21480
rect 19984 21360 20036 21412
rect 15384 21292 15436 21344
rect 15752 21292 15804 21344
rect 15936 21292 15988 21344
rect 19248 21292 19300 21344
rect 19524 21335 19576 21344
rect 19524 21301 19533 21335
rect 19533 21301 19567 21335
rect 19567 21301 19576 21335
rect 19524 21292 19576 21301
rect 19616 21335 19668 21344
rect 19616 21301 19625 21335
rect 19625 21301 19659 21335
rect 19659 21301 19668 21335
rect 19616 21292 19668 21301
rect 19800 21292 19852 21344
rect 21824 21335 21876 21344
rect 21824 21301 21833 21335
rect 21833 21301 21867 21335
rect 21867 21301 21876 21335
rect 21824 21292 21876 21301
rect 22836 21292 22888 21344
rect 3749 21190 3801 21242
rect 3813 21190 3865 21242
rect 3877 21190 3929 21242
rect 3941 21190 3993 21242
rect 4005 21190 4057 21242
rect 9347 21190 9399 21242
rect 9411 21190 9463 21242
rect 9475 21190 9527 21242
rect 9539 21190 9591 21242
rect 9603 21190 9655 21242
rect 14945 21190 14997 21242
rect 15009 21190 15061 21242
rect 15073 21190 15125 21242
rect 15137 21190 15189 21242
rect 15201 21190 15253 21242
rect 20543 21190 20595 21242
rect 20607 21190 20659 21242
rect 20671 21190 20723 21242
rect 20735 21190 20787 21242
rect 20799 21190 20851 21242
rect 2596 21088 2648 21140
rect 7656 21088 7708 21140
rect 7748 21088 7800 21140
rect 5356 21020 5408 21072
rect 5724 21063 5776 21072
rect 5724 21029 5733 21063
rect 5733 21029 5767 21063
rect 5767 21029 5776 21063
rect 5724 21020 5776 21029
rect 1768 20952 1820 21004
rect 7104 20952 7156 21004
rect 7656 20952 7708 21004
rect 9220 21088 9272 21140
rect 9404 21020 9456 21072
rect 9680 21020 9732 21072
rect 11336 21088 11388 21140
rect 11888 21088 11940 21140
rect 12164 21088 12216 21140
rect 12900 21088 12952 21140
rect 14004 21088 14056 21140
rect 14188 21088 14240 21140
rect 13912 21020 13964 21072
rect 19156 21088 19208 21140
rect 19248 21088 19300 21140
rect 20168 21088 20220 21140
rect 20352 21088 20404 21140
rect 21640 21088 21692 21140
rect 2228 20927 2280 20936
rect 2228 20893 2237 20927
rect 2237 20893 2271 20927
rect 2271 20893 2280 20927
rect 2228 20884 2280 20893
rect 2320 20884 2372 20936
rect 3608 20884 3660 20936
rect 4068 20884 4120 20936
rect 5908 20927 5960 20936
rect 5908 20893 5917 20927
rect 5917 20893 5951 20927
rect 5951 20893 5960 20927
rect 5908 20884 5960 20893
rect 2136 20791 2188 20800
rect 2136 20757 2145 20791
rect 2145 20757 2179 20791
rect 2179 20757 2188 20791
rect 2136 20748 2188 20757
rect 2596 20816 2648 20868
rect 3700 20748 3752 20800
rect 4804 20816 4856 20868
rect 7380 20884 7432 20936
rect 11520 20995 11572 21004
rect 11520 20961 11529 20995
rect 11529 20961 11563 20995
rect 11563 20961 11572 20995
rect 11520 20952 11572 20961
rect 12532 20995 12584 21004
rect 12532 20961 12541 20995
rect 12541 20961 12575 20995
rect 12575 20961 12584 20995
rect 12532 20952 12584 20961
rect 15568 20995 15620 21004
rect 15568 20961 15577 20995
rect 15577 20961 15611 20995
rect 15611 20961 15620 20995
rect 15568 20952 15620 20961
rect 19616 21020 19668 21072
rect 17224 20995 17276 21004
rect 17224 20961 17233 20995
rect 17233 20961 17267 20995
rect 17267 20961 17276 20995
rect 17224 20952 17276 20961
rect 18052 20995 18104 21004
rect 18052 20961 18061 20995
rect 18061 20961 18095 20995
rect 18095 20961 18104 20995
rect 18052 20952 18104 20961
rect 5540 20748 5592 20800
rect 6460 20748 6512 20800
rect 7104 20748 7156 20800
rect 7656 20816 7708 20868
rect 8116 20816 8168 20868
rect 8392 20816 8444 20868
rect 7472 20748 7524 20800
rect 9312 20884 9364 20936
rect 9496 20816 9548 20868
rect 9772 20816 9824 20868
rect 12072 20884 12124 20936
rect 14740 20884 14792 20936
rect 15384 20884 15436 20936
rect 9404 20748 9456 20800
rect 12624 20748 12676 20800
rect 13912 20791 13964 20800
rect 13912 20757 13921 20791
rect 13921 20757 13955 20791
rect 13955 20757 13964 20791
rect 13912 20748 13964 20757
rect 15660 20816 15712 20868
rect 15844 20927 15896 20936
rect 15844 20893 15878 20927
rect 15878 20893 15896 20927
rect 18880 20952 18932 21004
rect 15844 20884 15896 20893
rect 18420 20884 18472 20936
rect 19892 20927 19944 20936
rect 19892 20893 19901 20927
rect 19901 20893 19935 20927
rect 19935 20893 19944 20927
rect 19892 20884 19944 20893
rect 19984 20927 20036 20936
rect 19984 20893 19993 20927
rect 19993 20893 20027 20927
rect 20027 20893 20036 20927
rect 19984 20884 20036 20893
rect 20996 20884 21048 20936
rect 20720 20816 20772 20868
rect 21916 20816 21968 20868
rect 16396 20748 16448 20800
rect 17316 20791 17368 20800
rect 17316 20757 17325 20791
rect 17325 20757 17359 20791
rect 17359 20757 17368 20791
rect 17316 20748 17368 20757
rect 17408 20791 17460 20800
rect 17408 20757 17417 20791
rect 17417 20757 17451 20791
rect 17451 20757 17460 20791
rect 17408 20748 17460 20757
rect 18604 20791 18656 20800
rect 18604 20757 18613 20791
rect 18613 20757 18647 20791
rect 18647 20757 18656 20791
rect 18604 20748 18656 20757
rect 20812 20748 20864 20800
rect 21456 20748 21508 20800
rect 6548 20646 6600 20698
rect 6612 20646 6664 20698
rect 6676 20646 6728 20698
rect 6740 20646 6792 20698
rect 6804 20646 6856 20698
rect 12146 20646 12198 20698
rect 12210 20646 12262 20698
rect 12274 20646 12326 20698
rect 12338 20646 12390 20698
rect 12402 20646 12454 20698
rect 17744 20646 17796 20698
rect 17808 20646 17860 20698
rect 17872 20646 17924 20698
rect 17936 20646 17988 20698
rect 18000 20646 18052 20698
rect 1768 20587 1820 20596
rect 1768 20553 1777 20587
rect 1777 20553 1811 20587
rect 1811 20553 1820 20587
rect 1768 20544 1820 20553
rect 2228 20544 2280 20596
rect 2136 20476 2188 20528
rect 3240 20544 3292 20596
rect 4068 20544 4120 20596
rect 2596 20408 2648 20460
rect 2872 20451 2924 20460
rect 2872 20417 2890 20451
rect 2890 20417 2924 20451
rect 2872 20408 2924 20417
rect 3424 20476 3476 20528
rect 4712 20519 4764 20528
rect 4712 20485 4721 20519
rect 4721 20485 4755 20519
rect 4755 20485 4764 20519
rect 4712 20476 4764 20485
rect 5908 20544 5960 20596
rect 7748 20587 7800 20596
rect 7748 20553 7757 20587
rect 7757 20553 7791 20587
rect 7791 20553 7800 20587
rect 7748 20544 7800 20553
rect 3700 20408 3752 20460
rect 5080 20451 5132 20460
rect 5080 20417 5114 20451
rect 5114 20417 5132 20451
rect 5080 20408 5132 20417
rect 6460 20476 6512 20528
rect 8024 20476 8076 20528
rect 8576 20476 8628 20528
rect 8852 20544 8904 20596
rect 9496 20544 9548 20596
rect 7472 20408 7524 20460
rect 9680 20451 9732 20460
rect 4436 20340 4488 20392
rect 4712 20340 4764 20392
rect 8024 20340 8076 20392
rect 9680 20417 9689 20451
rect 9689 20417 9723 20451
rect 9723 20417 9732 20451
rect 9680 20408 9732 20417
rect 9956 20451 10008 20460
rect 9956 20417 9990 20451
rect 9990 20417 10008 20451
rect 9956 20408 10008 20417
rect 13636 20544 13688 20596
rect 15660 20587 15712 20596
rect 11980 20408 12032 20460
rect 12532 20476 12584 20528
rect 13452 20476 13504 20528
rect 15660 20553 15669 20587
rect 15669 20553 15703 20587
rect 15703 20553 15712 20587
rect 15660 20544 15712 20553
rect 18604 20544 18656 20596
rect 19708 20587 19760 20596
rect 19708 20553 19717 20587
rect 19717 20553 19751 20587
rect 19751 20553 19760 20587
rect 19708 20544 19760 20553
rect 7564 20272 7616 20324
rect 8484 20272 8536 20324
rect 3148 20204 3200 20256
rect 3240 20247 3292 20256
rect 3240 20213 3249 20247
rect 3249 20213 3283 20247
rect 3283 20213 3292 20247
rect 3240 20204 3292 20213
rect 4160 20204 4212 20256
rect 4988 20204 5040 20256
rect 6000 20204 6052 20256
rect 7840 20247 7892 20256
rect 7840 20213 7849 20247
rect 7849 20213 7883 20247
rect 7883 20213 7892 20247
rect 7840 20204 7892 20213
rect 8300 20204 8352 20256
rect 9220 20204 9272 20256
rect 9680 20272 9732 20324
rect 11152 20272 11204 20324
rect 10324 20204 10376 20256
rect 11244 20204 11296 20256
rect 12716 20408 12768 20460
rect 13820 20451 13872 20460
rect 13820 20417 13829 20451
rect 13829 20417 13863 20451
rect 13863 20417 13872 20451
rect 13820 20408 13872 20417
rect 13912 20408 13964 20460
rect 14556 20408 14608 20460
rect 15752 20476 15804 20528
rect 16304 20476 16356 20528
rect 17960 20476 18012 20528
rect 16948 20408 17000 20460
rect 17224 20451 17276 20460
rect 17224 20417 17233 20451
rect 17233 20417 17267 20451
rect 17267 20417 17276 20451
rect 17224 20408 17276 20417
rect 14280 20204 14332 20256
rect 14740 20340 14792 20392
rect 15936 20383 15988 20392
rect 15936 20349 15945 20383
rect 15945 20349 15979 20383
rect 15979 20349 15988 20383
rect 15936 20340 15988 20349
rect 17132 20340 17184 20392
rect 15292 20272 15344 20324
rect 17684 20340 17736 20392
rect 19064 20340 19116 20392
rect 19616 20408 19668 20460
rect 20352 20476 20404 20528
rect 21180 20544 21232 20596
rect 23388 20476 23440 20528
rect 20904 20408 20956 20460
rect 20996 20408 21048 20460
rect 19248 20383 19300 20392
rect 19248 20349 19257 20383
rect 19257 20349 19291 20383
rect 19291 20349 19300 20383
rect 19248 20340 19300 20349
rect 19984 20340 20036 20392
rect 21640 20408 21692 20460
rect 19524 20272 19576 20324
rect 16304 20204 16356 20256
rect 16488 20247 16540 20256
rect 16488 20213 16497 20247
rect 16497 20213 16531 20247
rect 16531 20213 16540 20247
rect 16488 20204 16540 20213
rect 19064 20204 19116 20256
rect 21640 20315 21692 20324
rect 21640 20281 21649 20315
rect 21649 20281 21683 20315
rect 21683 20281 21692 20315
rect 21640 20272 21692 20281
rect 22100 20383 22152 20392
rect 22100 20349 22109 20383
rect 22109 20349 22143 20383
rect 22143 20349 22152 20383
rect 22100 20340 22152 20349
rect 23020 20408 23072 20460
rect 23296 20408 23348 20460
rect 21180 20204 21232 20256
rect 21272 20204 21324 20256
rect 22008 20204 22060 20256
rect 22284 20204 22336 20256
rect 23020 20247 23072 20256
rect 23020 20213 23029 20247
rect 23029 20213 23063 20247
rect 23063 20213 23072 20247
rect 23020 20204 23072 20213
rect 3749 20102 3801 20154
rect 3813 20102 3865 20154
rect 3877 20102 3929 20154
rect 3941 20102 3993 20154
rect 4005 20102 4057 20154
rect 9347 20102 9399 20154
rect 9411 20102 9463 20154
rect 9475 20102 9527 20154
rect 9539 20102 9591 20154
rect 9603 20102 9655 20154
rect 14945 20102 14997 20154
rect 15009 20102 15061 20154
rect 15073 20102 15125 20154
rect 15137 20102 15189 20154
rect 15201 20102 15253 20154
rect 20543 20102 20595 20154
rect 20607 20102 20659 20154
rect 20671 20102 20723 20154
rect 20735 20102 20787 20154
rect 20799 20102 20851 20154
rect 2872 20000 2924 20052
rect 4620 20000 4672 20052
rect 7012 20000 7064 20052
rect 7196 20043 7248 20052
rect 7196 20009 7205 20043
rect 7205 20009 7239 20043
rect 7239 20009 7248 20043
rect 7196 20000 7248 20009
rect 8024 20043 8076 20052
rect 8024 20009 8033 20043
rect 8033 20009 8067 20043
rect 8067 20009 8076 20043
rect 8024 20000 8076 20009
rect 9772 20043 9824 20052
rect 9772 20009 9781 20043
rect 9781 20009 9815 20043
rect 9815 20009 9824 20043
rect 9772 20000 9824 20009
rect 11060 20000 11112 20052
rect 13544 20000 13596 20052
rect 14096 20043 14148 20052
rect 14096 20009 14105 20043
rect 14105 20009 14139 20043
rect 14139 20009 14148 20043
rect 14096 20000 14148 20009
rect 14832 20000 14884 20052
rect 2596 19932 2648 19984
rect 4896 19932 4948 19984
rect 5080 19975 5132 19984
rect 5080 19941 5089 19975
rect 5089 19941 5123 19975
rect 5123 19941 5132 19975
rect 5080 19932 5132 19941
rect 5540 19932 5592 19984
rect 3148 19864 3200 19916
rect 5264 19907 5316 19916
rect 1584 19796 1636 19848
rect 2228 19796 2280 19848
rect 2780 19796 2832 19848
rect 4620 19839 4672 19848
rect 2872 19703 2924 19712
rect 2872 19669 2881 19703
rect 2881 19669 2915 19703
rect 2915 19669 2924 19703
rect 4620 19805 4629 19839
rect 4629 19805 4663 19839
rect 4663 19805 4672 19839
rect 4620 19796 4672 19805
rect 4804 19796 4856 19848
rect 5264 19873 5273 19907
rect 5273 19873 5307 19907
rect 5307 19873 5316 19907
rect 5264 19864 5316 19873
rect 5908 19864 5960 19916
rect 7564 19932 7616 19984
rect 9680 19932 9732 19984
rect 7196 19864 7248 19916
rect 7748 19907 7800 19916
rect 6184 19796 6236 19848
rect 7288 19796 7340 19848
rect 7748 19873 7757 19907
rect 7757 19873 7791 19907
rect 7791 19873 7800 19907
rect 7748 19864 7800 19873
rect 8668 19907 8720 19916
rect 8668 19873 8677 19907
rect 8677 19873 8711 19907
rect 8711 19873 8720 19907
rect 8668 19864 8720 19873
rect 9220 19864 9272 19916
rect 11520 19932 11572 19984
rect 11336 19864 11388 19916
rect 11888 19907 11940 19916
rect 11888 19873 11897 19907
rect 11897 19873 11931 19907
rect 11931 19873 11940 19907
rect 11888 19864 11940 19873
rect 13084 19907 13136 19916
rect 13084 19873 13093 19907
rect 13093 19873 13127 19907
rect 13127 19873 13136 19907
rect 13084 19864 13136 19873
rect 12072 19796 12124 19848
rect 12808 19839 12860 19848
rect 12808 19805 12817 19839
rect 12817 19805 12851 19839
rect 12851 19805 12860 19839
rect 12808 19796 12860 19805
rect 13636 19796 13688 19848
rect 5080 19728 5132 19780
rect 2872 19660 2924 19669
rect 5816 19660 5868 19712
rect 6368 19703 6420 19712
rect 6368 19669 6377 19703
rect 6377 19669 6411 19703
rect 6411 19669 6420 19703
rect 6368 19660 6420 19669
rect 6920 19660 6972 19712
rect 7932 19728 7984 19780
rect 9772 19728 9824 19780
rect 10140 19728 10192 19780
rect 7564 19703 7616 19712
rect 7564 19669 7573 19703
rect 7573 19669 7607 19703
rect 7607 19669 7616 19703
rect 7564 19660 7616 19669
rect 8392 19703 8444 19712
rect 8392 19669 8401 19703
rect 8401 19669 8435 19703
rect 8435 19669 8444 19703
rect 8392 19660 8444 19669
rect 11152 19660 11204 19712
rect 11428 19660 11480 19712
rect 11796 19703 11848 19712
rect 11796 19669 11805 19703
rect 11805 19669 11839 19703
rect 11839 19669 11848 19703
rect 11796 19660 11848 19669
rect 12072 19660 12124 19712
rect 14004 19932 14056 19984
rect 14556 19907 14608 19916
rect 14556 19873 14565 19907
rect 14565 19873 14599 19907
rect 14599 19873 14608 19907
rect 14556 19864 14608 19873
rect 15016 19864 15068 19916
rect 14188 19796 14240 19848
rect 19156 20000 19208 20052
rect 18604 19864 18656 19916
rect 21456 20000 21508 20052
rect 22560 20000 22612 20052
rect 15660 19839 15712 19848
rect 15660 19805 15669 19839
rect 15669 19805 15703 19839
rect 15703 19805 15712 19839
rect 16396 19839 16448 19848
rect 15660 19796 15712 19805
rect 16396 19805 16405 19839
rect 16405 19805 16439 19839
rect 16439 19805 16448 19839
rect 16396 19796 16448 19805
rect 14372 19728 14424 19780
rect 17132 19796 17184 19848
rect 18144 19839 18196 19848
rect 18144 19805 18153 19839
rect 18153 19805 18187 19839
rect 18187 19805 18196 19839
rect 18144 19796 18196 19805
rect 14188 19660 14240 19712
rect 16304 19703 16356 19712
rect 16304 19669 16313 19703
rect 16313 19669 16347 19703
rect 16347 19669 16356 19703
rect 16304 19660 16356 19669
rect 17684 19728 17736 19780
rect 19708 19907 19760 19916
rect 19708 19873 19720 19907
rect 19720 19873 19754 19907
rect 19754 19873 19760 19907
rect 19708 19864 19760 19873
rect 20996 19864 21048 19916
rect 18972 19796 19024 19848
rect 19340 19796 19392 19848
rect 21180 19839 21232 19848
rect 21180 19805 21189 19839
rect 21189 19805 21223 19839
rect 21223 19805 21232 19839
rect 21180 19796 21232 19805
rect 20904 19728 20956 19780
rect 23572 19796 23624 19848
rect 17592 19660 17644 19712
rect 18236 19703 18288 19712
rect 18236 19669 18245 19703
rect 18245 19669 18279 19703
rect 18279 19669 18288 19703
rect 18236 19660 18288 19669
rect 18604 19703 18656 19712
rect 18604 19669 18613 19703
rect 18613 19669 18647 19703
rect 18647 19669 18656 19703
rect 18604 19660 18656 19669
rect 19616 19660 19668 19712
rect 21088 19703 21140 19712
rect 21088 19669 21097 19703
rect 21097 19669 21131 19703
rect 21131 19669 21140 19703
rect 21088 19660 21140 19669
rect 22100 19660 22152 19712
rect 22560 19703 22612 19712
rect 22560 19669 22569 19703
rect 22569 19669 22603 19703
rect 22603 19669 22612 19703
rect 22560 19660 22612 19669
rect 23020 19703 23072 19712
rect 23020 19669 23029 19703
rect 23029 19669 23063 19703
rect 23063 19669 23072 19703
rect 23020 19660 23072 19669
rect 6548 19558 6600 19610
rect 6612 19558 6664 19610
rect 6676 19558 6728 19610
rect 6740 19558 6792 19610
rect 6804 19558 6856 19610
rect 12146 19558 12198 19610
rect 12210 19558 12262 19610
rect 12274 19558 12326 19610
rect 12338 19558 12390 19610
rect 12402 19558 12454 19610
rect 17744 19558 17796 19610
rect 17808 19558 17860 19610
rect 17872 19558 17924 19610
rect 17936 19558 17988 19610
rect 18000 19558 18052 19610
rect 1492 19456 1544 19508
rect 2780 19456 2832 19508
rect 4160 19388 4212 19440
rect 4344 19431 4396 19440
rect 4344 19397 4353 19431
rect 4353 19397 4387 19431
rect 4387 19397 4396 19431
rect 4344 19388 4396 19397
rect 4896 19499 4948 19508
rect 4896 19465 4905 19499
rect 4905 19465 4939 19499
rect 4939 19465 4948 19499
rect 6368 19499 6420 19508
rect 4896 19456 4948 19465
rect 6368 19465 6377 19499
rect 6377 19465 6411 19499
rect 6411 19465 6420 19499
rect 6368 19456 6420 19465
rect 8116 19456 8168 19508
rect 8392 19456 8444 19508
rect 9772 19456 9824 19508
rect 10048 19499 10100 19508
rect 10048 19465 10057 19499
rect 10057 19465 10091 19499
rect 10091 19465 10100 19499
rect 10048 19456 10100 19465
rect 10324 19499 10376 19508
rect 10324 19465 10333 19499
rect 10333 19465 10367 19499
rect 10367 19465 10376 19499
rect 10324 19456 10376 19465
rect 11612 19456 11664 19508
rect 14096 19456 14148 19508
rect 14372 19499 14424 19508
rect 14372 19465 14381 19499
rect 14381 19465 14415 19499
rect 14415 19465 14424 19499
rect 14372 19456 14424 19465
rect 15200 19456 15252 19508
rect 1584 19320 1636 19372
rect 4436 19363 4488 19372
rect 4160 19295 4212 19304
rect 4160 19261 4169 19295
rect 4169 19261 4203 19295
rect 4203 19261 4212 19295
rect 4160 19252 4212 19261
rect 4436 19329 4445 19363
rect 4445 19329 4479 19363
rect 4479 19329 4488 19363
rect 4436 19320 4488 19329
rect 6000 19363 6052 19372
rect 6000 19329 6009 19363
rect 6009 19329 6043 19363
rect 6043 19329 6052 19363
rect 6000 19320 6052 19329
rect 7012 19388 7064 19440
rect 7196 19388 7248 19440
rect 8852 19388 8904 19440
rect 9220 19363 9272 19372
rect 4712 19252 4764 19304
rect 4804 19252 4856 19304
rect 3148 19184 3200 19236
rect 3424 19184 3476 19236
rect 4252 19184 4304 19236
rect 7012 19252 7064 19304
rect 7472 19252 7524 19304
rect 9220 19329 9229 19363
rect 9229 19329 9263 19363
rect 9263 19329 9272 19363
rect 9220 19320 9272 19329
rect 9864 19320 9916 19372
rect 11060 19388 11112 19440
rect 19248 19456 19300 19508
rect 21272 19456 21324 19508
rect 22284 19499 22336 19508
rect 20628 19388 20680 19440
rect 22284 19465 22293 19499
rect 22293 19465 22327 19499
rect 22327 19465 22336 19499
rect 22284 19456 22336 19465
rect 23204 19456 23256 19508
rect 7748 19295 7800 19304
rect 7748 19261 7760 19295
rect 7760 19261 7794 19295
rect 7794 19261 7800 19295
rect 7748 19252 7800 19261
rect 7932 19252 7984 19304
rect 8668 19252 8720 19304
rect 11152 19363 11204 19372
rect 11152 19329 11161 19363
rect 11161 19329 11195 19363
rect 11195 19329 11204 19363
rect 11152 19320 11204 19329
rect 11520 19363 11572 19372
rect 11520 19329 11529 19363
rect 11529 19329 11563 19363
rect 11563 19329 11572 19363
rect 11520 19320 11572 19329
rect 12440 19320 12492 19372
rect 13452 19363 13504 19372
rect 13452 19329 13461 19363
rect 13461 19329 13495 19363
rect 13495 19329 13504 19363
rect 13452 19320 13504 19329
rect 14004 19363 14056 19372
rect 14004 19329 14013 19363
rect 14013 19329 14047 19363
rect 14047 19329 14056 19363
rect 14004 19320 14056 19329
rect 14832 19363 14884 19372
rect 14832 19329 14841 19363
rect 14841 19329 14875 19363
rect 14875 19329 14884 19363
rect 14832 19320 14884 19329
rect 15660 19320 15712 19372
rect 10784 19295 10836 19304
rect 10784 19261 10793 19295
rect 10793 19261 10827 19295
rect 10827 19261 10836 19295
rect 10784 19252 10836 19261
rect 8852 19184 8904 19236
rect 9864 19184 9916 19236
rect 3516 19116 3568 19168
rect 4528 19116 4580 19168
rect 5816 19159 5868 19168
rect 5816 19125 5825 19159
rect 5825 19125 5859 19159
rect 5859 19125 5868 19159
rect 5816 19116 5868 19125
rect 6184 19159 6236 19168
rect 6184 19125 6193 19159
rect 6193 19125 6227 19159
rect 6227 19125 6236 19159
rect 6184 19116 6236 19125
rect 7012 19116 7064 19168
rect 8392 19116 8444 19168
rect 8668 19116 8720 19168
rect 9036 19116 9088 19168
rect 9128 19116 9180 19168
rect 9956 19116 10008 19168
rect 10508 19116 10560 19168
rect 11796 19184 11848 19236
rect 13820 19252 13872 19304
rect 15016 19295 15068 19304
rect 15016 19261 15025 19295
rect 15025 19261 15059 19295
rect 15059 19261 15068 19295
rect 15016 19252 15068 19261
rect 11244 19116 11296 19168
rect 11520 19116 11572 19168
rect 11704 19159 11756 19168
rect 11704 19125 11713 19159
rect 11713 19125 11747 19159
rect 11747 19125 11756 19159
rect 11704 19116 11756 19125
rect 11980 19116 12032 19168
rect 12440 19116 12492 19168
rect 14280 19184 14332 19236
rect 14464 19159 14516 19168
rect 14464 19125 14473 19159
rect 14473 19125 14507 19159
rect 14507 19125 14516 19159
rect 14832 19184 14884 19236
rect 16212 19252 16264 19304
rect 17040 19320 17092 19372
rect 20904 19363 20956 19372
rect 16856 19252 16908 19304
rect 14464 19116 14516 19125
rect 15292 19116 15344 19168
rect 16212 19159 16264 19168
rect 16212 19125 16221 19159
rect 16221 19125 16255 19159
rect 16255 19125 16264 19159
rect 16212 19116 16264 19125
rect 17500 19252 17552 19304
rect 17592 19295 17644 19304
rect 17592 19261 17604 19295
rect 17604 19261 17638 19295
rect 17638 19261 17644 19295
rect 17592 19252 17644 19261
rect 18604 19252 18656 19304
rect 19156 19252 19208 19304
rect 20904 19329 20913 19363
rect 20913 19329 20947 19363
rect 20947 19329 20956 19363
rect 20904 19320 20956 19329
rect 21364 19320 21416 19372
rect 23664 19388 23716 19440
rect 22192 19363 22244 19372
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 22836 19363 22888 19372
rect 19800 19227 19852 19236
rect 19800 19193 19809 19227
rect 19809 19193 19843 19227
rect 19843 19193 19852 19227
rect 19800 19184 19852 19193
rect 21456 19252 21508 19304
rect 22836 19329 22845 19363
rect 22845 19329 22879 19363
rect 22879 19329 22888 19363
rect 22836 19320 22888 19329
rect 19340 19116 19392 19168
rect 19524 19116 19576 19168
rect 20260 19159 20312 19168
rect 20260 19125 20269 19159
rect 20269 19125 20303 19159
rect 20303 19125 20312 19159
rect 20260 19116 20312 19125
rect 21640 19184 21692 19236
rect 22928 19116 22980 19168
rect 3749 19014 3801 19066
rect 3813 19014 3865 19066
rect 3877 19014 3929 19066
rect 3941 19014 3993 19066
rect 4005 19014 4057 19066
rect 9347 19014 9399 19066
rect 9411 19014 9463 19066
rect 9475 19014 9527 19066
rect 9539 19014 9591 19066
rect 9603 19014 9655 19066
rect 14945 19014 14997 19066
rect 15009 19014 15061 19066
rect 15073 19014 15125 19066
rect 15137 19014 15189 19066
rect 15201 19014 15253 19066
rect 20543 19014 20595 19066
rect 20607 19014 20659 19066
rect 20671 19014 20723 19066
rect 20735 19014 20787 19066
rect 20799 19014 20851 19066
rect 1676 18912 1728 18964
rect 4436 18912 4488 18964
rect 4804 18955 4856 18964
rect 4804 18921 4813 18955
rect 4813 18921 4847 18955
rect 4847 18921 4856 18955
rect 4804 18912 4856 18921
rect 6184 18912 6236 18964
rect 8668 18912 8720 18964
rect 1768 18844 1820 18896
rect 1308 18776 1360 18828
rect 3516 18776 3568 18828
rect 1400 18708 1452 18760
rect 3608 18751 3660 18760
rect 3608 18717 3617 18751
rect 3617 18717 3651 18751
rect 3651 18717 3660 18751
rect 3608 18708 3660 18717
rect 4160 18844 4212 18896
rect 7196 18887 7248 18896
rect 4620 18776 4672 18828
rect 7196 18853 7205 18887
rect 7205 18853 7239 18887
rect 7239 18853 7248 18887
rect 7196 18844 7248 18853
rect 8852 18776 8904 18828
rect 4436 18640 4488 18692
rect 5816 18708 5868 18760
rect 6184 18708 6236 18760
rect 6460 18708 6512 18760
rect 7932 18751 7984 18760
rect 7932 18717 7941 18751
rect 7941 18717 7975 18751
rect 7975 18717 7984 18751
rect 7932 18708 7984 18717
rect 8116 18708 8168 18760
rect 8300 18708 8352 18760
rect 8576 18708 8628 18760
rect 9312 18844 9364 18896
rect 9680 18844 9732 18896
rect 9220 18776 9272 18828
rect 10508 18844 10560 18896
rect 13820 18912 13872 18964
rect 14004 18912 14056 18964
rect 14832 18912 14884 18964
rect 15660 18912 15712 18964
rect 15936 18912 15988 18964
rect 14372 18844 14424 18896
rect 9680 18708 9732 18760
rect 11428 18776 11480 18828
rect 10508 18751 10560 18760
rect 10508 18717 10517 18751
rect 10517 18717 10551 18751
rect 10551 18717 10560 18751
rect 10508 18708 10560 18717
rect 10784 18708 10836 18760
rect 10324 18640 10376 18692
rect 2044 18572 2096 18624
rect 2228 18615 2280 18624
rect 2228 18581 2237 18615
rect 2237 18581 2271 18615
rect 2271 18581 2280 18615
rect 2228 18572 2280 18581
rect 2320 18572 2372 18624
rect 3424 18572 3476 18624
rect 4160 18615 4212 18624
rect 4160 18581 4169 18615
rect 4169 18581 4203 18615
rect 4203 18581 4212 18615
rect 4160 18572 4212 18581
rect 4252 18615 4304 18624
rect 4252 18581 4261 18615
rect 4261 18581 4295 18615
rect 4295 18581 4304 18615
rect 5264 18615 5316 18624
rect 4252 18572 4304 18581
rect 5264 18581 5273 18615
rect 5273 18581 5307 18615
rect 5307 18581 5316 18615
rect 5264 18572 5316 18581
rect 5356 18572 5408 18624
rect 5724 18572 5776 18624
rect 7196 18572 7248 18624
rect 8300 18572 8352 18624
rect 9496 18572 9548 18624
rect 10048 18615 10100 18624
rect 10048 18581 10057 18615
rect 10057 18581 10091 18615
rect 10091 18581 10100 18615
rect 10048 18572 10100 18581
rect 10876 18572 10928 18624
rect 10968 18615 11020 18624
rect 10968 18581 10983 18615
rect 10983 18581 11017 18615
rect 11017 18581 11020 18615
rect 12624 18751 12676 18760
rect 12624 18717 12633 18751
rect 12633 18717 12667 18751
rect 12667 18717 12676 18751
rect 12624 18708 12676 18717
rect 12900 18751 12952 18760
rect 12900 18717 12909 18751
rect 12909 18717 12943 18751
rect 12943 18717 12952 18751
rect 12900 18708 12952 18717
rect 12440 18640 12492 18692
rect 13268 18640 13320 18692
rect 13452 18776 13504 18828
rect 17592 18912 17644 18964
rect 17776 18912 17828 18964
rect 18236 18912 18288 18964
rect 19892 18912 19944 18964
rect 20444 18912 20496 18964
rect 17408 18844 17460 18896
rect 19340 18844 19392 18896
rect 20352 18844 20404 18896
rect 14096 18708 14148 18760
rect 17592 18776 17644 18828
rect 21916 18912 21968 18964
rect 23112 18912 23164 18964
rect 15476 18751 15528 18760
rect 15476 18717 15485 18751
rect 15485 18717 15519 18751
rect 15519 18717 15528 18751
rect 15476 18708 15528 18717
rect 17132 18708 17184 18760
rect 17776 18751 17828 18760
rect 17776 18717 17785 18751
rect 17785 18717 17819 18751
rect 17819 18717 17828 18751
rect 17776 18708 17828 18717
rect 10968 18572 11020 18581
rect 12532 18615 12584 18624
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 12992 18572 13044 18624
rect 16304 18640 16356 18692
rect 17868 18640 17920 18692
rect 17500 18572 17552 18624
rect 18696 18708 18748 18760
rect 19064 18751 19116 18760
rect 19064 18717 19073 18751
rect 19073 18717 19107 18751
rect 19107 18717 19116 18751
rect 19064 18708 19116 18717
rect 19892 18708 19944 18760
rect 18328 18640 18380 18692
rect 19524 18640 19576 18692
rect 19616 18640 19668 18692
rect 21180 18708 21232 18760
rect 22652 18751 22704 18760
rect 22652 18717 22661 18751
rect 22661 18717 22695 18751
rect 22695 18717 22704 18751
rect 22652 18708 22704 18717
rect 22836 18751 22888 18760
rect 22836 18717 22845 18751
rect 22845 18717 22879 18751
rect 22879 18717 22888 18751
rect 22836 18708 22888 18717
rect 21824 18640 21876 18692
rect 18236 18572 18288 18624
rect 18972 18572 19024 18624
rect 21272 18572 21324 18624
rect 22008 18615 22060 18624
rect 22008 18581 22017 18615
rect 22017 18581 22051 18615
rect 22051 18581 22060 18615
rect 22008 18572 22060 18581
rect 6548 18470 6600 18522
rect 6612 18470 6664 18522
rect 6676 18470 6728 18522
rect 6740 18470 6792 18522
rect 6804 18470 6856 18522
rect 12146 18470 12198 18522
rect 12210 18470 12262 18522
rect 12274 18470 12326 18522
rect 12338 18470 12390 18522
rect 12402 18470 12454 18522
rect 17744 18470 17796 18522
rect 17808 18470 17860 18522
rect 17872 18470 17924 18522
rect 17936 18470 17988 18522
rect 18000 18470 18052 18522
rect 1676 18411 1728 18420
rect 1676 18377 1685 18411
rect 1685 18377 1719 18411
rect 1719 18377 1728 18411
rect 1676 18368 1728 18377
rect 2228 18368 2280 18420
rect 1584 18300 1636 18352
rect 4712 18368 4764 18420
rect 6000 18368 6052 18420
rect 1768 18275 1820 18284
rect 1768 18241 1777 18275
rect 1777 18241 1811 18275
rect 1811 18241 1820 18275
rect 1768 18232 1820 18241
rect 2320 18275 2372 18284
rect 2320 18241 2354 18275
rect 2354 18241 2372 18275
rect 2320 18232 2372 18241
rect 6092 18300 6144 18352
rect 7104 18300 7156 18352
rect 8668 18300 8720 18352
rect 7012 18275 7064 18284
rect 1308 18096 1360 18148
rect 4620 18164 4672 18216
rect 6276 18164 6328 18216
rect 7012 18241 7021 18275
rect 7021 18241 7055 18275
rect 7055 18241 7064 18275
rect 7012 18232 7064 18241
rect 7380 18232 7432 18284
rect 10048 18368 10100 18420
rect 11704 18368 11756 18420
rect 12808 18411 12860 18420
rect 12808 18377 12817 18411
rect 12817 18377 12851 18411
rect 12851 18377 12860 18411
rect 12808 18368 12860 18377
rect 14464 18368 14516 18420
rect 13360 18300 13412 18352
rect 17040 18411 17092 18420
rect 17040 18377 17049 18411
rect 17049 18377 17083 18411
rect 17083 18377 17092 18411
rect 17040 18368 17092 18377
rect 17132 18368 17184 18420
rect 18512 18368 18564 18420
rect 10968 18232 11020 18284
rect 7104 18164 7156 18216
rect 9128 18164 9180 18216
rect 9496 18164 9548 18216
rect 9772 18164 9824 18216
rect 4528 18096 4580 18148
rect 10784 18139 10836 18148
rect 3240 18028 3292 18080
rect 4436 18028 4488 18080
rect 6368 18071 6420 18080
rect 6368 18037 6377 18071
rect 6377 18037 6411 18071
rect 6411 18037 6420 18071
rect 6368 18028 6420 18037
rect 10784 18105 10793 18139
rect 10793 18105 10827 18139
rect 10827 18105 10836 18139
rect 10784 18096 10836 18105
rect 11244 18096 11296 18148
rect 11704 18232 11756 18284
rect 11980 18275 12032 18284
rect 11980 18241 11989 18275
rect 11989 18241 12023 18275
rect 12023 18241 12032 18275
rect 12900 18275 12952 18284
rect 11980 18232 12032 18241
rect 12900 18241 12909 18275
rect 12909 18241 12943 18275
rect 12943 18241 12952 18275
rect 12900 18232 12952 18241
rect 14004 18275 14056 18284
rect 14004 18241 14013 18275
rect 14013 18241 14047 18275
rect 14047 18241 14056 18275
rect 14004 18232 14056 18241
rect 11520 18164 11572 18216
rect 13084 18164 13136 18216
rect 13268 18164 13320 18216
rect 15476 18300 15528 18352
rect 19248 18368 19300 18420
rect 20904 18368 20956 18420
rect 21548 18411 21600 18420
rect 21548 18377 21557 18411
rect 21557 18377 21591 18411
rect 21591 18377 21600 18411
rect 21548 18368 21600 18377
rect 19432 18300 19484 18352
rect 20260 18300 20312 18352
rect 20444 18300 20496 18352
rect 18512 18232 18564 18284
rect 17132 18207 17184 18216
rect 17132 18173 17141 18207
rect 17141 18173 17175 18207
rect 17175 18173 17184 18207
rect 17132 18164 17184 18173
rect 17224 18207 17276 18216
rect 17224 18173 17233 18207
rect 17233 18173 17267 18207
rect 17267 18173 17276 18207
rect 17224 18164 17276 18173
rect 17684 18164 17736 18216
rect 19708 18232 19760 18284
rect 21272 18275 21324 18284
rect 21272 18241 21281 18275
rect 21281 18241 21315 18275
rect 21315 18241 21324 18275
rect 21272 18232 21324 18241
rect 21456 18232 21508 18284
rect 19064 18207 19116 18216
rect 8208 18028 8260 18080
rect 8576 18028 8628 18080
rect 13268 18071 13320 18080
rect 13268 18037 13277 18071
rect 13277 18037 13311 18071
rect 13311 18037 13320 18071
rect 13268 18028 13320 18037
rect 13544 18028 13596 18080
rect 14188 18028 14240 18080
rect 14832 18028 14884 18080
rect 17040 18096 17092 18148
rect 18604 18028 18656 18080
rect 19064 18173 19073 18207
rect 19073 18173 19107 18207
rect 19107 18173 19116 18207
rect 19064 18164 19116 18173
rect 19432 18164 19484 18216
rect 19616 18207 19668 18216
rect 19616 18173 19625 18207
rect 19625 18173 19659 18207
rect 19659 18173 19668 18207
rect 19616 18164 19668 18173
rect 22468 18368 22520 18420
rect 22928 18368 22980 18420
rect 22928 18164 22980 18216
rect 19156 18028 19208 18080
rect 19524 18071 19576 18080
rect 19524 18037 19533 18071
rect 19533 18037 19567 18071
rect 19567 18037 19576 18071
rect 19524 18028 19576 18037
rect 19616 18028 19668 18080
rect 20352 18028 20404 18080
rect 21272 18028 21324 18080
rect 23020 18071 23072 18080
rect 23020 18037 23029 18071
rect 23029 18037 23063 18071
rect 23063 18037 23072 18071
rect 23020 18028 23072 18037
rect 3749 17926 3801 17978
rect 3813 17926 3865 17978
rect 3877 17926 3929 17978
rect 3941 17926 3993 17978
rect 4005 17926 4057 17978
rect 9347 17926 9399 17978
rect 9411 17926 9463 17978
rect 9475 17926 9527 17978
rect 9539 17926 9591 17978
rect 9603 17926 9655 17978
rect 14945 17926 14997 17978
rect 15009 17926 15061 17978
rect 15073 17926 15125 17978
rect 15137 17926 15189 17978
rect 15201 17926 15253 17978
rect 20543 17926 20595 17978
rect 20607 17926 20659 17978
rect 20671 17926 20723 17978
rect 20735 17926 20787 17978
rect 20799 17926 20851 17978
rect 2504 17824 2556 17876
rect 3608 17824 3660 17876
rect 5264 17824 5316 17876
rect 6460 17867 6512 17876
rect 6460 17833 6469 17867
rect 6469 17833 6503 17867
rect 6503 17833 6512 17867
rect 6460 17824 6512 17833
rect 6920 17824 6972 17876
rect 7380 17824 7432 17876
rect 2964 17756 3016 17808
rect 4528 17756 4580 17808
rect 8668 17799 8720 17808
rect 8668 17765 8677 17799
rect 8677 17765 8711 17799
rect 8711 17765 8720 17799
rect 8668 17756 8720 17765
rect 9036 17756 9088 17808
rect 1584 17688 1636 17740
rect 2044 17663 2096 17672
rect 2044 17629 2078 17663
rect 2078 17629 2096 17663
rect 2044 17620 2096 17629
rect 3424 17663 3476 17672
rect 3424 17629 3433 17663
rect 3433 17629 3467 17663
rect 3467 17629 3476 17663
rect 3424 17620 3476 17629
rect 3608 17620 3660 17672
rect 4528 17620 4580 17672
rect 8024 17688 8076 17740
rect 12716 17824 12768 17876
rect 12900 17867 12952 17876
rect 12900 17833 12909 17867
rect 12909 17833 12943 17867
rect 12943 17833 12952 17867
rect 12900 17824 12952 17833
rect 14096 17867 14148 17876
rect 14096 17833 14105 17867
rect 14105 17833 14139 17867
rect 14139 17833 14148 17867
rect 14096 17824 14148 17833
rect 14188 17824 14240 17876
rect 17316 17867 17368 17876
rect 12624 17756 12676 17808
rect 13360 17756 13412 17808
rect 6552 17663 6604 17672
rect 6552 17629 6561 17663
rect 6561 17629 6595 17663
rect 6595 17629 6604 17663
rect 6552 17620 6604 17629
rect 3148 17552 3200 17604
rect 4344 17552 4396 17604
rect 4804 17595 4856 17604
rect 4804 17561 4813 17595
rect 4813 17561 4847 17595
rect 4847 17561 4856 17595
rect 4804 17552 4856 17561
rect 6368 17552 6420 17604
rect 4896 17484 4948 17536
rect 7564 17620 7616 17672
rect 7840 17663 7892 17672
rect 7840 17629 7849 17663
rect 7849 17629 7883 17663
rect 7883 17629 7892 17663
rect 7840 17620 7892 17629
rect 9220 17620 9272 17672
rect 13268 17688 13320 17740
rect 14372 17756 14424 17808
rect 14556 17756 14608 17808
rect 11060 17620 11112 17672
rect 12072 17620 12124 17672
rect 17316 17833 17325 17867
rect 17325 17833 17359 17867
rect 17359 17833 17368 17867
rect 17316 17824 17368 17833
rect 19248 17867 19300 17876
rect 17684 17756 17736 17808
rect 19248 17833 19257 17867
rect 19257 17833 19291 17867
rect 19291 17833 19300 17867
rect 19248 17824 19300 17833
rect 19340 17756 19392 17808
rect 14832 17688 14884 17740
rect 15476 17688 15528 17740
rect 15200 17620 15252 17672
rect 16212 17688 16264 17740
rect 17224 17688 17276 17740
rect 18880 17688 18932 17740
rect 21180 17824 21232 17876
rect 22100 17824 22152 17876
rect 20628 17756 20680 17808
rect 21456 17731 21508 17740
rect 16488 17620 16540 17672
rect 9036 17552 9088 17604
rect 10324 17595 10376 17604
rect 10324 17561 10358 17595
rect 10358 17561 10376 17595
rect 10324 17552 10376 17561
rect 14832 17552 14884 17604
rect 16580 17552 16632 17604
rect 16948 17552 17000 17604
rect 19432 17620 19484 17672
rect 21456 17697 21465 17731
rect 21465 17697 21499 17731
rect 21499 17697 21508 17731
rect 21456 17688 21508 17697
rect 20720 17663 20772 17672
rect 20720 17629 20729 17663
rect 20729 17629 20763 17663
rect 20763 17629 20772 17663
rect 20720 17620 20772 17629
rect 21548 17620 21600 17672
rect 23296 17620 23348 17672
rect 8208 17484 8260 17536
rect 8668 17484 8720 17536
rect 10600 17484 10652 17536
rect 13360 17527 13412 17536
rect 13360 17493 13369 17527
rect 13369 17493 13403 17527
rect 13403 17493 13412 17527
rect 13360 17484 13412 17493
rect 14556 17527 14608 17536
rect 14556 17493 14565 17527
rect 14565 17493 14599 17527
rect 14599 17493 14608 17527
rect 14556 17484 14608 17493
rect 14740 17484 14792 17536
rect 16672 17527 16724 17536
rect 16672 17493 16681 17527
rect 16681 17493 16715 17527
rect 16715 17493 16724 17527
rect 16672 17484 16724 17493
rect 18144 17552 18196 17604
rect 20536 17552 20588 17604
rect 18236 17484 18288 17536
rect 19064 17527 19116 17536
rect 19064 17493 19073 17527
rect 19073 17493 19107 17527
rect 19107 17493 19116 17527
rect 19064 17484 19116 17493
rect 20720 17484 20772 17536
rect 22928 17527 22980 17536
rect 22928 17493 22937 17527
rect 22937 17493 22971 17527
rect 22971 17493 22980 17527
rect 22928 17484 22980 17493
rect 6548 17382 6600 17434
rect 6612 17382 6664 17434
rect 6676 17382 6728 17434
rect 6740 17382 6792 17434
rect 6804 17382 6856 17434
rect 12146 17382 12198 17434
rect 12210 17382 12262 17434
rect 12274 17382 12326 17434
rect 12338 17382 12390 17434
rect 12402 17382 12454 17434
rect 17744 17382 17796 17434
rect 17808 17382 17860 17434
rect 17872 17382 17924 17434
rect 17936 17382 17988 17434
rect 18000 17382 18052 17434
rect 1400 17280 1452 17332
rect 3516 17280 3568 17332
rect 4160 17280 4212 17332
rect 4988 17280 5040 17332
rect 6276 17280 6328 17332
rect 7104 17280 7156 17332
rect 8024 17280 8076 17332
rect 8208 17280 8260 17332
rect 8392 17280 8444 17332
rect 8852 17323 8904 17332
rect 1584 17212 1636 17264
rect 2596 17187 2648 17196
rect 4804 17212 4856 17264
rect 2596 17153 2614 17187
rect 2614 17153 2648 17187
rect 2596 17144 2648 17153
rect 4712 17144 4764 17196
rect 3148 17119 3200 17128
rect 3148 17085 3157 17119
rect 3157 17085 3191 17119
rect 3191 17085 3200 17119
rect 3884 17119 3936 17128
rect 3148 17076 3200 17085
rect 3884 17085 3893 17119
rect 3893 17085 3927 17119
rect 3927 17085 3936 17119
rect 3884 17076 3936 17085
rect 4436 17076 4488 17128
rect 5908 17212 5960 17264
rect 6644 17212 6696 17264
rect 5632 17144 5684 17196
rect 6736 17187 6788 17196
rect 6736 17153 6745 17187
rect 6745 17153 6779 17187
rect 6779 17153 6788 17187
rect 6736 17144 6788 17153
rect 7380 17212 7432 17264
rect 8852 17289 8861 17323
rect 8861 17289 8895 17323
rect 8895 17289 8904 17323
rect 8852 17280 8904 17289
rect 9680 17323 9732 17332
rect 9680 17289 9689 17323
rect 9689 17289 9723 17323
rect 9723 17289 9732 17323
rect 9680 17280 9732 17289
rect 6368 17076 6420 17128
rect 8300 17187 8352 17196
rect 11520 17280 11572 17332
rect 11612 17280 11664 17332
rect 8300 17153 8318 17187
rect 8318 17153 8352 17187
rect 8300 17144 8352 17153
rect 8852 17144 8904 17196
rect 9128 17144 9180 17196
rect 11060 17187 11112 17196
rect 11060 17153 11069 17187
rect 11069 17153 11103 17187
rect 11103 17153 11112 17187
rect 11060 17144 11112 17153
rect 11704 17187 11756 17196
rect 11704 17153 11713 17187
rect 11713 17153 11747 17187
rect 11747 17153 11756 17187
rect 11704 17144 11756 17153
rect 12992 17212 13044 17264
rect 13360 17280 13412 17332
rect 14004 17280 14056 17332
rect 14556 17280 14608 17332
rect 13820 17187 13872 17196
rect 8668 17076 8720 17128
rect 13820 17153 13829 17187
rect 13829 17153 13863 17187
rect 13863 17153 13872 17187
rect 13820 17144 13872 17153
rect 14372 17144 14424 17196
rect 14648 17187 14700 17196
rect 14648 17153 14657 17187
rect 14657 17153 14691 17187
rect 14691 17153 14700 17187
rect 14648 17144 14700 17153
rect 15476 17212 15528 17264
rect 17132 17280 17184 17332
rect 18696 17280 18748 17332
rect 19524 17280 19576 17332
rect 16764 17212 16816 17264
rect 18144 17212 18196 17264
rect 15200 17144 15252 17196
rect 16304 17144 16356 17196
rect 16948 17144 17000 17196
rect 4252 17008 4304 17060
rect 2596 16940 2648 16992
rect 7012 17008 7064 17060
rect 14556 17076 14608 17128
rect 5724 16940 5776 16992
rect 7932 16940 7984 16992
rect 9128 16940 9180 16992
rect 11520 16940 11572 16992
rect 11796 16940 11848 16992
rect 13912 16940 13964 16992
rect 16488 17008 16540 17060
rect 16396 16940 16448 16992
rect 17316 16983 17368 16992
rect 17316 16949 17325 16983
rect 17325 16949 17359 16983
rect 17359 16949 17368 16983
rect 17316 16940 17368 16949
rect 18420 16940 18472 16992
rect 18972 17076 19024 17128
rect 19800 17144 19852 17196
rect 22100 17280 22152 17332
rect 22284 17323 22336 17332
rect 22284 17289 22293 17323
rect 22293 17289 22327 17323
rect 22327 17289 22336 17323
rect 22284 17280 22336 17289
rect 21272 17255 21324 17264
rect 21272 17221 21281 17255
rect 21281 17221 21315 17255
rect 21315 17221 21324 17255
rect 21272 17212 21324 17221
rect 22836 17255 22888 17264
rect 22836 17221 22845 17255
rect 22845 17221 22879 17255
rect 22879 17221 22888 17255
rect 22836 17212 22888 17221
rect 19248 17008 19300 17060
rect 19800 17008 19852 17060
rect 19524 16940 19576 16992
rect 19708 16983 19760 16992
rect 19708 16949 19717 16983
rect 19717 16949 19751 16983
rect 19751 16949 19760 16983
rect 19708 16940 19760 16949
rect 20260 16940 20312 16992
rect 21088 17008 21140 17060
rect 22928 17076 22980 17128
rect 20904 16940 20956 16992
rect 23204 16940 23256 16992
rect 3749 16838 3801 16890
rect 3813 16838 3865 16890
rect 3877 16838 3929 16890
rect 3941 16838 3993 16890
rect 4005 16838 4057 16890
rect 9347 16838 9399 16890
rect 9411 16838 9463 16890
rect 9475 16838 9527 16890
rect 9539 16838 9591 16890
rect 9603 16838 9655 16890
rect 14945 16838 14997 16890
rect 15009 16838 15061 16890
rect 15073 16838 15125 16890
rect 15137 16838 15189 16890
rect 15201 16838 15253 16890
rect 20543 16838 20595 16890
rect 20607 16838 20659 16890
rect 20671 16838 20723 16890
rect 20735 16838 20787 16890
rect 20799 16838 20851 16890
rect 3608 16736 3660 16788
rect 3148 16600 3200 16652
rect 4528 16600 4580 16652
rect 4804 16736 4856 16788
rect 6184 16736 6236 16788
rect 6736 16736 6788 16788
rect 6920 16779 6972 16788
rect 6920 16745 6929 16779
rect 6929 16745 6963 16779
rect 6963 16745 6972 16779
rect 6920 16736 6972 16745
rect 7288 16736 7340 16788
rect 8668 16736 8720 16788
rect 10416 16736 10468 16788
rect 11520 16736 11572 16788
rect 7012 16668 7064 16720
rect 6644 16643 6696 16652
rect 6644 16609 6653 16643
rect 6653 16609 6687 16643
rect 6687 16609 6696 16643
rect 8576 16668 8628 16720
rect 6644 16600 6696 16609
rect 7656 16643 7708 16652
rect 7656 16609 7665 16643
rect 7665 16609 7699 16643
rect 7699 16609 7708 16643
rect 7656 16600 7708 16609
rect 8300 16600 8352 16652
rect 9220 16643 9272 16652
rect 9220 16609 9229 16643
rect 9229 16609 9263 16643
rect 9263 16609 9272 16643
rect 9220 16600 9272 16609
rect 15476 16736 15528 16788
rect 16304 16779 16356 16788
rect 16304 16745 16313 16779
rect 16313 16745 16347 16779
rect 16347 16745 16356 16779
rect 16304 16736 16356 16745
rect 18144 16736 18196 16788
rect 19248 16668 19300 16720
rect 19524 16668 19576 16720
rect 1860 16464 1912 16516
rect 2872 16575 2924 16584
rect 2872 16541 2881 16575
rect 2881 16541 2915 16575
rect 2915 16541 2924 16575
rect 2872 16532 2924 16541
rect 2964 16464 3016 16516
rect 1768 16439 1820 16448
rect 1768 16405 1777 16439
rect 1777 16405 1811 16439
rect 1811 16405 1820 16439
rect 1768 16396 1820 16405
rect 2320 16396 2372 16448
rect 5356 16532 5408 16584
rect 6460 16575 6512 16584
rect 6460 16541 6469 16575
rect 6469 16541 6503 16575
rect 6503 16541 6512 16575
rect 6460 16532 6512 16541
rect 7288 16532 7340 16584
rect 7840 16532 7892 16584
rect 8484 16575 8536 16584
rect 8484 16541 8493 16575
rect 8493 16541 8527 16575
rect 8527 16541 8536 16575
rect 8484 16532 8536 16541
rect 11244 16532 11296 16584
rect 8116 16464 8168 16516
rect 12072 16464 12124 16516
rect 3332 16396 3384 16448
rect 3700 16396 3752 16448
rect 6092 16439 6144 16448
rect 6092 16405 6101 16439
rect 6101 16405 6135 16439
rect 6135 16405 6144 16439
rect 7104 16439 7156 16448
rect 6092 16396 6144 16405
rect 7104 16405 7113 16439
rect 7113 16405 7147 16439
rect 7147 16405 7156 16439
rect 7104 16396 7156 16405
rect 8208 16439 8260 16448
rect 8208 16405 8217 16439
rect 8217 16405 8251 16439
rect 8251 16405 8260 16439
rect 8208 16396 8260 16405
rect 9496 16396 9548 16448
rect 9680 16439 9732 16448
rect 9680 16405 9689 16439
rect 9689 16405 9723 16439
rect 9723 16405 9732 16439
rect 9680 16396 9732 16405
rect 9864 16396 9916 16448
rect 10048 16396 10100 16448
rect 11704 16439 11756 16448
rect 11704 16405 11713 16439
rect 11713 16405 11747 16439
rect 11747 16405 11756 16439
rect 11704 16396 11756 16405
rect 13544 16575 13596 16584
rect 13544 16541 13562 16575
rect 13562 16541 13596 16575
rect 13544 16532 13596 16541
rect 14556 16532 14608 16584
rect 16672 16532 16724 16584
rect 17316 16532 17368 16584
rect 19708 16600 19760 16652
rect 21456 16643 21508 16652
rect 19248 16575 19300 16584
rect 19248 16541 19257 16575
rect 19257 16541 19291 16575
rect 19291 16541 19300 16575
rect 19984 16575 20036 16584
rect 19248 16532 19300 16541
rect 19984 16541 19993 16575
rect 19993 16541 20027 16575
rect 20027 16541 20036 16575
rect 19984 16532 20036 16541
rect 20536 16532 20588 16584
rect 20904 16532 20956 16584
rect 21456 16609 21465 16643
rect 21465 16609 21499 16643
rect 21499 16609 21508 16643
rect 21456 16600 21508 16609
rect 15752 16464 15804 16516
rect 13820 16396 13872 16448
rect 14096 16439 14148 16448
rect 14096 16405 14105 16439
rect 14105 16405 14139 16439
rect 14139 16405 14148 16439
rect 14096 16396 14148 16405
rect 17132 16507 17184 16516
rect 17132 16473 17141 16507
rect 17141 16473 17175 16507
rect 17175 16473 17184 16507
rect 17132 16464 17184 16473
rect 17592 16464 17644 16516
rect 16856 16396 16908 16448
rect 18880 16396 18932 16448
rect 21180 16507 21232 16516
rect 21180 16473 21189 16507
rect 21189 16473 21223 16507
rect 21223 16473 21232 16507
rect 21180 16464 21232 16473
rect 21732 16507 21784 16516
rect 21732 16473 21766 16507
rect 21766 16473 21784 16507
rect 21732 16464 21784 16473
rect 23388 16532 23440 16584
rect 20352 16396 20404 16448
rect 21088 16439 21140 16448
rect 21088 16405 21097 16439
rect 21097 16405 21131 16439
rect 21131 16405 21140 16439
rect 21088 16396 21140 16405
rect 22744 16396 22796 16448
rect 22928 16439 22980 16448
rect 22928 16405 22937 16439
rect 22937 16405 22971 16439
rect 22971 16405 22980 16439
rect 22928 16396 22980 16405
rect 6548 16294 6600 16346
rect 6612 16294 6664 16346
rect 6676 16294 6728 16346
rect 6740 16294 6792 16346
rect 6804 16294 6856 16346
rect 12146 16294 12198 16346
rect 12210 16294 12262 16346
rect 12274 16294 12326 16346
rect 12338 16294 12390 16346
rect 12402 16294 12454 16346
rect 17744 16294 17796 16346
rect 17808 16294 17860 16346
rect 17872 16294 17924 16346
rect 17936 16294 17988 16346
rect 18000 16294 18052 16346
rect 2872 16235 2924 16244
rect 2872 16201 2881 16235
rect 2881 16201 2915 16235
rect 2915 16201 2924 16235
rect 2872 16192 2924 16201
rect 3700 16235 3752 16244
rect 3700 16201 3709 16235
rect 3709 16201 3743 16235
rect 3743 16201 3752 16235
rect 3700 16192 3752 16201
rect 4252 16124 4304 16176
rect 5540 16192 5592 16244
rect 6368 16124 6420 16176
rect 2044 16056 2096 16108
rect 1492 16031 1544 16040
rect 1492 15997 1501 16031
rect 1501 15997 1535 16031
rect 1535 15997 1544 16031
rect 1492 15988 1544 15997
rect 3148 16056 3200 16108
rect 5172 16056 5224 16108
rect 3240 16031 3292 16040
rect 3240 15997 3249 16031
rect 3249 15997 3283 16031
rect 3283 15997 3292 16031
rect 3240 15988 3292 15997
rect 2872 15920 2924 15972
rect 5632 16056 5684 16108
rect 6184 16099 6236 16108
rect 6184 16065 6193 16099
rect 6193 16065 6227 16099
rect 6227 16065 6236 16099
rect 6184 16056 6236 16065
rect 8300 16192 8352 16244
rect 9496 16235 9548 16244
rect 9496 16201 9505 16235
rect 9505 16201 9539 16235
rect 9539 16201 9548 16235
rect 9496 16192 9548 16201
rect 9864 16192 9916 16244
rect 7748 16124 7800 16176
rect 9128 16099 9180 16108
rect 11244 16124 11296 16176
rect 5448 15988 5500 16040
rect 6460 15988 6512 16040
rect 9128 16065 9146 16099
rect 9146 16065 9180 16099
rect 9128 16056 9180 16065
rect 11060 16099 11112 16108
rect 12072 16192 12124 16244
rect 14556 16192 14608 16244
rect 14648 16192 14700 16244
rect 14096 16124 14148 16176
rect 11060 16065 11078 16099
rect 11078 16065 11112 16099
rect 11060 16056 11112 16065
rect 11704 15988 11756 16040
rect 13820 16056 13872 16108
rect 21732 16192 21784 16244
rect 17132 16124 17184 16176
rect 22744 16167 22796 16176
rect 22744 16133 22753 16167
rect 22753 16133 22787 16167
rect 22787 16133 22796 16167
rect 22744 16124 22796 16133
rect 16396 16056 16448 16108
rect 16764 16056 16816 16108
rect 18236 16056 18288 16108
rect 18788 16099 18840 16108
rect 18788 16065 18797 16099
rect 18797 16065 18831 16099
rect 18831 16065 18840 16099
rect 18788 16056 18840 16065
rect 19248 16099 19300 16108
rect 19248 16065 19257 16099
rect 19257 16065 19291 16099
rect 19291 16065 19300 16099
rect 19248 16056 19300 16065
rect 19340 16056 19392 16108
rect 21548 16056 21600 16108
rect 22468 16099 22520 16108
rect 18696 16031 18748 16040
rect 5632 15920 5684 15972
rect 16488 15963 16540 15972
rect 16488 15929 16497 15963
rect 16497 15929 16531 15963
rect 16531 15929 16540 15963
rect 16488 15920 16540 15929
rect 16856 15963 16908 15972
rect 16856 15929 16865 15963
rect 16865 15929 16899 15963
rect 16899 15929 16908 15963
rect 16856 15920 16908 15929
rect 18696 15997 18705 16031
rect 18705 15997 18739 16031
rect 18739 15997 18748 16031
rect 18696 15988 18748 15997
rect 19800 15988 19852 16040
rect 22468 16065 22477 16099
rect 22477 16065 22511 16099
rect 22511 16065 22520 16099
rect 22468 16056 22520 16065
rect 22560 16099 22612 16108
rect 22560 16065 22569 16099
rect 22569 16065 22603 16099
rect 22603 16065 22612 16099
rect 22560 16056 22612 16065
rect 19064 15920 19116 15972
rect 6920 15852 6972 15904
rect 7932 15895 7984 15904
rect 7932 15861 7941 15895
rect 7941 15861 7975 15895
rect 7975 15861 7984 15895
rect 7932 15852 7984 15861
rect 10416 15852 10468 15904
rect 11980 15852 12032 15904
rect 13452 15852 13504 15904
rect 15384 15852 15436 15904
rect 15844 15895 15896 15904
rect 15844 15861 15853 15895
rect 15853 15861 15887 15895
rect 15887 15861 15896 15895
rect 15844 15852 15896 15861
rect 16948 15895 17000 15904
rect 16948 15861 16957 15895
rect 16957 15861 16991 15895
rect 16991 15861 17000 15895
rect 16948 15852 17000 15861
rect 17684 15852 17736 15904
rect 17960 15852 18012 15904
rect 18512 15852 18564 15904
rect 18880 15852 18932 15904
rect 20444 15852 20496 15904
rect 21456 15895 21508 15904
rect 21456 15861 21465 15895
rect 21465 15861 21499 15895
rect 21499 15861 21508 15895
rect 21456 15852 21508 15861
rect 21548 15852 21600 15904
rect 23112 15895 23164 15904
rect 23112 15861 23121 15895
rect 23121 15861 23155 15895
rect 23155 15861 23164 15895
rect 23112 15852 23164 15861
rect 3749 15750 3801 15802
rect 3813 15750 3865 15802
rect 3877 15750 3929 15802
rect 3941 15750 3993 15802
rect 4005 15750 4057 15802
rect 9347 15750 9399 15802
rect 9411 15750 9463 15802
rect 9475 15750 9527 15802
rect 9539 15750 9591 15802
rect 9603 15750 9655 15802
rect 14945 15750 14997 15802
rect 15009 15750 15061 15802
rect 15073 15750 15125 15802
rect 15137 15750 15189 15802
rect 15201 15750 15253 15802
rect 20543 15750 20595 15802
rect 20607 15750 20659 15802
rect 20671 15750 20723 15802
rect 20735 15750 20787 15802
rect 20799 15750 20851 15802
rect 2044 15691 2096 15700
rect 2044 15657 2053 15691
rect 2053 15657 2087 15691
rect 2087 15657 2096 15691
rect 2044 15648 2096 15657
rect 2320 15648 2372 15700
rect 3056 15648 3108 15700
rect 3240 15648 3292 15700
rect 1492 15512 1544 15564
rect 2044 15512 2096 15564
rect 4896 15648 4948 15700
rect 5172 15648 5224 15700
rect 10140 15648 10192 15700
rect 6460 15555 6512 15564
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 6460 15521 6469 15555
rect 6469 15521 6503 15555
rect 6503 15521 6512 15555
rect 6460 15512 6512 15521
rect 7104 15512 7156 15564
rect 9864 15555 9916 15564
rect 9864 15521 9873 15555
rect 9873 15521 9907 15555
rect 9907 15521 9916 15555
rect 9864 15512 9916 15521
rect 11060 15648 11112 15700
rect 13452 15691 13504 15700
rect 13452 15657 13461 15691
rect 13461 15657 13495 15691
rect 13495 15657 13504 15691
rect 13452 15648 13504 15657
rect 13636 15691 13688 15700
rect 13636 15657 13645 15691
rect 13645 15657 13679 15691
rect 13679 15657 13688 15691
rect 13636 15648 13688 15657
rect 15752 15691 15804 15700
rect 10416 15623 10468 15632
rect 10416 15589 10425 15623
rect 10425 15589 10459 15623
rect 10459 15589 10468 15623
rect 10416 15580 10468 15589
rect 11428 15580 11480 15632
rect 15752 15657 15761 15691
rect 15761 15657 15795 15691
rect 15795 15657 15804 15691
rect 15752 15648 15804 15657
rect 17960 15648 18012 15700
rect 18052 15648 18104 15700
rect 18788 15648 18840 15700
rect 19984 15691 20036 15700
rect 19984 15657 19993 15691
rect 19993 15657 20027 15691
rect 20027 15657 20036 15691
rect 19984 15648 20036 15657
rect 22100 15648 22152 15700
rect 22652 15648 22704 15700
rect 11612 15512 11664 15564
rect 4160 15444 4212 15496
rect 4344 15444 4396 15496
rect 5448 15444 5500 15496
rect 7748 15444 7800 15496
rect 9772 15444 9824 15496
rect 10048 15487 10100 15496
rect 10048 15453 10057 15487
rect 10057 15453 10091 15487
rect 10091 15453 10100 15487
rect 10048 15444 10100 15453
rect 10140 15444 10192 15496
rect 11336 15487 11388 15496
rect 11336 15453 11345 15487
rect 11345 15453 11379 15487
rect 11379 15453 11388 15487
rect 11336 15444 11388 15453
rect 13820 15512 13872 15564
rect 18052 15555 18104 15564
rect 18052 15521 18061 15555
rect 18061 15521 18095 15555
rect 18095 15521 18104 15555
rect 18052 15512 18104 15521
rect 18328 15580 18380 15632
rect 18972 15580 19024 15632
rect 19248 15512 19300 15564
rect 19800 15512 19852 15564
rect 20904 15580 20956 15632
rect 21272 15580 21324 15632
rect 20352 15555 20404 15564
rect 20352 15521 20361 15555
rect 20361 15521 20395 15555
rect 20395 15521 20404 15555
rect 20352 15512 20404 15521
rect 20996 15512 21048 15564
rect 13636 15444 13688 15496
rect 15844 15444 15896 15496
rect 1768 15376 1820 15428
rect 7932 15376 7984 15428
rect 4896 15351 4948 15360
rect 4896 15317 4905 15351
rect 4905 15317 4939 15351
rect 4939 15317 4948 15351
rect 4896 15308 4948 15317
rect 5908 15308 5960 15360
rect 6000 15351 6052 15360
rect 6000 15317 6009 15351
rect 6009 15317 6043 15351
rect 6043 15317 6052 15351
rect 6000 15308 6052 15317
rect 6368 15308 6420 15360
rect 6920 15308 6972 15360
rect 8576 15351 8628 15360
rect 8576 15317 8585 15351
rect 8585 15317 8619 15351
rect 8619 15317 8628 15351
rect 8576 15308 8628 15317
rect 10876 15351 10928 15360
rect 10876 15317 10885 15351
rect 10885 15317 10919 15351
rect 10919 15317 10928 15351
rect 10876 15308 10928 15317
rect 14464 15376 14516 15428
rect 18144 15444 18196 15496
rect 18880 15487 18932 15496
rect 18880 15453 18889 15487
rect 18889 15453 18923 15487
rect 18923 15453 18932 15487
rect 18880 15444 18932 15453
rect 20904 15487 20956 15496
rect 20904 15453 20913 15487
rect 20913 15453 20947 15487
rect 20947 15453 20956 15487
rect 20904 15444 20956 15453
rect 15568 15308 15620 15360
rect 16580 15376 16632 15428
rect 17592 15376 17644 15428
rect 17684 15376 17736 15428
rect 21272 15444 21324 15496
rect 22744 15444 22796 15496
rect 22836 15444 22888 15496
rect 19524 15351 19576 15360
rect 19524 15317 19533 15351
rect 19533 15317 19567 15351
rect 19567 15317 19576 15351
rect 19524 15308 19576 15317
rect 19616 15351 19668 15360
rect 19616 15317 19625 15351
rect 19625 15317 19659 15351
rect 19659 15317 19668 15351
rect 19616 15308 19668 15317
rect 22376 15376 22428 15428
rect 21272 15308 21324 15360
rect 22192 15308 22244 15360
rect 22928 15351 22980 15360
rect 22928 15317 22937 15351
rect 22937 15317 22971 15351
rect 22971 15317 22980 15351
rect 22928 15308 22980 15317
rect 6548 15206 6600 15258
rect 6612 15206 6664 15258
rect 6676 15206 6728 15258
rect 6740 15206 6792 15258
rect 6804 15206 6856 15258
rect 12146 15206 12198 15258
rect 12210 15206 12262 15258
rect 12274 15206 12326 15258
rect 12338 15206 12390 15258
rect 12402 15206 12454 15258
rect 17744 15206 17796 15258
rect 17808 15206 17860 15258
rect 17872 15206 17924 15258
rect 17936 15206 17988 15258
rect 18000 15206 18052 15258
rect 1400 15147 1452 15156
rect 1400 15113 1409 15147
rect 1409 15113 1443 15147
rect 1443 15113 1452 15147
rect 1400 15104 1452 15113
rect 4252 15147 4304 15156
rect 4252 15113 4261 15147
rect 4261 15113 4295 15147
rect 4295 15113 4304 15147
rect 4252 15104 4304 15113
rect 5448 15104 5500 15156
rect 7564 15104 7616 15156
rect 8116 15104 8168 15156
rect 11612 15147 11664 15156
rect 11612 15113 11621 15147
rect 11621 15113 11655 15147
rect 11655 15113 11664 15147
rect 11612 15104 11664 15113
rect 16488 15104 16540 15156
rect 18696 15104 18748 15156
rect 19340 15147 19392 15156
rect 19340 15113 19349 15147
rect 19349 15113 19383 15147
rect 19383 15113 19392 15147
rect 19340 15104 19392 15113
rect 19616 15104 19668 15156
rect 20904 15147 20956 15156
rect 20904 15113 20913 15147
rect 20913 15113 20947 15147
rect 20947 15113 20956 15147
rect 20904 15104 20956 15113
rect 21272 15104 21324 15156
rect 22192 15147 22244 15156
rect 22192 15113 22201 15147
rect 22201 15113 22235 15147
rect 22235 15113 22244 15147
rect 22192 15104 22244 15113
rect 23480 15104 23532 15156
rect 2044 14968 2096 15020
rect 2872 15011 2924 15020
rect 2872 14977 2881 15011
rect 2881 14977 2915 15011
rect 2915 14977 2924 15011
rect 2872 14968 2924 14977
rect 2964 14968 3016 15020
rect 4436 15036 4488 15088
rect 4988 15036 5040 15088
rect 5172 15036 5224 15088
rect 7656 15036 7708 15088
rect 11244 15036 11296 15088
rect 14096 15079 14148 15088
rect 14096 15045 14105 15079
rect 14105 15045 14139 15079
rect 14139 15045 14148 15079
rect 14096 15036 14148 15045
rect 14832 15036 14884 15088
rect 22100 15079 22152 15088
rect 22100 15045 22109 15079
rect 22109 15045 22143 15079
rect 22143 15045 22152 15079
rect 22100 15036 22152 15045
rect 5632 14968 5684 15020
rect 5724 15011 5776 15020
rect 5724 14977 5733 15011
rect 5733 14977 5767 15011
rect 5767 14977 5776 15011
rect 5724 14968 5776 14977
rect 6920 14968 6972 15020
rect 7012 14968 7064 15020
rect 9036 14968 9088 15020
rect 11060 14968 11112 15020
rect 11980 14968 12032 15020
rect 12900 14968 12952 15020
rect 13820 14968 13872 15020
rect 15384 14968 15436 15020
rect 16488 15011 16540 15020
rect 2412 14764 2464 14816
rect 7748 14943 7800 14952
rect 4252 14832 4304 14884
rect 7748 14909 7757 14943
rect 7757 14909 7791 14943
rect 7791 14909 7800 14943
rect 7748 14900 7800 14909
rect 8760 14900 8812 14952
rect 9404 14943 9456 14952
rect 9404 14909 9410 14943
rect 9410 14909 9444 14943
rect 9444 14909 9456 14943
rect 9404 14900 9456 14909
rect 9680 14900 9732 14952
rect 14832 14900 14884 14952
rect 16488 14977 16497 15011
rect 16497 14977 16531 15011
rect 16531 14977 16540 15011
rect 16488 14968 16540 14977
rect 17040 14900 17092 14952
rect 18144 14968 18196 15020
rect 18512 15011 18564 15020
rect 18512 14977 18521 15011
rect 18521 14977 18555 15011
rect 18555 14977 18564 15011
rect 18512 14968 18564 14977
rect 19432 15011 19484 15020
rect 19432 14977 19441 15011
rect 19441 14977 19475 15011
rect 19475 14977 19484 15011
rect 19432 14968 19484 14977
rect 19892 15011 19944 15020
rect 19892 14977 19901 15011
rect 19901 14977 19935 15011
rect 19935 14977 19944 15011
rect 19892 14968 19944 14977
rect 21180 14968 21232 15020
rect 22376 14968 22428 15020
rect 23204 14968 23256 15020
rect 18328 14943 18380 14952
rect 6460 14832 6512 14884
rect 14188 14875 14240 14884
rect 4620 14764 4672 14816
rect 5632 14764 5684 14816
rect 11060 14807 11112 14816
rect 11060 14773 11069 14807
rect 11069 14773 11103 14807
rect 11103 14773 11112 14807
rect 11060 14764 11112 14773
rect 11152 14807 11204 14816
rect 11152 14773 11161 14807
rect 11161 14773 11195 14807
rect 11195 14773 11204 14807
rect 14188 14841 14197 14875
rect 14197 14841 14231 14875
rect 14231 14841 14240 14875
rect 14188 14832 14240 14841
rect 11152 14764 11204 14773
rect 13544 14764 13596 14816
rect 14004 14764 14056 14816
rect 15568 14807 15620 14816
rect 15568 14773 15577 14807
rect 15577 14773 15611 14807
rect 15611 14773 15620 14807
rect 15568 14764 15620 14773
rect 15844 14807 15896 14816
rect 15844 14773 15853 14807
rect 15853 14773 15887 14807
rect 15887 14773 15896 14807
rect 15844 14764 15896 14773
rect 18328 14909 18337 14943
rect 18337 14909 18371 14943
rect 18371 14909 18380 14943
rect 18328 14900 18380 14909
rect 19156 14943 19208 14952
rect 19156 14909 19165 14943
rect 19165 14909 19199 14943
rect 19199 14909 19208 14943
rect 19156 14900 19208 14909
rect 20996 14900 21048 14952
rect 21456 14943 21508 14952
rect 21456 14909 21465 14943
rect 21465 14909 21499 14943
rect 21499 14909 21508 14943
rect 21456 14900 21508 14909
rect 22652 14900 22704 14952
rect 18880 14832 18932 14884
rect 19616 14764 19668 14816
rect 22100 14764 22152 14816
rect 3749 14662 3801 14714
rect 3813 14662 3865 14714
rect 3877 14662 3929 14714
rect 3941 14662 3993 14714
rect 4005 14662 4057 14714
rect 9347 14662 9399 14714
rect 9411 14662 9463 14714
rect 9475 14662 9527 14714
rect 9539 14662 9591 14714
rect 9603 14662 9655 14714
rect 14945 14662 14997 14714
rect 15009 14662 15061 14714
rect 15073 14662 15125 14714
rect 15137 14662 15189 14714
rect 15201 14662 15253 14714
rect 20543 14662 20595 14714
rect 20607 14662 20659 14714
rect 20671 14662 20723 14714
rect 20735 14662 20787 14714
rect 20799 14662 20851 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 1952 14560 2004 14612
rect 2412 14603 2464 14612
rect 2412 14569 2421 14603
rect 2421 14569 2455 14603
rect 2455 14569 2464 14603
rect 2412 14560 2464 14569
rect 2688 14603 2740 14612
rect 2688 14569 2697 14603
rect 2697 14569 2731 14603
rect 2731 14569 2740 14603
rect 2688 14560 2740 14569
rect 2964 14603 3016 14612
rect 2964 14569 2973 14603
rect 2973 14569 3007 14603
rect 3007 14569 3016 14603
rect 2964 14560 3016 14569
rect 2136 14492 2188 14544
rect 1584 14356 1636 14408
rect 1952 14399 2004 14408
rect 1952 14365 1961 14399
rect 1961 14365 1995 14399
rect 1995 14365 2004 14399
rect 1952 14356 2004 14365
rect 5632 14560 5684 14612
rect 5724 14560 5776 14612
rect 4620 14467 4672 14476
rect 4620 14433 4629 14467
rect 4629 14433 4663 14467
rect 4663 14433 4672 14467
rect 4620 14424 4672 14433
rect 4988 14467 5040 14476
rect 3240 14356 3292 14408
rect 4160 14356 4212 14408
rect 4988 14433 4997 14467
rect 4997 14433 5031 14467
rect 5031 14433 5040 14467
rect 4988 14424 5040 14433
rect 7564 14467 7616 14476
rect 7564 14433 7573 14467
rect 7573 14433 7607 14467
rect 7607 14433 7616 14467
rect 7564 14424 7616 14433
rect 5724 14356 5776 14408
rect 6460 14356 6512 14408
rect 9220 14560 9272 14612
rect 10140 14603 10192 14612
rect 10140 14569 10149 14603
rect 10149 14569 10183 14603
rect 10183 14569 10192 14603
rect 10140 14560 10192 14569
rect 10876 14560 10928 14612
rect 12900 14560 12952 14612
rect 15936 14603 15988 14612
rect 15936 14569 15945 14603
rect 15945 14569 15979 14603
rect 15979 14569 15988 14603
rect 15936 14560 15988 14569
rect 17592 14603 17644 14612
rect 17592 14569 17601 14603
rect 17601 14569 17635 14603
rect 17635 14569 17644 14603
rect 17592 14560 17644 14569
rect 19524 14560 19576 14612
rect 19892 14560 19944 14612
rect 22192 14560 22244 14612
rect 23664 14560 23716 14612
rect 5632 14288 5684 14340
rect 6000 14220 6052 14272
rect 6276 14220 6328 14272
rect 7288 14220 7340 14272
rect 7840 14263 7892 14272
rect 7840 14229 7842 14263
rect 7842 14229 7876 14263
rect 7876 14229 7892 14263
rect 7840 14220 7892 14229
rect 8576 14424 8628 14476
rect 8852 14356 8904 14408
rect 9588 14356 9640 14408
rect 16028 14492 16080 14544
rect 11152 14467 11204 14476
rect 11152 14433 11161 14467
rect 11161 14433 11195 14467
rect 11195 14433 11204 14467
rect 11152 14424 11204 14433
rect 14832 14424 14884 14476
rect 10232 14399 10284 14408
rect 10232 14365 10241 14399
rect 10241 14365 10275 14399
rect 10275 14365 10284 14399
rect 10232 14356 10284 14365
rect 11336 14356 11388 14408
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12115 14399
rect 12115 14365 12124 14399
rect 12072 14356 12124 14365
rect 12624 14356 12676 14408
rect 12900 14399 12952 14408
rect 12900 14365 12909 14399
rect 12909 14365 12943 14399
rect 12943 14365 12952 14399
rect 12900 14356 12952 14365
rect 14740 14399 14792 14408
rect 14740 14365 14749 14399
rect 14749 14365 14783 14399
rect 14783 14365 14792 14399
rect 14740 14356 14792 14365
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 15844 14356 15896 14408
rect 19156 14424 19208 14476
rect 18512 14356 18564 14408
rect 20076 14356 20128 14408
rect 20352 14399 20404 14408
rect 20352 14365 20370 14399
rect 20370 14365 20404 14399
rect 20352 14356 20404 14365
rect 20720 14356 20772 14408
rect 20996 14424 21048 14476
rect 20904 14399 20956 14408
rect 20904 14365 20913 14399
rect 20913 14365 20947 14399
rect 20947 14365 20956 14399
rect 20904 14356 20956 14365
rect 22008 14356 22060 14408
rect 23112 14399 23164 14408
rect 23112 14365 23121 14399
rect 23121 14365 23155 14399
rect 23155 14365 23164 14399
rect 23112 14356 23164 14365
rect 11796 14288 11848 14340
rect 13912 14288 13964 14340
rect 14464 14288 14516 14340
rect 18880 14288 18932 14340
rect 19156 14288 19208 14340
rect 11428 14263 11480 14272
rect 11428 14229 11437 14263
rect 11437 14229 11471 14263
rect 11471 14229 11480 14263
rect 11428 14220 11480 14229
rect 12808 14263 12860 14272
rect 12808 14229 12817 14263
rect 12817 14229 12851 14263
rect 12851 14229 12860 14263
rect 12808 14220 12860 14229
rect 13728 14220 13780 14272
rect 14924 14220 14976 14272
rect 18604 14263 18656 14272
rect 18604 14229 18613 14263
rect 18613 14229 18647 14263
rect 18647 14229 18656 14263
rect 18604 14220 18656 14229
rect 19432 14220 19484 14272
rect 19984 14220 20036 14272
rect 20168 14220 20220 14272
rect 21732 14220 21784 14272
rect 22284 14220 22336 14272
rect 22652 14263 22704 14272
rect 22652 14229 22661 14263
rect 22661 14229 22695 14263
rect 22695 14229 22704 14263
rect 22652 14220 22704 14229
rect 6548 14118 6600 14170
rect 6612 14118 6664 14170
rect 6676 14118 6728 14170
rect 6740 14118 6792 14170
rect 6804 14118 6856 14170
rect 12146 14118 12198 14170
rect 12210 14118 12262 14170
rect 12274 14118 12326 14170
rect 12338 14118 12390 14170
rect 12402 14118 12454 14170
rect 17744 14118 17796 14170
rect 17808 14118 17860 14170
rect 17872 14118 17924 14170
rect 17936 14118 17988 14170
rect 18000 14118 18052 14170
rect 1952 14016 2004 14068
rect 5172 14016 5224 14068
rect 5724 14059 5776 14068
rect 5724 14025 5733 14059
rect 5733 14025 5767 14059
rect 5767 14025 5776 14059
rect 5724 14016 5776 14025
rect 6368 14016 6420 14068
rect 7288 14016 7340 14068
rect 8024 14016 8076 14068
rect 9128 14016 9180 14068
rect 2872 13948 2924 14000
rect 2504 13880 2556 13932
rect 3516 13880 3568 13932
rect 4252 13880 4304 13932
rect 4988 13948 5040 14000
rect 6092 13948 6144 14000
rect 8116 13948 8168 14000
rect 4896 13880 4948 13932
rect 5080 13880 5132 13932
rect 5816 13880 5868 13932
rect 6000 13923 6052 13932
rect 6000 13889 6009 13923
rect 6009 13889 6043 13923
rect 6043 13889 6052 13923
rect 6000 13880 6052 13889
rect 6460 13880 6512 13932
rect 7472 13923 7524 13932
rect 7472 13889 7481 13923
rect 7481 13889 7515 13923
rect 7515 13889 7524 13923
rect 7472 13880 7524 13889
rect 7840 13880 7892 13932
rect 8576 13923 8628 13932
rect 8576 13889 8585 13923
rect 8585 13889 8619 13923
rect 8619 13889 8628 13923
rect 8576 13880 8628 13889
rect 9128 13880 9180 13932
rect 11060 14016 11112 14068
rect 14096 14016 14148 14068
rect 15476 14016 15528 14068
rect 16672 14016 16724 14068
rect 11336 13948 11388 14000
rect 11428 13948 11480 14000
rect 9956 13923 10008 13932
rect 9956 13889 9965 13923
rect 9965 13889 9999 13923
rect 9999 13889 10008 13923
rect 9956 13880 10008 13889
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 11152 13923 11204 13932
rect 11152 13889 11161 13923
rect 11161 13889 11195 13923
rect 11195 13889 11204 13923
rect 11152 13880 11204 13889
rect 11244 13880 11296 13932
rect 13820 13948 13872 14000
rect 16488 13991 16540 14000
rect 16488 13957 16497 13991
rect 16497 13957 16531 13991
rect 16531 13957 16540 13991
rect 16488 13948 16540 13957
rect 13728 13880 13780 13932
rect 14924 13923 14976 13932
rect 14924 13889 14958 13923
rect 14958 13889 14976 13923
rect 14924 13880 14976 13889
rect 16304 13923 16356 13932
rect 16304 13889 16313 13923
rect 16313 13889 16347 13923
rect 16347 13889 16356 13923
rect 16304 13880 16356 13889
rect 16396 13880 16448 13932
rect 19156 14016 19208 14068
rect 19340 14016 19392 14068
rect 20076 14016 20128 14068
rect 17684 13880 17736 13932
rect 18144 13880 18196 13932
rect 19064 13880 19116 13932
rect 20720 13948 20772 14000
rect 21272 13948 21324 14000
rect 20076 13880 20128 13932
rect 22100 14059 22152 14068
rect 22100 14025 22109 14059
rect 22109 14025 22143 14059
rect 22143 14025 22152 14059
rect 22100 14016 22152 14025
rect 22652 14016 22704 14068
rect 22560 13948 22612 14000
rect 2872 13855 2924 13864
rect 2872 13821 2881 13855
rect 2881 13821 2915 13855
rect 2915 13821 2924 13855
rect 2872 13812 2924 13821
rect 1676 13744 1728 13796
rect 5448 13812 5500 13864
rect 1952 13719 2004 13728
rect 1952 13685 1961 13719
rect 1961 13685 1995 13719
rect 1995 13685 2004 13719
rect 1952 13676 2004 13685
rect 6184 13744 6236 13796
rect 6276 13744 6328 13796
rect 8024 13812 8076 13864
rect 9680 13744 9732 13796
rect 10876 13812 10928 13864
rect 15752 13812 15804 13864
rect 18420 13855 18472 13864
rect 18420 13821 18429 13855
rect 18429 13821 18463 13855
rect 18463 13821 18472 13855
rect 18420 13812 18472 13821
rect 21640 13880 21692 13932
rect 22192 13880 22244 13932
rect 22284 13880 22336 13932
rect 5816 13719 5868 13728
rect 5816 13685 5825 13719
rect 5825 13685 5859 13719
rect 5859 13685 5868 13719
rect 5816 13676 5868 13685
rect 10968 13676 11020 13728
rect 12440 13676 12492 13728
rect 12900 13719 12952 13728
rect 12900 13685 12909 13719
rect 12909 13685 12943 13719
rect 12943 13685 12952 13719
rect 12900 13676 12952 13685
rect 15384 13676 15436 13728
rect 22560 13812 22612 13864
rect 16028 13719 16080 13728
rect 16028 13685 16037 13719
rect 16037 13685 16071 13719
rect 16071 13685 16080 13719
rect 16028 13676 16080 13685
rect 16396 13676 16448 13728
rect 16580 13676 16632 13728
rect 21456 13676 21508 13728
rect 22836 13744 22888 13796
rect 22376 13676 22428 13728
rect 22744 13676 22796 13728
rect 22928 13719 22980 13728
rect 22928 13685 22937 13719
rect 22937 13685 22971 13719
rect 22971 13685 22980 13719
rect 22928 13676 22980 13685
rect 3749 13574 3801 13626
rect 3813 13574 3865 13626
rect 3877 13574 3929 13626
rect 3941 13574 3993 13626
rect 4005 13574 4057 13626
rect 9347 13574 9399 13626
rect 9411 13574 9463 13626
rect 9475 13574 9527 13626
rect 9539 13574 9591 13626
rect 9603 13574 9655 13626
rect 14945 13574 14997 13626
rect 15009 13574 15061 13626
rect 15073 13574 15125 13626
rect 15137 13574 15189 13626
rect 15201 13574 15253 13626
rect 20543 13574 20595 13626
rect 20607 13574 20659 13626
rect 20671 13574 20723 13626
rect 20735 13574 20787 13626
rect 20799 13574 20851 13626
rect 2504 13472 2556 13524
rect 5632 13515 5684 13524
rect 5080 13404 5132 13456
rect 3884 13379 3936 13388
rect 3884 13345 3893 13379
rect 3893 13345 3927 13379
rect 3927 13345 3936 13379
rect 3884 13336 3936 13345
rect 5632 13481 5641 13515
rect 5641 13481 5675 13515
rect 5675 13481 5684 13515
rect 5632 13472 5684 13481
rect 7012 13515 7064 13524
rect 7012 13481 7021 13515
rect 7021 13481 7055 13515
rect 7055 13481 7064 13515
rect 7012 13472 7064 13481
rect 10508 13472 10560 13524
rect 12072 13472 12124 13524
rect 14372 13472 14424 13524
rect 14740 13472 14792 13524
rect 16304 13472 16356 13524
rect 19616 13472 19668 13524
rect 9956 13404 10008 13456
rect 10232 13404 10284 13456
rect 11980 13404 12032 13456
rect 9496 13379 9548 13388
rect 9496 13345 9505 13379
rect 9505 13345 9539 13379
rect 9539 13345 9548 13379
rect 9496 13336 9548 13345
rect 9588 13336 9640 13388
rect 18788 13379 18840 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 2044 13268 2096 13320
rect 2872 13268 2924 13320
rect 4160 13311 4212 13320
rect 4160 13277 4169 13311
rect 4169 13277 4203 13311
rect 4203 13277 4212 13311
rect 4160 13268 4212 13277
rect 4252 13268 4304 13320
rect 6092 13268 6144 13320
rect 6368 13311 6420 13320
rect 6368 13277 6377 13311
rect 6377 13277 6411 13311
rect 6411 13277 6420 13311
rect 7104 13311 7156 13320
rect 6368 13268 6420 13277
rect 7104 13277 7113 13311
rect 7113 13277 7147 13311
rect 7147 13277 7156 13311
rect 7104 13268 7156 13277
rect 7196 13268 7248 13320
rect 8944 13268 8996 13320
rect 10140 13268 10192 13320
rect 18788 13345 18797 13379
rect 18797 13345 18831 13379
rect 18831 13345 18840 13379
rect 18788 13336 18840 13345
rect 19064 13379 19116 13388
rect 19064 13345 19073 13379
rect 19073 13345 19107 13379
rect 19107 13345 19116 13379
rect 19064 13336 19116 13345
rect 1952 13200 2004 13252
rect 2136 13132 2188 13184
rect 7748 13200 7800 13252
rect 11888 13268 11940 13320
rect 12440 13268 12492 13320
rect 13820 13268 13872 13320
rect 14740 13311 14792 13320
rect 14740 13277 14749 13311
rect 14749 13277 14783 13311
rect 14783 13277 14792 13311
rect 14740 13268 14792 13277
rect 15752 13268 15804 13320
rect 16304 13268 16356 13320
rect 16948 13268 17000 13320
rect 17132 13268 17184 13320
rect 10600 13200 10652 13252
rect 12808 13243 12860 13252
rect 4988 13175 5040 13184
rect 4988 13141 4997 13175
rect 4997 13141 5031 13175
rect 5031 13141 5040 13175
rect 4988 13132 5040 13141
rect 5816 13132 5868 13184
rect 8208 13132 8260 13184
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 9680 13175 9732 13184
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 9772 13175 9824 13184
rect 9772 13141 9781 13175
rect 9781 13141 9815 13175
rect 9815 13141 9824 13175
rect 9772 13132 9824 13141
rect 11152 13132 11204 13184
rect 11704 13132 11756 13184
rect 12808 13209 12842 13243
rect 12842 13209 12860 13243
rect 12808 13200 12860 13209
rect 19984 13311 20036 13320
rect 19984 13277 19993 13311
rect 19993 13277 20027 13311
rect 20027 13277 20036 13311
rect 19984 13268 20036 13277
rect 21180 13404 21232 13456
rect 22468 13472 22520 13524
rect 22836 13515 22888 13524
rect 22836 13481 22845 13515
rect 22845 13481 22879 13515
rect 22879 13481 22888 13515
rect 22836 13472 22888 13481
rect 23756 13472 23808 13524
rect 21088 13379 21140 13388
rect 21088 13345 21097 13379
rect 21097 13345 21131 13379
rect 21131 13345 21140 13379
rect 21088 13336 21140 13345
rect 21272 13379 21324 13388
rect 21272 13345 21281 13379
rect 21281 13345 21315 13379
rect 21315 13345 21324 13379
rect 21272 13336 21324 13345
rect 22652 13268 22704 13320
rect 23112 13311 23164 13320
rect 23112 13277 23121 13311
rect 23121 13277 23155 13311
rect 23155 13277 23164 13311
rect 23112 13268 23164 13277
rect 21364 13200 21416 13252
rect 22008 13200 22060 13252
rect 22928 13200 22980 13252
rect 16212 13175 16264 13184
rect 16212 13141 16221 13175
rect 16221 13141 16255 13175
rect 16255 13141 16264 13175
rect 16212 13132 16264 13141
rect 18236 13132 18288 13184
rect 18328 13132 18380 13184
rect 20260 13132 20312 13184
rect 20444 13175 20496 13184
rect 20444 13141 20453 13175
rect 20453 13141 20487 13175
rect 20487 13141 20496 13175
rect 20444 13132 20496 13141
rect 21824 13132 21876 13184
rect 6548 13030 6600 13082
rect 6612 13030 6664 13082
rect 6676 13030 6728 13082
rect 6740 13030 6792 13082
rect 6804 13030 6856 13082
rect 12146 13030 12198 13082
rect 12210 13030 12262 13082
rect 12274 13030 12326 13082
rect 12338 13030 12390 13082
rect 12402 13030 12454 13082
rect 17744 13030 17796 13082
rect 17808 13030 17860 13082
rect 17872 13030 17924 13082
rect 17936 13030 17988 13082
rect 18000 13030 18052 13082
rect 2504 12928 2556 12980
rect 3516 12971 3568 12980
rect 3516 12937 3525 12971
rect 3525 12937 3559 12971
rect 3559 12937 3568 12971
rect 3516 12928 3568 12937
rect 6000 12928 6052 12980
rect 6460 12928 6512 12980
rect 9956 12928 10008 12980
rect 10140 12971 10192 12980
rect 10140 12937 10149 12971
rect 10149 12937 10183 12971
rect 10183 12937 10192 12971
rect 10140 12928 10192 12937
rect 12072 12928 12124 12980
rect 12532 12928 12584 12980
rect 15292 12928 15344 12980
rect 2872 12860 2924 12912
rect 3148 12792 3200 12844
rect 4620 12860 4672 12912
rect 5816 12903 5868 12912
rect 5816 12869 5840 12903
rect 5840 12869 5868 12903
rect 5816 12860 5868 12869
rect 6184 12860 6236 12912
rect 3884 12792 3936 12844
rect 5356 12792 5408 12844
rect 7104 12860 7156 12912
rect 7748 12860 7800 12912
rect 4252 12724 4304 12776
rect 5724 12724 5776 12776
rect 8116 12835 8168 12844
rect 8576 12860 8628 12912
rect 9588 12860 9640 12912
rect 8116 12801 8134 12835
rect 8134 12801 8168 12835
rect 8116 12792 8168 12801
rect 8852 12835 8904 12844
rect 8852 12801 8861 12835
rect 8861 12801 8895 12835
rect 8895 12801 8904 12835
rect 8852 12792 8904 12801
rect 4344 12656 4396 12708
rect 8760 12724 8812 12776
rect 11612 12860 11664 12912
rect 14372 12903 14424 12912
rect 11520 12792 11572 12844
rect 13820 12792 13872 12844
rect 14372 12869 14381 12903
rect 14381 12869 14415 12903
rect 14415 12869 14424 12903
rect 14372 12860 14424 12869
rect 16028 12860 16080 12912
rect 14648 12792 14700 12844
rect 15476 12792 15528 12844
rect 18512 12928 18564 12980
rect 18604 12928 18656 12980
rect 16580 12792 16632 12844
rect 18144 12860 18196 12912
rect 20076 12928 20128 12980
rect 21088 12928 21140 12980
rect 21824 12971 21876 12980
rect 21824 12937 21833 12971
rect 21833 12937 21867 12971
rect 21867 12937 21876 12971
rect 21824 12928 21876 12937
rect 22652 12971 22704 12980
rect 22652 12937 22661 12971
rect 22661 12937 22695 12971
rect 22695 12937 22704 12971
rect 22652 12928 22704 12937
rect 21272 12860 21324 12912
rect 6368 12656 6420 12708
rect 4436 12631 4488 12640
rect 4436 12597 4445 12631
rect 4445 12597 4479 12631
rect 4479 12597 4488 12631
rect 4436 12588 4488 12597
rect 6460 12588 6512 12640
rect 7472 12588 7524 12640
rect 11980 12767 12032 12776
rect 9036 12656 9088 12708
rect 11980 12733 11989 12767
rect 11989 12733 12023 12767
rect 12023 12733 12032 12767
rect 11980 12724 12032 12733
rect 12072 12767 12124 12776
rect 12072 12733 12081 12767
rect 12081 12733 12115 12767
rect 12115 12733 12124 12767
rect 12072 12724 12124 12733
rect 14004 12724 14056 12776
rect 14188 12767 14240 12776
rect 14188 12733 14197 12767
rect 14197 12733 14231 12767
rect 14231 12733 14240 12767
rect 14188 12724 14240 12733
rect 15384 12767 15436 12776
rect 11152 12656 11204 12708
rect 12624 12656 12676 12708
rect 15384 12733 15393 12767
rect 15393 12733 15427 12767
rect 15427 12733 15436 12767
rect 15384 12724 15436 12733
rect 16856 12767 16908 12776
rect 16856 12733 16865 12767
rect 16865 12733 16899 12767
rect 16899 12733 16908 12767
rect 16856 12724 16908 12733
rect 17316 12724 17368 12776
rect 19708 12792 19760 12844
rect 21548 12792 21600 12844
rect 21732 12792 21784 12844
rect 22376 12792 22428 12844
rect 22836 12792 22888 12844
rect 19892 12724 19944 12776
rect 21824 12724 21876 12776
rect 22468 12767 22520 12776
rect 22468 12733 22477 12767
rect 22477 12733 22511 12767
rect 22511 12733 22520 12767
rect 22468 12724 22520 12733
rect 8944 12588 8996 12640
rect 14372 12588 14424 12640
rect 14832 12631 14884 12640
rect 14832 12597 14841 12631
rect 14841 12597 14875 12631
rect 14875 12597 14884 12631
rect 14832 12588 14884 12597
rect 17408 12631 17460 12640
rect 17408 12597 17417 12631
rect 17417 12597 17451 12631
rect 17451 12597 17460 12631
rect 17408 12588 17460 12597
rect 19248 12588 19300 12640
rect 19708 12588 19760 12640
rect 22560 12588 22612 12640
rect 22928 12631 22980 12640
rect 22928 12597 22937 12631
rect 22937 12597 22971 12631
rect 22971 12597 22980 12631
rect 22928 12588 22980 12597
rect 3749 12486 3801 12538
rect 3813 12486 3865 12538
rect 3877 12486 3929 12538
rect 3941 12486 3993 12538
rect 4005 12486 4057 12538
rect 9347 12486 9399 12538
rect 9411 12486 9463 12538
rect 9475 12486 9527 12538
rect 9539 12486 9591 12538
rect 9603 12486 9655 12538
rect 14945 12486 14997 12538
rect 15009 12486 15061 12538
rect 15073 12486 15125 12538
rect 15137 12486 15189 12538
rect 15201 12486 15253 12538
rect 20543 12486 20595 12538
rect 20607 12486 20659 12538
rect 20671 12486 20723 12538
rect 20735 12486 20787 12538
rect 20799 12486 20851 12538
rect 3148 12384 3200 12436
rect 9680 12384 9732 12436
rect 2044 12291 2096 12300
rect 2044 12257 2053 12291
rect 2053 12257 2087 12291
rect 2087 12257 2096 12291
rect 2044 12248 2096 12257
rect 9772 12316 9824 12368
rect 2136 12180 2188 12232
rect 4620 12248 4672 12300
rect 3700 12112 3752 12164
rect 4896 12180 4948 12232
rect 5540 12180 5592 12232
rect 4620 12112 4672 12164
rect 5908 12112 5960 12164
rect 4252 12044 4304 12096
rect 4528 12044 4580 12096
rect 5172 12087 5224 12096
rect 5172 12053 5181 12087
rect 5181 12053 5215 12087
rect 5215 12053 5224 12087
rect 5172 12044 5224 12053
rect 6000 12087 6052 12096
rect 6000 12053 6009 12087
rect 6009 12053 6043 12087
rect 6043 12053 6052 12087
rect 6000 12044 6052 12053
rect 8024 12180 8076 12232
rect 8392 12180 8444 12232
rect 8668 12180 8720 12232
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 11980 12384 12032 12436
rect 16856 12384 16908 12436
rect 17868 12384 17920 12436
rect 18144 12384 18196 12436
rect 19616 12427 19668 12436
rect 14096 12248 14148 12300
rect 14372 12291 14424 12300
rect 11520 12223 11572 12232
rect 11520 12189 11529 12223
rect 11529 12189 11563 12223
rect 11563 12189 11572 12223
rect 11520 12180 11572 12189
rect 10600 12112 10652 12164
rect 8484 12044 8536 12096
rect 11428 12112 11480 12164
rect 14372 12257 14381 12291
rect 14381 12257 14415 12291
rect 14415 12257 14424 12291
rect 14372 12248 14424 12257
rect 14740 12248 14792 12300
rect 19616 12393 19625 12427
rect 19625 12393 19659 12427
rect 19659 12393 19668 12427
rect 19616 12384 19668 12393
rect 18604 12316 18656 12368
rect 21456 12384 21508 12436
rect 22100 12384 22152 12436
rect 21640 12316 21692 12368
rect 20260 12248 20312 12300
rect 21548 12248 21600 12300
rect 21732 12291 21784 12300
rect 21732 12257 21741 12291
rect 21741 12257 21775 12291
rect 21775 12257 21784 12291
rect 21732 12248 21784 12257
rect 14832 12180 14884 12232
rect 15752 12180 15804 12232
rect 16212 12180 16264 12232
rect 19064 12223 19116 12232
rect 19064 12189 19073 12223
rect 19073 12189 19107 12223
rect 19107 12189 19116 12223
rect 19064 12180 19116 12189
rect 19800 12180 19852 12232
rect 21824 12180 21876 12232
rect 14740 12112 14792 12164
rect 18144 12112 18196 12164
rect 18512 12112 18564 12164
rect 11336 12044 11388 12096
rect 14464 12044 14516 12096
rect 14832 12087 14884 12096
rect 14832 12053 14841 12087
rect 14841 12053 14875 12087
rect 14875 12053 14884 12087
rect 14832 12044 14884 12053
rect 16948 12044 17000 12096
rect 17132 12087 17184 12096
rect 17132 12053 17141 12087
rect 17141 12053 17175 12087
rect 17175 12053 17184 12087
rect 17132 12044 17184 12053
rect 17224 12044 17276 12096
rect 19432 12087 19484 12096
rect 19432 12053 19441 12087
rect 19441 12053 19475 12087
rect 19475 12053 19484 12087
rect 19432 12044 19484 12053
rect 21732 12112 21784 12164
rect 22284 12180 22336 12232
rect 22468 12112 22520 12164
rect 19984 12044 20036 12096
rect 20076 12044 20128 12096
rect 20812 12044 20864 12096
rect 23020 12044 23072 12096
rect 6548 11942 6600 11994
rect 6612 11942 6664 11994
rect 6676 11942 6728 11994
rect 6740 11942 6792 11994
rect 6804 11942 6856 11994
rect 12146 11942 12198 11994
rect 12210 11942 12262 11994
rect 12274 11942 12326 11994
rect 12338 11942 12390 11994
rect 12402 11942 12454 11994
rect 17744 11942 17796 11994
rect 17808 11942 17860 11994
rect 17872 11942 17924 11994
rect 17936 11942 17988 11994
rect 18000 11942 18052 11994
rect 1400 11840 1452 11892
rect 3700 11883 3752 11892
rect 3700 11849 3709 11883
rect 3709 11849 3743 11883
rect 3743 11849 3752 11883
rect 3700 11840 3752 11849
rect 4988 11840 5040 11892
rect 5356 11883 5408 11892
rect 5356 11849 5365 11883
rect 5365 11849 5399 11883
rect 5399 11849 5408 11883
rect 5356 11840 5408 11849
rect 8484 11883 8536 11892
rect 5172 11772 5224 11824
rect 6000 11772 6052 11824
rect 8484 11849 8493 11883
rect 8493 11849 8527 11883
rect 8527 11849 8536 11883
rect 8484 11840 8536 11849
rect 8852 11840 8904 11892
rect 12072 11840 12124 11892
rect 17132 11840 17184 11892
rect 17500 11840 17552 11892
rect 17592 11840 17644 11892
rect 18604 11840 18656 11892
rect 4252 11704 4304 11756
rect 4620 11704 4672 11756
rect 4988 11747 5040 11756
rect 4988 11713 4997 11747
rect 4997 11713 5031 11747
rect 5031 11713 5040 11747
rect 4988 11704 5040 11713
rect 5448 11704 5500 11756
rect 6460 11704 6512 11756
rect 11520 11772 11572 11824
rect 14004 11815 14056 11824
rect 10048 11704 10100 11756
rect 11980 11704 12032 11756
rect 4344 11636 4396 11688
rect 4712 11679 4764 11688
rect 4712 11645 4721 11679
rect 4721 11645 4755 11679
rect 4755 11645 4764 11679
rect 4712 11636 4764 11645
rect 4804 11636 4856 11688
rect 6184 11636 6236 11688
rect 8576 11636 8628 11688
rect 10968 11636 11020 11688
rect 14004 11781 14013 11815
rect 14013 11781 14047 11815
rect 14047 11781 14056 11815
rect 14004 11772 14056 11781
rect 13820 11704 13872 11756
rect 13544 11636 13596 11688
rect 15568 11772 15620 11824
rect 18328 11772 18380 11824
rect 18420 11772 18472 11824
rect 19432 11840 19484 11892
rect 20812 11883 20864 11892
rect 20812 11849 20821 11883
rect 20821 11849 20855 11883
rect 20855 11849 20864 11883
rect 20812 11840 20864 11849
rect 22100 11840 22152 11892
rect 21180 11772 21232 11824
rect 14832 11704 14884 11756
rect 15476 11704 15528 11756
rect 16120 11747 16172 11756
rect 16120 11713 16129 11747
rect 16129 11713 16163 11747
rect 16163 11713 16172 11747
rect 16120 11704 16172 11713
rect 16672 11704 16724 11756
rect 17040 11704 17092 11756
rect 6276 11568 6328 11620
rect 11612 11611 11664 11620
rect 11612 11577 11621 11611
rect 11621 11577 11655 11611
rect 11655 11577 11664 11611
rect 11612 11568 11664 11577
rect 16028 11679 16080 11688
rect 16028 11645 16037 11679
rect 16037 11645 16071 11679
rect 16071 11645 16080 11679
rect 16028 11636 16080 11645
rect 16396 11636 16448 11688
rect 18604 11679 18656 11688
rect 18604 11645 18613 11679
rect 18613 11645 18647 11679
rect 18647 11645 18656 11679
rect 18604 11636 18656 11645
rect 19984 11636 20036 11688
rect 20352 11679 20404 11688
rect 20352 11645 20361 11679
rect 20361 11645 20395 11679
rect 20395 11645 20404 11679
rect 20352 11636 20404 11645
rect 21548 11704 21600 11756
rect 23112 11747 23164 11756
rect 23112 11713 23121 11747
rect 23121 11713 23155 11747
rect 23155 11713 23164 11747
rect 23112 11704 23164 11713
rect 22100 11636 22152 11688
rect 3240 11543 3292 11552
rect 3240 11509 3249 11543
rect 3249 11509 3283 11543
rect 3283 11509 3292 11543
rect 3240 11500 3292 11509
rect 4344 11543 4396 11552
rect 4344 11509 4353 11543
rect 4353 11509 4387 11543
rect 4387 11509 4396 11543
rect 4344 11500 4396 11509
rect 4528 11500 4580 11552
rect 9680 11543 9732 11552
rect 9680 11509 9689 11543
rect 9689 11509 9723 11543
rect 9723 11509 9732 11543
rect 9680 11500 9732 11509
rect 13728 11543 13780 11552
rect 13728 11509 13737 11543
rect 13737 11509 13771 11543
rect 13771 11509 13780 11543
rect 13728 11500 13780 11509
rect 14556 11500 14608 11552
rect 16120 11500 16172 11552
rect 17776 11500 17828 11552
rect 18972 11500 19024 11552
rect 21272 11568 21324 11620
rect 21640 11568 21692 11620
rect 23020 11636 23072 11688
rect 19984 11543 20036 11552
rect 19984 11509 19993 11543
rect 19993 11509 20027 11543
rect 20027 11509 20036 11543
rect 19984 11500 20036 11509
rect 20904 11543 20956 11552
rect 20904 11509 20913 11543
rect 20913 11509 20947 11543
rect 20947 11509 20956 11543
rect 20904 11500 20956 11509
rect 22652 11500 22704 11552
rect 3749 11398 3801 11450
rect 3813 11398 3865 11450
rect 3877 11398 3929 11450
rect 3941 11398 3993 11450
rect 4005 11398 4057 11450
rect 9347 11398 9399 11450
rect 9411 11398 9463 11450
rect 9475 11398 9527 11450
rect 9539 11398 9591 11450
rect 9603 11398 9655 11450
rect 14945 11398 14997 11450
rect 15009 11398 15061 11450
rect 15073 11398 15125 11450
rect 15137 11398 15189 11450
rect 15201 11398 15253 11450
rect 20543 11398 20595 11450
rect 20607 11398 20659 11450
rect 20671 11398 20723 11450
rect 20735 11398 20787 11450
rect 20799 11398 20851 11450
rect 3516 11296 3568 11348
rect 4160 11296 4212 11348
rect 4988 11296 5040 11348
rect 9128 11339 9180 11348
rect 9128 11305 9137 11339
rect 9137 11305 9171 11339
rect 9171 11305 9180 11339
rect 9128 11296 9180 11305
rect 10048 11296 10100 11348
rect 4804 11228 4856 11280
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 3424 11135 3476 11144
rect 3424 11101 3433 11135
rect 3433 11101 3467 11135
rect 3467 11101 3476 11135
rect 3424 11092 3476 11101
rect 4436 11160 4488 11212
rect 4712 11160 4764 11212
rect 6368 11228 6420 11280
rect 10968 11296 11020 11348
rect 11336 11296 11388 11348
rect 13820 11296 13872 11348
rect 13912 11296 13964 11348
rect 14188 11296 14240 11348
rect 15476 11296 15528 11348
rect 3148 11024 3200 11076
rect 3516 11024 3568 11076
rect 4620 11092 4672 11144
rect 5448 11092 5500 11144
rect 6460 11092 6512 11144
rect 8392 11135 8444 11144
rect 4712 11067 4764 11076
rect 4712 11033 4721 11067
rect 4721 11033 4755 11067
rect 4755 11033 4764 11067
rect 4712 11024 4764 11033
rect 4528 10956 4580 11008
rect 5172 10999 5224 11008
rect 5172 10965 5181 10999
rect 5181 10965 5215 10999
rect 5215 10965 5224 10999
rect 5172 10956 5224 10965
rect 6092 10956 6144 11008
rect 7012 10999 7064 11008
rect 7012 10965 7021 10999
rect 7021 10965 7055 10999
rect 7055 10965 7064 10999
rect 7012 10956 7064 10965
rect 8392 11101 8401 11135
rect 8401 11101 8435 11135
rect 8435 11101 8444 11135
rect 8392 11092 8444 11101
rect 8576 11092 8628 11144
rect 8944 11135 8996 11144
rect 8944 11101 8953 11135
rect 8953 11101 8987 11135
rect 8987 11101 8996 11135
rect 8944 11092 8996 11101
rect 10508 11092 10560 11144
rect 11520 11160 11572 11212
rect 12072 11135 12124 11144
rect 12072 11101 12081 11135
rect 12081 11101 12115 11135
rect 12115 11101 12124 11135
rect 12072 11092 12124 11101
rect 13912 11160 13964 11212
rect 14280 11203 14332 11212
rect 14280 11169 14289 11203
rect 14289 11169 14323 11203
rect 14323 11169 14332 11203
rect 14280 11160 14332 11169
rect 14740 11160 14792 11212
rect 15568 11160 15620 11212
rect 9680 11024 9732 11076
rect 10692 11024 10744 11076
rect 8300 10956 8352 11008
rect 12072 10956 12124 11008
rect 13728 11092 13780 11144
rect 16028 11296 16080 11348
rect 16580 11228 16632 11280
rect 17040 11296 17092 11348
rect 17316 11296 17368 11348
rect 20352 11296 20404 11348
rect 20996 11339 21048 11348
rect 20996 11305 21005 11339
rect 21005 11305 21039 11339
rect 21039 11305 21048 11339
rect 20996 11296 21048 11305
rect 17500 11271 17552 11280
rect 17500 11237 17509 11271
rect 17509 11237 17543 11271
rect 17543 11237 17552 11271
rect 18972 11271 19024 11280
rect 17500 11228 17552 11237
rect 16948 11203 17000 11212
rect 16948 11169 16957 11203
rect 16957 11169 16991 11203
rect 16991 11169 17000 11203
rect 16948 11160 17000 11169
rect 17408 11160 17460 11212
rect 17592 11160 17644 11212
rect 17224 11092 17276 11144
rect 17776 11135 17828 11144
rect 17776 11101 17785 11135
rect 17785 11101 17819 11135
rect 17819 11101 17828 11135
rect 17776 11092 17828 11101
rect 18972 11237 18981 11271
rect 18981 11237 19015 11271
rect 19015 11237 19024 11271
rect 18972 11228 19024 11237
rect 20444 11228 20496 11280
rect 23112 11296 23164 11348
rect 22100 11228 22152 11280
rect 18604 11160 18656 11212
rect 23204 11228 23256 11280
rect 18972 11092 19024 11144
rect 23572 11160 23624 11212
rect 21180 11092 21232 11144
rect 22192 11092 22244 11144
rect 23112 11135 23164 11144
rect 23112 11101 23121 11135
rect 23121 11101 23155 11135
rect 23155 11101 23164 11135
rect 23112 11092 23164 11101
rect 13636 11024 13688 11076
rect 13360 10956 13412 11008
rect 14372 10999 14424 11008
rect 14372 10965 14381 10999
rect 14381 10965 14415 10999
rect 14415 10965 14424 10999
rect 14372 10956 14424 10965
rect 15384 10956 15436 11008
rect 18696 11024 18748 11076
rect 19064 10956 19116 11008
rect 19248 11024 19300 11076
rect 23020 10956 23072 11008
rect 6548 10854 6600 10906
rect 6612 10854 6664 10906
rect 6676 10854 6728 10906
rect 6740 10854 6792 10906
rect 6804 10854 6856 10906
rect 12146 10854 12198 10906
rect 12210 10854 12262 10906
rect 12274 10854 12326 10906
rect 12338 10854 12390 10906
rect 12402 10854 12454 10906
rect 17744 10854 17796 10906
rect 17808 10854 17860 10906
rect 17872 10854 17924 10906
rect 17936 10854 17988 10906
rect 18000 10854 18052 10906
rect 3424 10752 3476 10804
rect 5172 10752 5224 10804
rect 7012 10752 7064 10804
rect 8668 10795 8720 10804
rect 8668 10761 8677 10795
rect 8677 10761 8711 10795
rect 8711 10761 8720 10795
rect 8668 10752 8720 10761
rect 8944 10752 8996 10804
rect 10968 10752 11020 10804
rect 11980 10752 12032 10804
rect 14372 10795 14424 10804
rect 14372 10761 14381 10795
rect 14381 10761 14415 10795
rect 14415 10761 14424 10795
rect 14372 10752 14424 10761
rect 14648 10752 14700 10804
rect 17500 10752 17552 10804
rect 6920 10684 6972 10736
rect 9772 10684 9824 10736
rect 10508 10684 10560 10736
rect 13912 10684 13964 10736
rect 16120 10684 16172 10736
rect 1860 10616 1912 10668
rect 4804 10616 4856 10668
rect 5356 10616 5408 10668
rect 6184 10659 6236 10668
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 7288 10616 7340 10668
rect 8944 10616 8996 10668
rect 1768 10591 1820 10600
rect 1768 10557 1777 10591
rect 1777 10557 1811 10591
rect 1811 10557 1820 10591
rect 1768 10548 1820 10557
rect 4436 10591 4488 10600
rect 4436 10557 4445 10591
rect 4445 10557 4479 10591
rect 4479 10557 4488 10591
rect 4436 10548 4488 10557
rect 4896 10548 4948 10600
rect 4160 10480 4212 10532
rect 8760 10548 8812 10600
rect 9680 10480 9732 10532
rect 4620 10412 4672 10464
rect 5448 10412 5500 10464
rect 7472 10412 7524 10464
rect 11336 10616 11388 10668
rect 12072 10616 12124 10668
rect 12716 10616 12768 10668
rect 13820 10616 13872 10668
rect 10876 10548 10928 10600
rect 13912 10591 13964 10600
rect 13544 10523 13596 10532
rect 13544 10489 13553 10523
rect 13553 10489 13587 10523
rect 13587 10489 13596 10523
rect 13544 10480 13596 10489
rect 13912 10557 13921 10591
rect 13921 10557 13955 10591
rect 13955 10557 13964 10591
rect 13912 10548 13964 10557
rect 14004 10480 14056 10532
rect 11520 10455 11572 10464
rect 11520 10421 11529 10455
rect 11529 10421 11563 10455
rect 11563 10421 11572 10455
rect 11520 10412 11572 10421
rect 17408 10616 17460 10668
rect 19708 10752 19760 10804
rect 22468 10795 22520 10804
rect 22468 10761 22477 10795
rect 22477 10761 22511 10795
rect 22511 10761 22520 10795
rect 22468 10752 22520 10761
rect 23296 10752 23348 10804
rect 21180 10684 21232 10736
rect 16672 10548 16724 10600
rect 17224 10548 17276 10600
rect 18328 10548 18380 10600
rect 18972 10616 19024 10668
rect 18512 10548 18564 10600
rect 18696 10591 18748 10600
rect 18696 10557 18705 10591
rect 18705 10557 18739 10591
rect 18739 10557 18748 10591
rect 18696 10548 18748 10557
rect 19064 10548 19116 10600
rect 21088 10616 21140 10668
rect 22560 10591 22612 10600
rect 22560 10557 22569 10591
rect 22569 10557 22603 10591
rect 22603 10557 22612 10591
rect 22560 10548 22612 10557
rect 21272 10480 21324 10532
rect 23940 10616 23992 10668
rect 16948 10412 17000 10464
rect 18512 10412 18564 10464
rect 19064 10412 19116 10464
rect 20260 10412 20312 10464
rect 21640 10455 21692 10464
rect 21640 10421 21649 10455
rect 21649 10421 21683 10455
rect 21683 10421 21692 10455
rect 21640 10412 21692 10421
rect 3749 10310 3801 10362
rect 3813 10310 3865 10362
rect 3877 10310 3929 10362
rect 3941 10310 3993 10362
rect 4005 10310 4057 10362
rect 9347 10310 9399 10362
rect 9411 10310 9463 10362
rect 9475 10310 9527 10362
rect 9539 10310 9591 10362
rect 9603 10310 9655 10362
rect 14945 10310 14997 10362
rect 15009 10310 15061 10362
rect 15073 10310 15125 10362
rect 15137 10310 15189 10362
rect 15201 10310 15253 10362
rect 20543 10310 20595 10362
rect 20607 10310 20659 10362
rect 20671 10310 20723 10362
rect 20735 10310 20787 10362
rect 20799 10310 20851 10362
rect 1768 10208 1820 10260
rect 4436 10208 4488 10260
rect 7288 10208 7340 10260
rect 8944 10251 8996 10260
rect 8944 10217 8953 10251
rect 8953 10217 8987 10251
rect 8987 10217 8996 10251
rect 8944 10208 8996 10217
rect 4528 10140 4580 10192
rect 6092 10183 6144 10192
rect 6092 10149 6101 10183
rect 6101 10149 6135 10183
rect 6135 10149 6144 10183
rect 6092 10140 6144 10149
rect 3424 10047 3476 10056
rect 3424 10013 3433 10047
rect 3433 10013 3467 10047
rect 3467 10013 3476 10047
rect 3424 10004 3476 10013
rect 3884 10072 3936 10124
rect 4436 10115 4488 10124
rect 4436 10081 4445 10115
rect 4445 10081 4479 10115
rect 4479 10081 4488 10115
rect 4436 10072 4488 10081
rect 6460 10072 6512 10124
rect 9680 10072 9732 10124
rect 10876 10208 10928 10260
rect 11980 10251 12032 10260
rect 11980 10217 11989 10251
rect 11989 10217 12023 10251
rect 12023 10217 12032 10251
rect 11980 10208 12032 10217
rect 13636 10251 13688 10260
rect 13636 10217 13645 10251
rect 13645 10217 13679 10251
rect 13679 10217 13688 10251
rect 13636 10208 13688 10217
rect 15384 10208 15436 10260
rect 16764 10208 16816 10260
rect 19892 10251 19944 10260
rect 5356 10004 5408 10056
rect 8300 10047 8352 10056
rect 8300 10013 8318 10047
rect 8318 10013 8352 10047
rect 8300 10004 8352 10013
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 9588 10004 9640 10056
rect 10508 10004 10560 10056
rect 13360 10047 13412 10056
rect 13360 10013 13369 10047
rect 13369 10013 13403 10047
rect 13403 10013 13412 10047
rect 13360 10004 13412 10013
rect 13452 10047 13504 10056
rect 13452 10013 13461 10047
rect 13461 10013 13495 10047
rect 13495 10013 13504 10047
rect 13452 10004 13504 10013
rect 14004 10004 14056 10056
rect 15660 10004 15712 10056
rect 16396 10004 16448 10056
rect 16488 10004 16540 10056
rect 18144 10004 18196 10056
rect 4160 9979 4212 9988
rect 2596 9868 2648 9920
rect 3608 9868 3660 9920
rect 3792 9911 3844 9920
rect 3792 9877 3801 9911
rect 3801 9877 3835 9911
rect 3835 9877 3844 9911
rect 3792 9868 3844 9877
rect 4160 9945 4169 9979
rect 4169 9945 4203 9979
rect 4203 9945 4212 9979
rect 4160 9936 4212 9945
rect 4344 9936 4396 9988
rect 4620 9936 4672 9988
rect 9680 9936 9732 9988
rect 15384 9936 15436 9988
rect 4804 9868 4856 9920
rect 6920 9868 6972 9920
rect 8760 9868 8812 9920
rect 9404 9911 9456 9920
rect 9404 9877 9413 9911
rect 9413 9877 9447 9911
rect 9447 9877 9456 9911
rect 9404 9868 9456 9877
rect 11336 9868 11388 9920
rect 13912 9868 13964 9920
rect 15936 9868 15988 9920
rect 18972 10004 19024 10056
rect 18420 9979 18472 9988
rect 18420 9945 18460 9979
rect 18460 9945 18472 9979
rect 18880 9979 18932 9988
rect 18420 9936 18472 9945
rect 18880 9945 18889 9979
rect 18889 9945 18923 9979
rect 18923 9945 18932 9979
rect 18880 9936 18932 9945
rect 17132 9868 17184 9920
rect 17224 9911 17276 9920
rect 17224 9877 17233 9911
rect 17233 9877 17267 9911
rect 17267 9877 17276 9911
rect 17224 9868 17276 9877
rect 18604 9868 18656 9920
rect 19892 10217 19901 10251
rect 19901 10217 19935 10251
rect 19935 10217 19944 10251
rect 19892 10208 19944 10217
rect 20904 10208 20956 10260
rect 21824 10251 21876 10260
rect 21824 10217 21833 10251
rect 21833 10217 21867 10251
rect 21867 10217 21876 10251
rect 21824 10208 21876 10217
rect 21916 10208 21968 10260
rect 21640 10140 21692 10192
rect 22836 10183 22888 10192
rect 21824 10072 21876 10124
rect 22376 10115 22428 10124
rect 22376 10081 22385 10115
rect 22385 10081 22419 10115
rect 22419 10081 22428 10115
rect 22376 10072 22428 10081
rect 22836 10149 22845 10183
rect 22845 10149 22879 10183
rect 22879 10149 22888 10183
rect 22836 10140 22888 10149
rect 19708 10004 19760 10056
rect 20260 10004 20312 10056
rect 23020 10004 23072 10056
rect 19984 9868 20036 9920
rect 22100 9868 22152 9920
rect 6548 9766 6600 9818
rect 6612 9766 6664 9818
rect 6676 9766 6728 9818
rect 6740 9766 6792 9818
rect 6804 9766 6856 9818
rect 12146 9766 12198 9818
rect 12210 9766 12262 9818
rect 12274 9766 12326 9818
rect 12338 9766 12390 9818
rect 12402 9766 12454 9818
rect 17744 9766 17796 9818
rect 17808 9766 17860 9818
rect 17872 9766 17924 9818
rect 17936 9766 17988 9818
rect 18000 9766 18052 9818
rect 3792 9664 3844 9716
rect 4804 9707 4856 9716
rect 4804 9673 4813 9707
rect 4813 9673 4847 9707
rect 4847 9673 4856 9707
rect 4804 9664 4856 9673
rect 3240 9596 3292 9648
rect 5356 9596 5408 9648
rect 1400 9571 1452 9580
rect 1400 9537 1409 9571
rect 1409 9537 1443 9571
rect 1443 9537 1452 9571
rect 1400 9528 1452 9537
rect 3332 9528 3384 9580
rect 4528 9528 4580 9580
rect 5540 9528 5592 9580
rect 9404 9664 9456 9716
rect 10968 9707 11020 9716
rect 10968 9673 10977 9707
rect 10977 9673 11011 9707
rect 11011 9673 11020 9707
rect 10968 9664 11020 9673
rect 11520 9664 11572 9716
rect 8576 9596 8628 9648
rect 9680 9596 9732 9648
rect 12716 9639 12768 9648
rect 12716 9605 12725 9639
rect 12725 9605 12759 9639
rect 12759 9605 12768 9639
rect 12716 9596 12768 9605
rect 14096 9596 14148 9648
rect 15660 9639 15712 9648
rect 15660 9605 15669 9639
rect 15669 9605 15703 9639
rect 15703 9605 15712 9639
rect 15660 9596 15712 9605
rect 18328 9664 18380 9716
rect 18696 9664 18748 9716
rect 21824 9707 21876 9716
rect 21824 9673 21833 9707
rect 21833 9673 21867 9707
rect 21867 9673 21876 9707
rect 21824 9664 21876 9673
rect 22560 9664 22612 9716
rect 2872 9503 2924 9512
rect 2872 9469 2881 9503
rect 2881 9469 2915 9503
rect 2915 9469 2924 9503
rect 2872 9460 2924 9469
rect 7472 9528 7524 9580
rect 7196 9460 7248 9512
rect 3516 9392 3568 9444
rect 4712 9392 4764 9444
rect 1492 9324 1544 9376
rect 2504 9324 2556 9376
rect 6644 9367 6696 9376
rect 6644 9333 6653 9367
rect 6653 9333 6687 9367
rect 6687 9333 6696 9367
rect 6644 9324 6696 9333
rect 9588 9571 9640 9580
rect 9588 9537 9597 9571
rect 9597 9537 9631 9571
rect 9631 9537 9640 9571
rect 9588 9528 9640 9537
rect 9864 9571 9916 9580
rect 9864 9537 9898 9571
rect 9898 9537 9916 9571
rect 9864 9528 9916 9537
rect 11980 9528 12032 9580
rect 13268 9571 13320 9580
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 14372 9571 14424 9580
rect 14372 9537 14381 9571
rect 14381 9537 14415 9571
rect 14415 9537 14424 9571
rect 14372 9528 14424 9537
rect 18880 9596 18932 9648
rect 21180 9639 21232 9648
rect 21180 9605 21189 9639
rect 21189 9605 21223 9639
rect 21223 9605 21232 9639
rect 21180 9596 21232 9605
rect 22100 9596 22152 9648
rect 23112 9639 23164 9648
rect 23112 9605 23121 9639
rect 23121 9605 23155 9639
rect 23155 9605 23164 9639
rect 23112 9596 23164 9605
rect 15936 9528 15988 9580
rect 17408 9571 17460 9580
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 14004 9435 14056 9444
rect 14004 9401 14013 9435
rect 14013 9401 14047 9435
rect 14047 9401 14056 9435
rect 14004 9392 14056 9401
rect 14280 9392 14332 9444
rect 14832 9460 14884 9512
rect 15384 9460 15436 9512
rect 14740 9392 14792 9444
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 18604 9571 18656 9580
rect 18604 9537 18613 9571
rect 18613 9537 18647 9571
rect 18647 9537 18656 9571
rect 18604 9528 18656 9537
rect 18972 9528 19024 9580
rect 21548 9528 21600 9580
rect 22836 9571 22888 9580
rect 22836 9537 22845 9571
rect 22845 9537 22879 9571
rect 22879 9537 22888 9571
rect 22836 9528 22888 9537
rect 16856 9460 16908 9512
rect 17316 9460 17368 9512
rect 18420 9460 18472 9512
rect 21180 9460 21232 9512
rect 21364 9392 21416 9444
rect 23112 9460 23164 9512
rect 21732 9392 21784 9444
rect 10968 9324 11020 9376
rect 13912 9367 13964 9376
rect 13912 9333 13921 9367
rect 13921 9333 13955 9367
rect 13955 9333 13964 9367
rect 13912 9324 13964 9333
rect 16304 9324 16356 9376
rect 17040 9324 17092 9376
rect 20996 9324 21048 9376
rect 21456 9324 21508 9376
rect 3749 9222 3801 9274
rect 3813 9222 3865 9274
rect 3877 9222 3929 9274
rect 3941 9222 3993 9274
rect 4005 9222 4057 9274
rect 9347 9222 9399 9274
rect 9411 9222 9463 9274
rect 9475 9222 9527 9274
rect 9539 9222 9591 9274
rect 9603 9222 9655 9274
rect 14945 9222 14997 9274
rect 15009 9222 15061 9274
rect 15073 9222 15125 9274
rect 15137 9222 15189 9274
rect 15201 9222 15253 9274
rect 20543 9222 20595 9274
rect 20607 9222 20659 9274
rect 20671 9222 20723 9274
rect 20735 9222 20787 9274
rect 20799 9222 20851 9274
rect 1768 9120 1820 9172
rect 3424 9120 3476 9172
rect 4528 9163 4580 9172
rect 4528 9129 4537 9163
rect 4537 9129 4571 9163
rect 4571 9129 4580 9163
rect 4528 9120 4580 9129
rect 5540 9120 5592 9172
rect 3148 9052 3200 9104
rect 2872 8984 2924 9036
rect 4896 8984 4948 9036
rect 5356 8984 5408 9036
rect 1492 8916 1544 8968
rect 4160 8916 4212 8968
rect 11428 9120 11480 9172
rect 13452 9163 13504 9172
rect 13452 9129 13461 9163
rect 13461 9129 13495 9163
rect 13495 9129 13504 9163
rect 13452 9120 13504 9129
rect 14096 9120 14148 9172
rect 19432 9120 19484 9172
rect 21548 9163 21600 9172
rect 8392 9052 8444 9104
rect 8760 9095 8812 9104
rect 8760 9061 8769 9095
rect 8769 9061 8803 9095
rect 8803 9061 8812 9095
rect 8760 9052 8812 9061
rect 16856 9052 16908 9104
rect 10508 8984 10560 9036
rect 4344 8848 4396 8900
rect 4712 8848 4764 8900
rect 8392 8916 8444 8968
rect 14280 8984 14332 9036
rect 15384 8984 15436 9036
rect 16764 9027 16816 9036
rect 11980 8916 12032 8968
rect 13452 8916 13504 8968
rect 15660 8916 15712 8968
rect 16764 8993 16773 9027
rect 16773 8993 16807 9027
rect 16807 8993 16816 9027
rect 16764 8984 16816 8993
rect 16948 9027 17000 9036
rect 16948 8993 16957 9027
rect 16957 8993 16991 9027
rect 16991 8993 17000 9027
rect 16948 8984 17000 8993
rect 17316 9052 17368 9104
rect 19708 9052 19760 9104
rect 16672 8916 16724 8968
rect 18972 8984 19024 9036
rect 19616 8984 19668 9036
rect 20444 9052 20496 9104
rect 19248 8916 19300 8968
rect 21548 9129 21557 9163
rect 21557 9129 21591 9163
rect 21591 9129 21600 9163
rect 21548 9120 21600 9129
rect 21732 9120 21784 9172
rect 21088 9052 21140 9104
rect 2780 8823 2832 8832
rect 2780 8789 2789 8823
rect 2789 8789 2823 8823
rect 2823 8789 2832 8823
rect 2780 8780 2832 8789
rect 3516 8780 3568 8832
rect 4896 8823 4948 8832
rect 4896 8789 4905 8823
rect 4905 8789 4939 8823
rect 4939 8789 4948 8823
rect 4896 8780 4948 8789
rect 4988 8823 5040 8832
rect 4988 8789 4997 8823
rect 4997 8789 5031 8823
rect 5031 8789 5040 8823
rect 4988 8780 5040 8789
rect 5264 8780 5316 8832
rect 6644 8848 6696 8900
rect 8576 8848 8628 8900
rect 11060 8848 11112 8900
rect 6920 8823 6972 8832
rect 6920 8789 6929 8823
rect 6929 8789 6963 8823
rect 6963 8789 6972 8823
rect 10508 8823 10560 8832
rect 6920 8780 6972 8789
rect 10508 8789 10517 8823
rect 10517 8789 10551 8823
rect 10551 8789 10560 8823
rect 10508 8780 10560 8789
rect 14648 8891 14700 8900
rect 14648 8857 14682 8891
rect 14682 8857 14700 8891
rect 14648 8848 14700 8857
rect 15292 8848 15344 8900
rect 19524 8848 19576 8900
rect 12992 8823 13044 8832
rect 12992 8789 13001 8823
rect 13001 8789 13035 8823
rect 13035 8789 13044 8823
rect 12992 8780 13044 8789
rect 13084 8823 13136 8832
rect 13084 8789 13093 8823
rect 13093 8789 13127 8823
rect 13127 8789 13136 8823
rect 13084 8780 13136 8789
rect 13636 8780 13688 8832
rect 15384 8780 15436 8832
rect 15752 8823 15804 8832
rect 15752 8789 15761 8823
rect 15761 8789 15795 8823
rect 15795 8789 15804 8823
rect 15752 8780 15804 8789
rect 15844 8780 15896 8832
rect 21824 8848 21876 8900
rect 22560 8780 22612 8832
rect 23112 8823 23164 8832
rect 23112 8789 23121 8823
rect 23121 8789 23155 8823
rect 23155 8789 23164 8823
rect 23112 8780 23164 8789
rect 6548 8678 6600 8730
rect 6612 8678 6664 8730
rect 6676 8678 6728 8730
rect 6740 8678 6792 8730
rect 6804 8678 6856 8730
rect 12146 8678 12198 8730
rect 12210 8678 12262 8730
rect 12274 8678 12326 8730
rect 12338 8678 12390 8730
rect 12402 8678 12454 8730
rect 17744 8678 17796 8730
rect 17808 8678 17860 8730
rect 17872 8678 17924 8730
rect 17936 8678 17988 8730
rect 18000 8678 18052 8730
rect 3516 8619 3568 8628
rect 3516 8585 3525 8619
rect 3525 8585 3559 8619
rect 3559 8585 3568 8619
rect 3516 8576 3568 8585
rect 3608 8576 3660 8628
rect 4344 8619 4396 8628
rect 4344 8585 4353 8619
rect 4353 8585 4387 8619
rect 4387 8585 4396 8619
rect 4344 8576 4396 8585
rect 4896 8576 4948 8628
rect 7012 8619 7064 8628
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 9772 8619 9824 8628
rect 9772 8585 9781 8619
rect 9781 8585 9815 8619
rect 9815 8585 9824 8619
rect 9772 8576 9824 8585
rect 10140 8619 10192 8628
rect 10140 8585 10149 8619
rect 10149 8585 10183 8619
rect 10183 8585 10192 8619
rect 10140 8576 10192 8585
rect 10508 8576 10560 8628
rect 10692 8619 10744 8628
rect 10692 8585 10701 8619
rect 10701 8585 10735 8619
rect 10735 8585 10744 8619
rect 10692 8576 10744 8585
rect 13268 8576 13320 8628
rect 2780 8508 2832 8560
rect 3240 8508 3292 8560
rect 13912 8508 13964 8560
rect 14372 8576 14424 8628
rect 17132 8576 17184 8628
rect 19340 8576 19392 8628
rect 20260 8576 20312 8628
rect 21180 8576 21232 8628
rect 15752 8508 15804 8560
rect 1768 8440 1820 8492
rect 2320 8483 2372 8492
rect 2320 8449 2354 8483
rect 2354 8449 2372 8483
rect 2320 8440 2372 8449
rect 2688 8440 2740 8492
rect 5724 8483 5776 8492
rect 5724 8449 5733 8483
rect 5733 8449 5767 8483
rect 5767 8449 5776 8483
rect 5724 8440 5776 8449
rect 6092 8440 6144 8492
rect 8208 8483 8260 8492
rect 8208 8449 8217 8483
rect 8217 8449 8251 8483
rect 8251 8449 8260 8483
rect 8208 8440 8260 8449
rect 8392 8440 8444 8492
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 11980 8483 12032 8492
rect 11980 8449 11989 8483
rect 11989 8449 12023 8483
rect 12023 8449 12032 8483
rect 11980 8440 12032 8449
rect 12072 8440 12124 8492
rect 13452 8483 13504 8492
rect 13452 8449 13461 8483
rect 13461 8449 13495 8483
rect 13495 8449 13504 8483
rect 13452 8440 13504 8449
rect 14556 8440 14608 8492
rect 16120 8483 16172 8492
rect 5816 8415 5868 8424
rect 3332 8304 3384 8356
rect 5816 8381 5825 8415
rect 5825 8381 5859 8415
rect 5859 8381 5868 8415
rect 5816 8372 5868 8381
rect 5172 8304 5224 8356
rect 6276 8372 6328 8424
rect 9680 8347 9732 8356
rect 9680 8313 9689 8347
rect 9689 8313 9723 8347
rect 9723 8313 9732 8347
rect 10876 8372 10928 8424
rect 15384 8415 15436 8424
rect 15384 8381 15393 8415
rect 15393 8381 15427 8415
rect 15427 8381 15436 8415
rect 15384 8372 15436 8381
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 22744 8508 22796 8560
rect 17500 8440 17552 8492
rect 18972 8440 19024 8492
rect 19064 8440 19116 8492
rect 21364 8483 21416 8492
rect 21364 8449 21373 8483
rect 21373 8449 21407 8483
rect 21407 8449 21416 8483
rect 21364 8440 21416 8449
rect 21732 8440 21784 8492
rect 22560 8483 22612 8492
rect 22560 8449 22569 8483
rect 22569 8449 22603 8483
rect 22603 8449 22612 8483
rect 22560 8440 22612 8449
rect 20444 8372 20496 8424
rect 20812 8372 20864 8424
rect 20904 8372 20956 8424
rect 21548 8372 21600 8424
rect 9680 8304 9732 8313
rect 10692 8304 10744 8356
rect 11704 8304 11756 8356
rect 14464 8304 14516 8356
rect 17592 8304 17644 8356
rect 21180 8304 21232 8356
rect 16120 8236 16172 8288
rect 20260 8236 20312 8288
rect 21732 8236 21784 8288
rect 3749 8134 3801 8186
rect 3813 8134 3865 8186
rect 3877 8134 3929 8186
rect 3941 8134 3993 8186
rect 4005 8134 4057 8186
rect 9347 8134 9399 8186
rect 9411 8134 9463 8186
rect 9475 8134 9527 8186
rect 9539 8134 9591 8186
rect 9603 8134 9655 8186
rect 14945 8134 14997 8186
rect 15009 8134 15061 8186
rect 15073 8134 15125 8186
rect 15137 8134 15189 8186
rect 15201 8134 15253 8186
rect 20543 8134 20595 8186
rect 20607 8134 20659 8186
rect 20671 8134 20723 8186
rect 20735 8134 20787 8186
rect 20799 8134 20851 8186
rect 4988 8032 5040 8084
rect 5264 7964 5316 8016
rect 1768 7896 1820 7948
rect 5172 7939 5224 7948
rect 5172 7905 5181 7939
rect 5181 7905 5215 7939
rect 5215 7905 5224 7939
rect 5172 7896 5224 7905
rect 2136 7871 2188 7880
rect 2136 7837 2145 7871
rect 2145 7837 2179 7871
rect 2179 7837 2188 7871
rect 2136 7828 2188 7837
rect 2504 7871 2556 7880
rect 2504 7837 2538 7871
rect 2538 7837 2556 7871
rect 2504 7828 2556 7837
rect 5724 8032 5776 8084
rect 7196 8032 7248 8084
rect 8576 8032 8628 8084
rect 9864 8032 9916 8084
rect 13084 8032 13136 8084
rect 19156 8032 19208 8084
rect 20904 8032 20956 8084
rect 21364 8075 21416 8084
rect 21364 8041 21373 8075
rect 21373 8041 21407 8075
rect 21407 8041 21416 8075
rect 21364 8032 21416 8041
rect 22836 8032 22888 8084
rect 9956 7896 10008 7948
rect 13452 7896 13504 7948
rect 13636 7939 13688 7948
rect 13636 7905 13645 7939
rect 13645 7905 13679 7939
rect 13679 7905 13688 7939
rect 13636 7896 13688 7905
rect 13820 7896 13872 7948
rect 14464 7896 14516 7948
rect 15660 7896 15712 7948
rect 18604 7896 18656 7948
rect 4252 7760 4304 7812
rect 6920 7871 6972 7880
rect 6920 7837 6929 7871
rect 6929 7837 6963 7871
rect 6963 7837 6972 7871
rect 6920 7828 6972 7837
rect 9680 7828 9732 7880
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 15844 7828 15896 7880
rect 16764 7828 16816 7880
rect 18972 7896 19024 7948
rect 20168 7896 20220 7948
rect 3608 7735 3660 7744
rect 3608 7701 3617 7735
rect 3617 7701 3651 7735
rect 3651 7701 3660 7735
rect 3608 7692 3660 7701
rect 4988 7735 5040 7744
rect 4988 7701 4997 7735
rect 4997 7701 5031 7735
rect 5031 7701 5040 7735
rect 4988 7692 5040 7701
rect 5080 7735 5132 7744
rect 5080 7701 5089 7735
rect 5089 7701 5123 7735
rect 5123 7701 5132 7735
rect 8024 7760 8076 7812
rect 8576 7760 8628 7812
rect 11980 7760 12032 7812
rect 15200 7803 15252 7812
rect 15200 7769 15218 7803
rect 15218 7769 15252 7803
rect 15200 7760 15252 7769
rect 16304 7803 16356 7812
rect 16304 7769 16338 7803
rect 16338 7769 16356 7803
rect 16304 7760 16356 7769
rect 16396 7760 16448 7812
rect 16672 7760 16724 7812
rect 19156 7760 19208 7812
rect 19340 7828 19392 7880
rect 21180 7871 21232 7880
rect 21180 7837 21189 7871
rect 21189 7837 21223 7871
rect 21223 7837 21232 7871
rect 21180 7828 21232 7837
rect 21272 7828 21324 7880
rect 23296 7828 23348 7880
rect 21364 7760 21416 7812
rect 22284 7760 22336 7812
rect 5080 7692 5132 7701
rect 7012 7692 7064 7744
rect 9220 7735 9272 7744
rect 9220 7701 9229 7735
rect 9229 7701 9263 7735
rect 9263 7701 9272 7735
rect 9220 7692 9272 7701
rect 11336 7692 11388 7744
rect 12716 7692 12768 7744
rect 15384 7692 15436 7744
rect 17500 7692 17552 7744
rect 18972 7692 19024 7744
rect 19984 7692 20036 7744
rect 20812 7692 20864 7744
rect 22744 7692 22796 7744
rect 6548 7590 6600 7642
rect 6612 7590 6664 7642
rect 6676 7590 6728 7642
rect 6740 7590 6792 7642
rect 6804 7590 6856 7642
rect 12146 7590 12198 7642
rect 12210 7590 12262 7642
rect 12274 7590 12326 7642
rect 12338 7590 12390 7642
rect 12402 7590 12454 7642
rect 17744 7590 17796 7642
rect 17808 7590 17860 7642
rect 17872 7590 17924 7642
rect 17936 7590 17988 7642
rect 18000 7590 18052 7642
rect 1584 7488 1636 7540
rect 2136 7488 2188 7540
rect 5080 7488 5132 7540
rect 5540 7488 5592 7540
rect 11520 7531 11572 7540
rect 1676 7420 1728 7472
rect 2780 7395 2832 7404
rect 2780 7361 2798 7395
rect 2798 7361 2832 7395
rect 2780 7352 2832 7361
rect 4344 7395 4396 7404
rect 4344 7361 4362 7395
rect 4362 7361 4396 7395
rect 4344 7352 4396 7361
rect 4528 7352 4580 7404
rect 8024 7420 8076 7472
rect 9036 7395 9088 7404
rect 11520 7497 11529 7531
rect 11529 7497 11563 7531
rect 11563 7497 11572 7531
rect 11520 7488 11572 7497
rect 11888 7488 11940 7540
rect 12992 7488 13044 7540
rect 14648 7488 14700 7540
rect 15200 7488 15252 7540
rect 11060 7420 11112 7472
rect 19340 7488 19392 7540
rect 17592 7420 17644 7472
rect 18972 7420 19024 7472
rect 20168 7488 20220 7540
rect 20812 7531 20864 7540
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 21364 7488 21416 7540
rect 22192 7488 22244 7540
rect 3056 7327 3108 7336
rect 3056 7293 3065 7327
rect 3065 7293 3099 7327
rect 3099 7293 3108 7327
rect 3056 7284 3108 7293
rect 4620 7327 4672 7336
rect 4620 7293 4629 7327
rect 4629 7293 4663 7327
rect 4663 7293 4672 7327
rect 4620 7284 4672 7293
rect 5816 7216 5868 7268
rect 6368 7216 6420 7268
rect 1768 7148 1820 7200
rect 2688 7148 2740 7200
rect 9036 7361 9054 7395
rect 9054 7361 9088 7395
rect 9036 7352 9088 7361
rect 10600 7395 10652 7404
rect 7380 7284 7432 7336
rect 7840 7284 7892 7336
rect 10600 7361 10609 7395
rect 10609 7361 10643 7395
rect 10643 7361 10652 7395
rect 10600 7352 10652 7361
rect 11336 7395 11388 7404
rect 11336 7361 11345 7395
rect 11345 7361 11379 7395
rect 11379 7361 11388 7395
rect 11336 7352 11388 7361
rect 15384 7352 15436 7404
rect 16120 7352 16172 7404
rect 9956 7284 10008 7336
rect 12164 7327 12216 7336
rect 12164 7293 12173 7327
rect 12173 7293 12207 7327
rect 12207 7293 12216 7327
rect 12164 7284 12216 7293
rect 12808 7284 12860 7336
rect 16856 7284 16908 7336
rect 18236 7284 18288 7336
rect 19800 7352 19852 7404
rect 21548 7420 21600 7472
rect 22928 7420 22980 7472
rect 22192 7352 22244 7404
rect 23020 7395 23072 7404
rect 23020 7361 23029 7395
rect 23029 7361 23063 7395
rect 23063 7361 23072 7395
rect 23020 7352 23072 7361
rect 20168 7327 20220 7336
rect 20168 7293 20177 7327
rect 20177 7293 20211 7327
rect 20211 7293 20220 7327
rect 20168 7284 20220 7293
rect 20352 7327 20404 7336
rect 20352 7293 20361 7327
rect 20361 7293 20395 7327
rect 20395 7293 20404 7327
rect 20352 7284 20404 7293
rect 22376 7327 22428 7336
rect 13820 7216 13872 7268
rect 16212 7259 16264 7268
rect 16212 7225 16221 7259
rect 16221 7225 16255 7259
rect 16255 7225 16264 7259
rect 16212 7216 16264 7225
rect 16764 7216 16816 7268
rect 7564 7191 7616 7200
rect 7564 7157 7573 7191
rect 7573 7157 7607 7191
rect 7607 7157 7616 7191
rect 7564 7148 7616 7157
rect 8116 7148 8168 7200
rect 8576 7148 8628 7200
rect 12992 7191 13044 7200
rect 12992 7157 13001 7191
rect 13001 7157 13035 7191
rect 13035 7157 13044 7191
rect 12992 7148 13044 7157
rect 18604 7148 18656 7200
rect 19616 7216 19668 7268
rect 19800 7216 19852 7268
rect 20260 7216 20312 7268
rect 22376 7293 22385 7327
rect 22385 7293 22419 7327
rect 22419 7293 22428 7327
rect 22376 7284 22428 7293
rect 22744 7284 22796 7336
rect 19340 7148 19392 7200
rect 21732 7148 21784 7200
rect 22100 7216 22152 7268
rect 22744 7148 22796 7200
rect 3749 7046 3801 7098
rect 3813 7046 3865 7098
rect 3877 7046 3929 7098
rect 3941 7046 3993 7098
rect 4005 7046 4057 7098
rect 9347 7046 9399 7098
rect 9411 7046 9463 7098
rect 9475 7046 9527 7098
rect 9539 7046 9591 7098
rect 9603 7046 9655 7098
rect 14945 7046 14997 7098
rect 15009 7046 15061 7098
rect 15073 7046 15125 7098
rect 15137 7046 15189 7098
rect 15201 7046 15253 7098
rect 20543 7046 20595 7098
rect 20607 7046 20659 7098
rect 20671 7046 20723 7098
rect 20735 7046 20787 7098
rect 20799 7046 20851 7098
rect 1676 6987 1728 6996
rect 1676 6953 1685 6987
rect 1685 6953 1719 6987
rect 1719 6953 1728 6987
rect 1676 6944 1728 6953
rect 1860 6851 1912 6860
rect 1860 6817 1869 6851
rect 1869 6817 1903 6851
rect 1903 6817 1912 6851
rect 1860 6808 1912 6817
rect 3056 6808 3108 6860
rect 4620 6944 4672 6996
rect 5448 6944 5500 6996
rect 7564 6944 7616 6996
rect 12164 6987 12216 6996
rect 12164 6953 12173 6987
rect 12173 6953 12207 6987
rect 12207 6953 12216 6987
rect 12164 6944 12216 6953
rect 20168 6944 20220 6996
rect 22100 6944 22152 6996
rect 22192 6944 22244 6996
rect 6184 6851 6236 6860
rect 6184 6817 6193 6851
rect 6193 6817 6227 6851
rect 6227 6817 6236 6851
rect 6184 6808 6236 6817
rect 8300 6808 8352 6860
rect 8576 6851 8628 6860
rect 8576 6817 8585 6851
rect 8585 6817 8619 6851
rect 8619 6817 8628 6851
rect 8576 6808 8628 6817
rect 12072 6808 12124 6860
rect 2596 6740 2648 6792
rect 2964 6715 3016 6724
rect 2964 6681 2973 6715
rect 2973 6681 3007 6715
rect 3007 6681 3016 6715
rect 2964 6672 3016 6681
rect 4252 6783 4304 6792
rect 4252 6749 4286 6783
rect 4286 6749 4304 6783
rect 4252 6740 4304 6749
rect 5540 6740 5592 6792
rect 8668 6740 8720 6792
rect 8116 6672 8168 6724
rect 4988 6604 5040 6656
rect 7196 6604 7248 6656
rect 7472 6604 7524 6656
rect 8576 6604 8628 6656
rect 9956 6672 10008 6724
rect 10416 6672 10468 6724
rect 11888 6740 11940 6792
rect 12164 6740 12216 6792
rect 12716 6740 12768 6792
rect 17500 6851 17552 6860
rect 17500 6817 17509 6851
rect 17509 6817 17543 6851
rect 17543 6817 17552 6851
rect 17500 6808 17552 6817
rect 18420 6851 18472 6860
rect 13636 6740 13688 6792
rect 13176 6672 13228 6724
rect 9036 6604 9088 6656
rect 11980 6604 12032 6656
rect 14832 6647 14884 6656
rect 14832 6613 14841 6647
rect 14841 6613 14875 6647
rect 14875 6613 14884 6647
rect 16396 6740 16448 6792
rect 17316 6740 17368 6792
rect 18420 6817 18429 6851
rect 18429 6817 18463 6851
rect 18463 6817 18472 6851
rect 18420 6808 18472 6817
rect 18604 6876 18656 6928
rect 19156 6876 19208 6928
rect 20812 6876 20864 6928
rect 19432 6808 19484 6860
rect 18236 6740 18288 6792
rect 20812 6783 20864 6792
rect 20812 6749 20821 6783
rect 20821 6749 20855 6783
rect 20855 6749 20864 6783
rect 20812 6740 20864 6749
rect 21180 6740 21232 6792
rect 16672 6715 16724 6724
rect 16672 6681 16690 6715
rect 16690 6681 16724 6715
rect 16672 6672 16724 6681
rect 18144 6715 18196 6724
rect 18144 6681 18153 6715
rect 18153 6681 18187 6715
rect 18187 6681 18196 6715
rect 18144 6672 18196 6681
rect 19432 6672 19484 6724
rect 22192 6740 22244 6792
rect 14832 6604 14884 6613
rect 16580 6604 16632 6656
rect 16764 6604 16816 6656
rect 16948 6604 17000 6656
rect 18604 6647 18656 6656
rect 18604 6613 18613 6647
rect 18613 6613 18647 6647
rect 18647 6613 18656 6647
rect 18604 6604 18656 6613
rect 18696 6647 18748 6656
rect 18696 6613 18705 6647
rect 18705 6613 18739 6647
rect 18739 6613 18748 6647
rect 18696 6604 18748 6613
rect 21456 6672 21508 6724
rect 21548 6672 21600 6724
rect 21916 6672 21968 6724
rect 22652 6740 22704 6792
rect 23388 6808 23440 6860
rect 23020 6647 23072 6656
rect 23020 6613 23029 6647
rect 23029 6613 23063 6647
rect 23063 6613 23072 6647
rect 23020 6604 23072 6613
rect 6548 6502 6600 6554
rect 6612 6502 6664 6554
rect 6676 6502 6728 6554
rect 6740 6502 6792 6554
rect 6804 6502 6856 6554
rect 12146 6502 12198 6554
rect 12210 6502 12262 6554
rect 12274 6502 12326 6554
rect 12338 6502 12390 6554
rect 12402 6502 12454 6554
rect 17744 6502 17796 6554
rect 17808 6502 17860 6554
rect 17872 6502 17924 6554
rect 17936 6502 17988 6554
rect 18000 6502 18052 6554
rect 2320 6400 2372 6452
rect 2780 6443 2832 6452
rect 2780 6409 2789 6443
rect 2789 6409 2823 6443
rect 2823 6409 2832 6443
rect 2780 6400 2832 6409
rect 2964 6400 3016 6452
rect 4528 6400 4580 6452
rect 1768 6307 1820 6316
rect 1768 6273 1777 6307
rect 1777 6273 1811 6307
rect 1811 6273 1820 6307
rect 1768 6264 1820 6273
rect 3332 6264 3384 6316
rect 5540 6400 5592 6452
rect 7012 6443 7064 6452
rect 7012 6409 7021 6443
rect 7021 6409 7055 6443
rect 7055 6409 7064 6443
rect 7012 6400 7064 6409
rect 7472 6443 7524 6452
rect 7472 6409 7481 6443
rect 7481 6409 7515 6443
rect 7515 6409 7524 6443
rect 7472 6400 7524 6409
rect 7564 6400 7616 6452
rect 6184 6307 6236 6316
rect 6184 6273 6193 6307
rect 6193 6273 6227 6307
rect 6227 6273 6236 6307
rect 6184 6264 6236 6273
rect 6368 6307 6420 6316
rect 6368 6273 6377 6307
rect 6377 6273 6411 6307
rect 6411 6273 6420 6307
rect 6368 6264 6420 6273
rect 7196 6332 7248 6384
rect 7472 6264 7524 6316
rect 7840 6264 7892 6316
rect 8024 6307 8076 6316
rect 8024 6273 8033 6307
rect 8033 6273 8067 6307
rect 8067 6273 8076 6307
rect 8024 6264 8076 6273
rect 9036 6332 9088 6384
rect 9220 6332 9272 6384
rect 13084 6400 13136 6452
rect 13176 6400 13228 6452
rect 14740 6400 14792 6452
rect 16764 6400 16816 6452
rect 16948 6443 17000 6452
rect 16948 6409 16957 6443
rect 16957 6409 16991 6443
rect 16991 6409 17000 6443
rect 16948 6400 17000 6409
rect 19984 6400 20036 6452
rect 22376 6400 22428 6452
rect 12072 6332 12124 6384
rect 7748 6196 7800 6248
rect 8576 6264 8628 6316
rect 9956 6307 10008 6316
rect 5172 6128 5224 6180
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 10968 6264 11020 6316
rect 11980 6239 12032 6248
rect 11980 6205 11989 6239
rect 11989 6205 12023 6239
rect 12023 6205 12032 6239
rect 11980 6196 12032 6205
rect 12808 6307 12860 6316
rect 12808 6273 12817 6307
rect 12817 6273 12851 6307
rect 12851 6273 12860 6307
rect 12808 6264 12860 6273
rect 14832 6332 14884 6384
rect 18144 6375 18196 6384
rect 18144 6341 18153 6375
rect 18153 6341 18187 6375
rect 18187 6341 18196 6375
rect 18144 6332 18196 6341
rect 22284 6332 22336 6384
rect 13636 6264 13688 6316
rect 15108 6307 15160 6316
rect 15108 6273 15117 6307
rect 15117 6273 15151 6307
rect 15151 6273 15160 6307
rect 15108 6264 15160 6273
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 17500 6307 17552 6316
rect 17500 6273 17509 6307
rect 17509 6273 17543 6307
rect 17543 6273 17552 6307
rect 17500 6264 17552 6273
rect 18236 6307 18288 6316
rect 18236 6273 18245 6307
rect 18245 6273 18279 6307
rect 18279 6273 18288 6307
rect 18236 6264 18288 6273
rect 18328 6264 18380 6316
rect 19340 6264 19392 6316
rect 9772 6128 9824 6180
rect 13176 6196 13228 6248
rect 13268 6239 13320 6248
rect 13268 6205 13280 6239
rect 13280 6205 13314 6239
rect 13314 6205 13320 6239
rect 13268 6196 13320 6205
rect 13452 6196 13504 6248
rect 17132 6196 17184 6248
rect 19708 6239 19760 6248
rect 19708 6205 19717 6239
rect 19717 6205 19751 6239
rect 19751 6205 19760 6239
rect 19708 6196 19760 6205
rect 20904 6264 20956 6316
rect 23112 6264 23164 6316
rect 21916 6239 21968 6248
rect 21916 6205 21925 6239
rect 21925 6205 21959 6239
rect 21959 6205 21968 6239
rect 21916 6196 21968 6205
rect 8392 6060 8444 6112
rect 9864 6060 9916 6112
rect 11888 6060 11940 6112
rect 13636 6060 13688 6112
rect 14648 6103 14700 6112
rect 14648 6069 14657 6103
rect 14657 6069 14691 6103
rect 14691 6069 14700 6103
rect 14648 6060 14700 6069
rect 16948 6060 17000 6112
rect 17408 6103 17460 6112
rect 17408 6069 17417 6103
rect 17417 6069 17451 6103
rect 17451 6069 17460 6103
rect 17408 6060 17460 6069
rect 19432 6060 19484 6112
rect 20168 6060 20220 6112
rect 20260 6060 20312 6112
rect 23020 6103 23072 6112
rect 23020 6069 23029 6103
rect 23029 6069 23063 6103
rect 23063 6069 23072 6103
rect 23020 6060 23072 6069
rect 3749 5958 3801 6010
rect 3813 5958 3865 6010
rect 3877 5958 3929 6010
rect 3941 5958 3993 6010
rect 4005 5958 4057 6010
rect 9347 5958 9399 6010
rect 9411 5958 9463 6010
rect 9475 5958 9527 6010
rect 9539 5958 9591 6010
rect 9603 5958 9655 6010
rect 14945 5958 14997 6010
rect 15009 5958 15061 6010
rect 15073 5958 15125 6010
rect 15137 5958 15189 6010
rect 15201 5958 15253 6010
rect 20543 5958 20595 6010
rect 20607 5958 20659 6010
rect 20671 5958 20723 6010
rect 20735 5958 20787 6010
rect 20799 5958 20851 6010
rect 4344 5856 4396 5908
rect 4620 5899 4672 5908
rect 4620 5865 4629 5899
rect 4629 5865 4663 5899
rect 4663 5865 4672 5899
rect 4620 5856 4672 5865
rect 4804 5856 4856 5908
rect 5356 5856 5408 5908
rect 6368 5856 6420 5908
rect 8024 5856 8076 5908
rect 3700 5652 3752 5704
rect 4804 5720 4856 5772
rect 5448 5763 5500 5772
rect 5448 5729 5464 5763
rect 5464 5729 5498 5763
rect 5498 5729 5500 5763
rect 5448 5720 5500 5729
rect 8484 5720 8536 5772
rect 10324 5720 10376 5772
rect 12808 5856 12860 5908
rect 13636 5856 13688 5908
rect 14096 5856 14148 5908
rect 11888 5763 11940 5772
rect 11888 5729 11900 5763
rect 11900 5729 11934 5763
rect 11934 5729 11940 5763
rect 11888 5720 11940 5729
rect 5264 5652 5316 5704
rect 5356 5695 5408 5704
rect 5356 5661 5365 5695
rect 5365 5661 5399 5695
rect 5399 5661 5408 5695
rect 5356 5652 5408 5661
rect 3516 5584 3568 5636
rect 4528 5516 4580 5568
rect 5080 5516 5132 5568
rect 5172 5516 5224 5568
rect 5816 5584 5868 5636
rect 8392 5652 8444 5704
rect 12992 5720 13044 5772
rect 20260 5856 20312 5908
rect 15200 5788 15252 5840
rect 16672 5831 16724 5840
rect 16672 5797 16681 5831
rect 16681 5797 16715 5831
rect 16715 5797 16724 5831
rect 19892 5831 19944 5840
rect 16672 5788 16724 5797
rect 19892 5797 19901 5831
rect 19901 5797 19935 5831
rect 19935 5797 19944 5831
rect 19892 5788 19944 5797
rect 21456 5856 21508 5908
rect 12624 5652 12676 5704
rect 13728 5627 13780 5636
rect 13728 5593 13737 5627
rect 13737 5593 13771 5627
rect 13771 5593 13780 5627
rect 13728 5584 13780 5593
rect 6460 5516 6512 5568
rect 10692 5516 10744 5568
rect 12072 5516 12124 5568
rect 13360 5516 13412 5568
rect 15292 5652 15344 5704
rect 16764 5720 16816 5772
rect 18696 5720 18748 5772
rect 19432 5720 19484 5772
rect 22928 5763 22980 5772
rect 22928 5729 22937 5763
rect 22937 5729 22971 5763
rect 22971 5729 22980 5763
rect 22928 5720 22980 5729
rect 15384 5584 15436 5636
rect 17408 5695 17460 5704
rect 17408 5661 17417 5695
rect 17417 5661 17451 5695
rect 17451 5661 17460 5695
rect 17408 5652 17460 5661
rect 18236 5652 18288 5704
rect 20720 5652 20772 5704
rect 21180 5652 21232 5704
rect 21548 5652 21600 5704
rect 16396 5584 16448 5636
rect 17224 5627 17276 5636
rect 15200 5516 15252 5568
rect 17224 5593 17233 5627
rect 17233 5593 17267 5627
rect 17267 5593 17276 5627
rect 17224 5584 17276 5593
rect 18144 5584 18196 5636
rect 18880 5584 18932 5636
rect 20260 5584 20312 5636
rect 16764 5516 16816 5568
rect 17592 5559 17644 5568
rect 17592 5525 17601 5559
rect 17601 5525 17635 5559
rect 17635 5525 17644 5559
rect 17592 5516 17644 5525
rect 18420 5516 18472 5568
rect 19708 5559 19760 5568
rect 19708 5525 19717 5559
rect 19717 5525 19751 5559
rect 19751 5525 19760 5559
rect 19708 5516 19760 5525
rect 22100 5584 22152 5636
rect 22376 5516 22428 5568
rect 6548 5414 6600 5466
rect 6612 5414 6664 5466
rect 6676 5414 6728 5466
rect 6740 5414 6792 5466
rect 6804 5414 6856 5466
rect 12146 5414 12198 5466
rect 12210 5414 12262 5466
rect 12274 5414 12326 5466
rect 12338 5414 12390 5466
rect 12402 5414 12454 5466
rect 17744 5414 17796 5466
rect 17808 5414 17860 5466
rect 17872 5414 17924 5466
rect 17936 5414 17988 5466
rect 18000 5414 18052 5466
rect 5172 5312 5224 5364
rect 5264 5312 5316 5364
rect 6184 5355 6236 5364
rect 6184 5321 6193 5355
rect 6193 5321 6227 5355
rect 6227 5321 6236 5355
rect 6184 5312 6236 5321
rect 6460 5312 6512 5364
rect 7840 5312 7892 5364
rect 8852 5312 8904 5364
rect 10692 5355 10744 5364
rect 10692 5321 10701 5355
rect 10701 5321 10735 5355
rect 10735 5321 10744 5355
rect 10692 5312 10744 5321
rect 11980 5312 12032 5364
rect 12624 5312 12676 5364
rect 5080 5287 5132 5296
rect 4620 5176 4672 5228
rect 4804 5219 4856 5228
rect 4804 5185 4813 5219
rect 4813 5185 4847 5219
rect 4847 5185 4856 5219
rect 4804 5176 4856 5185
rect 5080 5253 5114 5287
rect 5114 5253 5132 5287
rect 5080 5244 5132 5253
rect 5540 5244 5592 5296
rect 7380 5244 7432 5296
rect 6368 5108 6420 5160
rect 6920 5176 6972 5228
rect 7748 5151 7800 5160
rect 7380 5040 7432 5092
rect 5448 4972 5500 5024
rect 7104 4972 7156 5024
rect 7748 5117 7757 5151
rect 7757 5117 7791 5151
rect 7791 5117 7800 5151
rect 7748 5108 7800 5117
rect 8668 5244 8720 5296
rect 9680 5244 9732 5296
rect 12808 5244 12860 5296
rect 12992 5287 13044 5296
rect 12992 5253 13001 5287
rect 13001 5253 13035 5287
rect 13035 5253 13044 5287
rect 12992 5244 13044 5253
rect 8300 5176 8352 5228
rect 10324 5219 10376 5228
rect 10324 5185 10333 5219
rect 10333 5185 10367 5219
rect 10367 5185 10376 5219
rect 10324 5176 10376 5185
rect 11336 5176 11388 5228
rect 16120 5176 16172 5228
rect 16488 5312 16540 5364
rect 16580 5312 16632 5364
rect 17040 5312 17092 5364
rect 17592 5312 17644 5364
rect 18604 5355 18656 5364
rect 18604 5321 18613 5355
rect 18613 5321 18647 5355
rect 18647 5321 18656 5355
rect 18604 5312 18656 5321
rect 18880 5312 18932 5364
rect 19340 5312 19392 5364
rect 20260 5355 20312 5364
rect 20260 5321 20269 5355
rect 20269 5321 20303 5355
rect 20303 5321 20312 5355
rect 20260 5312 20312 5321
rect 21824 5312 21876 5364
rect 22192 5355 22244 5364
rect 22192 5321 22201 5355
rect 22201 5321 22235 5355
rect 22235 5321 22244 5355
rect 22192 5312 22244 5321
rect 16948 5176 17000 5228
rect 17684 5176 17736 5228
rect 19524 5244 19576 5296
rect 18972 5219 19024 5228
rect 18972 5185 18981 5219
rect 18981 5185 19015 5219
rect 19015 5185 19024 5219
rect 18972 5176 19024 5185
rect 19432 5176 19484 5228
rect 21732 5244 21784 5296
rect 23204 5244 23256 5296
rect 21640 5219 21692 5228
rect 21640 5185 21649 5219
rect 21649 5185 21683 5219
rect 21683 5185 21692 5219
rect 21640 5176 21692 5185
rect 22836 5219 22888 5228
rect 22836 5185 22845 5219
rect 22845 5185 22879 5219
rect 22879 5185 22888 5219
rect 22836 5176 22888 5185
rect 9220 5108 9272 5160
rect 10508 5151 10560 5160
rect 10508 5117 10517 5151
rect 10517 5117 10551 5151
rect 10551 5117 10560 5151
rect 10508 5108 10560 5117
rect 12624 5108 12676 5160
rect 14740 5151 14792 5160
rect 14464 5040 14516 5092
rect 14740 5117 14749 5151
rect 14749 5117 14783 5151
rect 14783 5117 14792 5151
rect 14740 5108 14792 5117
rect 16396 5108 16448 5160
rect 17316 5108 17368 5160
rect 17592 5151 17644 5160
rect 17592 5117 17601 5151
rect 17601 5117 17635 5151
rect 17635 5117 17644 5151
rect 17592 5108 17644 5117
rect 11428 4972 11480 5024
rect 13268 4972 13320 5024
rect 13452 4972 13504 5024
rect 18788 5040 18840 5092
rect 19248 5040 19300 5092
rect 19800 5040 19852 5092
rect 21824 5108 21876 5160
rect 22284 5108 22336 5160
rect 19984 5040 20036 5092
rect 21732 5040 21784 5092
rect 17500 4972 17552 5024
rect 19892 4972 19944 5024
rect 21640 4972 21692 5024
rect 23112 4972 23164 5024
rect 3749 4870 3801 4922
rect 3813 4870 3865 4922
rect 3877 4870 3929 4922
rect 3941 4870 3993 4922
rect 4005 4870 4057 4922
rect 9347 4870 9399 4922
rect 9411 4870 9463 4922
rect 9475 4870 9527 4922
rect 9539 4870 9591 4922
rect 9603 4870 9655 4922
rect 14945 4870 14997 4922
rect 15009 4870 15061 4922
rect 15073 4870 15125 4922
rect 15137 4870 15189 4922
rect 15201 4870 15253 4922
rect 20543 4870 20595 4922
rect 20607 4870 20659 4922
rect 20671 4870 20723 4922
rect 20735 4870 20787 4922
rect 20799 4870 20851 4922
rect 2872 4607 2924 4616
rect 2872 4573 2881 4607
rect 2881 4573 2915 4607
rect 2915 4573 2924 4607
rect 2872 4564 2924 4573
rect 4160 4768 4212 4820
rect 5816 4768 5868 4820
rect 6184 4768 6236 4820
rect 6552 4768 6604 4820
rect 6920 4811 6972 4820
rect 6920 4777 6929 4811
rect 6929 4777 6963 4811
rect 6963 4777 6972 4811
rect 6920 4768 6972 4777
rect 7472 4768 7524 4820
rect 6368 4675 6420 4684
rect 6368 4641 6377 4675
rect 6377 4641 6411 4675
rect 6411 4641 6420 4675
rect 6368 4632 6420 4641
rect 5356 4607 5408 4616
rect 2964 4539 3016 4548
rect 2964 4505 2973 4539
rect 2973 4505 3007 4539
rect 3007 4505 3016 4539
rect 2964 4496 3016 4505
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 6460 4564 6512 4616
rect 6552 4607 6604 4616
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 6184 4496 6236 4548
rect 7196 4496 7248 4548
rect 9864 4768 9916 4820
rect 10416 4811 10468 4820
rect 10416 4777 10425 4811
rect 10425 4777 10459 4811
rect 10459 4777 10468 4811
rect 10416 4768 10468 4777
rect 10600 4811 10652 4820
rect 10600 4777 10609 4811
rect 10609 4777 10643 4811
rect 10643 4777 10652 4811
rect 10600 4768 10652 4777
rect 10232 4700 10284 4752
rect 7840 4607 7892 4616
rect 7840 4573 7849 4607
rect 7849 4573 7883 4607
rect 7883 4573 7892 4607
rect 7840 4564 7892 4573
rect 10508 4632 10560 4684
rect 11796 4768 11848 4820
rect 8852 4564 8904 4616
rect 9220 4564 9272 4616
rect 9772 4607 9824 4616
rect 2228 4471 2280 4480
rect 2228 4437 2237 4471
rect 2237 4437 2271 4471
rect 2271 4437 2280 4471
rect 2228 4428 2280 4437
rect 5080 4428 5132 4480
rect 6276 4428 6328 4480
rect 7012 4471 7064 4480
rect 7012 4437 7021 4471
rect 7021 4437 7055 4471
rect 7055 4437 7064 4471
rect 7380 4471 7432 4480
rect 7012 4428 7064 4437
rect 7380 4437 7389 4471
rect 7389 4437 7423 4471
rect 7423 4437 7432 4471
rect 7380 4428 7432 4437
rect 9772 4573 9781 4607
rect 9781 4573 9815 4607
rect 9815 4573 9824 4607
rect 9772 4564 9824 4573
rect 16488 4768 16540 4820
rect 18052 4811 18104 4820
rect 18052 4777 18061 4811
rect 18061 4777 18095 4811
rect 18095 4777 18104 4811
rect 18052 4768 18104 4777
rect 18880 4768 18932 4820
rect 19248 4811 19300 4820
rect 19248 4777 19257 4811
rect 19257 4777 19291 4811
rect 19291 4777 19300 4811
rect 19248 4768 19300 4777
rect 19432 4811 19484 4820
rect 19432 4777 19441 4811
rect 19441 4777 19475 4811
rect 19475 4777 19484 4811
rect 19432 4768 19484 4777
rect 19524 4768 19576 4820
rect 21548 4811 21600 4820
rect 15016 4743 15068 4752
rect 15016 4709 15025 4743
rect 15025 4709 15059 4743
rect 15059 4709 15068 4743
rect 15016 4700 15068 4709
rect 15476 4632 15528 4684
rect 17132 4700 17184 4752
rect 18236 4700 18288 4752
rect 18972 4700 19024 4752
rect 16948 4632 17000 4684
rect 12532 4564 12584 4616
rect 11060 4496 11112 4548
rect 13452 4496 13504 4548
rect 8392 4428 8444 4480
rect 11336 4471 11388 4480
rect 11336 4437 11345 4471
rect 11345 4437 11379 4471
rect 11379 4437 11388 4471
rect 11336 4428 11388 4437
rect 11428 4471 11480 4480
rect 11428 4437 11437 4471
rect 11437 4437 11471 4471
rect 11471 4437 11480 4471
rect 11428 4428 11480 4437
rect 12624 4428 12676 4480
rect 14280 4428 14332 4480
rect 14648 4428 14700 4480
rect 16396 4564 16448 4616
rect 17224 4564 17276 4616
rect 17592 4632 17644 4684
rect 21548 4777 21557 4811
rect 21557 4777 21591 4811
rect 21591 4777 21600 4811
rect 21548 4768 21600 4777
rect 21088 4632 21140 4684
rect 21180 4632 21232 4684
rect 19432 4564 19484 4616
rect 19892 4564 19944 4616
rect 20904 4564 20956 4616
rect 21272 4564 21324 4616
rect 21456 4564 21508 4616
rect 16580 4428 16632 4480
rect 16856 4471 16908 4480
rect 16856 4437 16865 4471
rect 16865 4437 16899 4471
rect 16899 4437 16908 4471
rect 16856 4428 16908 4437
rect 16948 4471 17000 4480
rect 16948 4437 16957 4471
rect 16957 4437 16991 4471
rect 16991 4437 17000 4471
rect 16948 4428 17000 4437
rect 17500 4428 17552 4480
rect 18236 4428 18288 4480
rect 19524 4428 19576 4480
rect 19800 4471 19852 4480
rect 19800 4437 19809 4471
rect 19809 4437 19843 4471
rect 19843 4437 19852 4471
rect 19800 4428 19852 4437
rect 21088 4496 21140 4548
rect 20996 4428 21048 4480
rect 21732 4496 21784 4548
rect 23020 4428 23072 4480
rect 6548 4326 6600 4378
rect 6612 4326 6664 4378
rect 6676 4326 6728 4378
rect 6740 4326 6792 4378
rect 6804 4326 6856 4378
rect 12146 4326 12198 4378
rect 12210 4326 12262 4378
rect 12274 4326 12326 4378
rect 12338 4326 12390 4378
rect 12402 4326 12454 4378
rect 17744 4326 17796 4378
rect 17808 4326 17860 4378
rect 17872 4326 17924 4378
rect 17936 4326 17988 4378
rect 18000 4326 18052 4378
rect 2872 4224 2924 4276
rect 5172 4224 5224 4276
rect 4528 4088 4580 4140
rect 7012 4224 7064 4276
rect 7288 4267 7340 4276
rect 7288 4233 7297 4267
rect 7297 4233 7331 4267
rect 7331 4233 7340 4267
rect 7288 4224 7340 4233
rect 7840 4224 7892 4276
rect 8944 4224 8996 4276
rect 12808 4224 12860 4276
rect 13452 4267 13504 4276
rect 13452 4233 13461 4267
rect 13461 4233 13495 4267
rect 13495 4233 13504 4267
rect 13452 4224 13504 4233
rect 16856 4224 16908 4276
rect 9036 4156 9088 4208
rect 7196 4088 7248 4140
rect 7288 4088 7340 4140
rect 7748 4088 7800 4140
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 3976 3995 4028 4004
rect 3976 3961 3985 3995
rect 3985 3961 4019 3995
rect 4019 3961 4028 3995
rect 3976 3952 4028 3961
rect 5816 3952 5868 4004
rect 6184 3995 6236 4004
rect 6184 3961 6193 3995
rect 6193 3961 6227 3995
rect 6227 3961 6236 3995
rect 6184 3952 6236 3961
rect 7012 4020 7064 4072
rect 8208 4063 8260 4072
rect 8208 4029 8217 4063
rect 8217 4029 8251 4063
rect 8251 4029 8260 4063
rect 8208 4020 8260 4029
rect 8484 4088 8536 4140
rect 11428 4156 11480 4208
rect 16580 4156 16632 4208
rect 10600 4088 10652 4140
rect 11336 4088 11388 4140
rect 13360 4131 13412 4140
rect 13360 4097 13369 4131
rect 13369 4097 13403 4131
rect 13403 4097 13412 4131
rect 13360 4088 13412 4097
rect 13820 4088 13872 4140
rect 14280 4088 14332 4140
rect 17592 4224 17644 4276
rect 19156 4267 19208 4276
rect 17868 4156 17920 4208
rect 17500 4131 17552 4140
rect 8392 3952 8444 4004
rect 3424 3884 3476 3936
rect 6092 3884 6144 3936
rect 6920 3884 6972 3936
rect 10876 4063 10928 4072
rect 10508 3952 10560 4004
rect 10876 4029 10885 4063
rect 10885 4029 10919 4063
rect 10919 4029 10928 4063
rect 10876 4020 10928 4029
rect 14004 4020 14056 4072
rect 14096 4020 14148 4072
rect 9864 3884 9916 3936
rect 11244 3884 11296 3936
rect 11520 3927 11572 3936
rect 11520 3893 11529 3927
rect 11529 3893 11563 3927
rect 11563 3893 11572 3927
rect 11520 3884 11572 3893
rect 12532 3884 12584 3936
rect 17500 4097 17509 4131
rect 17509 4097 17543 4131
rect 17543 4097 17552 4131
rect 17500 4088 17552 4097
rect 18328 4088 18380 4140
rect 18420 4131 18472 4140
rect 18420 4097 18429 4131
rect 18429 4097 18463 4131
rect 18463 4097 18472 4131
rect 19156 4233 19165 4267
rect 19165 4233 19199 4267
rect 19199 4233 19208 4267
rect 19156 4224 19208 4233
rect 19616 4224 19668 4276
rect 19800 4224 19852 4276
rect 18420 4088 18472 4097
rect 17316 4063 17368 4072
rect 17316 4029 17325 4063
rect 17325 4029 17359 4063
rect 17359 4029 17368 4063
rect 17316 4020 17368 4029
rect 17684 4020 17736 4072
rect 18972 4088 19024 4140
rect 19248 4131 19300 4140
rect 19248 4097 19257 4131
rect 19257 4097 19291 4131
rect 19291 4097 19300 4131
rect 19248 4088 19300 4097
rect 19064 4063 19116 4072
rect 13912 3884 13964 3936
rect 14556 3927 14608 3936
rect 14556 3893 14565 3927
rect 14565 3893 14599 3927
rect 14599 3893 14608 3927
rect 14556 3884 14608 3893
rect 14832 3884 14884 3936
rect 15292 3884 15344 3936
rect 19064 4029 19073 4063
rect 19073 4029 19107 4063
rect 19107 4029 19116 4063
rect 19064 4020 19116 4029
rect 20076 4088 20128 4140
rect 20352 4156 20404 4208
rect 20996 4156 21048 4208
rect 21364 4156 21416 4208
rect 21456 4156 21508 4208
rect 21640 4156 21692 4208
rect 22468 4156 22520 4208
rect 22744 4199 22796 4208
rect 22744 4165 22753 4199
rect 22753 4165 22787 4199
rect 22787 4165 22796 4199
rect 22744 4156 22796 4165
rect 23020 4088 23072 4140
rect 20260 4063 20312 4072
rect 17868 3952 17920 4004
rect 20260 4029 20269 4063
rect 20269 4029 20303 4063
rect 20303 4029 20312 4063
rect 20260 4020 20312 4029
rect 21272 4020 21324 4072
rect 19984 3995 20036 4004
rect 19984 3961 19993 3995
rect 19993 3961 20027 3995
rect 20027 3961 20036 3995
rect 19984 3952 20036 3961
rect 19064 3884 19116 3936
rect 19616 3927 19668 3936
rect 19616 3893 19625 3927
rect 19625 3893 19659 3927
rect 19659 3893 19668 3927
rect 19616 3884 19668 3893
rect 19800 3884 19852 3936
rect 21732 3884 21784 3936
rect 22008 3952 22060 4004
rect 3749 3782 3801 3834
rect 3813 3782 3865 3834
rect 3877 3782 3929 3834
rect 3941 3782 3993 3834
rect 4005 3782 4057 3834
rect 9347 3782 9399 3834
rect 9411 3782 9463 3834
rect 9475 3782 9527 3834
rect 9539 3782 9591 3834
rect 9603 3782 9655 3834
rect 14945 3782 14997 3834
rect 15009 3782 15061 3834
rect 15073 3782 15125 3834
rect 15137 3782 15189 3834
rect 15201 3782 15253 3834
rect 20543 3782 20595 3834
rect 20607 3782 20659 3834
rect 20671 3782 20723 3834
rect 20735 3782 20787 3834
rect 20799 3782 20851 3834
rect 2044 3476 2096 3528
rect 1400 3383 1452 3392
rect 1400 3349 1409 3383
rect 1409 3349 1443 3383
rect 1443 3349 1452 3383
rect 1400 3340 1452 3349
rect 2964 3383 3016 3392
rect 2964 3349 2973 3383
rect 2973 3349 3007 3383
rect 3007 3349 3016 3383
rect 2964 3340 3016 3349
rect 7196 3612 7248 3664
rect 11060 3612 11112 3664
rect 12072 3612 12124 3664
rect 12440 3655 12492 3664
rect 12440 3621 12449 3655
rect 12449 3621 12483 3655
rect 12483 3621 12492 3655
rect 12440 3612 12492 3621
rect 13820 3680 13872 3732
rect 15292 3680 15344 3732
rect 15476 3723 15528 3732
rect 15476 3689 15485 3723
rect 15485 3689 15519 3723
rect 15519 3689 15528 3723
rect 15476 3680 15528 3689
rect 16948 3680 17000 3732
rect 19800 3680 19852 3732
rect 22652 3680 22704 3732
rect 22836 3680 22888 3732
rect 3516 3544 3568 3596
rect 4712 3544 4764 3596
rect 4804 3544 4856 3596
rect 7104 3519 7156 3528
rect 7104 3485 7113 3519
rect 7113 3485 7147 3519
rect 7147 3485 7156 3519
rect 7104 3476 7156 3485
rect 8484 3476 8536 3528
rect 9220 3476 9272 3528
rect 10600 3476 10652 3528
rect 12532 3519 12584 3528
rect 12532 3485 12541 3519
rect 12541 3485 12575 3519
rect 12575 3485 12584 3519
rect 12532 3476 12584 3485
rect 16396 3476 16448 3528
rect 5908 3408 5960 3460
rect 6184 3340 6236 3392
rect 6460 3340 6512 3392
rect 6920 3340 6972 3392
rect 9680 3408 9732 3460
rect 11152 3408 11204 3460
rect 12072 3408 12124 3460
rect 14188 3408 14240 3460
rect 14556 3408 14608 3460
rect 17684 3587 17736 3596
rect 17684 3553 17693 3587
rect 17693 3553 17727 3587
rect 17727 3553 17736 3587
rect 17684 3544 17736 3553
rect 19432 3587 19484 3596
rect 18236 3476 18288 3528
rect 19432 3553 19441 3587
rect 19441 3553 19475 3587
rect 19475 3553 19484 3587
rect 19432 3544 19484 3553
rect 20260 3587 20312 3596
rect 20260 3553 20269 3587
rect 20269 3553 20303 3587
rect 20303 3553 20312 3587
rect 20260 3544 20312 3553
rect 18972 3476 19024 3528
rect 19616 3519 19668 3528
rect 19616 3485 19625 3519
rect 19625 3485 19659 3519
rect 19659 3485 19668 3519
rect 19616 3476 19668 3485
rect 21272 3476 21324 3528
rect 8392 3340 8444 3392
rect 10876 3340 10928 3392
rect 10968 3340 11020 3392
rect 13636 3340 13688 3392
rect 13728 3340 13780 3392
rect 16764 3340 16816 3392
rect 17684 3408 17736 3460
rect 17408 3383 17460 3392
rect 17408 3349 17417 3383
rect 17417 3349 17451 3383
rect 17451 3349 17460 3383
rect 17408 3340 17460 3349
rect 18144 3383 18196 3392
rect 18144 3349 18153 3383
rect 18153 3349 18187 3383
rect 18187 3349 18196 3383
rect 18144 3340 18196 3349
rect 18328 3340 18380 3392
rect 20536 3451 20588 3460
rect 20536 3417 20570 3451
rect 20570 3417 20588 3451
rect 20536 3408 20588 3417
rect 20720 3408 20772 3460
rect 21272 3340 21324 3392
rect 21640 3383 21692 3392
rect 21640 3349 21649 3383
rect 21649 3349 21683 3383
rect 21683 3349 21692 3383
rect 21640 3340 21692 3349
rect 6548 3238 6600 3290
rect 6612 3238 6664 3290
rect 6676 3238 6728 3290
rect 6740 3238 6792 3290
rect 6804 3238 6856 3290
rect 12146 3238 12198 3290
rect 12210 3238 12262 3290
rect 12274 3238 12326 3290
rect 12338 3238 12390 3290
rect 12402 3238 12454 3290
rect 17744 3238 17796 3290
rect 17808 3238 17860 3290
rect 17872 3238 17924 3290
rect 17936 3238 17988 3290
rect 18000 3238 18052 3290
rect 2504 3179 2556 3188
rect 2504 3145 2513 3179
rect 2513 3145 2547 3179
rect 2547 3145 2556 3179
rect 2504 3136 2556 3145
rect 3240 3179 3292 3188
rect 3240 3145 3249 3179
rect 3249 3145 3283 3179
rect 3283 3145 3292 3179
rect 3240 3136 3292 3145
rect 5908 3136 5960 3188
rect 6000 3136 6052 3188
rect 6184 3179 6236 3188
rect 6184 3145 6193 3179
rect 6193 3145 6227 3179
rect 6227 3145 6236 3179
rect 6184 3136 6236 3145
rect 6460 3136 6512 3188
rect 2044 3111 2096 3120
rect 2044 3077 2053 3111
rect 2053 3077 2087 3111
rect 2087 3077 2096 3111
rect 2044 3068 2096 3077
rect 1584 3043 1636 3052
rect 1584 3009 1593 3043
rect 1593 3009 1627 3043
rect 1627 3009 1636 3043
rect 1584 3000 1636 3009
rect 3516 3068 3568 3120
rect 10968 3136 11020 3188
rect 11336 3179 11388 3188
rect 11336 3145 11345 3179
rect 11345 3145 11379 3179
rect 11379 3145 11388 3179
rect 11336 3136 11388 3145
rect 12072 3136 12124 3188
rect 2504 3000 2556 3052
rect 7196 3068 7248 3120
rect 8944 3111 8996 3120
rect 8944 3077 8953 3111
rect 8953 3077 8987 3111
rect 8987 3077 8996 3111
rect 8944 3068 8996 3077
rect 1860 2796 1912 2848
rect 3332 2839 3384 2848
rect 3332 2805 3341 2839
rect 3341 2805 3375 2839
rect 3375 2805 3384 2839
rect 4804 3043 4856 3052
rect 4804 3009 4813 3043
rect 4813 3009 4847 3043
rect 4847 3009 4856 3043
rect 5080 3043 5132 3052
rect 4804 3000 4856 3009
rect 5080 3009 5114 3043
rect 5114 3009 5132 3043
rect 5080 3000 5132 3009
rect 8392 3000 8444 3052
rect 10324 3043 10376 3052
rect 10324 3009 10342 3043
rect 10342 3009 10376 3043
rect 10324 3000 10376 3009
rect 10600 3043 10652 3052
rect 10600 3009 10609 3043
rect 10609 3009 10643 3043
rect 10643 3009 10652 3043
rect 10600 3000 10652 3009
rect 11060 3000 11112 3052
rect 6368 2932 6420 2984
rect 9128 2975 9180 2984
rect 9128 2941 9137 2975
rect 9137 2941 9171 2975
rect 9171 2941 9180 2975
rect 9128 2932 9180 2941
rect 6828 2864 6880 2916
rect 3332 2796 3384 2805
rect 6276 2796 6328 2848
rect 8300 2796 8352 2848
rect 9680 2796 9732 2848
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 12532 3136 12584 3188
rect 13912 3179 13964 3188
rect 13912 3145 13921 3179
rect 13921 3145 13955 3179
rect 13955 3145 13964 3179
rect 13912 3136 13964 3145
rect 14556 3179 14608 3188
rect 14556 3145 14565 3179
rect 14565 3145 14599 3179
rect 14599 3145 14608 3179
rect 14556 3136 14608 3145
rect 14740 3136 14792 3188
rect 20812 3136 20864 3188
rect 21364 3136 21416 3188
rect 12624 3068 12676 3120
rect 13820 3111 13872 3120
rect 13820 3077 13829 3111
rect 13829 3077 13863 3111
rect 13863 3077 13872 3111
rect 13820 3068 13872 3077
rect 14096 3111 14148 3120
rect 14096 3077 14105 3111
rect 14105 3077 14139 3111
rect 14139 3077 14148 3111
rect 14096 3068 14148 3077
rect 14096 2932 14148 2984
rect 14648 3000 14700 3052
rect 15660 3000 15712 3052
rect 16212 3043 16264 3052
rect 16212 3009 16230 3043
rect 16230 3009 16264 3043
rect 16212 3000 16264 3009
rect 16396 3000 16448 3052
rect 16580 3000 16632 3052
rect 16764 3000 16816 3052
rect 19340 3068 19392 3120
rect 14464 2932 14516 2984
rect 14004 2864 14056 2916
rect 14280 2864 14332 2916
rect 13728 2796 13780 2848
rect 14372 2839 14424 2848
rect 14372 2805 14381 2839
rect 14381 2805 14415 2839
rect 14415 2805 14424 2839
rect 14372 2796 14424 2805
rect 17408 2796 17460 2848
rect 18420 3043 18472 3052
rect 18420 3009 18454 3043
rect 18454 3009 18472 3043
rect 18420 3000 18472 3009
rect 20444 3000 20496 3052
rect 21180 3068 21232 3120
rect 21548 3068 21600 3120
rect 21272 3043 21324 3052
rect 21272 3009 21281 3043
rect 21281 3009 21315 3043
rect 21315 3009 21324 3043
rect 21272 3000 21324 3009
rect 21364 3043 21416 3052
rect 21364 3009 21373 3043
rect 21373 3009 21407 3043
rect 21407 3009 21416 3043
rect 21364 3000 21416 3009
rect 22652 3043 22704 3052
rect 18144 2864 18196 2916
rect 19248 2864 19300 2916
rect 19156 2796 19208 2848
rect 22100 2932 22152 2984
rect 22652 3009 22661 3043
rect 22661 3009 22695 3043
rect 22695 3009 22704 3043
rect 22652 3000 22704 3009
rect 22468 2975 22520 2984
rect 22468 2941 22477 2975
rect 22477 2941 22511 2975
rect 22511 2941 22520 2975
rect 22468 2932 22520 2941
rect 22836 2975 22888 2984
rect 22836 2941 22845 2975
rect 22845 2941 22879 2975
rect 22879 2941 22888 2975
rect 22836 2932 22888 2941
rect 21088 2839 21140 2848
rect 21088 2805 21097 2839
rect 21097 2805 21131 2839
rect 21131 2805 21140 2839
rect 21548 2839 21600 2848
rect 21088 2796 21140 2805
rect 21548 2805 21557 2839
rect 21557 2805 21591 2839
rect 21591 2805 21600 2839
rect 21548 2796 21600 2805
rect 3749 2694 3801 2746
rect 3813 2694 3865 2746
rect 3877 2694 3929 2746
rect 3941 2694 3993 2746
rect 4005 2694 4057 2746
rect 9347 2694 9399 2746
rect 9411 2694 9463 2746
rect 9475 2694 9527 2746
rect 9539 2694 9591 2746
rect 9603 2694 9655 2746
rect 14945 2694 14997 2746
rect 15009 2694 15061 2746
rect 15073 2694 15125 2746
rect 15137 2694 15189 2746
rect 15201 2694 15253 2746
rect 20543 2694 20595 2746
rect 20607 2694 20659 2746
rect 20671 2694 20723 2746
rect 20735 2694 20787 2746
rect 20799 2694 20851 2746
rect 4804 2592 4856 2644
rect 5908 2524 5960 2576
rect 5816 2456 5868 2508
rect 7012 2592 7064 2644
rect 7104 2592 7156 2644
rect 7380 2592 7432 2644
rect 8208 2592 8260 2644
rect 9036 2592 9088 2644
rect 9956 2592 10008 2644
rect 10324 2592 10376 2644
rect 11152 2592 11204 2644
rect 13452 2592 13504 2644
rect 14188 2592 14240 2644
rect 17500 2592 17552 2644
rect 6368 2499 6420 2508
rect 6368 2465 6377 2499
rect 6377 2465 6411 2499
rect 6411 2465 6420 2499
rect 6368 2456 6420 2465
rect 8300 2456 8352 2508
rect 9864 2499 9916 2508
rect 1860 2431 1912 2440
rect 1860 2397 1869 2431
rect 1869 2397 1903 2431
rect 1903 2397 1912 2431
rect 1860 2388 1912 2397
rect 3608 2431 3660 2440
rect 2044 2295 2096 2304
rect 2044 2261 2053 2295
rect 2053 2261 2087 2295
rect 2087 2261 2096 2295
rect 2044 2252 2096 2261
rect 2228 2295 2280 2304
rect 2228 2261 2237 2295
rect 2237 2261 2271 2295
rect 2271 2261 2280 2295
rect 2228 2252 2280 2261
rect 3608 2397 3617 2431
rect 3617 2397 3651 2431
rect 3651 2397 3660 2431
rect 3608 2388 3660 2397
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5356 2431 5408 2440
rect 5356 2397 5365 2431
rect 5365 2397 5399 2431
rect 5399 2397 5408 2431
rect 5356 2388 5408 2397
rect 3792 2295 3844 2304
rect 3792 2261 3801 2295
rect 3801 2261 3835 2295
rect 3835 2261 3844 2295
rect 3792 2252 3844 2261
rect 3976 2295 4028 2304
rect 3976 2261 3985 2295
rect 3985 2261 4019 2295
rect 4019 2261 4028 2295
rect 3976 2252 4028 2261
rect 8208 2388 8260 2440
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 5816 2363 5868 2372
rect 5816 2329 5825 2363
rect 5825 2329 5859 2363
rect 5859 2329 5868 2363
rect 5816 2320 5868 2329
rect 6092 2320 6144 2372
rect 6828 2320 6880 2372
rect 8116 2320 8168 2372
rect 9864 2465 9873 2499
rect 9873 2465 9907 2499
rect 9907 2465 9916 2499
rect 9864 2456 9916 2465
rect 9956 2499 10008 2508
rect 9956 2465 9965 2499
rect 9965 2465 9999 2499
rect 9999 2465 10008 2499
rect 10232 2524 10284 2576
rect 11244 2524 11296 2576
rect 9956 2456 10008 2465
rect 9680 2388 9732 2440
rect 11704 2456 11756 2508
rect 9128 2363 9180 2372
rect 9128 2329 9137 2363
rect 9137 2329 9171 2363
rect 9171 2329 9180 2363
rect 9128 2320 9180 2329
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 11704 2320 11756 2372
rect 12072 2456 12124 2508
rect 14096 2524 14148 2576
rect 15292 2567 15344 2576
rect 15292 2533 15301 2567
rect 15301 2533 15335 2567
rect 15335 2533 15344 2567
rect 15292 2524 15344 2533
rect 15384 2524 15436 2576
rect 16396 2567 16448 2576
rect 16396 2533 16405 2567
rect 16405 2533 16439 2567
rect 16439 2533 16448 2567
rect 16396 2524 16448 2533
rect 12716 2388 12768 2440
rect 14280 2456 14332 2508
rect 14372 2456 14424 2508
rect 14004 2388 14056 2440
rect 16580 2456 16632 2508
rect 15476 2431 15528 2440
rect 15476 2397 15485 2431
rect 15485 2397 15519 2431
rect 15519 2397 15528 2431
rect 15476 2388 15528 2397
rect 16212 2431 16264 2440
rect 16212 2397 16221 2431
rect 16221 2397 16255 2431
rect 16255 2397 16264 2431
rect 16212 2388 16264 2397
rect 22836 2592 22888 2644
rect 20720 2567 20772 2576
rect 20720 2533 20729 2567
rect 20729 2533 20763 2567
rect 20763 2533 20772 2567
rect 20720 2524 20772 2533
rect 20904 2524 20956 2576
rect 22376 2524 22428 2576
rect 22744 2567 22796 2576
rect 22744 2533 22753 2567
rect 22753 2533 22787 2567
rect 22787 2533 22796 2567
rect 22744 2524 22796 2533
rect 19340 2499 19392 2508
rect 19340 2465 19349 2499
rect 19349 2465 19383 2499
rect 19383 2465 19392 2499
rect 19340 2456 19392 2465
rect 20352 2456 20404 2508
rect 18236 2431 18288 2440
rect 18236 2397 18245 2431
rect 18245 2397 18279 2431
rect 18279 2397 18288 2431
rect 18236 2388 18288 2397
rect 18972 2388 19024 2440
rect 20444 2388 20496 2440
rect 22008 2456 22060 2508
rect 21916 2388 21968 2440
rect 23112 2431 23164 2440
rect 23112 2397 23121 2431
rect 23121 2397 23155 2431
rect 23155 2397 23164 2431
rect 23112 2388 23164 2397
rect 12900 2252 12952 2304
rect 17040 2363 17092 2372
rect 17040 2329 17074 2363
rect 17074 2329 17092 2363
rect 17040 2320 17092 2329
rect 18236 2252 18288 2304
rect 18880 2295 18932 2304
rect 18880 2261 18889 2295
rect 18889 2261 18923 2295
rect 18923 2261 18932 2295
rect 18880 2252 18932 2261
rect 18972 2295 19024 2304
rect 18972 2261 18981 2295
rect 18981 2261 19015 2295
rect 19015 2261 19024 2295
rect 19340 2320 19392 2372
rect 20812 2320 20864 2372
rect 18972 2252 19024 2261
rect 21640 2252 21692 2304
rect 21824 2252 21876 2304
rect 6548 2150 6600 2202
rect 6612 2150 6664 2202
rect 6676 2150 6728 2202
rect 6740 2150 6792 2202
rect 6804 2150 6856 2202
rect 12146 2150 12198 2202
rect 12210 2150 12262 2202
rect 12274 2150 12326 2202
rect 12338 2150 12390 2202
rect 12402 2150 12454 2202
rect 17744 2150 17796 2202
rect 17808 2150 17860 2202
rect 17872 2150 17924 2202
rect 17936 2150 17988 2202
rect 18000 2150 18052 2202
rect 3792 2048 3844 2100
rect 9312 2048 9364 2100
rect 2228 1980 2280 2032
rect 4620 1912 4672 1964
rect 7932 1912 7984 1964
rect 8208 1980 8260 2032
rect 17040 1980 17092 2032
rect 17500 2048 17552 2100
rect 22468 2048 22520 2100
rect 20720 1980 20772 2032
rect 14832 1912 14884 1964
rect 16396 1912 16448 1964
rect 20260 1912 20312 1964
rect 3608 1844 3660 1896
rect 7380 1844 7432 1896
rect 16304 1844 16356 1896
rect 18880 1844 18932 1896
rect 3424 1776 3476 1828
rect 9128 1776 9180 1828
rect 15292 1776 15344 1828
rect 20168 1776 20220 1828
rect 7932 1572 7984 1624
rect 18236 1708 18288 1760
<< metal2 >>
rect 294 23800 350 24600
rect 938 23800 994 24600
rect 1582 23800 1638 24600
rect 2226 23800 2282 24600
rect 2870 23800 2926 24600
rect 3514 23800 3570 24600
rect 4158 23800 4214 24600
rect 4802 23800 4858 24600
rect 5446 23800 5502 24600
rect 6090 23800 6146 24600
rect 6734 23800 6790 24600
rect 7378 23800 7434 24600
rect 8022 23800 8078 24600
rect 8666 23800 8722 24600
rect 9048 23854 9260 23882
rect 308 21894 336 23800
rect 296 21888 348 21894
rect 296 21830 348 21836
rect 952 21690 980 23800
rect 1596 21894 1624 23800
rect 1952 22092 2004 22098
rect 1952 22034 2004 22040
rect 1860 22024 1912 22030
rect 1860 21966 1912 21972
rect 1584 21888 1636 21894
rect 1584 21830 1636 21836
rect 940 21684 992 21690
rect 940 21626 992 21632
rect 1768 21548 1820 21554
rect 1768 21490 1820 21496
rect 1780 21010 1808 21490
rect 1768 21004 1820 21010
rect 1768 20946 1820 20952
rect 1780 20602 1808 20946
rect 1768 20596 1820 20602
rect 1768 20538 1820 20544
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 1492 19508 1544 19514
rect 1492 19450 1544 19456
rect 1308 18828 1360 18834
rect 1308 18770 1360 18776
rect 1320 18154 1348 18770
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1308 18148 1360 18154
rect 1308 18090 1360 18096
rect 1412 17338 1440 18702
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1504 16574 1532 19450
rect 1596 19378 1624 19790
rect 1584 19372 1636 19378
rect 1584 19314 1636 19320
rect 1596 18358 1624 19314
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 1688 18426 1716 18906
rect 1768 18896 1820 18902
rect 1768 18838 1820 18844
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 1584 18352 1636 18358
rect 1584 18294 1636 18300
rect 1596 17746 1624 18294
rect 1780 18290 1808 18838
rect 1768 18284 1820 18290
rect 1768 18226 1820 18232
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1596 17270 1624 17682
rect 1584 17264 1636 17270
rect 1584 17206 1636 17212
rect 1504 16546 1716 16574
rect 1492 16040 1544 16046
rect 1492 15982 1544 15988
rect 1504 15570 1532 15982
rect 1492 15564 1544 15570
rect 1492 15506 1544 15512
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1412 15162 1440 15438
rect 1582 15328 1638 15337
rect 1582 15263 1638 15272
rect 1400 15156 1452 15162
rect 1400 15098 1452 15104
rect 1596 14618 1624 15263
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1584 14408 1636 14414
rect 1584 14350 1636 14356
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 11898 1440 13262
rect 1400 11892 1452 11898
rect 1400 11834 1452 11840
rect 1400 9580 1452 9586
rect 1400 9522 1452 9528
rect 1412 9217 1440 9522
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 1504 8974 1532 9318
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1596 7546 1624 14350
rect 1688 13802 1716 16546
rect 1872 16522 1900 21966
rect 1860 16516 1912 16522
rect 1860 16458 1912 16464
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1780 15434 1808 16390
rect 1768 15428 1820 15434
rect 1768 15370 1820 15376
rect 1964 14618 1992 22034
rect 2044 21956 2096 21962
rect 2044 21898 2096 21904
rect 2056 18714 2084 21898
rect 2240 21894 2268 23800
rect 2884 22094 2912 23800
rect 2884 22066 3004 22094
rect 2976 21894 3004 22066
rect 3056 22024 3108 22030
rect 3056 21966 3108 21972
rect 3332 22024 3384 22030
rect 3332 21966 3384 21972
rect 2228 21888 2280 21894
rect 2228 21830 2280 21836
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 2964 21888 3016 21894
rect 2964 21830 3016 21836
rect 2884 21690 2912 21830
rect 2872 21684 2924 21690
rect 2872 21626 2924 21632
rect 2504 21616 2556 21622
rect 2504 21558 2556 21564
rect 2320 21344 2372 21350
rect 2320 21286 2372 21292
rect 2332 20942 2360 21286
rect 2228 20936 2280 20942
rect 2228 20878 2280 20884
rect 2320 20936 2372 20942
rect 2320 20878 2372 20884
rect 2136 20800 2188 20806
rect 2136 20742 2188 20748
rect 2148 20534 2176 20742
rect 2240 20602 2268 20878
rect 2228 20596 2280 20602
rect 2228 20538 2280 20544
rect 2136 20528 2188 20534
rect 2136 20470 2188 20476
rect 2240 19854 2268 20538
rect 2228 19848 2280 19854
rect 2228 19790 2280 19796
rect 2056 18686 2176 18714
rect 2044 18624 2096 18630
rect 2044 18566 2096 18572
rect 2056 17678 2084 18566
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 2044 16108 2096 16114
rect 2044 16050 2096 16056
rect 2056 15706 2084 16050
rect 2044 15700 2096 15706
rect 2044 15642 2096 15648
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 2056 15026 2084 15506
rect 2044 15020 2096 15026
rect 2044 14962 2096 14968
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2148 14550 2176 18686
rect 2228 18624 2280 18630
rect 2228 18566 2280 18572
rect 2320 18624 2372 18630
rect 2320 18566 2372 18572
rect 2240 18426 2268 18566
rect 2228 18420 2280 18426
rect 2228 18362 2280 18368
rect 2332 18290 2360 18566
rect 2320 18284 2372 18290
rect 2320 18226 2372 18232
rect 2516 17882 2544 21558
rect 2964 21548 3016 21554
rect 2964 21490 3016 21496
rect 2596 21480 2648 21486
rect 2596 21422 2648 21428
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2608 21146 2636 21422
rect 2688 21412 2740 21418
rect 2688 21354 2740 21360
rect 2596 21140 2648 21146
rect 2596 21082 2648 21088
rect 2608 20874 2636 21082
rect 2596 20868 2648 20874
rect 2596 20810 2648 20816
rect 2596 20460 2648 20466
rect 2596 20402 2648 20408
rect 2608 19990 2636 20402
rect 2596 19984 2648 19990
rect 2596 19926 2648 19932
rect 2504 17876 2556 17882
rect 2504 17818 2556 17824
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 2608 16998 2636 17138
rect 2596 16992 2648 16998
rect 2596 16934 2648 16940
rect 2320 16448 2372 16454
rect 2320 16390 2372 16396
rect 2332 15706 2360 16390
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 2412 14816 2464 14822
rect 2412 14758 2464 14764
rect 2424 14618 2452 14758
rect 2700 14618 2728 21354
rect 2792 19854 2820 21422
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 2884 20058 2912 20402
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2780 19848 2832 19854
rect 2976 19802 3004 21490
rect 2780 19790 2832 19796
rect 2792 19514 2820 19790
rect 2884 19774 3004 19802
rect 2884 19718 2912 19774
rect 2872 19712 2924 19718
rect 2872 19654 2924 19660
rect 2780 19508 2832 19514
rect 2780 19450 2832 19456
rect 2964 17808 3016 17814
rect 2964 17750 3016 17756
rect 2872 16584 2924 16590
rect 2872 16526 2924 16532
rect 2884 16250 2912 16526
rect 2976 16522 3004 17750
rect 2964 16516 3016 16522
rect 2964 16458 3016 16464
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2872 15972 2924 15978
rect 2872 15914 2924 15920
rect 2884 15026 2912 15914
rect 3068 15706 3096 21966
rect 3240 21344 3292 21350
rect 3240 21286 3292 21292
rect 3252 20602 3280 21286
rect 3240 20596 3292 20602
rect 3240 20538 3292 20544
rect 3148 20256 3200 20262
rect 3148 20198 3200 20204
rect 3240 20256 3292 20262
rect 3240 20198 3292 20204
rect 3160 19922 3188 20198
rect 3148 19916 3200 19922
rect 3148 19858 3200 19864
rect 3148 19236 3200 19242
rect 3148 19178 3200 19184
rect 3160 17610 3188 19178
rect 3252 18086 3280 20198
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3148 17604 3200 17610
rect 3148 17546 3200 17552
rect 3148 17128 3200 17134
rect 3148 17070 3200 17076
rect 3160 16658 3188 17070
rect 3148 16652 3200 16658
rect 3148 16594 3200 16600
rect 3160 16114 3188 16594
rect 3344 16454 3372 21966
rect 3528 21894 3556 23800
rect 3749 22332 4057 22352
rect 3749 22330 3755 22332
rect 3811 22330 3835 22332
rect 3891 22330 3915 22332
rect 3971 22330 3995 22332
rect 4051 22330 4057 22332
rect 3811 22278 3813 22330
rect 3993 22278 3995 22330
rect 3749 22276 3755 22278
rect 3811 22276 3835 22278
rect 3891 22276 3915 22278
rect 3971 22276 3995 22278
rect 4051 22276 4057 22278
rect 3749 22256 4057 22276
rect 4068 22024 4120 22030
rect 4068 21966 4120 21972
rect 3516 21888 3568 21894
rect 3516 21830 3568 21836
rect 4080 21622 4108 21966
rect 4172 21894 4200 23800
rect 4816 22094 4844 23800
rect 4724 22066 4844 22094
rect 4988 22092 5040 22098
rect 4528 22024 4580 22030
rect 4528 21966 4580 21972
rect 4160 21888 4212 21894
rect 4160 21830 4212 21836
rect 4252 21684 4304 21690
rect 4252 21626 4304 21632
rect 4068 21616 4120 21622
rect 4068 21558 4120 21564
rect 3424 21480 3476 21486
rect 3424 21422 3476 21428
rect 3436 20534 3464 21422
rect 3749 21244 4057 21264
rect 3749 21242 3755 21244
rect 3811 21242 3835 21244
rect 3891 21242 3915 21244
rect 3971 21242 3995 21244
rect 4051 21242 4057 21244
rect 3811 21190 3813 21242
rect 3993 21190 3995 21242
rect 3749 21188 3755 21190
rect 3811 21188 3835 21190
rect 3891 21188 3915 21190
rect 3971 21188 3995 21190
rect 4051 21188 4057 21190
rect 3749 21168 4057 21188
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 4068 20936 4120 20942
rect 4068 20878 4120 20884
rect 3424 20528 3476 20534
rect 3424 20470 3476 20476
rect 3422 19272 3478 19281
rect 3422 19207 3424 19216
rect 3476 19207 3478 19216
rect 3424 19178 3476 19184
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3528 18834 3556 19110
rect 3620 18850 3648 20878
rect 3700 20800 3752 20806
rect 3700 20742 3752 20748
rect 3712 20466 3740 20742
rect 4080 20602 4108 20878
rect 4068 20596 4120 20602
rect 4068 20538 4120 20544
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 4160 20256 4212 20262
rect 4160 20198 4212 20204
rect 3749 20156 4057 20176
rect 3749 20154 3755 20156
rect 3811 20154 3835 20156
rect 3891 20154 3915 20156
rect 3971 20154 3995 20156
rect 4051 20154 4057 20156
rect 3811 20102 3813 20154
rect 3993 20102 3995 20154
rect 3749 20100 3755 20102
rect 3811 20100 3835 20102
rect 3891 20100 3915 20102
rect 3971 20100 3995 20102
rect 4051 20100 4057 20102
rect 3749 20080 4057 20100
rect 4172 19446 4200 20198
rect 4160 19440 4212 19446
rect 4160 19382 4212 19388
rect 4160 19304 4212 19310
rect 4160 19246 4212 19252
rect 3749 19068 4057 19088
rect 3749 19066 3755 19068
rect 3811 19066 3835 19068
rect 3891 19066 3915 19068
rect 3971 19066 3995 19068
rect 4051 19066 4057 19068
rect 3811 19014 3813 19066
rect 3993 19014 3995 19066
rect 3749 19012 3755 19014
rect 3811 19012 3835 19014
rect 3891 19012 3915 19014
rect 3971 19012 3995 19014
rect 4051 19012 4057 19014
rect 3749 18992 4057 19012
rect 4172 18902 4200 19246
rect 4264 19242 4292 21626
rect 4436 21480 4488 21486
rect 4436 21422 4488 21428
rect 4448 20398 4476 21422
rect 4436 20392 4488 20398
rect 4436 20334 4488 20340
rect 4344 19440 4396 19446
rect 4344 19382 4396 19388
rect 4252 19236 4304 19242
rect 4252 19178 4304 19184
rect 4160 18896 4212 18902
rect 3516 18828 3568 18834
rect 3620 18822 3740 18850
rect 4160 18838 4212 18844
rect 3516 18770 3568 18776
rect 3608 18760 3660 18766
rect 3608 18702 3660 18708
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3436 17678 3464 18566
rect 3620 17882 3648 18702
rect 3712 18193 3740 18822
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 3698 18184 3754 18193
rect 3698 18119 3754 18128
rect 3749 17980 4057 18000
rect 3749 17978 3755 17980
rect 3811 17978 3835 17980
rect 3891 17978 3915 17980
rect 3971 17978 3995 17980
rect 4051 17978 4057 17980
rect 3811 17926 3813 17978
rect 3993 17926 3995 17978
rect 3749 17924 3755 17926
rect 3811 17924 3835 17926
rect 3891 17924 3915 17926
rect 3971 17924 3995 17926
rect 4051 17924 4057 17926
rect 3749 17904 4057 17924
rect 3608 17876 3660 17882
rect 3528 17836 3608 17864
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3528 17338 3556 17836
rect 3608 17818 3660 17824
rect 3882 17776 3938 17785
rect 3882 17711 3938 17720
rect 3608 17672 3660 17678
rect 3608 17614 3660 17620
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3620 16794 3648 17614
rect 3896 17134 3924 17711
rect 4172 17338 4200 18566
rect 4160 17332 4212 17338
rect 4160 17274 4212 17280
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 4264 17066 4292 18566
rect 4356 17610 4384 19382
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4448 18970 4476 19314
rect 4540 19174 4568 21966
rect 4724 21894 4752 22066
rect 4988 22034 5040 22040
rect 4712 21888 4764 21894
rect 4712 21830 4764 21836
rect 4804 21888 4856 21894
rect 4804 21830 4856 21836
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 4724 20534 4752 21490
rect 4816 20874 4844 21830
rect 5000 21622 5028 22034
rect 5172 22024 5224 22030
rect 5172 21966 5224 21972
rect 5184 21622 5212 21966
rect 4988 21616 5040 21622
rect 4988 21558 5040 21564
rect 5172 21616 5224 21622
rect 5172 21558 5224 21564
rect 5080 21344 5132 21350
rect 5080 21286 5132 21292
rect 4804 20868 4856 20874
rect 4804 20810 4856 20816
rect 4712 20528 4764 20534
rect 4712 20470 4764 20476
rect 5092 20466 5120 21286
rect 5356 21072 5408 21078
rect 5276 21032 5356 21060
rect 5080 20460 5132 20466
rect 5080 20402 5132 20408
rect 4712 20392 4764 20398
rect 4712 20334 4764 20340
rect 4620 20052 4672 20058
rect 4620 19994 4672 20000
rect 4632 19854 4660 19994
rect 4620 19848 4672 19854
rect 4620 19790 4672 19796
rect 4724 19394 4752 20334
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 4896 19984 4948 19990
rect 4896 19926 4948 19932
rect 4804 19848 4856 19854
rect 4804 19790 4856 19796
rect 4632 19366 4752 19394
rect 4528 19168 4580 19174
rect 4528 19110 4580 19116
rect 4436 18964 4488 18970
rect 4436 18906 4488 18912
rect 4632 18834 4660 19366
rect 4816 19310 4844 19790
rect 4908 19514 4936 19926
rect 4896 19508 4948 19514
rect 4896 19450 4948 19456
rect 4712 19304 4764 19310
rect 4712 19246 4764 19252
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4620 18828 4672 18834
rect 4620 18770 4672 18776
rect 4436 18692 4488 18698
rect 4436 18634 4488 18640
rect 4448 18086 4476 18634
rect 4632 18222 4660 18770
rect 4724 18426 4752 19246
rect 4816 18970 4844 19246
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4712 18420 4764 18426
rect 4712 18362 4764 18368
rect 4620 18216 4672 18222
rect 4620 18158 4672 18164
rect 4528 18148 4580 18154
rect 4528 18090 4580 18096
rect 4436 18080 4488 18086
rect 4436 18022 4488 18028
rect 4344 17604 4396 17610
rect 4344 17546 4396 17552
rect 4448 17134 4476 18022
rect 4540 17814 4568 18090
rect 4528 17808 4580 17814
rect 4528 17750 4580 17756
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4252 17060 4304 17066
rect 4252 17002 4304 17008
rect 3749 16892 4057 16912
rect 3749 16890 3755 16892
rect 3811 16890 3835 16892
rect 3891 16890 3915 16892
rect 3971 16890 3995 16892
rect 4051 16890 4057 16892
rect 3811 16838 3813 16890
rect 3993 16838 3995 16890
rect 3749 16836 3755 16838
rect 3811 16836 3835 16838
rect 3891 16836 3915 16838
rect 3971 16836 3995 16838
rect 4051 16836 4057 16838
rect 3749 16816 4057 16836
rect 3608 16788 3660 16794
rect 4540 16776 4568 17614
rect 3608 16730 3660 16736
rect 4448 16748 4568 16776
rect 3332 16448 3384 16454
rect 3332 16390 3384 16396
rect 3700 16448 3752 16454
rect 3700 16390 3752 16396
rect 3712 16250 3740 16390
rect 3700 16244 3752 16250
rect 3700 16186 3752 16192
rect 4252 16176 4304 16182
rect 4252 16118 4304 16124
rect 3148 16108 3200 16114
rect 3148 16050 3200 16056
rect 3240 16040 3292 16046
rect 3240 15982 3292 15988
rect 3252 15706 3280 15982
rect 3749 15804 4057 15824
rect 3749 15802 3755 15804
rect 3811 15802 3835 15804
rect 3891 15802 3915 15804
rect 3971 15802 3995 15804
rect 4051 15802 4057 15804
rect 3811 15750 3813 15802
rect 3993 15750 3995 15802
rect 3749 15748 3755 15750
rect 3811 15748 3835 15750
rect 3891 15748 3915 15750
rect 3971 15748 3995 15750
rect 4051 15748 4057 15750
rect 3749 15728 4057 15748
rect 3056 15700 3108 15706
rect 3056 15642 3108 15648
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 2412 14612 2464 14618
rect 2412 14554 2464 14560
rect 2688 14612 2740 14618
rect 2688 14554 2740 14560
rect 2136 14544 2188 14550
rect 2136 14486 2188 14492
rect 1952 14408 2004 14414
rect 1952 14350 2004 14356
rect 1964 14074 1992 14350
rect 1952 14068 2004 14074
rect 1952 14010 2004 14016
rect 2884 14006 2912 14962
rect 2976 14618 3004 14962
rect 2964 14612 3016 14618
rect 2964 14554 3016 14560
rect 3252 14414 3280 15642
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 4264 15450 4292 16118
rect 4344 15496 4396 15502
rect 4264 15444 4344 15450
rect 4264 15438 4396 15444
rect 4172 15042 4200 15438
rect 4264 15422 4384 15438
rect 4264 15162 4292 15422
rect 4252 15156 4304 15162
rect 4252 15098 4304 15104
rect 4448 15094 4476 16748
rect 4632 16674 4660 18158
rect 4724 17202 4752 18362
rect 4804 17604 4856 17610
rect 4804 17546 4856 17552
rect 4816 17270 4844 17546
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4712 17196 4764 17202
rect 4712 17138 4764 17144
rect 4816 16794 4844 17206
rect 4804 16788 4856 16794
rect 4804 16730 4856 16736
rect 4540 16658 4660 16674
rect 4528 16652 4660 16658
rect 4580 16646 4660 16652
rect 4528 16594 4580 16600
rect 4908 15706 4936 17478
rect 5000 17338 5028 20198
rect 5080 19984 5132 19990
rect 5080 19926 5132 19932
rect 5092 19786 5120 19926
rect 5276 19922 5304 21032
rect 5356 21014 5408 21020
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 5080 19780 5132 19786
rect 5080 19722 5132 19728
rect 5264 18624 5316 18630
rect 5264 18566 5316 18572
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5276 17882 5304 18566
rect 5264 17876 5316 17882
rect 5264 17818 5316 17824
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 5368 16590 5396 18566
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5172 16108 5224 16114
rect 5172 16050 5224 16056
rect 5184 15706 5212 16050
rect 5460 16046 5488 23800
rect 6000 22976 6052 22982
rect 6000 22918 6052 22924
rect 5540 21888 5592 21894
rect 5540 21830 5592 21836
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 5552 21622 5580 21830
rect 5644 21690 5672 21830
rect 5632 21684 5684 21690
rect 5632 21626 5684 21632
rect 5540 21616 5592 21622
rect 5540 21558 5592 21564
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5736 21078 5764 21490
rect 5724 21072 5776 21078
rect 5724 21014 5776 21020
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 5540 20800 5592 20806
rect 5540 20742 5592 20748
rect 5552 19990 5580 20742
rect 5920 20602 5948 20878
rect 5908 20596 5960 20602
rect 5908 20538 5960 20544
rect 5540 19984 5592 19990
rect 5540 19926 5592 19932
rect 5920 19922 5948 20538
rect 6012 20262 6040 22918
rect 6104 22094 6132 23800
rect 6748 22982 6776 23800
rect 6736 22976 6788 22982
rect 6736 22918 6788 22924
rect 7392 22094 7420 23800
rect 6104 22066 6224 22094
rect 7392 22066 7604 22094
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 5908 19916 5960 19922
rect 5908 19858 5960 19864
rect 6196 19854 6224 22066
rect 6460 22024 6512 22030
rect 6460 21966 6512 21972
rect 7380 22024 7432 22030
rect 7380 21966 7432 21972
rect 6368 21956 6420 21962
rect 6368 21898 6420 21904
rect 6380 21690 6408 21898
rect 6368 21684 6420 21690
rect 6368 21626 6420 21632
rect 6472 21486 6500 21966
rect 6736 21956 6788 21962
rect 6788 21916 6960 21944
rect 6736 21898 6788 21904
rect 6548 21788 6856 21808
rect 6548 21786 6554 21788
rect 6610 21786 6634 21788
rect 6690 21786 6714 21788
rect 6770 21786 6794 21788
rect 6850 21786 6856 21788
rect 6610 21734 6612 21786
rect 6792 21734 6794 21786
rect 6548 21732 6554 21734
rect 6610 21732 6634 21734
rect 6690 21732 6714 21734
rect 6770 21732 6794 21734
rect 6850 21732 6856 21734
rect 6548 21712 6856 21732
rect 6932 21690 6960 21916
rect 6920 21684 6972 21690
rect 6920 21626 6972 21632
rect 7392 21554 7420 21966
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 6460 21480 6512 21486
rect 6460 21422 6512 21428
rect 7196 21480 7248 21486
rect 7196 21422 7248 21428
rect 7104 21344 7156 21350
rect 7104 21286 7156 21292
rect 7116 21010 7144 21286
rect 7104 21004 7156 21010
rect 7104 20946 7156 20952
rect 6460 20800 6512 20806
rect 6460 20742 6512 20748
rect 7104 20800 7156 20806
rect 7104 20742 7156 20748
rect 6472 20534 6500 20742
rect 6548 20700 6856 20720
rect 6548 20698 6554 20700
rect 6610 20698 6634 20700
rect 6690 20698 6714 20700
rect 6770 20698 6794 20700
rect 6850 20698 6856 20700
rect 6610 20646 6612 20698
rect 6792 20646 6794 20698
rect 6548 20644 6554 20646
rect 6610 20644 6634 20646
rect 6690 20644 6714 20646
rect 6770 20644 6794 20646
rect 6850 20644 6856 20646
rect 6548 20624 6856 20644
rect 6460 20528 6512 20534
rect 6460 20470 6512 20476
rect 7012 20052 7064 20058
rect 7012 19994 7064 20000
rect 6184 19848 6236 19854
rect 6184 19790 6236 19796
rect 5816 19712 5868 19718
rect 5816 19654 5868 19660
rect 6368 19712 6420 19718
rect 6368 19654 6420 19660
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 5828 19258 5856 19654
rect 6380 19514 6408 19654
rect 6548 19612 6856 19632
rect 6548 19610 6554 19612
rect 6610 19610 6634 19612
rect 6690 19610 6714 19612
rect 6770 19610 6794 19612
rect 6850 19610 6856 19612
rect 6610 19558 6612 19610
rect 6792 19558 6794 19610
rect 6548 19556 6554 19558
rect 6610 19556 6634 19558
rect 6690 19556 6714 19558
rect 6770 19556 6794 19558
rect 6850 19556 6856 19558
rect 6548 19536 6856 19556
rect 6368 19508 6420 19514
rect 6368 19450 6420 19456
rect 6000 19372 6052 19378
rect 6000 19314 6052 19320
rect 5828 19230 5948 19258
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5828 18766 5856 19110
rect 5816 18760 5868 18766
rect 5816 18702 5868 18708
rect 5724 18624 5776 18630
rect 5724 18566 5776 18572
rect 5632 17196 5684 17202
rect 5632 17138 5684 17144
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 4896 15700 4948 15706
rect 4896 15642 4948 15648
rect 5172 15700 5224 15706
rect 5172 15642 5224 15648
rect 5460 15502 5488 15982
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 4896 15360 4948 15366
rect 4896 15302 4948 15308
rect 4436 15088 4488 15094
rect 4172 15014 4292 15042
rect 4436 15030 4488 15036
rect 4264 14890 4292 15014
rect 4252 14884 4304 14890
rect 4252 14826 4304 14832
rect 3749 14716 4057 14736
rect 3749 14714 3755 14716
rect 3811 14714 3835 14716
rect 3891 14714 3915 14716
rect 3971 14714 3995 14716
rect 4051 14714 4057 14716
rect 3811 14662 3813 14714
rect 3993 14662 3995 14714
rect 3749 14660 3755 14662
rect 3811 14660 3835 14662
rect 3891 14660 3915 14662
rect 3971 14660 3995 14662
rect 4051 14660 4057 14662
rect 3749 14640 4057 14660
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 4160 14408 4212 14414
rect 4160 14350 4212 14356
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 1676 13796 1728 13802
rect 1676 13738 1728 13744
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 13258 1992 13670
rect 2516 13530 2544 13874
rect 2884 13870 2912 13942
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2504 13524 2556 13530
rect 2504 13466 2556 13472
rect 2044 13320 2096 13326
rect 2044 13262 2096 13268
rect 1952 13252 2004 13258
rect 1952 13194 2004 13200
rect 2056 12306 2084 13262
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2044 12300 2096 12306
rect 2044 12242 2096 12248
rect 2148 12238 2176 13126
rect 2516 12986 2544 13466
rect 2884 13326 2912 13806
rect 2872 13320 2924 13326
rect 2872 13262 2924 13268
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2884 12918 2912 13262
rect 3528 12986 3556 13874
rect 3749 13628 4057 13648
rect 3749 13626 3755 13628
rect 3811 13626 3835 13628
rect 3891 13626 3915 13628
rect 3971 13626 3995 13628
rect 4051 13626 4057 13628
rect 3811 13574 3813 13626
rect 3993 13574 3995 13626
rect 3749 13572 3755 13574
rect 3811 13572 3835 13574
rect 3891 13572 3915 13574
rect 3971 13572 3995 13574
rect 4051 13572 4057 13574
rect 3749 13552 4057 13572
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3516 12980 3568 12986
rect 3516 12922 3568 12928
rect 2872 12912 2924 12918
rect 2872 12854 2924 12860
rect 3896 12850 3924 13330
rect 4172 13326 4200 14350
rect 4264 13938 4292 14826
rect 4620 14816 4672 14822
rect 4620 14758 4672 14764
rect 4632 14482 4660 14758
rect 4620 14476 4672 14482
rect 4620 14418 4672 14424
rect 4908 13938 4936 15302
rect 5448 15156 5500 15162
rect 5448 15098 5500 15104
rect 4988 15088 5040 15094
rect 4988 15030 5040 15036
rect 5172 15088 5224 15094
rect 5172 15030 5224 15036
rect 5000 14482 5028 15030
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 5000 14006 5028 14418
rect 5184 14074 5212 15030
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 4988 14000 5040 14006
rect 4988 13942 5040 13948
rect 4252 13932 4304 13938
rect 4252 13874 4304 13880
rect 4896 13932 4948 13938
rect 4896 13874 4948 13880
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5092 13462 5120 13874
rect 5460 13870 5488 15098
rect 5448 13864 5500 13870
rect 5448 13806 5500 13812
rect 5080 13456 5132 13462
rect 5080 13398 5132 13404
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4264 12866 4292 13262
rect 4988 13184 5040 13190
rect 4988 13126 5040 13132
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 4172 12838 4292 12866
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 3160 12442 3188 12786
rect 3749 12540 4057 12560
rect 3749 12538 3755 12540
rect 3811 12538 3835 12540
rect 3891 12538 3915 12540
rect 3971 12538 3995 12540
rect 4051 12538 4057 12540
rect 3811 12486 3813 12538
rect 3993 12486 3995 12538
rect 3749 12484 3755 12486
rect 3811 12484 3835 12486
rect 3891 12484 3915 12486
rect 3971 12484 3995 12486
rect 4051 12484 4057 12486
rect 3749 12464 4057 12484
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 2136 12232 2188 12238
rect 2136 12174 2188 12180
rect 3700 12164 3752 12170
rect 3700 12106 3752 12112
rect 3712 11898 3740 12106
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3712 11642 3740 11834
rect 3528 11614 3740 11642
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10606 1808 11086
rect 3148 11076 3200 11082
rect 3148 11018 3200 11024
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1768 10600 1820 10606
rect 1768 10542 1820 10548
rect 1780 10266 1808 10542
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1780 9178 1808 10202
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 1780 8498 1808 9114
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1780 7954 1808 8434
rect 1768 7948 1820 7954
rect 1768 7890 1820 7896
rect 1584 7540 1636 7546
rect 1584 7482 1636 7488
rect 1676 7472 1728 7478
rect 1676 7414 1728 7420
rect 1688 7002 1716 7414
rect 1768 7200 1820 7206
rect 1768 7142 1820 7148
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1780 6322 1808 7142
rect 1872 6866 1900 10610
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2136 7880 2188 7886
rect 2136 7822 2188 7828
rect 2148 7546 2176 7822
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 1860 6860 1912 6866
rect 1860 6802 1912 6808
rect 2332 6458 2360 8434
rect 2516 7886 2544 9318
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2608 6798 2636 9862
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2884 9042 2912 9454
rect 3160 9110 3188 11018
rect 3252 9654 3280 11494
rect 3528 11354 3556 11614
rect 3749 11452 4057 11472
rect 3749 11450 3755 11452
rect 3811 11450 3835 11452
rect 3891 11450 3915 11452
rect 3971 11450 3995 11452
rect 4051 11450 4057 11452
rect 3811 11398 3813 11450
rect 3993 11398 3995 11450
rect 3749 11396 3755 11398
rect 3811 11396 3835 11398
rect 3891 11396 3915 11398
rect 3971 11396 3995 11398
rect 4051 11396 4057 11398
rect 3749 11376 4057 11396
rect 4172 11354 4200 12838
rect 4252 12776 4304 12782
rect 4252 12718 4304 12724
rect 4264 12102 4292 12718
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 4264 11762 4292 12038
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4356 11694 4384 12650
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4356 11558 4384 11630
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 3516 11348 3568 11354
rect 3516 11290 3568 11296
rect 4160 11348 4212 11354
rect 4160 11290 4212 11296
rect 4356 11234 4384 11494
rect 4264 11206 4384 11234
rect 4448 11218 4476 12582
rect 4632 12306 4660 12854
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4896 12232 4948 12238
rect 4896 12174 4948 12180
rect 4620 12164 4672 12170
rect 4620 12106 4672 12112
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4540 11642 4568 12038
rect 4632 11762 4660 12106
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4712 11688 4764 11694
rect 4540 11614 4660 11642
rect 4712 11630 4764 11636
rect 4804 11688 4856 11694
rect 4804 11630 4856 11636
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4436 11212 4488 11218
rect 3424 11144 3476 11150
rect 3424 11086 3476 11092
rect 3436 10810 3464 11086
rect 3516 11076 3568 11082
rect 3516 11018 3568 11024
rect 3424 10804 3476 10810
rect 3424 10746 3476 10752
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3240 9648 3292 9654
rect 3240 9590 3292 9596
rect 3332 9580 3384 9586
rect 3332 9522 3384 9528
rect 3148 9104 3200 9110
rect 3148 9046 3200 9052
rect 2872 9036 2924 9042
rect 2872 8978 2924 8984
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2792 8566 2820 8774
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2700 7206 2728 8434
rect 2780 7404 2832 7410
rect 2780 7346 2832 7352
rect 2688 7200 2740 7206
rect 2688 7142 2740 7148
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2792 6458 2820 7346
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 3068 6866 3096 7278
rect 3252 6914 3280 8502
rect 3344 8362 3372 9522
rect 3436 9178 3464 9998
rect 3528 9450 3556 11018
rect 4160 10532 4212 10538
rect 4160 10474 4212 10480
rect 3749 10364 4057 10384
rect 3749 10362 3755 10364
rect 3811 10362 3835 10364
rect 3891 10362 3915 10364
rect 3971 10362 3995 10364
rect 4051 10362 4057 10364
rect 3811 10310 3813 10362
rect 3993 10310 3995 10362
rect 3749 10308 3755 10310
rect 3811 10308 3835 10310
rect 3891 10308 3915 10310
rect 3971 10308 3995 10310
rect 4051 10308 4057 10310
rect 3749 10288 4057 10308
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3896 10010 3924 10066
rect 3620 9982 3924 10010
rect 4172 9994 4200 10474
rect 4160 9988 4212 9994
rect 3620 9926 3648 9982
rect 4160 9930 4212 9936
rect 3608 9920 3660 9926
rect 3608 9862 3660 9868
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3804 9722 3832 9862
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3516 9444 3568 9450
rect 3516 9386 3568 9392
rect 3749 9276 4057 9296
rect 3749 9274 3755 9276
rect 3811 9274 3835 9276
rect 3891 9274 3915 9276
rect 3971 9274 3995 9276
rect 4051 9274 4057 9276
rect 3811 9222 3813 9274
rect 3993 9222 3995 9274
rect 3749 9220 3755 9222
rect 3811 9220 3835 9222
rect 3891 9220 3915 9222
rect 3971 9220 3995 9222
rect 4051 9220 4057 9222
rect 3749 9200 4057 9220
rect 3424 9172 3476 9178
rect 3424 9114 3476 9120
rect 4172 8974 4200 9930
rect 4264 9874 4292 11206
rect 4436 11154 4488 11160
rect 4540 11098 4568 11494
rect 4632 11150 4660 11614
rect 4724 11218 4752 11630
rect 4816 11286 4844 11630
rect 4804 11280 4856 11286
rect 4804 11222 4856 11228
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4356 11070 4568 11098
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4712 11076 4764 11082
rect 4356 9994 4384 11070
rect 4712 11018 4764 11024
rect 4528 11008 4580 11014
rect 4528 10950 4580 10956
rect 4436 10600 4488 10606
rect 4436 10542 4488 10548
rect 4448 10266 4476 10542
rect 4436 10260 4488 10266
rect 4436 10202 4488 10208
rect 4540 10198 4568 10950
rect 4620 10464 4672 10470
rect 4620 10406 4672 10412
rect 4528 10192 4580 10198
rect 4528 10134 4580 10140
rect 4436 10124 4488 10130
rect 4436 10066 4488 10072
rect 4344 9988 4396 9994
rect 4344 9930 4396 9936
rect 4448 9874 4476 10066
rect 4632 9994 4660 10406
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 4264 9846 4476 9874
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4540 9178 4568 9522
rect 4724 9450 4752 11018
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4816 9926 4844 10610
rect 4908 10606 4936 12174
rect 5000 11898 5028 13126
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5172 12096 5224 12102
rect 5172 12038 5224 12044
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 5184 11830 5212 12038
rect 5368 11898 5396 12786
rect 5552 12238 5580 16186
rect 5644 16114 5672 17138
rect 5736 16998 5764 18566
rect 5920 17270 5948 19230
rect 6012 18426 6040 19314
rect 6184 19168 6236 19174
rect 6184 19110 6236 19116
rect 6196 18970 6224 19110
rect 6184 18964 6236 18970
rect 6184 18906 6236 18912
rect 6184 18760 6236 18766
rect 6184 18702 6236 18708
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6092 18352 6144 18358
rect 6092 18294 6144 18300
rect 5908 17264 5960 17270
rect 5908 17206 5960 17212
rect 5724 16992 5776 16998
rect 5724 16934 5776 16940
rect 6104 16454 6132 18294
rect 6196 17218 6224 18702
rect 6276 18216 6328 18222
rect 6276 18158 6328 18164
rect 6288 17338 6316 18158
rect 6368 18080 6420 18086
rect 6368 18022 6420 18028
rect 6380 17610 6408 18022
rect 6472 17882 6500 18702
rect 6548 18524 6856 18544
rect 6548 18522 6554 18524
rect 6610 18522 6634 18524
rect 6690 18522 6714 18524
rect 6770 18522 6794 18524
rect 6850 18522 6856 18524
rect 6610 18470 6612 18522
rect 6792 18470 6794 18522
rect 6548 18468 6554 18470
rect 6610 18468 6634 18470
rect 6690 18468 6714 18470
rect 6770 18468 6794 18470
rect 6850 18468 6856 18470
rect 6548 18448 6856 18468
rect 6932 17882 6960 19654
rect 7024 19553 7052 19994
rect 7010 19544 7066 19553
rect 7010 19479 7066 19488
rect 7012 19440 7064 19446
rect 7010 19408 7012 19417
rect 7064 19408 7066 19417
rect 7010 19343 7066 19352
rect 7012 19304 7064 19310
rect 7012 19246 7064 19252
rect 7024 19174 7052 19246
rect 7012 19168 7064 19174
rect 7012 19110 7064 19116
rect 7116 18358 7144 20742
rect 7208 20058 7236 21422
rect 7392 20942 7420 21490
rect 7380 20936 7432 20942
rect 7380 20878 7432 20884
rect 7196 20052 7248 20058
rect 7196 19994 7248 20000
rect 7196 19916 7248 19922
rect 7196 19858 7248 19864
rect 7208 19446 7236 19858
rect 7288 19848 7340 19854
rect 7288 19790 7340 19796
rect 7196 19440 7248 19446
rect 7196 19382 7248 19388
rect 7300 19292 7328 19790
rect 7208 19264 7328 19292
rect 7208 18986 7236 19264
rect 7208 18958 7328 18986
rect 7196 18896 7248 18902
rect 7194 18864 7196 18873
rect 7248 18864 7250 18873
rect 7194 18799 7250 18808
rect 7196 18624 7248 18630
rect 7196 18566 7248 18572
rect 7104 18352 7156 18358
rect 7104 18294 7156 18300
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 6460 17876 6512 17882
rect 6460 17818 6512 17824
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6368 17604 6420 17610
rect 6368 17546 6420 17552
rect 6276 17332 6328 17338
rect 6276 17274 6328 17280
rect 6196 17190 6408 17218
rect 6380 17134 6408 17190
rect 6368 17128 6420 17134
rect 6368 17070 6420 17076
rect 6184 16788 6236 16794
rect 6184 16730 6236 16736
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 6196 16114 6224 16730
rect 6380 16182 6408 17070
rect 6472 16590 6500 17818
rect 6550 17776 6606 17785
rect 6550 17711 6606 17720
rect 6564 17678 6592 17711
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6548 17436 6856 17456
rect 6548 17434 6554 17436
rect 6610 17434 6634 17436
rect 6690 17434 6714 17436
rect 6770 17434 6794 17436
rect 6850 17434 6856 17436
rect 6610 17382 6612 17434
rect 6792 17382 6794 17434
rect 6548 17380 6554 17382
rect 6610 17380 6634 17382
rect 6690 17380 6714 17382
rect 6770 17380 6794 17382
rect 6850 17380 6856 17382
rect 6548 17360 6856 17380
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6656 16658 6684 17206
rect 6736 17196 6788 17202
rect 6736 17138 6788 17144
rect 6748 16794 6776 17138
rect 7024 17066 7052 18226
rect 7116 18222 7144 18253
rect 7104 18216 7156 18222
rect 7102 18184 7104 18193
rect 7156 18184 7158 18193
rect 7102 18119 7158 18128
rect 7116 17338 7144 18119
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7012 17060 7064 17066
rect 7012 17002 7064 17008
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6644 16652 6696 16658
rect 6644 16594 6696 16600
rect 6460 16584 6512 16590
rect 6460 16526 6512 16532
rect 6548 16348 6856 16368
rect 6548 16346 6554 16348
rect 6610 16346 6634 16348
rect 6690 16346 6714 16348
rect 6770 16346 6794 16348
rect 6850 16346 6856 16348
rect 6610 16294 6612 16346
rect 6792 16294 6794 16346
rect 6548 16292 6554 16294
rect 6610 16292 6634 16294
rect 6690 16292 6714 16294
rect 6770 16292 6794 16294
rect 6850 16292 6856 16294
rect 6548 16272 6856 16292
rect 6368 16176 6420 16182
rect 6368 16118 6420 16124
rect 5632 16108 5684 16114
rect 5632 16050 5684 16056
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 6460 16040 6512 16046
rect 6460 15982 6512 15988
rect 5632 15972 5684 15978
rect 5632 15914 5684 15920
rect 5644 15026 5672 15914
rect 6472 15570 6500 15982
rect 6932 15910 6960 16730
rect 7024 16726 7052 17002
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 6920 15904 6972 15910
rect 6920 15846 6972 15852
rect 7116 15570 7144 16390
rect 6460 15564 6512 15570
rect 6460 15506 6512 15512
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 5908 15360 5960 15366
rect 5908 15302 5960 15308
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 6368 15360 6420 15366
rect 6368 15302 6420 15308
rect 5632 15020 5684 15026
rect 5632 14962 5684 14968
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5632 14816 5684 14822
rect 5632 14758 5684 14764
rect 5644 14618 5672 14758
rect 5736 14618 5764 14962
rect 5632 14612 5684 14618
rect 5632 14554 5684 14560
rect 5724 14612 5776 14618
rect 5776 14572 5856 14600
rect 5724 14554 5776 14560
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5632 14340 5684 14346
rect 5632 14282 5684 14288
rect 5644 13530 5672 14282
rect 5736 14074 5764 14350
rect 5724 14068 5776 14074
rect 5724 14010 5776 14016
rect 5828 13938 5856 14572
rect 5816 13932 5868 13938
rect 5816 13874 5868 13880
rect 5816 13728 5868 13734
rect 5736 13688 5816 13716
rect 5632 13524 5684 13530
rect 5632 13466 5684 13472
rect 5736 12782 5764 13688
rect 5816 13670 5868 13676
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5828 12918 5856 13126
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 5724 12776 5776 12782
rect 5724 12718 5776 12724
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5920 12170 5948 15302
rect 6012 14278 6040 15302
rect 6000 14272 6052 14278
rect 6000 14214 6052 14220
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 6092 14000 6144 14006
rect 6092 13942 6144 13948
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 6012 12986 6040 13874
rect 6104 13326 6132 13942
rect 6288 13802 6316 14214
rect 6380 14074 6408 15302
rect 6472 14890 6500 15506
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6548 15260 6856 15280
rect 6548 15258 6554 15260
rect 6610 15258 6634 15260
rect 6690 15258 6714 15260
rect 6770 15258 6794 15260
rect 6850 15258 6856 15260
rect 6610 15206 6612 15258
rect 6792 15206 6794 15258
rect 6548 15204 6554 15206
rect 6610 15204 6634 15206
rect 6690 15204 6714 15206
rect 6770 15204 6794 15206
rect 6850 15204 6856 15206
rect 6548 15184 6856 15204
rect 6932 15026 6960 15302
rect 6920 15020 6972 15026
rect 6920 14962 6972 14968
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 6460 14884 6512 14890
rect 6460 14826 6512 14832
rect 6460 14408 6512 14414
rect 6460 14350 6512 14356
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6472 13938 6500 14350
rect 6548 14172 6856 14192
rect 6548 14170 6554 14172
rect 6610 14170 6634 14172
rect 6690 14170 6714 14172
rect 6770 14170 6794 14172
rect 6850 14170 6856 14172
rect 6610 14118 6612 14170
rect 6792 14118 6794 14170
rect 6548 14116 6554 14118
rect 6610 14116 6634 14118
rect 6690 14116 6714 14118
rect 6770 14116 6794 14118
rect 6850 14116 6856 14118
rect 6548 14096 6856 14116
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6184 13796 6236 13802
rect 6184 13738 6236 13744
rect 6276 13796 6328 13802
rect 6276 13738 6328 13744
rect 6092 13320 6144 13326
rect 6092 13262 6144 13268
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6196 12918 6224 13738
rect 6288 13308 6316 13738
rect 6368 13320 6420 13326
rect 6288 13280 6368 13308
rect 6368 13262 6420 13268
rect 6472 12986 6500 13874
rect 7024 13530 7052 14962
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 7208 13326 7236 18566
rect 7300 16794 7328 18958
rect 7392 18290 7420 20878
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 7484 20466 7512 20742
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7576 20330 7604 22066
rect 7654 21448 7710 21457
rect 7654 21383 7710 21392
rect 7668 21146 7696 21383
rect 7656 21140 7708 21146
rect 7656 21082 7708 21088
rect 7748 21140 7800 21146
rect 7748 21082 7800 21088
rect 7656 21004 7708 21010
rect 7656 20946 7708 20952
rect 7668 20874 7696 20946
rect 7656 20868 7708 20874
rect 7656 20810 7708 20816
rect 7760 20602 7788 21082
rect 7748 20596 7800 20602
rect 7748 20538 7800 20544
rect 7564 20324 7616 20330
rect 7564 20266 7616 20272
rect 7564 19984 7616 19990
rect 7564 19926 7616 19932
rect 7576 19718 7604 19926
rect 7760 19922 7788 20538
rect 8036 20534 8064 23800
rect 8484 22228 8536 22234
rect 8484 22170 8536 22176
rect 8496 22030 8524 22170
rect 8680 22094 8708 23800
rect 8680 22066 8892 22094
rect 8484 22024 8536 22030
rect 8668 22024 8720 22030
rect 8536 21984 8616 22012
rect 8484 21966 8536 21972
rect 8116 21956 8168 21962
rect 8116 21898 8168 21904
rect 8392 21956 8444 21962
rect 8392 21898 8444 21904
rect 8128 21622 8156 21898
rect 8116 21616 8168 21622
rect 8116 21558 8168 21564
rect 8404 20874 8432 21898
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8496 21593 8524 21830
rect 8482 21584 8538 21593
rect 8482 21519 8538 21528
rect 8588 21049 8616 21984
rect 8668 21966 8720 21972
rect 8680 21350 8708 21966
rect 8760 21888 8812 21894
rect 8760 21830 8812 21836
rect 8668 21344 8720 21350
rect 8668 21286 8720 21292
rect 8574 21040 8630 21049
rect 8574 20975 8630 20984
rect 8116 20868 8168 20874
rect 8116 20810 8168 20816
rect 8392 20868 8444 20874
rect 8392 20810 8444 20816
rect 8024 20528 8076 20534
rect 8024 20470 8076 20476
rect 8128 20482 8156 20810
rect 8576 20528 8628 20534
rect 8128 20454 8248 20482
rect 8576 20470 8628 20476
rect 8024 20392 8076 20398
rect 8024 20334 8076 20340
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7852 20097 7880 20198
rect 7838 20088 7894 20097
rect 7894 20046 7972 20074
rect 8036 20058 8064 20334
rect 7838 20023 7894 20032
rect 7748 19916 7800 19922
rect 7944 19904 7972 20046
rect 8024 20052 8076 20058
rect 8024 19994 8076 20000
rect 7944 19876 8064 19904
rect 7748 19858 7800 19864
rect 7932 19780 7984 19786
rect 7932 19722 7984 19728
rect 7564 19712 7616 19718
rect 7564 19654 7616 19660
rect 7472 19304 7524 19310
rect 7472 19246 7524 19252
rect 7576 19258 7604 19654
rect 7838 19408 7894 19417
rect 7838 19343 7894 19352
rect 7748 19304 7800 19310
rect 7380 18284 7432 18290
rect 7380 18226 7432 18232
rect 7392 17882 7420 18226
rect 7484 18193 7512 19246
rect 7576 19230 7651 19258
rect 7852 19292 7880 19343
rect 7944 19310 7972 19722
rect 7800 19264 7880 19292
rect 7932 19304 7984 19310
rect 7748 19246 7800 19252
rect 7932 19246 7984 19252
rect 7623 19224 7651 19230
rect 7623 19196 7696 19224
rect 7470 18184 7526 18193
rect 7470 18119 7526 18128
rect 7380 17876 7432 17882
rect 7380 17818 7432 17824
rect 7392 17270 7420 17818
rect 7564 17672 7616 17678
rect 7562 17640 7564 17649
rect 7616 17640 7618 17649
rect 7562 17575 7618 17584
rect 7380 17264 7432 17270
rect 7380 17206 7432 17212
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7668 16658 7696 19196
rect 8036 19156 8064 19876
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8128 19417 8156 19450
rect 8114 19408 8170 19417
rect 8114 19343 8170 19352
rect 7760 19128 8064 19156
rect 7656 16652 7708 16658
rect 7656 16594 7708 16600
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7300 14278 7328 16526
rect 7760 16266 7788 19128
rect 7932 18760 7984 18766
rect 7932 18702 7984 18708
rect 8116 18760 8168 18766
rect 8116 18702 8168 18708
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 7852 16590 7880 17614
rect 7944 16998 7972 18702
rect 8022 17912 8078 17921
rect 8022 17847 8078 17856
rect 8036 17746 8064 17847
rect 8024 17740 8076 17746
rect 8024 17682 8076 17688
rect 8024 17332 8076 17338
rect 8024 17274 8076 17280
rect 7932 16992 7984 16998
rect 7932 16934 7984 16940
rect 7840 16584 7892 16590
rect 7840 16526 7892 16532
rect 7668 16238 7788 16266
rect 7564 15156 7616 15162
rect 7564 15098 7616 15104
rect 7576 14482 7604 15098
rect 7668 15094 7696 16238
rect 7748 16176 7800 16182
rect 7748 16118 7800 16124
rect 7760 15502 7788 16118
rect 7932 15904 7984 15910
rect 7932 15846 7984 15852
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 7760 14958 7788 15438
rect 7944 15434 7972 15846
rect 7932 15428 7984 15434
rect 7932 15370 7984 15376
rect 8036 15144 8064 17274
rect 8128 16522 8156 18702
rect 8220 18329 8248 20454
rect 8484 20324 8536 20330
rect 8484 20266 8536 20272
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8312 18766 8340 20198
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 8404 19514 8432 19654
rect 8392 19508 8444 19514
rect 8392 19450 8444 19456
rect 8392 19168 8444 19174
rect 8392 19110 8444 19116
rect 8300 18760 8352 18766
rect 8300 18702 8352 18708
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8206 18320 8262 18329
rect 8206 18255 8262 18264
rect 8220 18086 8248 18255
rect 8208 18080 8260 18086
rect 8208 18022 8260 18028
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 8220 17338 8248 17478
rect 8208 17332 8260 17338
rect 8208 17274 8260 17280
rect 8312 17202 8340 18566
rect 8404 17338 8432 19110
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8300 16652 8352 16658
rect 8300 16594 8352 16600
rect 8116 16516 8168 16522
rect 8116 16458 8168 16464
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8116 15156 8168 15162
rect 8036 15116 8116 15144
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7564 14476 7616 14482
rect 7564 14418 7616 14424
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 14074 7328 14214
rect 7288 14068 7340 14074
rect 7288 14010 7340 14016
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 6548 13084 6856 13104
rect 6548 13082 6554 13084
rect 6610 13082 6634 13084
rect 6690 13082 6714 13084
rect 6770 13082 6794 13084
rect 6850 13082 6856 13084
rect 6610 13030 6612 13082
rect 6792 13030 6794 13082
rect 6548 13028 6554 13030
rect 6610 13028 6634 13030
rect 6690 13028 6714 13030
rect 6770 13028 6794 13030
rect 6850 13028 6856 13030
rect 6548 13008 6856 13028
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 7116 12918 7144 13262
rect 6184 12912 6236 12918
rect 6184 12854 6236 12860
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 6368 12708 6420 12714
rect 6368 12650 6420 12656
rect 5908 12164 5960 12170
rect 5908 12106 5960 12112
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5356 11892 5408 11898
rect 5356 11834 5408 11840
rect 6012 11830 6040 12038
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5000 11354 5028 11698
rect 4988 11348 5040 11354
rect 4988 11290 5040 11296
rect 5460 11150 5488 11698
rect 6184 11688 6236 11694
rect 6184 11630 6236 11636
rect 5448 11144 5500 11150
rect 5448 11086 5500 11092
rect 5172 11008 5224 11014
rect 5172 10950 5224 10956
rect 5184 10810 5212 10950
rect 5172 10804 5224 10810
rect 5172 10746 5224 10752
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4804 9920 4856 9926
rect 4804 9862 4856 9868
rect 4816 9722 4844 9862
rect 4804 9716 4856 9722
rect 4804 9658 4856 9664
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4908 9042 4936 10542
rect 5368 10062 5396 10610
rect 5460 10470 5488 11086
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 6104 10198 6132 10950
rect 6196 10674 6224 11630
rect 6276 11620 6328 11626
rect 6276 11562 6328 11568
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6092 10192 6144 10198
rect 6092 10134 6144 10140
rect 5356 10056 5408 10062
rect 5356 9998 5408 10004
rect 5368 9654 5396 9998
rect 5356 9648 5408 9654
rect 5356 9590 5408 9596
rect 5368 9042 5396 9590
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5552 9178 5580 9522
rect 5540 9172 5592 9178
rect 5540 9114 5592 9120
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 5356 9036 5408 9042
rect 5356 8978 5408 8984
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 3516 8832 3568 8838
rect 3516 8774 3568 8780
rect 3528 8634 3556 8774
rect 4356 8634 4384 8842
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 3332 8356 3384 8362
rect 3332 8298 3384 8304
rect 3620 7750 3648 8570
rect 3749 8188 4057 8208
rect 3749 8186 3755 8188
rect 3811 8186 3835 8188
rect 3891 8186 3915 8188
rect 3971 8186 3995 8188
rect 4051 8186 4057 8188
rect 3811 8134 3813 8186
rect 3993 8134 3995 8186
rect 3749 8132 3755 8134
rect 3811 8132 3835 8134
rect 3891 8132 3915 8134
rect 3971 8132 3995 8134
rect 4051 8132 4057 8134
rect 3749 8112 4057 8132
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 3608 7744 3660 7750
rect 3608 7686 3660 7692
rect 3252 6886 3372 6914
rect 3056 6860 3108 6866
rect 3056 6802 3108 6808
rect 2964 6724 3016 6730
rect 2964 6666 3016 6672
rect 2976 6458 3004 6666
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 3344 6322 3372 6886
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 3332 6316 3384 6322
rect 3332 6258 3384 6264
rect 2870 6216 2926 6225
rect 2870 6151 2926 6160
rect 2502 5672 2558 5681
rect 2502 5607 2558 5616
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 2240 4185 2268 4422
rect 2226 4176 2282 4185
rect 2226 4111 2282 4120
rect 2044 3528 2096 3534
rect 2044 3470 2096 3476
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1412 3097 1440 3334
rect 2056 3126 2084 3470
rect 2516 3194 2544 5607
rect 2884 4622 2912 6151
rect 3620 5794 3648 7686
rect 3749 7100 4057 7120
rect 3749 7098 3755 7100
rect 3811 7098 3835 7100
rect 3891 7098 3915 7100
rect 3971 7098 3995 7100
rect 4051 7098 4057 7100
rect 3811 7046 3813 7098
rect 3993 7046 3995 7098
rect 3749 7044 3755 7046
rect 3811 7044 3835 7046
rect 3891 7044 3915 7046
rect 3971 7044 3995 7046
rect 4051 7044 4057 7046
rect 3749 7024 4057 7044
rect 4158 6896 4214 6905
rect 4158 6831 4214 6840
rect 3749 6012 4057 6032
rect 3749 6010 3755 6012
rect 3811 6010 3835 6012
rect 3891 6010 3915 6012
rect 3971 6010 3995 6012
rect 4051 6010 4057 6012
rect 3811 5958 3813 6010
rect 3993 5958 3995 6010
rect 3749 5956 3755 5958
rect 3811 5956 3835 5958
rect 3891 5956 3915 5958
rect 3971 5956 3995 5958
rect 4051 5956 4057 5958
rect 3749 5936 4057 5956
rect 3620 5766 3740 5794
rect 3712 5710 3740 5766
rect 3700 5704 3752 5710
rect 3700 5646 3752 5652
rect 3516 5636 3568 5642
rect 3516 5578 3568 5584
rect 2872 4616 2924 4622
rect 2872 4558 2924 4564
rect 2962 4584 3018 4593
rect 2884 4282 2912 4558
rect 2962 4519 2964 4528
rect 3016 4519 3018 4528
rect 2964 4490 3016 4496
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 3424 3936 3476 3942
rect 3424 3878 3476 3884
rect 3238 3496 3294 3505
rect 3238 3431 3294 3440
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2044 3120 2096 3126
rect 1398 3088 1454 3097
rect 2044 3062 2096 3068
rect 2516 3058 2544 3130
rect 1398 3023 1454 3032
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 2504 3052 2556 3058
rect 2504 2994 2556 3000
rect 1596 2961 1624 2994
rect 1582 2952 1638 2961
rect 1582 2887 1638 2896
rect 1860 2848 1912 2854
rect 1860 2790 1912 2796
rect 1872 2446 1900 2790
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 2044 2304 2096 2310
rect 2044 2246 2096 2252
rect 2228 2304 2280 2310
rect 2228 2246 2280 2252
rect 2056 800 2084 2246
rect 2240 2038 2268 2246
rect 2228 2032 2280 2038
rect 2228 1974 2280 1980
rect 2976 1737 3004 3334
rect 3252 3194 3280 3431
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3332 2848 3384 2854
rect 3332 2790 3384 2796
rect 3344 2417 3372 2790
rect 3330 2408 3386 2417
rect 3330 2343 3386 2352
rect 3436 1834 3464 3878
rect 3528 3602 3556 5578
rect 3749 4924 4057 4944
rect 3749 4922 3755 4924
rect 3811 4922 3835 4924
rect 3891 4922 3915 4924
rect 3971 4922 3995 4924
rect 4051 4922 4057 4924
rect 3811 4870 3813 4922
rect 3993 4870 3995 4922
rect 3749 4868 3755 4870
rect 3811 4868 3835 4870
rect 3891 4868 3915 4870
rect 3971 4868 3995 4870
rect 4051 4868 4057 4870
rect 3749 4848 4057 4868
rect 4172 4826 4200 6831
rect 4264 6798 4292 7754
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4528 7404 4580 7410
rect 4528 7346 4580 7352
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 4356 5914 4384 7346
rect 4540 6458 4568 7346
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4632 7002 4660 7278
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4620 5908 4672 5914
rect 4620 5850 4672 5856
rect 4528 5568 4580 5574
rect 4528 5510 4580 5516
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4540 4146 4568 5510
rect 4632 5234 4660 5850
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 3974 4040 4030 4049
rect 3974 3975 3976 3984
rect 4028 3975 4030 3984
rect 3976 3946 4028 3952
rect 3749 3836 4057 3856
rect 3749 3834 3755 3836
rect 3811 3834 3835 3836
rect 3891 3834 3915 3836
rect 3971 3834 3995 3836
rect 4051 3834 4057 3836
rect 3811 3782 3813 3834
rect 3993 3782 3995 3834
rect 3749 3780 3755 3782
rect 3811 3780 3835 3782
rect 3891 3780 3915 3782
rect 3971 3780 3995 3782
rect 4051 3780 4057 3782
rect 3749 3760 4057 3780
rect 4724 3602 4752 8842
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 5264 8832 5316 8838
rect 5264 8774 5316 8780
rect 4908 8634 4936 8774
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5000 8090 5028 8774
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5184 7954 5212 8298
rect 5276 8022 5304 8774
rect 5264 8016 5316 8022
rect 5264 7958 5316 7964
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 4988 7744 5040 7750
rect 4988 7686 5040 7692
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4802 7304 4858 7313
rect 4802 7239 4858 7248
rect 4816 5914 4844 7239
rect 5000 6662 5028 7686
rect 5092 7546 5120 7686
rect 5552 7546 5580 9114
rect 6104 8498 6132 10134
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 5736 8090 5764 8434
rect 6288 8430 6316 11562
rect 6380 11286 6408 12650
rect 7484 12646 7512 13874
rect 7760 13258 7788 14894
rect 7840 14272 7892 14278
rect 7840 14214 7892 14220
rect 7852 13938 7880 14214
rect 8036 14074 8064 15116
rect 8116 15098 8168 15104
rect 8024 14068 8076 14074
rect 8024 14010 8076 14016
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 7748 13252 7800 13258
rect 7748 13194 7800 13200
rect 7760 12918 7788 13194
rect 7748 12912 7800 12918
rect 7748 12854 7800 12860
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 6472 11762 6500 12582
rect 6548 11996 6856 12016
rect 6548 11994 6554 11996
rect 6610 11994 6634 11996
rect 6690 11994 6714 11996
rect 6770 11994 6794 11996
rect 6850 11994 6856 11996
rect 6610 11942 6612 11994
rect 6792 11942 6794 11994
rect 6548 11940 6554 11942
rect 6610 11940 6634 11942
rect 6690 11940 6714 11942
rect 6770 11940 6794 11942
rect 6850 11940 6856 11942
rect 6548 11920 6856 11940
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6368 11280 6420 11286
rect 6368 11222 6420 11228
rect 6472 11150 6500 11698
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6472 10130 6500 11086
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 6548 10908 6856 10928
rect 6548 10906 6554 10908
rect 6610 10906 6634 10908
rect 6690 10906 6714 10908
rect 6770 10906 6794 10908
rect 6850 10906 6856 10908
rect 6610 10854 6612 10906
rect 6792 10854 6794 10906
rect 6548 10852 6554 10854
rect 6610 10852 6634 10854
rect 6690 10852 6714 10854
rect 6770 10852 6794 10854
rect 6850 10852 6856 10854
rect 6548 10832 6856 10852
rect 7024 10810 7052 10950
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6932 10010 6960 10678
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7300 10266 7328 10610
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 6932 9982 7052 10010
rect 6920 9920 6972 9926
rect 6920 9862 6972 9868
rect 6548 9820 6856 9840
rect 6548 9818 6554 9820
rect 6610 9818 6634 9820
rect 6690 9818 6714 9820
rect 6770 9818 6794 9820
rect 6850 9818 6856 9820
rect 6610 9766 6612 9818
rect 6792 9766 6794 9818
rect 6548 9764 6554 9766
rect 6610 9764 6634 9766
rect 6690 9764 6714 9766
rect 6770 9764 6794 9766
rect 6850 9764 6856 9766
rect 6548 9744 6856 9764
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6656 8906 6684 9318
rect 6644 8900 6696 8906
rect 6644 8842 6696 8848
rect 6932 8838 6960 9862
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6548 8732 6856 8752
rect 6548 8730 6554 8732
rect 6610 8730 6634 8732
rect 6690 8730 6714 8732
rect 6770 8730 6794 8732
rect 6850 8730 6856 8732
rect 6610 8678 6612 8730
rect 6792 8678 6794 8730
rect 6548 8676 6554 8678
rect 6610 8676 6634 8678
rect 6690 8676 6714 8678
rect 6770 8676 6794 8678
rect 6850 8676 6856 8678
rect 6548 8656 6856 8676
rect 5816 8424 5868 8430
rect 5816 8366 5868 8372
rect 6276 8424 6328 8430
rect 6276 8366 6328 8372
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5080 7540 5132 7546
rect 5080 7482 5132 7488
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 4804 5908 4856 5914
rect 4804 5850 4856 5856
rect 4804 5772 4856 5778
rect 4804 5714 4856 5720
rect 4816 5234 4844 5714
rect 5184 5574 5212 6122
rect 5356 5908 5408 5914
rect 5356 5850 5408 5856
rect 5368 5710 5396 5850
rect 5460 5778 5488 6938
rect 5552 6798 5580 7482
rect 5828 7274 5856 8366
rect 6932 7886 6960 8774
rect 7024 8634 7052 9982
rect 7484 9586 7512 10406
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7012 8628 7064 8634
rect 7012 8570 7064 8576
rect 7208 8090 7236 9454
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 6920 7880 6972 7886
rect 6920 7822 6972 7828
rect 7012 7744 7064 7750
rect 7012 7686 7064 7692
rect 6548 7644 6856 7664
rect 6548 7642 6554 7644
rect 6610 7642 6634 7644
rect 6690 7642 6714 7644
rect 6770 7642 6794 7644
rect 6850 7642 6856 7644
rect 6610 7590 6612 7642
rect 6792 7590 6794 7642
rect 6548 7588 6554 7590
rect 6610 7588 6634 7590
rect 6690 7588 6714 7590
rect 6770 7588 6794 7590
rect 6850 7588 6856 7590
rect 6548 7568 6856 7588
rect 5816 7268 5868 7274
rect 5816 7210 5868 7216
rect 6368 7268 6420 7274
rect 6368 7210 6420 7216
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5448 5772 5500 5778
rect 5448 5714 5500 5720
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5080 5568 5132 5574
rect 5080 5510 5132 5516
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 5092 5302 5120 5510
rect 5276 5370 5304 5646
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 5264 5364 5316 5370
rect 5264 5306 5316 5312
rect 5080 5296 5132 5302
rect 5080 5238 5132 5244
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4816 4078 4844 5170
rect 5080 4480 5132 4486
rect 5080 4422 5132 4428
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4816 3602 4844 4014
rect 3516 3596 3568 3602
rect 3516 3538 3568 3544
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4804 3596 4856 3602
rect 4804 3538 4856 3544
rect 3528 3126 3556 3538
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 4816 3058 4844 3538
rect 5092 3058 5120 4422
rect 5184 4282 5212 5306
rect 5552 5302 5580 6394
rect 6196 6322 6224 6802
rect 6380 6322 6408 7210
rect 6548 6556 6856 6576
rect 6548 6554 6554 6556
rect 6610 6554 6634 6556
rect 6690 6554 6714 6556
rect 6770 6554 6794 6556
rect 6850 6554 6856 6556
rect 6610 6502 6612 6554
rect 6792 6502 6794 6554
rect 6548 6500 6554 6502
rect 6610 6500 6634 6502
rect 6690 6500 6714 6502
rect 6770 6500 6794 6502
rect 6850 6500 6856 6502
rect 6548 6480 6856 6500
rect 7024 6458 7052 7686
rect 7852 7342 7880 13874
rect 8024 13864 8076 13870
rect 8024 13806 8076 13812
rect 8036 12238 8064 13806
rect 8128 12850 8156 13942
rect 8220 13190 8248 16390
rect 8312 16250 8340 16594
rect 8496 16590 8524 20266
rect 8588 19258 8616 20470
rect 8680 19922 8708 21286
rect 8668 19916 8720 19922
rect 8668 19858 8720 19864
rect 8668 19304 8720 19310
rect 8588 19252 8668 19258
rect 8588 19246 8720 19252
rect 8588 19230 8708 19246
rect 8588 18850 8616 19230
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8680 18970 8708 19110
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 8588 18822 8708 18850
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8588 18086 8616 18702
rect 8680 18358 8708 18822
rect 8668 18352 8720 18358
rect 8668 18294 8720 18300
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8588 16726 8616 18022
rect 8668 17808 8720 17814
rect 8666 17776 8668 17785
rect 8720 17776 8722 17785
rect 8666 17711 8722 17720
rect 8666 17640 8722 17649
rect 8666 17575 8722 17584
rect 8680 17542 8708 17575
rect 8668 17536 8720 17542
rect 8668 17478 8720 17484
rect 8668 17128 8720 17134
rect 8668 17070 8720 17076
rect 8680 16794 8708 17070
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8576 16720 8628 16726
rect 8576 16662 8628 16668
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8300 16244 8352 16250
rect 8300 16186 8352 16192
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8588 14482 8616 15302
rect 8772 14958 8800 21830
rect 8864 20602 8892 22066
rect 8944 21684 8996 21690
rect 8944 21626 8996 21632
rect 8852 20596 8904 20602
rect 8852 20538 8904 20544
rect 8864 19446 8892 20538
rect 8852 19440 8904 19446
rect 8852 19382 8904 19388
rect 8852 19236 8904 19242
rect 8852 19178 8904 19184
rect 8864 18834 8892 19178
rect 8852 18828 8904 18834
rect 8852 18770 8904 18776
rect 8850 17912 8906 17921
rect 8850 17847 8906 17856
rect 8864 17338 8892 17847
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8588 13938 8616 14418
rect 8864 14414 8892 17138
rect 8852 14408 8904 14414
rect 8852 14350 8904 14356
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8956 13326 8984 21626
rect 9048 21554 9076 23854
rect 9232 23746 9260 23854
rect 9310 23800 9366 24600
rect 9954 23800 10010 24600
rect 10598 23800 10654 24600
rect 11242 23800 11298 24600
rect 11886 23800 11942 24600
rect 12530 23800 12586 24600
rect 13174 23800 13230 24600
rect 13818 23800 13874 24600
rect 14462 23800 14518 24600
rect 14660 23854 15056 23882
rect 9324 23746 9352 23800
rect 9232 23718 9352 23746
rect 9347 22332 9655 22352
rect 9347 22330 9353 22332
rect 9409 22330 9433 22332
rect 9489 22330 9513 22332
rect 9569 22330 9593 22332
rect 9649 22330 9655 22332
rect 9409 22278 9411 22330
rect 9591 22278 9593 22330
rect 9347 22276 9353 22278
rect 9409 22276 9433 22278
rect 9489 22276 9513 22278
rect 9569 22276 9593 22278
rect 9649 22276 9655 22278
rect 9347 22256 9655 22276
rect 9968 22094 9996 23800
rect 9876 22066 9996 22094
rect 9128 22024 9180 22030
rect 9126 21992 9128 22001
rect 9180 21992 9182 22001
rect 9126 21927 9182 21936
rect 9876 21690 9904 22066
rect 10324 22024 10376 22030
rect 10138 21992 10194 22001
rect 10324 21966 10376 21972
rect 10138 21927 10194 21936
rect 9956 21888 10008 21894
rect 9956 21830 10008 21836
rect 9864 21684 9916 21690
rect 9864 21626 9916 21632
rect 9220 21616 9272 21622
rect 9220 21558 9272 21564
rect 9036 21548 9088 21554
rect 9036 21490 9088 21496
rect 9128 21548 9180 21554
rect 9128 21490 9180 21496
rect 9048 20913 9076 21490
rect 9034 20904 9090 20913
rect 9034 20839 9090 20848
rect 9140 20788 9168 21490
rect 9232 21146 9260 21558
rect 9680 21548 9732 21554
rect 9680 21490 9732 21496
rect 9692 21457 9720 21490
rect 9678 21448 9734 21457
rect 9678 21383 9734 21392
rect 9772 21412 9824 21418
rect 9824 21372 9904 21400
rect 9772 21354 9824 21360
rect 9347 21244 9655 21264
rect 9347 21242 9353 21244
rect 9409 21242 9433 21244
rect 9489 21242 9513 21244
rect 9569 21242 9593 21244
rect 9649 21242 9655 21244
rect 9409 21190 9411 21242
rect 9591 21190 9593 21242
rect 9347 21188 9353 21190
rect 9409 21188 9433 21190
rect 9489 21188 9513 21190
rect 9569 21188 9593 21190
rect 9649 21188 9655 21190
rect 9347 21168 9655 21188
rect 9220 21140 9272 21146
rect 9220 21082 9272 21088
rect 9404 21072 9456 21078
rect 9404 21014 9456 21020
rect 9680 21072 9732 21078
rect 9680 21014 9732 21020
rect 9312 20936 9364 20942
rect 9310 20904 9312 20913
rect 9364 20904 9366 20913
rect 9310 20839 9366 20848
rect 9416 20806 9444 21014
rect 9496 20868 9548 20874
rect 9496 20810 9548 20816
rect 9048 20760 9168 20788
rect 9404 20800 9456 20806
rect 9048 19174 9076 20760
rect 9404 20742 9456 20748
rect 9508 20602 9536 20810
rect 9496 20596 9548 20602
rect 9496 20538 9548 20544
rect 9692 20466 9720 21014
rect 9772 20868 9824 20874
rect 9772 20810 9824 20816
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9218 20360 9274 20369
rect 9218 20295 9274 20304
rect 9680 20324 9732 20330
rect 9232 20262 9260 20295
rect 9680 20266 9732 20272
rect 9220 20256 9272 20262
rect 9220 20198 9272 20204
rect 9347 20156 9655 20176
rect 9347 20154 9353 20156
rect 9409 20154 9433 20156
rect 9489 20154 9513 20156
rect 9569 20154 9593 20156
rect 9649 20154 9655 20156
rect 9409 20102 9411 20154
rect 9591 20102 9593 20154
rect 9347 20100 9353 20102
rect 9409 20100 9433 20102
rect 9489 20100 9513 20102
rect 9569 20100 9593 20102
rect 9649 20100 9655 20102
rect 9347 20080 9655 20100
rect 9692 19990 9720 20266
rect 9784 20058 9812 20810
rect 9772 20052 9824 20058
rect 9772 19994 9824 20000
rect 9680 19984 9732 19990
rect 9680 19926 9732 19932
rect 9220 19916 9272 19922
rect 9220 19858 9272 19864
rect 9232 19378 9260 19858
rect 9678 19816 9734 19825
rect 9678 19751 9734 19760
rect 9772 19780 9824 19786
rect 9220 19372 9272 19378
rect 9220 19314 9272 19320
rect 9036 19168 9088 19174
rect 9036 19110 9088 19116
rect 9128 19168 9180 19174
rect 9128 19110 9180 19116
rect 9140 18222 9168 19110
rect 9232 18834 9260 19314
rect 9347 19068 9655 19088
rect 9347 19066 9353 19068
rect 9409 19066 9433 19068
rect 9489 19066 9513 19068
rect 9569 19066 9593 19068
rect 9649 19066 9655 19068
rect 9409 19014 9411 19066
rect 9591 19014 9593 19066
rect 9347 19012 9353 19014
rect 9409 19012 9433 19014
rect 9489 19012 9513 19014
rect 9569 19012 9593 19014
rect 9649 19012 9655 19014
rect 9347 18992 9655 19012
rect 9692 18902 9720 19751
rect 9772 19722 9824 19728
rect 9784 19514 9812 19722
rect 9772 19508 9824 19514
rect 9772 19450 9824 19456
rect 9312 18896 9364 18902
rect 9310 18864 9312 18873
rect 9680 18896 9732 18902
rect 9364 18864 9366 18873
rect 9220 18828 9272 18834
rect 9680 18838 9732 18844
rect 9310 18799 9366 18808
rect 9220 18770 9272 18776
rect 9128 18216 9180 18222
rect 9128 18158 9180 18164
rect 9036 17808 9088 17814
rect 9036 17750 9088 17756
rect 9048 17610 9076 17750
rect 9036 17604 9088 17610
rect 9036 17546 9088 17552
rect 9048 15026 9076 17546
rect 9140 17202 9168 18158
rect 9232 17678 9260 18770
rect 9680 18760 9732 18766
rect 9680 18702 9732 18708
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9508 18222 9536 18566
rect 9496 18216 9548 18222
rect 9496 18158 9548 18164
rect 9347 17980 9655 18000
rect 9347 17978 9353 17980
rect 9409 17978 9433 17980
rect 9489 17978 9513 17980
rect 9569 17978 9593 17980
rect 9649 17978 9655 17980
rect 9409 17926 9411 17978
rect 9591 17926 9593 17978
rect 9347 17924 9353 17926
rect 9409 17924 9433 17926
rect 9489 17924 9513 17926
rect 9569 17924 9593 17926
rect 9649 17924 9655 17926
rect 9347 17904 9655 17924
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9692 17338 9720 18702
rect 9784 18222 9812 19450
rect 9876 19378 9904 21372
rect 9968 20466 9996 21830
rect 10048 21480 10100 21486
rect 10048 21422 10100 21428
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 10060 19666 10088 21422
rect 10152 20369 10180 21927
rect 10336 21690 10364 21966
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10324 21684 10376 21690
rect 10324 21626 10376 21632
rect 10232 21616 10284 21622
rect 10232 21558 10284 21564
rect 10138 20360 10194 20369
rect 10138 20295 10194 20304
rect 10244 19825 10272 21558
rect 10416 21344 10468 21350
rect 10416 21286 10468 21292
rect 10324 20256 10376 20262
rect 10324 20198 10376 20204
rect 10230 19816 10286 19825
rect 10140 19780 10192 19786
rect 10230 19751 10286 19760
rect 10140 19722 10192 19728
rect 9968 19638 10088 19666
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9864 19236 9916 19242
rect 9864 19178 9916 19184
rect 9772 18216 9824 18222
rect 9770 18184 9772 18193
rect 9824 18184 9826 18193
rect 9770 18119 9826 18128
rect 9680 17332 9732 17338
rect 9680 17274 9732 17280
rect 9128 17196 9180 17202
rect 9128 17138 9180 17144
rect 9126 17096 9182 17105
rect 9126 17031 9182 17040
rect 9140 16998 9168 17031
rect 9128 16992 9180 16998
rect 9128 16934 9180 16940
rect 9347 16892 9655 16912
rect 9347 16890 9353 16892
rect 9409 16890 9433 16892
rect 9489 16890 9513 16892
rect 9569 16890 9593 16892
rect 9649 16890 9655 16892
rect 9409 16838 9411 16890
rect 9591 16838 9593 16890
rect 9347 16836 9353 16838
rect 9409 16836 9433 16838
rect 9489 16836 9513 16838
rect 9569 16836 9593 16838
rect 9649 16836 9655 16838
rect 9347 16816 9655 16836
rect 9220 16652 9272 16658
rect 9220 16594 9272 16600
rect 9128 16108 9180 16114
rect 9128 16050 9180 16056
rect 9036 15020 9088 15026
rect 9036 14962 9088 14968
rect 9140 14074 9168 16050
rect 9232 14618 9260 16594
rect 9876 16454 9904 19178
rect 9968 19174 9996 19638
rect 10046 19544 10102 19553
rect 10046 19479 10048 19488
rect 10100 19479 10102 19488
rect 10048 19450 10100 19456
rect 9956 19168 10008 19174
rect 9956 19110 10008 19116
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 10060 18426 10088 18566
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9680 16448 9732 16454
rect 9864 16448 9916 16454
rect 9680 16390 9732 16396
rect 9784 16408 9864 16436
rect 9508 16250 9536 16390
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9347 15804 9655 15824
rect 9347 15802 9353 15804
rect 9409 15802 9433 15804
rect 9489 15802 9513 15804
rect 9569 15802 9593 15804
rect 9649 15802 9655 15804
rect 9409 15750 9411 15802
rect 9591 15750 9593 15802
rect 9347 15748 9353 15750
rect 9409 15748 9433 15750
rect 9489 15748 9513 15750
rect 9569 15748 9593 15750
rect 9649 15748 9655 15750
rect 9347 15728 9655 15748
rect 9692 15042 9720 16390
rect 9784 15502 9812 16408
rect 9864 16390 9916 16396
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 9864 16244 9916 16250
rect 9864 16186 9916 16192
rect 9876 15570 9904 16186
rect 9864 15564 9916 15570
rect 9864 15506 9916 15512
rect 10060 15502 10088 16390
rect 10152 15706 10180 19722
rect 10336 19514 10364 20198
rect 10324 19508 10376 19514
rect 10324 19450 10376 19456
rect 10324 18692 10376 18698
rect 10324 18634 10376 18640
rect 10336 17610 10364 18634
rect 10324 17604 10376 17610
rect 10324 17546 10376 17552
rect 10428 16794 10456 21286
rect 10520 20913 10548 21830
rect 10612 21622 10640 23800
rect 11060 21888 11112 21894
rect 11060 21830 11112 21836
rect 10600 21616 10652 21622
rect 10600 21558 10652 21564
rect 10506 20904 10562 20913
rect 10562 20862 10640 20890
rect 10506 20839 10562 20848
rect 10508 19168 10560 19174
rect 10508 19110 10560 19116
rect 10520 18902 10548 19110
rect 10508 18896 10560 18902
rect 10508 18838 10560 18844
rect 10520 18766 10548 18838
rect 10508 18760 10560 18766
rect 10508 18702 10560 18708
rect 10612 17542 10640 20862
rect 11072 20058 11100 21830
rect 11256 21554 11284 23800
rect 11900 22094 11928 23800
rect 12544 22234 12572 23800
rect 12532 22228 12584 22234
rect 12532 22170 12584 22176
rect 13084 22160 13136 22166
rect 13084 22102 13136 22108
rect 11900 22066 12020 22094
rect 11520 21956 11572 21962
rect 11520 21898 11572 21904
rect 11244 21548 11296 21554
rect 11244 21490 11296 21496
rect 11336 21480 11388 21486
rect 11336 21422 11388 21428
rect 11348 21146 11376 21422
rect 11336 21140 11388 21146
rect 11336 21082 11388 21088
rect 11152 20324 11204 20330
rect 11152 20266 11204 20272
rect 11060 20052 11112 20058
rect 11060 19994 11112 20000
rect 11164 19938 11192 20266
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 11072 19910 11192 19938
rect 11072 19530 11100 19910
rect 11150 19816 11206 19825
rect 11150 19751 11206 19760
rect 11164 19718 11192 19751
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 10980 19502 11100 19530
rect 10784 19304 10836 19310
rect 10784 19246 10836 19252
rect 10796 18766 10824 19246
rect 10980 19156 11008 19502
rect 11060 19440 11112 19446
rect 11060 19382 11112 19388
rect 11072 19224 11100 19382
rect 11164 19378 11192 19654
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11072 19196 11192 19224
rect 10980 19128 11100 19156
rect 10784 18760 10836 18766
rect 10784 18702 10836 18708
rect 10796 18154 10824 18702
rect 10876 18624 10928 18630
rect 10874 18592 10876 18601
rect 10968 18624 11020 18630
rect 10928 18592 10930 18601
rect 10968 18566 11020 18572
rect 10874 18527 10930 18536
rect 10980 18290 11008 18566
rect 10968 18284 11020 18290
rect 10968 18226 11020 18232
rect 10784 18148 10836 18154
rect 10784 18090 10836 18096
rect 11072 17762 11100 19128
rect 11164 18465 11192 19196
rect 11256 19174 11284 20198
rect 11348 19922 11376 21082
rect 11532 21010 11560 21898
rect 11796 21888 11848 21894
rect 11796 21830 11848 21836
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11520 19984 11572 19990
rect 11520 19926 11572 19932
rect 11336 19916 11388 19922
rect 11336 19858 11388 19864
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 11244 19168 11296 19174
rect 11244 19110 11296 19116
rect 11440 18834 11468 19654
rect 11532 19378 11560 19926
rect 11808 19802 11836 21830
rect 11888 21140 11940 21146
rect 11888 21082 11940 21088
rect 11900 19922 11928 21082
rect 11992 20466 12020 22066
rect 12164 22024 12216 22030
rect 12162 21992 12164 22001
rect 12216 21992 12218 22001
rect 12162 21927 12218 21936
rect 12438 21992 12494 22001
rect 12438 21927 12440 21936
rect 12492 21927 12494 21936
rect 12992 21956 13044 21962
rect 12440 21898 12492 21904
rect 12992 21898 13044 21904
rect 12072 21888 12124 21894
rect 12072 21830 12124 21836
rect 12084 21418 12112 21830
rect 12146 21788 12454 21808
rect 12146 21786 12152 21788
rect 12208 21786 12232 21788
rect 12288 21786 12312 21788
rect 12368 21786 12392 21788
rect 12448 21786 12454 21788
rect 12208 21734 12210 21786
rect 12390 21734 12392 21786
rect 12146 21732 12152 21734
rect 12208 21732 12232 21734
rect 12288 21732 12312 21734
rect 12368 21732 12392 21734
rect 12448 21732 12454 21734
rect 12146 21712 12454 21732
rect 13004 21690 13032 21898
rect 12992 21684 13044 21690
rect 12992 21626 13044 21632
rect 12532 21616 12584 21622
rect 12532 21558 12584 21564
rect 12164 21548 12216 21554
rect 12164 21490 12216 21496
rect 12072 21412 12124 21418
rect 12072 21354 12124 21360
rect 12176 21146 12204 21490
rect 12164 21140 12216 21146
rect 12164 21082 12216 21088
rect 12544 21010 12572 21558
rect 12900 21412 12952 21418
rect 12900 21354 12952 21360
rect 12912 21146 12940 21354
rect 12900 21140 12952 21146
rect 12900 21082 12952 21088
rect 12532 21004 12584 21010
rect 12532 20946 12584 20952
rect 12072 20936 12124 20942
rect 12072 20878 12124 20884
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 11888 19916 11940 19922
rect 11888 19858 11940 19864
rect 12084 19854 12112 20878
rect 12146 20700 12454 20720
rect 12146 20698 12152 20700
rect 12208 20698 12232 20700
rect 12288 20698 12312 20700
rect 12368 20698 12392 20700
rect 12448 20698 12454 20700
rect 12208 20646 12210 20698
rect 12390 20646 12392 20698
rect 12146 20644 12152 20646
rect 12208 20644 12232 20646
rect 12288 20644 12312 20646
rect 12368 20644 12392 20646
rect 12448 20644 12454 20646
rect 12146 20624 12454 20644
rect 12544 20534 12572 20946
rect 12624 20800 12676 20806
rect 12624 20742 12676 20748
rect 12532 20528 12584 20534
rect 12532 20470 12584 20476
rect 12636 20448 12664 20742
rect 12716 20460 12768 20466
rect 12636 20420 12716 20448
rect 12716 20402 12768 20408
rect 13096 19922 13124 22102
rect 13188 21418 13216 23800
rect 13360 22024 13412 22030
rect 13360 21966 13412 21972
rect 13268 21548 13320 21554
rect 13268 21490 13320 21496
rect 13176 21412 13228 21418
rect 13176 21354 13228 21360
rect 13280 20505 13308 21490
rect 13372 21486 13400 21966
rect 13636 21956 13688 21962
rect 13636 21898 13688 21904
rect 13360 21480 13412 21486
rect 13360 21422 13412 21428
rect 13544 21480 13596 21486
rect 13544 21422 13596 21428
rect 13266 20496 13322 20505
rect 13266 20431 13322 20440
rect 13084 19916 13136 19922
rect 13084 19858 13136 19864
rect 12072 19848 12124 19854
rect 11992 19808 12072 19836
rect 11808 19774 11928 19802
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11612 19508 11664 19514
rect 11612 19450 11664 19456
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11520 19168 11572 19174
rect 11520 19110 11572 19116
rect 11428 18828 11480 18834
rect 11428 18770 11480 18776
rect 11150 18456 11206 18465
rect 11150 18391 11206 18400
rect 11244 18148 11296 18154
rect 11244 18090 11296 18096
rect 10980 17734 11100 17762
rect 10600 17536 10652 17542
rect 10600 17478 10652 17484
rect 10416 16788 10468 16794
rect 10416 16730 10468 16736
rect 10416 15904 10468 15910
rect 10416 15846 10468 15852
rect 10140 15700 10192 15706
rect 10140 15642 10192 15648
rect 10428 15638 10456 15846
rect 10416 15632 10468 15638
rect 10416 15574 10468 15580
rect 9772 15496 9824 15502
rect 9772 15438 9824 15444
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 9416 15014 9720 15042
rect 9416 14958 9444 15014
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 9680 14952 9732 14958
rect 9680 14894 9732 14900
rect 9347 14716 9655 14736
rect 9347 14714 9353 14716
rect 9409 14714 9433 14716
rect 9489 14714 9513 14716
rect 9569 14714 9593 14716
rect 9649 14714 9655 14716
rect 9409 14662 9411 14714
rect 9591 14662 9593 14714
rect 9347 14660 9353 14662
rect 9409 14660 9433 14662
rect 9489 14660 9513 14662
rect 9569 14660 9593 14662
rect 9649 14660 9655 14662
rect 9347 14640 9655 14660
rect 9220 14612 9272 14618
rect 9692 14600 9720 14894
rect 10152 14618 10180 15438
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10888 14618 10916 15302
rect 9220 14554 9272 14560
rect 9600 14572 9720 14600
rect 10140 14612 10192 14618
rect 9600 14414 9628 14572
rect 10140 14554 10192 14560
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 9588 14408 9640 14414
rect 9588 14350 9640 14356
rect 10232 14408 10284 14414
rect 10232 14350 10284 14356
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 9128 13932 9180 13938
rect 9128 13874 9180 13880
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 8944 13320 8996 13326
rect 8944 13262 8996 13268
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8588 12918 8616 13126
rect 8772 12940 9076 12968
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 8392 12232 8444 12238
rect 8392 12174 8444 12180
rect 8404 11150 8432 12174
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11898 8524 12038
rect 8484 11892 8536 11898
rect 8484 11834 8536 11840
rect 8588 11694 8616 12854
rect 8772 12782 8800 12940
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8760 12776 8812 12782
rect 8760 12718 8812 12724
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8300 11008 8352 11014
rect 8300 10950 8352 10956
rect 8312 10062 8340 10950
rect 8588 10062 8616 11086
rect 8680 10810 8708 12174
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 8772 10606 8800 12718
rect 8864 11898 8892 12786
rect 9048 12714 9076 12940
rect 9036 12708 9088 12714
rect 9036 12650 9088 12656
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8956 12238 8984 12582
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 9140 11354 9168 13874
rect 9680 13796 9732 13802
rect 9680 13738 9732 13744
rect 9347 13628 9655 13648
rect 9347 13626 9353 13628
rect 9409 13626 9433 13628
rect 9489 13626 9513 13628
rect 9569 13626 9593 13628
rect 9649 13626 9655 13628
rect 9409 13574 9411 13626
rect 9591 13574 9593 13626
rect 9347 13572 9353 13574
rect 9409 13572 9433 13574
rect 9489 13572 9513 13574
rect 9569 13572 9593 13574
rect 9649 13572 9655 13574
rect 9347 13552 9655 13572
rect 9692 13512 9720 13738
rect 9508 13484 9720 13512
rect 9508 13394 9536 13484
rect 9968 13462 9996 13874
rect 10244 13462 10272 14350
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10520 13530 10548 13874
rect 10876 13864 10928 13870
rect 10876 13806 10928 13812
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 9496 13388 9548 13394
rect 9496 13330 9548 13336
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9600 12918 9628 13330
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9347 12540 9655 12560
rect 9347 12538 9353 12540
rect 9409 12538 9433 12540
rect 9489 12538 9513 12540
rect 9569 12538 9593 12540
rect 9649 12538 9655 12540
rect 9409 12486 9411 12538
rect 9591 12486 9593 12538
rect 9347 12484 9353 12486
rect 9409 12484 9433 12486
rect 9489 12484 9513 12486
rect 9569 12484 9593 12486
rect 9649 12484 9655 12486
rect 9347 12464 9655 12484
rect 9692 12442 9720 13126
rect 9680 12436 9732 12442
rect 9680 12378 9732 12384
rect 9784 12374 9812 13126
rect 9968 12986 9996 13398
rect 10140 13320 10192 13326
rect 10140 13262 10192 13268
rect 10152 12986 10180 13262
rect 10600 13252 10652 13258
rect 10600 13194 10652 13200
rect 9956 12980 10008 12986
rect 9956 12922 10008 12928
rect 10140 12980 10192 12986
rect 10140 12922 10192 12928
rect 9772 12368 9824 12374
rect 9772 12310 9824 12316
rect 10612 12170 10640 13194
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9347 11452 9655 11472
rect 9347 11450 9353 11452
rect 9409 11450 9433 11452
rect 9489 11450 9513 11452
rect 9569 11450 9593 11452
rect 9649 11450 9655 11452
rect 9409 11398 9411 11450
rect 9591 11398 9593 11450
rect 9347 11396 9353 11398
rect 9409 11396 9433 11398
rect 9489 11396 9513 11398
rect 9569 11396 9593 11398
rect 9649 11396 9655 11398
rect 9347 11376 9655 11396
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8956 10810 8984 11086
rect 9692 11082 9720 11494
rect 10060 11354 10088 11698
rect 10048 11348 10100 11354
rect 10048 11290 10100 11296
rect 10508 11144 10560 11150
rect 10508 11086 10560 11092
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 10520 10742 10548 11086
rect 10692 11076 10744 11082
rect 10692 11018 10744 11024
rect 9772 10736 9824 10742
rect 9772 10678 9824 10684
rect 10508 10736 10560 10742
rect 10508 10678 10560 10684
rect 8944 10668 8996 10674
rect 8944 10610 8996 10616
rect 8760 10600 8812 10606
rect 8760 10542 8812 10548
rect 8956 10266 8984 10610
rect 9680 10532 9732 10538
rect 9680 10474 9732 10480
rect 9347 10364 9655 10384
rect 9347 10362 9353 10364
rect 9409 10362 9433 10364
rect 9489 10362 9513 10364
rect 9569 10362 9593 10364
rect 9649 10362 9655 10364
rect 9409 10310 9411 10362
rect 9591 10310 9593 10362
rect 9347 10308 9353 10310
rect 9409 10308 9433 10310
rect 9489 10308 9513 10310
rect 9569 10308 9593 10310
rect 9649 10308 9655 10310
rect 9347 10288 9655 10308
rect 8944 10260 8996 10266
rect 8944 10202 8996 10208
rect 9692 10130 9720 10474
rect 9680 10124 9732 10130
rect 9680 10066 9732 10072
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 9588 10056 9640 10062
rect 9588 9998 9640 10004
rect 8588 9654 8616 9998
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 9404 9920 9456 9926
rect 9404 9862 9456 9868
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8772 9110 8800 9862
rect 9416 9722 9444 9862
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9600 9586 9628 9998
rect 9680 9988 9732 9994
rect 9680 9930 9732 9936
rect 9692 9654 9720 9930
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9347 9276 9655 9296
rect 9347 9274 9353 9276
rect 9409 9274 9433 9276
rect 9489 9274 9513 9276
rect 9569 9274 9593 9276
rect 9649 9274 9655 9276
rect 9409 9222 9411 9274
rect 9591 9222 9593 9274
rect 9347 9220 9353 9222
rect 9409 9220 9433 9222
rect 9489 9220 9513 9222
rect 9569 9220 9593 9222
rect 9649 9220 9655 9222
rect 9347 9200 9655 9220
rect 8392 9104 8444 9110
rect 8312 9064 8392 9092
rect 8312 8514 8340 9064
rect 8392 9046 8444 9052
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8220 8498 8340 8514
rect 8404 8498 8432 8910
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8208 8492 8340 8498
rect 8260 8486 8340 8492
rect 8392 8492 8444 8498
rect 8208 8434 8260 8440
rect 8392 8434 8444 8440
rect 8588 8090 8616 8842
rect 9784 8634 9812 10678
rect 10520 10062 10548 10678
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9680 8356 9732 8362
rect 9680 8298 9732 8304
rect 9347 8188 9655 8208
rect 9347 8186 9353 8188
rect 9409 8186 9433 8188
rect 9489 8186 9513 8188
rect 9569 8186 9593 8188
rect 9649 8186 9655 8188
rect 9409 8134 9411 8186
rect 9591 8134 9593 8186
rect 9347 8132 9353 8134
rect 9409 8132 9433 8134
rect 9489 8132 9513 8134
rect 9569 8132 9593 8134
rect 9649 8132 9655 8134
rect 9347 8112 9655 8132
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 9692 7886 9720 8298
rect 9876 8090 9904 9522
rect 10520 9042 10548 9998
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10520 8634 10548 8774
rect 10704 8634 10732 11018
rect 10888 10606 10916 13806
rect 10980 13734 11008 17734
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 11072 17202 11100 17614
rect 11256 17241 11284 18090
rect 11242 17232 11298 17241
rect 11060 17196 11112 17202
rect 11242 17167 11298 17176
rect 11060 17138 11112 17144
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11256 16182 11284 16526
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11072 15706 11100 16050
rect 11060 15700 11112 15706
rect 11060 15642 11112 15648
rect 11256 15094 11284 16118
rect 11440 15638 11468 18770
rect 11532 18222 11560 19110
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11532 17338 11560 18158
rect 11624 17338 11652 19450
rect 11808 19242 11836 19654
rect 11796 19236 11848 19242
rect 11796 19178 11848 19184
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11716 18873 11744 19110
rect 11702 18864 11758 18873
rect 11702 18799 11758 18808
rect 11702 18592 11758 18601
rect 11702 18527 11758 18536
rect 11716 18426 11744 18527
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11716 18193 11744 18226
rect 11702 18184 11758 18193
rect 11702 18119 11758 18128
rect 11520 17332 11572 17338
rect 11520 17274 11572 17280
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11704 17196 11756 17202
rect 11704 17138 11756 17144
rect 11520 16992 11572 16998
rect 11716 16980 11744 17138
rect 11796 16992 11848 16998
rect 11572 16952 11652 16980
rect 11716 16952 11796 16980
rect 11520 16934 11572 16940
rect 11520 16788 11572 16794
rect 11520 16730 11572 16736
rect 11428 15632 11480 15638
rect 11428 15574 11480 15580
rect 11336 15496 11388 15502
rect 11336 15438 11388 15444
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 11072 14822 11100 14962
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 11152 14816 11204 14822
rect 11152 14758 11204 14764
rect 11072 14074 11100 14758
rect 11164 14482 11192 14758
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11256 13938 11284 15030
rect 11348 14414 11376 15438
rect 11336 14408 11388 14414
rect 11336 14350 11388 14356
rect 11348 14006 11376 14350
rect 11428 14272 11480 14278
rect 11428 14214 11480 14220
rect 11440 14006 11468 14214
rect 11336 14000 11388 14006
rect 11336 13942 11388 13948
rect 11428 14000 11480 14006
rect 11428 13942 11480 13948
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11244 13932 11296 13938
rect 11244 13874 11296 13880
rect 10968 13728 11020 13734
rect 10968 13670 11020 13676
rect 11164 13190 11192 13874
rect 11152 13184 11204 13190
rect 11152 13126 11204 13132
rect 11164 12714 11192 13126
rect 11532 12850 11560 16730
rect 11624 15858 11652 16952
rect 11796 16934 11848 16940
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11716 16046 11744 16390
rect 11704 16040 11756 16046
rect 11704 15982 11756 15988
rect 11624 15830 11744 15858
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 11624 15162 11652 15506
rect 11612 15156 11664 15162
rect 11612 15098 11664 15104
rect 11716 14226 11744 15830
rect 11808 14346 11836 16934
rect 11796 14340 11848 14346
rect 11796 14282 11848 14288
rect 11716 14198 11836 14226
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11152 12708 11204 12714
rect 11152 12650 11204 12656
rect 11520 12232 11572 12238
rect 11520 12174 11572 12180
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11336 12096 11388 12102
rect 11336 12038 11388 12044
rect 10968 11688 11020 11694
rect 10968 11630 11020 11636
rect 10980 11354 11008 11630
rect 11348 11354 11376 12038
rect 10968 11348 11020 11354
rect 10968 11290 11020 11296
rect 11336 11348 11388 11354
rect 11336 11290 11388 11296
rect 10968 10804 11020 10810
rect 10968 10746 11020 10752
rect 10876 10600 10928 10606
rect 10876 10542 10928 10548
rect 10888 10266 10916 10542
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10508 8628 10560 8634
rect 10508 8570 10560 8576
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9680 7880 9732 7886
rect 9034 7848 9090 7857
rect 8024 7812 8076 7818
rect 8024 7754 8076 7760
rect 8576 7812 8628 7818
rect 9680 7822 9732 7828
rect 9034 7783 9090 7792
rect 8576 7754 8628 7760
rect 8036 7478 8064 7754
rect 8024 7472 8076 7478
rect 8024 7414 8076 7420
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7392 6746 7420 7278
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7576 7002 7604 7142
rect 7564 6996 7616 7002
rect 7564 6938 7616 6944
rect 7392 6718 7604 6746
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7208 6390 7236 6598
rect 7484 6458 7512 6598
rect 7576 6458 7604 6718
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7196 6384 7248 6390
rect 7196 6326 7248 6332
rect 8036 6322 8064 7414
rect 8588 7206 8616 7754
rect 9048 7410 9076 7783
rect 9220 7744 9272 7750
rect 9220 7686 9272 7692
rect 9036 7404 9088 7410
rect 9036 7346 9088 7352
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8128 6730 8156 7142
rect 8588 6866 8616 7142
rect 8300 6860 8352 6866
rect 8300 6802 8352 6808
rect 8576 6860 8628 6866
rect 8576 6802 8628 6808
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6368 6316 6420 6322
rect 6368 6258 6420 6264
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7840 6316 7892 6322
rect 7840 6258 7892 6264
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 5816 5636 5868 5642
rect 5816 5578 5868 5584
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5446 5128 5502 5137
rect 5446 5063 5502 5072
rect 5460 5030 5488 5063
rect 5448 5024 5500 5030
rect 5448 4966 5500 4972
rect 5828 4826 5856 5578
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6196 4826 6224 5306
rect 6380 5250 6408 5850
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6472 5370 6500 5510
rect 6548 5468 6856 5488
rect 6548 5466 6554 5468
rect 6610 5466 6634 5468
rect 6690 5466 6714 5468
rect 6770 5466 6794 5468
rect 6850 5466 6856 5468
rect 6610 5414 6612 5466
rect 6792 5414 6794 5466
rect 6548 5412 6554 5414
rect 6610 5412 6634 5414
rect 6690 5412 6714 5414
rect 6770 5412 6794 5414
rect 6850 5412 6856 5414
rect 6548 5392 6856 5412
rect 6460 5364 6512 5370
rect 6460 5306 6512 5312
rect 6288 5222 6408 5250
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 6184 4820 6236 4826
rect 6184 4762 6236 4768
rect 5354 4720 5410 4729
rect 5354 4655 5410 4664
rect 5368 4622 5396 4655
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 6184 4548 6236 4554
rect 6184 4490 6236 4496
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 6196 4010 6224 4490
rect 6288 4486 6316 5222
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6380 4690 6408 5102
rect 6368 4684 6420 4690
rect 6368 4626 6420 4632
rect 6472 4622 6500 5306
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 6920 5228 6972 5234
rect 6920 5170 6972 5176
rect 6932 4826 6960 5170
rect 7392 5098 7420 5238
rect 7380 5092 7432 5098
rect 7380 5034 7432 5040
rect 7104 5024 7156 5030
rect 7104 4966 7156 4972
rect 6552 4820 6604 4826
rect 6552 4762 6604 4768
rect 6920 4820 6972 4826
rect 6920 4762 6972 4768
rect 6564 4622 6592 4762
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6276 4480 6328 4486
rect 6276 4422 6328 4428
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6548 4380 6856 4400
rect 6548 4378 6554 4380
rect 6610 4378 6634 4380
rect 6690 4378 6714 4380
rect 6770 4378 6794 4380
rect 6850 4378 6856 4380
rect 6610 4326 6612 4378
rect 6792 4326 6794 4378
rect 6548 4324 6554 4326
rect 6610 4324 6634 4326
rect 6690 4324 6714 4326
rect 6770 4324 6794 4326
rect 6850 4324 6856 4326
rect 6548 4304 6856 4324
rect 7024 4282 7052 4422
rect 7012 4276 7064 4282
rect 7012 4218 7064 4224
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 5816 4004 5868 4010
rect 5816 3946 5868 3952
rect 6184 4004 6236 4010
rect 6184 3946 6236 3952
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 5080 3052 5132 3058
rect 5080 2994 5132 3000
rect 3749 2748 4057 2768
rect 3749 2746 3755 2748
rect 3811 2746 3835 2748
rect 3891 2746 3915 2748
rect 3971 2746 3995 2748
rect 4051 2746 4057 2748
rect 3811 2694 3813 2746
rect 3993 2694 3995 2746
rect 3749 2692 3755 2694
rect 3811 2692 3835 2694
rect 3891 2692 3915 2694
rect 3971 2692 3995 2694
rect 4051 2692 4057 2694
rect 3749 2672 4057 2692
rect 4816 2650 4844 2994
rect 4804 2644 4856 2650
rect 4804 2586 4856 2592
rect 5828 2514 5856 3946
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 5920 3194 5948 3402
rect 5908 3188 5960 3194
rect 5908 3130 5960 3136
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 5908 2576 5960 2582
rect 5906 2544 5908 2553
rect 5960 2544 5962 2553
rect 5816 2508 5868 2514
rect 5906 2479 5962 2488
rect 5816 2450 5868 2456
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 5356 2440 5408 2446
rect 6012 2394 6040 3130
rect 5356 2382 5408 2388
rect 3620 1902 3648 2382
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 3976 2304 4028 2310
rect 3976 2246 4028 2252
rect 3804 2106 3832 2246
rect 3792 2100 3844 2106
rect 3792 2042 3844 2048
rect 3608 1896 3660 1902
rect 3988 1873 4016 2246
rect 4632 1970 4660 2382
rect 5368 2009 5396 2382
rect 5828 2378 6040 2394
rect 6104 2378 6132 3878
rect 6932 3398 6960 3878
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 6460 3392 6512 3398
rect 6460 3334 6512 3340
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6196 3194 6224 3334
rect 6472 3194 6500 3334
rect 6548 3292 6856 3312
rect 6548 3290 6554 3292
rect 6610 3290 6634 3292
rect 6690 3290 6714 3292
rect 6770 3290 6794 3292
rect 6850 3290 6856 3292
rect 6610 3238 6612 3290
rect 6792 3238 6794 3290
rect 6548 3236 6554 3238
rect 6610 3236 6634 3238
rect 6690 3236 6714 3238
rect 6770 3236 6794 3238
rect 6850 3236 6856 3238
rect 6548 3216 6856 3236
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6368 2984 6420 2990
rect 6368 2926 6420 2932
rect 6276 2848 6328 2854
rect 6276 2790 6328 2796
rect 5816 2372 6040 2378
rect 5868 2366 6040 2372
rect 6092 2372 6144 2378
rect 5816 2314 5868 2320
rect 6092 2314 6144 2320
rect 5354 2000 5410 2009
rect 4620 1964 4672 1970
rect 5354 1935 5410 1944
rect 4620 1906 4672 1912
rect 3608 1838 3660 1844
rect 3974 1864 4030 1873
rect 3424 1828 3476 1834
rect 3974 1799 4030 1808
rect 3424 1770 3476 1776
rect 2962 1728 3018 1737
rect 2962 1663 3018 1672
rect 6288 1442 6316 2790
rect 6380 2514 6408 2926
rect 6828 2916 6880 2922
rect 6828 2858 6880 2864
rect 6840 2825 6868 2858
rect 6826 2816 6882 2825
rect 6826 2751 6882 2760
rect 7024 2650 7052 4014
rect 7116 3534 7144 4966
rect 7484 4826 7512 6258
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7760 5166 7788 6190
rect 7852 5370 7880 6258
rect 8036 5914 8064 6258
rect 8024 5908 8076 5914
rect 8024 5850 8076 5856
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 8312 5234 8340 6802
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8576 6656 8628 6662
rect 8576 6598 8628 6604
rect 8588 6322 8616 6598
rect 8576 6316 8628 6322
rect 8576 6258 8628 6264
rect 8392 6112 8444 6118
rect 8392 6054 8444 6060
rect 8404 5710 8432 6054
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7472 4820 7524 4826
rect 7472 4762 7524 4768
rect 7196 4548 7248 4554
rect 7196 4490 7248 4496
rect 7208 4146 7236 4490
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7288 4276 7340 4282
rect 7288 4218 7340 4224
rect 7300 4146 7328 4218
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7208 3670 7236 4082
rect 7196 3664 7248 3670
rect 7196 3606 7248 3612
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7196 3120 7248 3126
rect 7196 3062 7248 3068
rect 7012 2644 7064 2650
rect 7012 2586 7064 2592
rect 7104 2644 7156 2650
rect 7104 2586 7156 2592
rect 7116 2553 7144 2586
rect 7102 2544 7158 2553
rect 6368 2508 6420 2514
rect 7102 2479 7158 2488
rect 6368 2450 6420 2456
rect 7208 2394 7236 3062
rect 7392 2650 7420 4422
rect 7760 4146 7788 5102
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7852 4282 7880 4558
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 7840 4276 7892 4282
rect 7840 4218 7892 4224
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 8208 4072 8260 4078
rect 8208 4014 8260 4020
rect 8114 2952 8170 2961
rect 8114 2887 8170 2896
rect 7380 2644 7432 2650
rect 7380 2586 7432 2592
rect 6840 2378 7236 2394
rect 6828 2372 7236 2378
rect 6880 2366 7236 2372
rect 6828 2314 6880 2320
rect 6548 2204 6856 2224
rect 6548 2202 6554 2204
rect 6610 2202 6634 2204
rect 6690 2202 6714 2204
rect 6770 2202 6794 2204
rect 6850 2202 6856 2204
rect 6610 2150 6612 2202
rect 6792 2150 6794 2202
rect 6548 2148 6554 2150
rect 6610 2148 6634 2150
rect 6690 2148 6714 2150
rect 6770 2148 6794 2150
rect 6850 2148 6856 2150
rect 6548 2128 6856 2148
rect 7392 1902 7420 2586
rect 8128 2378 8156 2887
rect 8220 2650 8248 4014
rect 8404 4010 8432 4422
rect 8496 4146 8524 5714
rect 8680 5302 8708 6734
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 6390 9076 6598
rect 9232 6390 9260 7686
rect 9968 7342 9996 7890
rect 10152 7886 10180 8570
rect 10888 8430 10916 10202
rect 10980 9722 11008 10746
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11348 9926 11376 10610
rect 11336 9920 11388 9926
rect 11336 9862 11388 9868
rect 10968 9716 11020 9722
rect 10968 9658 11020 9664
rect 10980 9382 11008 9658
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 11060 8900 11112 8906
rect 11060 8842 11112 8848
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10692 8356 10744 8362
rect 10692 8298 10744 8304
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10598 7440 10654 7449
rect 10598 7375 10600 7384
rect 10652 7375 10654 7384
rect 10600 7346 10652 7352
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9347 7100 9655 7120
rect 9347 7098 9353 7100
rect 9409 7098 9433 7100
rect 9489 7098 9513 7100
rect 9569 7098 9593 7100
rect 9649 7098 9655 7100
rect 9409 7046 9411 7098
rect 9591 7046 9593 7098
rect 9347 7044 9353 7046
rect 9409 7044 9433 7046
rect 9489 7044 9513 7046
rect 9569 7044 9593 7046
rect 9649 7044 9655 7046
rect 9347 7024 9655 7044
rect 9968 6730 9996 7278
rect 10704 6914 10732 8298
rect 11072 7478 11100 8842
rect 11348 8498 11376 9862
rect 11440 9178 11468 12106
rect 11532 11830 11560 12174
rect 11520 11824 11572 11830
rect 11520 11766 11572 11772
rect 11532 11218 11560 11766
rect 11624 11626 11652 12854
rect 11612 11620 11664 11626
rect 11612 11562 11664 11568
rect 11520 11212 11572 11218
rect 11520 11154 11572 11160
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11532 9722 11560 10406
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 11336 7744 11388 7750
rect 11336 7686 11388 7692
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 11348 7410 11376 7686
rect 11532 7546 11560 9658
rect 11716 8362 11744 13126
rect 11808 12889 11836 14198
rect 11900 13326 11928 19774
rect 11992 19174 12020 19808
rect 12072 19790 12124 19796
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12072 19712 12124 19718
rect 12072 19654 12124 19660
rect 11980 19168 12032 19174
rect 11980 19110 12032 19116
rect 11978 18456 12034 18465
rect 11978 18391 12034 18400
rect 11992 18290 12020 18391
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 11992 15910 12020 18226
rect 12084 17678 12112 19654
rect 12146 19612 12454 19632
rect 12146 19610 12152 19612
rect 12208 19610 12232 19612
rect 12288 19610 12312 19612
rect 12368 19610 12392 19612
rect 12448 19610 12454 19612
rect 12208 19558 12210 19610
rect 12390 19558 12392 19610
rect 12146 19556 12152 19558
rect 12208 19556 12232 19558
rect 12288 19556 12312 19558
rect 12368 19556 12392 19558
rect 12448 19556 12454 19558
rect 12146 19536 12454 19556
rect 12440 19372 12492 19378
rect 12492 19332 12572 19360
rect 12440 19314 12492 19320
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12452 18698 12480 19110
rect 12440 18692 12492 18698
rect 12440 18634 12492 18640
rect 12544 18630 12572 19332
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12146 18524 12454 18544
rect 12146 18522 12152 18524
rect 12208 18522 12232 18524
rect 12288 18522 12312 18524
rect 12368 18522 12392 18524
rect 12448 18522 12454 18524
rect 12208 18470 12210 18522
rect 12390 18470 12392 18522
rect 12146 18468 12152 18470
rect 12208 18468 12232 18470
rect 12288 18468 12312 18470
rect 12368 18468 12392 18470
rect 12448 18468 12454 18470
rect 12146 18448 12454 18468
rect 12072 17672 12124 17678
rect 12072 17614 12124 17620
rect 12146 17436 12454 17456
rect 12146 17434 12152 17436
rect 12208 17434 12232 17436
rect 12288 17434 12312 17436
rect 12368 17434 12392 17436
rect 12448 17434 12454 17436
rect 12208 17382 12210 17434
rect 12390 17382 12392 17434
rect 12146 17380 12152 17382
rect 12208 17380 12232 17382
rect 12288 17380 12312 17382
rect 12368 17380 12392 17382
rect 12448 17380 12454 17382
rect 12146 17360 12454 17380
rect 12072 16516 12124 16522
rect 12072 16458 12124 16464
rect 12084 16250 12112 16458
rect 12146 16348 12454 16368
rect 12146 16346 12152 16348
rect 12208 16346 12232 16348
rect 12288 16346 12312 16348
rect 12368 16346 12392 16348
rect 12448 16346 12454 16348
rect 12208 16294 12210 16346
rect 12390 16294 12392 16346
rect 12146 16292 12152 16294
rect 12208 16292 12232 16294
rect 12288 16292 12312 16294
rect 12368 16292 12392 16294
rect 12448 16292 12454 16294
rect 12146 16272 12454 16292
rect 12072 16244 12124 16250
rect 12072 16186 12124 16192
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 12146 15260 12454 15280
rect 12146 15258 12152 15260
rect 12208 15258 12232 15260
rect 12288 15258 12312 15260
rect 12368 15258 12392 15260
rect 12448 15258 12454 15260
rect 12208 15206 12210 15258
rect 12390 15206 12392 15258
rect 12146 15204 12152 15206
rect 12208 15204 12232 15206
rect 12288 15204 12312 15206
rect 12368 15204 12392 15206
rect 12448 15204 12454 15206
rect 12146 15184 12454 15204
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11992 13462 12020 14962
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 12084 13530 12112 14350
rect 12146 14172 12454 14192
rect 12146 14170 12152 14172
rect 12208 14170 12232 14172
rect 12288 14170 12312 14172
rect 12368 14170 12392 14172
rect 12448 14170 12454 14172
rect 12208 14118 12210 14170
rect 12390 14118 12392 14170
rect 12146 14116 12152 14118
rect 12208 14116 12232 14118
rect 12288 14116 12312 14118
rect 12368 14116 12392 14118
rect 12448 14116 12454 14118
rect 12146 14096 12454 14116
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 11980 13456 12032 13462
rect 11980 13398 12032 13404
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 12084 12986 12112 13466
rect 12452 13326 12480 13670
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12146 13084 12454 13104
rect 12146 13082 12152 13084
rect 12208 13082 12232 13084
rect 12288 13082 12312 13084
rect 12368 13082 12392 13084
rect 12448 13082 12454 13084
rect 12208 13030 12210 13082
rect 12390 13030 12392 13082
rect 12146 13028 12152 13030
rect 12208 13028 12232 13030
rect 12288 13028 12312 13030
rect 12368 13028 12392 13030
rect 12448 13028 12454 13030
rect 12146 13008 12454 13028
rect 12544 12986 12572 18566
rect 12636 17814 12664 18702
rect 12820 18426 12848 19790
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 12808 18420 12860 18426
rect 12728 18380 12808 18408
rect 12728 17882 12756 18380
rect 12808 18362 12860 18368
rect 12912 18290 12940 18702
rect 12992 18624 13044 18630
rect 12992 18566 13044 18572
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 12912 17882 12940 18226
rect 12716 17876 12768 17882
rect 12716 17818 12768 17824
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12624 17808 12676 17814
rect 12624 17750 12676 17756
rect 13004 17270 13032 18566
rect 13096 18222 13124 19858
rect 13268 18692 13320 18698
rect 13268 18634 13320 18640
rect 13280 18222 13308 18634
rect 13372 18358 13400 21422
rect 13452 20528 13504 20534
rect 13452 20470 13504 20476
rect 13464 19378 13492 20470
rect 13556 20058 13584 21422
rect 13648 20602 13676 21898
rect 13832 21894 13860 23800
rect 13912 22024 13964 22030
rect 13912 21966 13964 21972
rect 13728 21888 13780 21894
rect 13728 21830 13780 21836
rect 13820 21888 13872 21894
rect 13820 21830 13872 21836
rect 13740 21486 13768 21830
rect 13728 21480 13780 21486
rect 13728 21422 13780 21428
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13820 21344 13872 21350
rect 13820 21286 13872 21292
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13648 19854 13676 20538
rect 13636 19848 13688 19854
rect 13636 19790 13688 19796
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13464 18834 13492 19314
rect 13452 18828 13504 18834
rect 13452 18770 13504 18776
rect 13360 18352 13412 18358
rect 13740 18306 13768 21286
rect 13832 20466 13860 21286
rect 13924 21078 13952 21966
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 14096 21548 14148 21554
rect 14096 21490 14148 21496
rect 14004 21140 14056 21146
rect 14004 21082 14056 21088
rect 13912 21072 13964 21078
rect 13912 21014 13964 21020
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 13924 20466 13952 20742
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 13912 20460 13964 20466
rect 13912 20402 13964 20408
rect 14016 19990 14044 21082
rect 14108 20058 14136 21490
rect 14200 21146 14228 21626
rect 14476 21457 14504 23800
rect 14660 21729 14688 23854
rect 15028 23746 15056 23854
rect 15106 23800 15162 24600
rect 15488 23854 15700 23882
rect 15120 23746 15148 23800
rect 15028 23718 15148 23746
rect 14945 22332 15253 22352
rect 14945 22330 14951 22332
rect 15007 22330 15031 22332
rect 15087 22330 15111 22332
rect 15167 22330 15191 22332
rect 15247 22330 15253 22332
rect 15007 22278 15009 22330
rect 15189 22278 15191 22330
rect 14945 22276 14951 22278
rect 15007 22276 15031 22278
rect 15087 22276 15111 22278
rect 15167 22276 15191 22278
rect 15247 22276 15253 22278
rect 14945 22256 15253 22276
rect 14740 21888 14792 21894
rect 14740 21830 14792 21836
rect 14832 21888 14884 21894
rect 14832 21830 14884 21836
rect 14646 21720 14702 21729
rect 14646 21655 14702 21664
rect 14462 21448 14518 21457
rect 14462 21383 14518 21392
rect 14188 21140 14240 21146
rect 14188 21082 14240 21088
rect 14096 20052 14148 20058
rect 14096 19994 14148 20000
rect 14004 19984 14056 19990
rect 14004 19926 14056 19932
rect 14094 19952 14150 19961
rect 14094 19887 14150 19896
rect 14108 19514 14136 19887
rect 14200 19854 14228 21082
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14188 19848 14240 19854
rect 14188 19790 14240 19796
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14096 19508 14148 19514
rect 14096 19450 14148 19456
rect 14004 19372 14056 19378
rect 14004 19314 14056 19320
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 13832 18970 13860 19246
rect 14016 18970 14044 19314
rect 14200 19122 14228 19654
rect 14292 19242 14320 20198
rect 14476 19802 14504 21383
rect 14556 20460 14608 20466
rect 14556 20402 14608 20408
rect 14568 19922 14596 20402
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14372 19780 14424 19786
rect 14476 19774 14596 19802
rect 14372 19722 14424 19728
rect 14384 19514 14412 19722
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14280 19236 14332 19242
rect 14280 19178 14332 19184
rect 14464 19168 14516 19174
rect 14200 19094 14320 19122
rect 14464 19110 14516 19116
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 14004 18964 14056 18970
rect 14004 18906 14056 18912
rect 14096 18760 14148 18766
rect 14096 18702 14148 18708
rect 13360 18294 13412 18300
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13268 18216 13320 18222
rect 13268 18158 13320 18164
rect 13268 18080 13320 18086
rect 13268 18022 13320 18028
rect 13280 17746 13308 18022
rect 13372 17814 13400 18294
rect 13648 18278 13768 18306
rect 14004 18284 14056 18290
rect 13544 18080 13596 18086
rect 13544 18022 13596 18028
rect 13360 17808 13412 17814
rect 13360 17750 13412 17756
rect 13268 17740 13320 17746
rect 13268 17682 13320 17688
rect 13360 17536 13412 17542
rect 13360 17478 13412 17484
rect 13372 17338 13400 17478
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 12992 17264 13044 17270
rect 12992 17206 13044 17212
rect 13556 16590 13584 18022
rect 13648 17785 13676 18278
rect 14004 18226 14056 18232
rect 13634 17776 13690 17785
rect 13634 17711 13690 17720
rect 14016 17338 14044 18226
rect 14108 17882 14136 18702
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14200 17882 14228 18022
rect 14096 17876 14148 17882
rect 14096 17818 14148 17824
rect 14188 17876 14240 17882
rect 14188 17818 14240 17824
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 13820 17196 13872 17202
rect 13820 17138 13872 17144
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 13832 16454 13860 17138
rect 13912 16992 13964 16998
rect 14016 16946 14044 17274
rect 13964 16940 14044 16946
rect 13912 16934 14044 16940
rect 13924 16918 14044 16934
rect 13820 16448 13872 16454
rect 13820 16390 13872 16396
rect 14096 16448 14148 16454
rect 14096 16390 14148 16396
rect 14108 16182 14136 16390
rect 14096 16176 14148 16182
rect 14096 16118 14148 16124
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13634 16008 13690 16017
rect 13634 15943 13690 15952
rect 13452 15904 13504 15910
rect 13452 15846 13504 15852
rect 13464 15706 13492 15846
rect 13648 15706 13676 15943
rect 13452 15700 13504 15706
rect 13636 15700 13688 15706
rect 13452 15642 13504 15648
rect 13556 15660 13636 15688
rect 12900 15020 12952 15026
rect 12900 14962 12952 14968
rect 12912 14618 12940 14962
rect 13556 14822 13584 15660
rect 13636 15642 13688 15648
rect 13832 15570 13860 16050
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13636 15496 13688 15502
rect 13636 15438 13688 15444
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 12624 14408 12676 14414
rect 12624 14350 12676 14356
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12532 12980 12584 12986
rect 12532 12922 12584 12928
rect 11794 12880 11850 12889
rect 11794 12815 11850 12824
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 12072 12776 12124 12782
rect 12072 12718 12124 12724
rect 11992 12442 12020 12718
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 12084 12322 12112 12718
rect 12636 12714 12664 14350
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12820 13258 12848 14214
rect 12912 13734 12940 14350
rect 12900 13728 12952 13734
rect 12900 13670 12952 13676
rect 12808 13252 12860 13258
rect 12808 13194 12860 13200
rect 12624 12708 12676 12714
rect 12624 12650 12676 12656
rect 11992 12294 12112 12322
rect 11992 11762 12020 12294
rect 12146 11996 12454 12016
rect 12146 11994 12152 11996
rect 12208 11994 12232 11996
rect 12288 11994 12312 11996
rect 12368 11994 12392 11996
rect 12448 11994 12454 11996
rect 12208 11942 12210 11994
rect 12390 11942 12392 11994
rect 12146 11940 12152 11942
rect 12208 11940 12232 11942
rect 12288 11940 12312 11942
rect 12368 11940 12392 11942
rect 12448 11940 12454 11942
rect 12146 11920 12454 11940
rect 12072 11892 12124 11898
rect 12072 11834 12124 11840
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 12084 11150 12112 11834
rect 13544 11688 13596 11694
rect 13544 11630 13596 11636
rect 12072 11144 12124 11150
rect 12072 11086 12124 11092
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 13360 11008 13412 11014
rect 13360 10950 13412 10956
rect 11980 10804 12032 10810
rect 11980 10746 12032 10752
rect 11794 10568 11850 10577
rect 11794 10503 11850 10512
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11520 7540 11572 7546
rect 11520 7482 11572 7488
rect 11336 7404 11388 7410
rect 11336 7346 11388 7352
rect 10612 6886 10732 6914
rect 10230 6760 10286 6769
rect 9956 6724 10008 6730
rect 10230 6695 10286 6704
rect 10416 6724 10468 6730
rect 9956 6666 10008 6672
rect 9036 6384 9088 6390
rect 9036 6326 9088 6332
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 8864 4622 8892 5306
rect 9232 5166 9260 6326
rect 9968 6322 9996 6666
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9347 6012 9655 6032
rect 9347 6010 9353 6012
rect 9409 6010 9433 6012
rect 9489 6010 9513 6012
rect 9569 6010 9593 6012
rect 9649 6010 9655 6012
rect 9409 5958 9411 6010
rect 9591 5958 9593 6010
rect 9347 5956 9353 5958
rect 9409 5956 9433 5958
rect 9489 5956 9513 5958
rect 9569 5956 9593 5958
rect 9649 5956 9655 5958
rect 9347 5936 9655 5956
rect 9680 5296 9732 5302
rect 9680 5238 9732 5244
rect 9220 5160 9272 5166
rect 9220 5102 9272 5108
rect 9347 4924 9655 4944
rect 9347 4922 9353 4924
rect 9409 4922 9433 4924
rect 9489 4922 9513 4924
rect 9569 4922 9593 4924
rect 9649 4922 9655 4924
rect 9409 4870 9411 4922
rect 9591 4870 9593 4922
rect 9347 4868 9353 4870
rect 9409 4868 9433 4870
rect 9489 4868 9513 4870
rect 9569 4868 9593 4870
rect 9649 4868 9655 4870
rect 9347 4848 9655 4868
rect 8852 4616 8904 4622
rect 8852 4558 8904 4564
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8392 4004 8444 4010
rect 8392 3946 8444 3952
rect 8496 3534 8524 4082
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8404 3058 8432 3334
rect 8956 3126 8984 4218
rect 9036 4208 9088 4214
rect 9036 4150 9088 4156
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 8300 2848 8352 2854
rect 8298 2816 8300 2825
rect 8352 2816 8354 2825
rect 8298 2751 8354 2760
rect 8208 2644 8260 2650
rect 8208 2586 8260 2592
rect 8312 2514 8340 2751
rect 8300 2508 8352 2514
rect 8300 2450 8352 2456
rect 8404 2446 8432 2994
rect 9048 2650 9076 4150
rect 9232 3534 9260 4558
rect 9347 3836 9655 3856
rect 9347 3834 9353 3836
rect 9409 3834 9433 3836
rect 9489 3834 9513 3836
rect 9569 3834 9593 3836
rect 9649 3834 9655 3836
rect 9409 3782 9411 3834
rect 9591 3782 9593 3834
rect 9347 3780 9353 3782
rect 9409 3780 9433 3782
rect 9489 3780 9513 3782
rect 9569 3780 9593 3782
rect 9649 3780 9655 3782
rect 9347 3760 9655 3780
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9692 3466 9720 5238
rect 9784 4622 9812 6122
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9876 4826 9904 6054
rect 9864 4820 9916 4826
rect 9916 4780 9996 4808
rect 9864 4762 9916 4768
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9864 3936 9916 3942
rect 9864 3878 9916 3884
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9128 2984 9180 2990
rect 9126 2952 9128 2961
rect 9180 2952 9182 2961
rect 9126 2887 9182 2896
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9347 2748 9655 2768
rect 9347 2746 9353 2748
rect 9409 2746 9433 2748
rect 9489 2746 9513 2748
rect 9569 2746 9593 2748
rect 9649 2746 9655 2748
rect 9409 2694 9411 2746
rect 9591 2694 9593 2746
rect 9347 2692 9353 2694
rect 9409 2692 9433 2694
rect 9489 2692 9513 2694
rect 9569 2692 9593 2694
rect 9649 2692 9655 2694
rect 9347 2672 9655 2692
rect 9036 2644 9088 2650
rect 9036 2586 9088 2592
rect 9692 2446 9720 2790
rect 9876 2514 9904 3878
rect 9968 2650 9996 4780
rect 10244 4758 10272 6695
rect 10416 6666 10468 6672
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10336 5234 10364 5714
rect 10324 5228 10376 5234
rect 10324 5170 10376 5176
rect 10428 4826 10456 6666
rect 10508 5160 10560 5166
rect 10508 5102 10560 5108
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10232 4752 10284 4758
rect 10232 4694 10284 4700
rect 10520 4690 10548 5102
rect 10612 4826 10640 6886
rect 10966 6352 11022 6361
rect 10966 6287 10968 6296
rect 11020 6287 11022 6296
rect 10968 6258 11020 6264
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10704 5370 10732 5510
rect 10692 5364 10744 5370
rect 10692 5306 10744 5312
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 10600 4820 10652 4826
rect 10600 4762 10652 4768
rect 10508 4684 10560 4690
rect 10508 4626 10560 4632
rect 10520 4010 10548 4626
rect 10612 4146 10640 4762
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10508 4004 10560 4010
rect 10508 3946 10560 3952
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10612 3058 10640 3470
rect 10888 3398 10916 4014
rect 11072 3670 11100 4490
rect 11348 4486 11376 5170
rect 11428 5024 11480 5030
rect 11428 4966 11480 4972
rect 11440 4486 11468 4966
rect 11808 4826 11836 10503
rect 11992 10266 12020 10746
rect 12084 10674 12112 10950
rect 12146 10908 12454 10928
rect 12146 10906 12152 10908
rect 12208 10906 12232 10908
rect 12288 10906 12312 10908
rect 12368 10906 12392 10908
rect 12448 10906 12454 10908
rect 12208 10854 12210 10906
rect 12390 10854 12392 10906
rect 12146 10852 12152 10854
rect 12208 10852 12232 10854
rect 12288 10852 12312 10854
rect 12368 10852 12392 10854
rect 12448 10852 12454 10854
rect 12146 10832 12454 10852
rect 12072 10668 12124 10674
rect 12072 10610 12124 10616
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11992 9586 12020 10202
rect 12146 9820 12454 9840
rect 12146 9818 12152 9820
rect 12208 9818 12232 9820
rect 12288 9818 12312 9820
rect 12368 9818 12392 9820
rect 12448 9818 12454 9820
rect 12208 9766 12210 9818
rect 12390 9766 12392 9818
rect 12146 9764 12152 9766
rect 12208 9764 12232 9766
rect 12288 9764 12312 9766
rect 12368 9764 12392 9766
rect 12448 9764 12454 9766
rect 12146 9744 12454 9764
rect 12728 9654 12756 10610
rect 13372 10062 13400 10950
rect 13556 10538 13584 11630
rect 13648 11257 13676 15438
rect 13832 15026 13860 15506
rect 14096 15088 14148 15094
rect 14096 15030 14148 15036
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 13728 14272 13780 14278
rect 13728 14214 13780 14220
rect 13740 13938 13768 14214
rect 13832 14006 13860 14962
rect 14004 14816 14056 14822
rect 14004 14758 14056 14764
rect 13912 14340 13964 14346
rect 13912 14282 13964 14288
rect 13820 14000 13872 14006
rect 13820 13942 13872 13948
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13832 13326 13860 13942
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13832 12850 13860 13262
rect 13820 12844 13872 12850
rect 13820 12786 13872 12792
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13634 11248 13690 11257
rect 13634 11183 13690 11192
rect 13740 11150 13768 11494
rect 13832 11354 13860 11698
rect 13924 11354 13952 14282
rect 14016 13841 14044 14758
rect 14108 14074 14136 15030
rect 14188 14884 14240 14890
rect 14188 14826 14240 14832
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14002 13832 14058 13841
rect 14002 13767 14058 13776
rect 14004 12776 14056 12782
rect 14004 12718 14056 12724
rect 14016 11830 14044 12718
rect 14108 12306 14136 14010
rect 14200 12782 14228 14826
rect 14188 12776 14240 12782
rect 14188 12718 14240 12724
rect 14096 12300 14148 12306
rect 14096 12242 14148 12248
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 13820 11348 13872 11354
rect 13820 11290 13872 11296
rect 13912 11348 13964 11354
rect 13912 11290 13964 11296
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13636 11076 13688 11082
rect 13636 11018 13688 11024
rect 13544 10532 13596 10538
rect 13544 10474 13596 10480
rect 13648 10266 13676 11018
rect 13832 10674 13860 11290
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13924 10742 13952 11154
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 12716 9648 12768 9654
rect 12716 9590 12768 9596
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 12898 9480 12954 9489
rect 12898 9415 12954 9424
rect 11980 8968 12032 8974
rect 11886 8936 11942 8945
rect 11980 8910 12032 8916
rect 11886 8871 11942 8880
rect 11900 7546 11928 8871
rect 11992 8498 12020 8910
rect 12146 8732 12454 8752
rect 12146 8730 12152 8732
rect 12208 8730 12232 8732
rect 12288 8730 12312 8732
rect 12368 8730 12392 8732
rect 12448 8730 12454 8732
rect 12208 8678 12210 8730
rect 12390 8678 12392 8730
rect 12146 8676 12152 8678
rect 12208 8676 12232 8678
rect 12288 8676 12312 8678
rect 12368 8676 12392 8678
rect 12448 8676 12454 8678
rect 12146 8656 12454 8676
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 11980 7812 12032 7818
rect 11980 7754 12032 7760
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 11900 6798 11928 7482
rect 11888 6792 11940 6798
rect 11888 6734 11940 6740
rect 11992 6662 12020 7754
rect 12084 6866 12112 8434
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12146 7644 12454 7664
rect 12146 7642 12152 7644
rect 12208 7642 12232 7644
rect 12288 7642 12312 7644
rect 12368 7642 12392 7644
rect 12448 7642 12454 7644
rect 12208 7590 12210 7642
rect 12390 7590 12392 7642
rect 12146 7588 12152 7590
rect 12208 7588 12232 7590
rect 12288 7588 12312 7590
rect 12368 7588 12392 7590
rect 12448 7588 12454 7590
rect 12146 7568 12454 7588
rect 12164 7336 12216 7342
rect 12164 7278 12216 7284
rect 12176 7002 12204 7278
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12072 6860 12124 6866
rect 12072 6802 12124 6808
rect 12176 6798 12204 6938
rect 12728 6798 12756 7686
rect 12808 7336 12860 7342
rect 12808 7278 12860 7284
rect 12164 6792 12216 6798
rect 12164 6734 12216 6740
rect 12716 6792 12768 6798
rect 12716 6734 12768 6740
rect 11980 6656 12032 6662
rect 11980 6598 12032 6604
rect 12146 6556 12454 6576
rect 12146 6554 12152 6556
rect 12208 6554 12232 6556
rect 12288 6554 12312 6556
rect 12368 6554 12392 6556
rect 12448 6554 12454 6556
rect 12208 6502 12210 6554
rect 12390 6502 12392 6554
rect 12146 6500 12152 6502
rect 12208 6500 12232 6502
rect 12288 6500 12312 6502
rect 12368 6500 12392 6502
rect 12448 6500 12454 6502
rect 12146 6480 12454 6500
rect 12072 6384 12124 6390
rect 12072 6326 12124 6332
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11900 5778 11928 6054
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11992 5370 12020 6190
rect 12084 5574 12112 6326
rect 12820 6322 12848 7278
rect 12808 6316 12860 6322
rect 12808 6258 12860 6264
rect 12820 5914 12848 6258
rect 12808 5908 12860 5914
rect 12808 5850 12860 5856
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12072 5568 12124 5574
rect 12072 5510 12124 5516
rect 12146 5468 12454 5488
rect 12146 5466 12152 5468
rect 12208 5466 12232 5468
rect 12288 5466 12312 5468
rect 12368 5466 12392 5468
rect 12448 5466 12454 5468
rect 12208 5414 12210 5466
rect 12390 5414 12392 5466
rect 12146 5412 12152 5414
rect 12208 5412 12232 5414
rect 12288 5412 12312 5414
rect 12368 5412 12392 5414
rect 12448 5412 12454 5414
rect 12146 5392 12454 5412
rect 12636 5370 12664 5646
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12808 5296 12860 5302
rect 12808 5238 12860 5244
rect 12624 5160 12676 5166
rect 12676 5120 12756 5148
rect 12624 5102 12676 5108
rect 11796 4820 11848 4826
rect 11796 4762 11848 4768
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 11440 4214 11468 4422
rect 12146 4380 12454 4400
rect 12146 4378 12152 4380
rect 12208 4378 12232 4380
rect 12288 4378 12312 4380
rect 12368 4378 12392 4380
rect 12448 4378 12454 4380
rect 12208 4326 12210 4378
rect 12390 4326 12392 4378
rect 12146 4324 12152 4326
rect 12208 4324 12232 4326
rect 12288 4324 12312 4326
rect 12368 4324 12392 4326
rect 12448 4324 12454 4326
rect 12146 4304 12454 4324
rect 11428 4208 11480 4214
rect 11428 4150 11480 4156
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 10876 3392 10928 3398
rect 10876 3334 10928 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 10980 3194 11008 3334
rect 10968 3188 11020 3194
rect 10968 3130 11020 3136
rect 11072 3058 11100 3606
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 10336 2650 10364 2994
rect 11164 2650 11192 3402
rect 9956 2644 10008 2650
rect 9956 2586 10008 2592
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 11152 2644 11204 2650
rect 11152 2586 11204 2592
rect 9968 2514 9996 2586
rect 11256 2582 11284 3878
rect 11348 3194 11376 4082
rect 12544 4026 12572 4558
rect 12624 4480 12676 4486
rect 12624 4422 12676 4428
rect 12452 3998 12572 4026
rect 11520 3936 11572 3942
rect 11520 3878 11572 3884
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11532 3058 11560 3878
rect 12452 3670 12480 3998
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 12072 3664 12124 3670
rect 11992 3624 12072 3652
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 10232 2576 10284 2582
rect 10232 2518 10284 2524
rect 11244 2576 11296 2582
rect 11244 2518 11296 2524
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 9956 2508 10008 2514
rect 9956 2450 10008 2456
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 8116 2372 8168 2378
rect 8116 2314 8168 2320
rect 8220 2038 8248 2382
rect 9128 2372 9180 2378
rect 9128 2314 9180 2320
rect 8208 2032 8260 2038
rect 8208 1974 8260 1980
rect 7932 1964 7984 1970
rect 7932 1906 7984 1912
rect 7380 1896 7432 1902
rect 7380 1838 7432 1844
rect 7944 1630 7972 1906
rect 9140 1834 9168 2314
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9324 2106 9352 2246
rect 9312 2100 9364 2106
rect 9312 2042 9364 2048
rect 9128 1828 9180 1834
rect 9128 1770 9180 1776
rect 7932 1624 7984 1630
rect 7932 1566 7984 1572
rect 6104 1414 6316 1442
rect 6104 800 6132 1414
rect 10244 800 10272 2518
rect 11704 2508 11756 2514
rect 11992 2496 12020 3624
rect 12072 3606 12124 3612
rect 12440 3664 12492 3670
rect 12440 3606 12492 3612
rect 12544 3534 12572 3878
rect 12532 3528 12584 3534
rect 12532 3470 12584 3476
rect 12072 3460 12124 3466
rect 12072 3402 12124 3408
rect 12084 3194 12112 3402
rect 12146 3292 12454 3312
rect 12146 3290 12152 3292
rect 12208 3290 12232 3292
rect 12288 3290 12312 3292
rect 12368 3290 12392 3292
rect 12448 3290 12454 3292
rect 12208 3238 12210 3290
rect 12390 3238 12392 3290
rect 12146 3236 12152 3238
rect 12208 3236 12232 3238
rect 12288 3236 12312 3238
rect 12368 3236 12392 3238
rect 12448 3236 12454 3238
rect 12146 3216 12454 3236
rect 12544 3194 12572 3470
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 12636 3126 12664 4422
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 12072 2508 12124 2514
rect 11992 2468 12072 2496
rect 11704 2450 11756 2456
rect 12072 2450 12124 2456
rect 11716 2378 11744 2450
rect 12728 2446 12756 5120
rect 12820 4282 12848 5238
rect 12808 4276 12860 4282
rect 12808 4218 12860 4224
rect 12716 2440 12768 2446
rect 12716 2382 12768 2388
rect 11704 2372 11756 2378
rect 11704 2314 11756 2320
rect 12912 2310 12940 9415
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 13004 7546 13032 8774
rect 13096 8090 13124 8774
rect 13280 8634 13308 9522
rect 13372 8956 13400 9998
rect 13464 9178 13492 9998
rect 13924 9926 13952 10542
rect 14016 10538 14044 11766
rect 14004 10532 14056 10538
rect 14004 10474 14056 10480
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 13912 9920 13964 9926
rect 13912 9862 13964 9868
rect 13542 9752 13598 9761
rect 13542 9687 13598 9696
rect 13452 9172 13504 9178
rect 13452 9114 13504 9120
rect 13452 8968 13504 8974
rect 13372 8928 13452 8956
rect 13452 8910 13504 8916
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13464 8498 13492 8910
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 13464 7954 13492 8434
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 13004 5778 13032 7142
rect 13176 6724 13228 6730
rect 13176 6666 13228 6672
rect 13188 6610 13216 6666
rect 13096 6582 13216 6610
rect 13096 6458 13124 6582
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 13188 6254 13216 6394
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13268 6248 13320 6254
rect 13452 6248 13504 6254
rect 13268 6190 13320 6196
rect 13372 6208 13452 6236
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 13004 5302 13032 5714
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 13280 5030 13308 6190
rect 13372 5574 13400 6208
rect 13452 6190 13504 6196
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13268 5024 13320 5030
rect 13268 4966 13320 4972
rect 13372 4146 13400 5510
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 13464 4554 13492 4966
rect 13452 4548 13504 4554
rect 13452 4490 13504 4496
rect 13452 4276 13504 4282
rect 13452 4218 13504 4224
rect 13360 4140 13412 4146
rect 13360 4082 13412 4088
rect 13464 2650 13492 4218
rect 13556 2961 13584 9687
rect 14016 9450 14044 9998
rect 14108 9654 14136 12242
rect 14292 11642 14320 19094
rect 14372 18896 14424 18902
rect 14372 18838 14424 18844
rect 14384 18465 14412 18838
rect 14370 18456 14426 18465
rect 14476 18426 14504 19110
rect 14370 18391 14426 18400
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14568 18306 14596 19774
rect 14476 18278 14596 18306
rect 14372 17808 14424 17814
rect 14372 17750 14424 17756
rect 14384 17202 14412 17750
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14476 15434 14504 18278
rect 14660 17898 14688 21655
rect 14752 20942 14780 21830
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 14740 20392 14792 20398
rect 14844 20369 14872 21830
rect 15384 21344 15436 21350
rect 15488 21321 15516 23854
rect 15672 23746 15700 23854
rect 15750 23800 15806 24600
rect 16394 23800 16450 24600
rect 17038 23800 17094 24600
rect 17682 23800 17738 24600
rect 18326 23800 18382 24600
rect 18970 23800 19026 24600
rect 19614 23800 19670 24600
rect 20258 23800 20314 24600
rect 20902 23800 20958 24600
rect 21008 23854 21220 23882
rect 15764 23746 15792 23800
rect 15672 23718 15792 23746
rect 15660 22024 15712 22030
rect 16304 22024 16356 22030
rect 15712 21984 15976 22012
rect 15660 21966 15712 21972
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 15568 21480 15620 21486
rect 15568 21422 15620 21428
rect 15384 21286 15436 21292
rect 15474 21312 15530 21321
rect 14945 21244 15253 21264
rect 14945 21242 14951 21244
rect 15007 21242 15031 21244
rect 15087 21242 15111 21244
rect 15167 21242 15191 21244
rect 15247 21242 15253 21244
rect 15007 21190 15009 21242
rect 15189 21190 15191 21242
rect 14945 21188 14951 21190
rect 15007 21188 15031 21190
rect 15087 21188 15111 21190
rect 15167 21188 15191 21190
rect 15247 21188 15253 21190
rect 14945 21168 15253 21188
rect 15396 20942 15424 21286
rect 15474 21247 15530 21256
rect 15384 20936 15436 20942
rect 14922 20904 14978 20913
rect 15384 20878 15436 20884
rect 14922 20839 14978 20848
rect 14740 20334 14792 20340
rect 14830 20360 14886 20369
rect 14568 17870 14688 17898
rect 14568 17814 14596 17870
rect 14556 17808 14608 17814
rect 14556 17750 14608 17756
rect 14752 17542 14780 20334
rect 14830 20295 14886 20304
rect 14936 20244 14964 20839
rect 15488 20754 15516 21247
rect 15580 21010 15608 21422
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15568 21004 15620 21010
rect 15568 20946 15620 20952
rect 15660 20868 15712 20874
rect 15660 20810 15712 20816
rect 15396 20726 15516 20754
rect 15292 20324 15344 20330
rect 15292 20266 15344 20272
rect 14844 20216 14964 20244
rect 14844 20058 14872 20216
rect 14945 20156 15253 20176
rect 14945 20154 14951 20156
rect 15007 20154 15031 20156
rect 15087 20154 15111 20156
rect 15167 20154 15191 20156
rect 15247 20154 15253 20156
rect 15007 20102 15009 20154
rect 15189 20102 15191 20154
rect 14945 20100 14951 20102
rect 15007 20100 15031 20102
rect 15087 20100 15111 20102
rect 15167 20100 15191 20102
rect 15247 20100 15253 20102
rect 14945 20080 15253 20100
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 15016 19916 15068 19922
rect 15016 19858 15068 19864
rect 15028 19394 15056 19858
rect 15200 19508 15252 19514
rect 15200 19450 15252 19456
rect 15212 19394 15240 19450
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 15028 19366 15240 19394
rect 14844 19242 14872 19314
rect 15028 19310 15056 19366
rect 15016 19304 15068 19310
rect 15016 19246 15068 19252
rect 14832 19236 14884 19242
rect 14832 19178 14884 19184
rect 14844 18970 14872 19178
rect 15304 19174 15332 20266
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 14945 19068 15253 19088
rect 14945 19066 14951 19068
rect 15007 19066 15031 19068
rect 15087 19066 15111 19068
rect 15167 19066 15191 19068
rect 15247 19066 15253 19068
rect 15007 19014 15009 19066
rect 15189 19014 15191 19066
rect 14945 19012 14951 19014
rect 15007 19012 15031 19014
rect 15087 19012 15111 19014
rect 15167 19012 15191 19014
rect 15247 19012 15253 19014
rect 14945 18992 15253 19012
rect 14832 18964 14884 18970
rect 14832 18906 14884 18912
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 14844 17746 14872 18022
rect 14945 17980 15253 18000
rect 14945 17978 14951 17980
rect 15007 17978 15031 17980
rect 15087 17978 15111 17980
rect 15167 17978 15191 17980
rect 15247 17978 15253 17980
rect 15007 17926 15009 17978
rect 15189 17926 15191 17978
rect 14945 17924 14951 17926
rect 15007 17924 15031 17926
rect 15087 17924 15111 17926
rect 15167 17924 15191 17926
rect 15247 17924 15253 17926
rect 14945 17904 15253 17924
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 14832 17604 14884 17610
rect 14832 17546 14884 17552
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14740 17536 14792 17542
rect 14740 17478 14792 17484
rect 14568 17338 14596 17478
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 14568 16590 14596 17070
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14568 16250 14596 16526
rect 14660 16250 14688 17138
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14648 16244 14700 16250
rect 14648 16186 14700 16192
rect 14464 15428 14516 15434
rect 14464 15370 14516 15376
rect 14844 15094 14872 17546
rect 15212 17202 15240 17614
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 14945 16892 15253 16912
rect 14945 16890 14951 16892
rect 15007 16890 15031 16892
rect 15087 16890 15111 16892
rect 15167 16890 15191 16892
rect 15247 16890 15253 16892
rect 15007 16838 15009 16890
rect 15189 16838 15191 16890
rect 14945 16836 14951 16838
rect 15007 16836 15031 16838
rect 15087 16836 15111 16838
rect 15167 16836 15191 16838
rect 15247 16836 15253 16838
rect 14945 16816 15253 16836
rect 15396 15910 15424 20726
rect 15672 20602 15700 20810
rect 15660 20596 15712 20602
rect 15660 20538 15712 20544
rect 15764 20534 15792 21286
rect 15856 20942 15884 21830
rect 15948 21554 15976 21984
rect 16304 21966 16356 21972
rect 16118 21720 16174 21729
rect 16118 21655 16174 21664
rect 15936 21548 15988 21554
rect 15936 21490 15988 21496
rect 16132 21457 16160 21655
rect 15934 21448 15990 21457
rect 15934 21383 15990 21392
rect 16118 21448 16174 21457
rect 16118 21383 16174 21392
rect 15948 21350 15976 21383
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 15844 20936 15896 20942
rect 15844 20878 15896 20884
rect 16210 20632 16266 20641
rect 16210 20567 16266 20576
rect 15752 20528 15804 20534
rect 15752 20470 15804 20476
rect 15936 20392 15988 20398
rect 15936 20334 15988 20340
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15672 19378 15700 19790
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15672 18970 15700 19314
rect 15948 18970 15976 20334
rect 16224 19310 16252 20567
rect 16316 20534 16344 21966
rect 16580 21956 16632 21962
rect 16580 21898 16632 21904
rect 16396 21888 16448 21894
rect 16396 21830 16448 21836
rect 16408 20806 16436 21830
rect 16592 21690 16620 21898
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16948 21888 17000 21894
rect 16948 21830 17000 21836
rect 16580 21684 16632 21690
rect 16580 21626 16632 21632
rect 16396 20800 16448 20806
rect 16396 20742 16448 20748
rect 16304 20528 16356 20534
rect 16304 20470 16356 20476
rect 16684 20346 16712 21830
rect 16960 21622 16988 21830
rect 16948 21616 17000 21622
rect 16948 21558 17000 21564
rect 17052 21049 17080 23800
rect 17696 22234 17724 23800
rect 17684 22228 17736 22234
rect 17684 22170 17736 22176
rect 17224 22024 17276 22030
rect 17684 22024 17736 22030
rect 17224 21966 17276 21972
rect 17604 21984 17684 22012
rect 17038 21040 17094 21049
rect 17236 21010 17264 21966
rect 17604 21593 17632 21984
rect 17684 21966 17736 21972
rect 18144 22024 18196 22030
rect 18144 21966 18196 21972
rect 17744 21788 18052 21808
rect 17744 21786 17750 21788
rect 17806 21786 17830 21788
rect 17886 21786 17910 21788
rect 17966 21786 17990 21788
rect 18046 21786 18052 21788
rect 17806 21734 17808 21786
rect 17988 21734 17990 21786
rect 17744 21732 17750 21734
rect 17806 21732 17830 21734
rect 17886 21732 17910 21734
rect 17966 21732 17990 21734
rect 18046 21732 18052 21734
rect 17744 21712 18052 21732
rect 18156 21690 18184 21966
rect 18144 21684 18196 21690
rect 18064 21644 18144 21672
rect 17590 21584 17646 21593
rect 17590 21519 17646 21528
rect 18064 21010 18092 21644
rect 18144 21626 18196 21632
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 17038 20975 17094 20984
rect 17224 21004 17276 21010
rect 17224 20946 17276 20952
rect 18052 21004 18104 21010
rect 18052 20946 18104 20952
rect 17316 20800 17368 20806
rect 17316 20742 17368 20748
rect 17408 20800 17460 20806
rect 17408 20742 17460 20748
rect 16316 20318 16712 20346
rect 16868 20590 17264 20618
rect 16316 20262 16344 20318
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16488 20256 16540 20262
rect 16488 20198 16540 20204
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 16212 19168 16264 19174
rect 16212 19110 16264 19116
rect 15660 18964 15712 18970
rect 15660 18906 15712 18912
rect 15936 18964 15988 18970
rect 15936 18906 15988 18912
rect 15476 18760 15528 18766
rect 15476 18702 15528 18708
rect 15488 18358 15516 18702
rect 15476 18352 15528 18358
rect 15476 18294 15528 18300
rect 15488 17746 15516 18294
rect 16224 17746 16252 19110
rect 16316 18698 16344 19654
rect 16304 18692 16356 18698
rect 16304 18634 16356 18640
rect 15476 17740 15528 17746
rect 15476 17682 15528 17688
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 15488 17270 15516 17682
rect 16026 17640 16082 17649
rect 16026 17575 16082 17584
rect 15476 17264 15528 17270
rect 15476 17206 15528 17212
rect 15488 16794 15516 17206
rect 15476 16788 15528 16794
rect 15476 16730 15528 16736
rect 15752 16516 15804 16522
rect 15752 16458 15804 16464
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 14945 15804 15253 15824
rect 14945 15802 14951 15804
rect 15007 15802 15031 15804
rect 15087 15802 15111 15804
rect 15167 15802 15191 15804
rect 15247 15802 15253 15804
rect 15007 15750 15009 15802
rect 15189 15750 15191 15802
rect 14945 15748 14951 15750
rect 15007 15748 15031 15750
rect 15087 15748 15111 15750
rect 15167 15748 15191 15750
rect 15247 15748 15253 15750
rect 14945 15728 15253 15748
rect 15764 15706 15792 16458
rect 15844 15904 15896 15910
rect 15844 15846 15896 15852
rect 15752 15700 15804 15706
rect 15752 15642 15804 15648
rect 15856 15502 15884 15846
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 14832 15088 14884 15094
rect 14832 15030 14884 15036
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14844 14482 14872 14894
rect 14945 14716 15253 14736
rect 14945 14714 14951 14716
rect 15007 14714 15031 14716
rect 15087 14714 15111 14716
rect 15167 14714 15191 14716
rect 15247 14714 15253 14716
rect 15007 14662 15009 14714
rect 15189 14662 15191 14714
rect 14945 14660 14951 14662
rect 15007 14660 15031 14662
rect 15087 14660 15111 14662
rect 15167 14660 15191 14662
rect 15247 14660 15253 14662
rect 14945 14640 15253 14660
rect 14832 14476 14884 14482
rect 14832 14418 14884 14424
rect 14740 14408 14792 14414
rect 14740 14350 14792 14356
rect 14464 14340 14516 14346
rect 14464 14282 14516 14288
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14384 12918 14412 13466
rect 14372 12912 14424 12918
rect 14372 12854 14424 12860
rect 14372 12640 14424 12646
rect 14372 12582 14424 12588
rect 14384 12306 14412 12582
rect 14372 12300 14424 12306
rect 14372 12242 14424 12248
rect 14476 12102 14504 14282
rect 14752 13530 14780 14350
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 13938 14964 14214
rect 14924 13932 14976 13938
rect 14924 13874 14976 13880
rect 15396 13734 15424 14962
rect 15580 14929 15608 15302
rect 15566 14920 15622 14929
rect 15566 14855 15622 14864
rect 15934 14920 15990 14929
rect 15934 14855 15990 14864
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15844 14816 15896 14822
rect 15844 14758 15896 14764
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15488 14074 15516 14350
rect 15476 14068 15528 14074
rect 15476 14010 15528 14016
rect 15384 13728 15436 13734
rect 15384 13670 15436 13676
rect 14945 13628 15253 13648
rect 14945 13626 14951 13628
rect 15007 13626 15031 13628
rect 15087 13626 15111 13628
rect 15167 13626 15191 13628
rect 15247 13626 15253 13628
rect 15007 13574 15009 13626
rect 15189 13574 15191 13626
rect 14945 13572 14951 13574
rect 15007 13572 15031 13574
rect 15087 13572 15111 13574
rect 15167 13572 15191 13574
rect 15247 13572 15253 13574
rect 14945 13552 15253 13572
rect 14740 13524 14792 13530
rect 14740 13466 14792 13472
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14292 11614 14504 11642
rect 14188 11348 14240 11354
rect 14188 11290 14240 11296
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 14004 9444 14056 9450
rect 14004 9386 14056 9392
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13648 7954 13676 8774
rect 13924 8566 13952 9318
rect 14108 9178 14136 9590
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 13912 8560 13964 8566
rect 13912 8502 13964 8508
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 13832 7274 13860 7890
rect 13820 7268 13872 7274
rect 13820 7210 13872 7216
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13648 6322 13676 6734
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13634 6216 13690 6225
rect 13634 6151 13690 6160
rect 13648 6118 13676 6151
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13648 5914 13676 6054
rect 14108 5914 14136 9114
rect 13636 5908 13688 5914
rect 13636 5850 13688 5856
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 13634 5808 13690 5817
rect 13634 5743 13690 5752
rect 13648 4729 13676 5743
rect 13726 5672 13782 5681
rect 13726 5607 13728 5616
rect 13780 5607 13782 5616
rect 13728 5578 13780 5584
rect 14200 5250 14228 11290
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14292 9450 14320 11154
rect 14372 11008 14424 11014
rect 14372 10950 14424 10956
rect 14384 10810 14412 10950
rect 14372 10804 14424 10810
rect 14372 10746 14424 10752
rect 14476 9761 14504 11614
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14462 9752 14518 9761
rect 14462 9687 14518 9696
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14280 9444 14332 9450
rect 14280 9386 14332 9392
rect 14292 9042 14320 9386
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14384 8634 14412 9522
rect 14464 9512 14516 9518
rect 14464 9454 14516 9460
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14476 8362 14504 9454
rect 14568 8498 14596 11494
rect 14660 10810 14688 12786
rect 14752 12306 14780 13262
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14844 12238 14872 12582
rect 14945 12540 15253 12560
rect 14945 12538 14951 12540
rect 15007 12538 15031 12540
rect 15087 12538 15111 12540
rect 15167 12538 15191 12540
rect 15247 12538 15253 12540
rect 15007 12486 15009 12538
rect 15189 12486 15191 12538
rect 14945 12484 14951 12486
rect 15007 12484 15031 12486
rect 15087 12484 15111 12486
rect 15167 12484 15191 12486
rect 15247 12484 15253 12486
rect 14945 12464 15253 12484
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14752 11218 14780 12106
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14844 11762 14872 12038
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14945 11452 15253 11472
rect 14945 11450 14951 11452
rect 15007 11450 15031 11452
rect 15087 11450 15111 11452
rect 15167 11450 15191 11452
rect 15247 11450 15253 11452
rect 15007 11398 15009 11450
rect 15189 11398 15191 11450
rect 14945 11396 14951 11398
rect 15007 11396 15031 11398
rect 15087 11396 15111 11398
rect 15167 11396 15191 11398
rect 15247 11396 15253 11398
rect 14945 11376 15253 11396
rect 14740 11212 14792 11218
rect 14740 11154 14792 11160
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14945 10364 15253 10384
rect 14945 10362 14951 10364
rect 15007 10362 15031 10364
rect 15087 10362 15111 10364
rect 15167 10362 15191 10364
rect 15247 10362 15253 10364
rect 15007 10310 15009 10362
rect 15189 10310 15191 10362
rect 14945 10308 14951 10310
rect 15007 10308 15031 10310
rect 15087 10308 15111 10310
rect 15167 10308 15191 10310
rect 15247 10308 15253 10310
rect 14945 10288 15253 10308
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 14740 9444 14792 9450
rect 14740 9386 14792 9392
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14464 8356 14516 8362
rect 14464 8298 14516 8304
rect 14568 7970 14596 8434
rect 14476 7954 14596 7970
rect 14464 7948 14596 7954
rect 14516 7942 14596 7948
rect 14464 7890 14516 7896
rect 14660 7546 14688 8842
rect 14648 7540 14700 7546
rect 14648 7482 14700 7488
rect 14752 7426 14780 9386
rect 14660 7398 14780 7426
rect 14660 6118 14688 7398
rect 14844 7324 14872 9454
rect 14945 9276 15253 9296
rect 14945 9274 14951 9276
rect 15007 9274 15031 9276
rect 15087 9274 15111 9276
rect 15167 9274 15191 9276
rect 15247 9274 15253 9276
rect 15007 9222 15009 9274
rect 15189 9222 15191 9274
rect 14945 9220 14951 9222
rect 15007 9220 15031 9222
rect 15087 9220 15111 9222
rect 15167 9220 15191 9222
rect 15247 9220 15253 9222
rect 14945 9200 15253 9220
rect 15304 8906 15332 12922
rect 15396 12782 15424 13670
rect 15488 12850 15516 14010
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15580 11830 15608 14758
rect 15856 14414 15884 14758
rect 15948 14618 15976 14855
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 16040 14550 16068 17575
rect 16304 17196 16356 17202
rect 16304 17138 16356 17144
rect 16316 16794 16344 17138
rect 16408 16998 16436 19790
rect 16500 17678 16528 20198
rect 16868 19310 16896 20590
rect 17236 20466 17264 20590
rect 16948 20460 17000 20466
rect 16948 20402 17000 20408
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 16856 19304 16908 19310
rect 16856 19246 16908 19252
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16960 17610 16988 20402
rect 17132 20392 17184 20398
rect 17132 20334 17184 20340
rect 17144 19854 17172 20334
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17040 19372 17092 19378
rect 17040 19314 17092 19320
rect 17052 18426 17080 19314
rect 17144 18766 17172 19790
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17130 18456 17186 18465
rect 17040 18420 17092 18426
rect 17130 18391 17132 18400
rect 17040 18362 17092 18368
rect 17184 18391 17186 18400
rect 17132 18362 17184 18368
rect 17052 18154 17080 18362
rect 17132 18216 17184 18222
rect 17132 18158 17184 18164
rect 17224 18216 17276 18222
rect 17224 18158 17276 18164
rect 17040 18148 17092 18154
rect 17040 18090 17092 18096
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 16948 17604 17000 17610
rect 16948 17546 17000 17552
rect 16488 17060 16540 17066
rect 16488 17002 16540 17008
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16028 14544 16080 14550
rect 16028 14486 16080 14492
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 16408 14090 16436 16050
rect 16500 15978 16528 17002
rect 16488 15972 16540 15978
rect 16488 15914 16540 15920
rect 16592 15434 16620 17546
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16684 16590 16712 17478
rect 17144 17338 17172 18158
rect 17236 17746 17264 18158
rect 17328 17882 17356 20742
rect 17420 18902 17448 20742
rect 17744 20700 18052 20720
rect 17744 20698 17750 20700
rect 17806 20698 17830 20700
rect 17886 20698 17910 20700
rect 17966 20698 17990 20700
rect 18046 20698 18052 20700
rect 17806 20646 17808 20698
rect 17988 20646 17990 20698
rect 17744 20644 17750 20646
rect 17806 20644 17830 20646
rect 17886 20644 17910 20646
rect 17966 20644 17990 20646
rect 18046 20644 18052 20646
rect 17744 20624 18052 20644
rect 17960 20528 18012 20534
rect 17590 20496 17646 20505
rect 17590 20431 17646 20440
rect 17958 20496 17960 20505
rect 18012 20496 18014 20505
rect 17958 20431 18014 20440
rect 17604 20097 17632 20431
rect 17684 20392 17736 20398
rect 17684 20334 17736 20340
rect 17590 20088 17646 20097
rect 17590 20023 17646 20032
rect 17696 19786 17724 20334
rect 18156 19854 18184 21422
rect 18144 19848 18196 19854
rect 18340 19825 18368 23800
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18420 20936 18472 20942
rect 18420 20878 18472 20884
rect 18144 19790 18196 19796
rect 18326 19816 18382 19825
rect 17684 19780 17736 19786
rect 17684 19722 17736 19728
rect 17592 19712 17644 19718
rect 17592 19654 17644 19660
rect 17604 19496 17632 19654
rect 17744 19612 18052 19632
rect 17744 19610 17750 19612
rect 17806 19610 17830 19612
rect 17886 19610 17910 19612
rect 17966 19610 17990 19612
rect 18046 19610 18052 19612
rect 17806 19558 17808 19610
rect 17988 19558 17990 19610
rect 17744 19556 17750 19558
rect 17806 19556 17830 19558
rect 17886 19556 17910 19558
rect 17966 19556 17990 19558
rect 18046 19556 18052 19558
rect 17744 19536 18052 19556
rect 17604 19468 17724 19496
rect 17498 19408 17554 19417
rect 17498 19343 17554 19352
rect 17512 19310 17540 19343
rect 17500 19304 17552 19310
rect 17500 19246 17552 19252
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17408 18896 17460 18902
rect 17408 18838 17460 18844
rect 17512 18630 17540 19246
rect 17604 18970 17632 19246
rect 17592 18964 17644 18970
rect 17592 18906 17644 18912
rect 17696 18850 17724 19468
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17604 18834 17724 18850
rect 17592 18828 17724 18834
rect 17644 18822 17724 18828
rect 17592 18770 17644 18776
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17604 18442 17632 18770
rect 17788 18766 17816 18906
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17866 18728 17922 18737
rect 17866 18663 17868 18672
rect 17920 18663 17922 18672
rect 17868 18634 17920 18640
rect 17744 18524 18052 18544
rect 17744 18522 17750 18524
rect 17806 18522 17830 18524
rect 17886 18522 17910 18524
rect 17966 18522 17990 18524
rect 18046 18522 18052 18524
rect 17806 18470 17808 18522
rect 17988 18470 17990 18522
rect 17744 18468 17750 18470
rect 17806 18468 17830 18470
rect 17886 18468 17910 18470
rect 17966 18468 17990 18470
rect 18046 18468 18052 18470
rect 17744 18448 18052 18468
rect 17512 18414 17632 18442
rect 17316 17876 17368 17882
rect 17316 17818 17368 17824
rect 17224 17740 17276 17746
rect 17224 17682 17276 17688
rect 17132 17332 17184 17338
rect 17132 17274 17184 17280
rect 16764 17264 16816 17270
rect 16764 17206 16816 17212
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16776 16114 16804 17206
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16856 16448 16908 16454
rect 16856 16390 16908 16396
rect 16764 16108 16816 16114
rect 16764 16050 16816 16056
rect 16868 15978 16896 16390
rect 16856 15972 16908 15978
rect 16856 15914 16908 15920
rect 16960 15910 16988 17138
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17328 16590 17356 16934
rect 17316 16584 17368 16590
rect 17316 16526 17368 16532
rect 17132 16516 17184 16522
rect 17132 16458 17184 16464
rect 17144 16182 17172 16458
rect 17132 16176 17184 16182
rect 17038 16144 17094 16153
rect 17132 16118 17184 16124
rect 17038 16079 17094 16088
rect 16948 15904 17000 15910
rect 16948 15846 17000 15852
rect 16580 15428 16632 15434
rect 16580 15370 16632 15376
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16500 15026 16528 15098
rect 16488 15020 16540 15026
rect 16488 14962 16540 14968
rect 17052 14958 17080 16079
rect 17040 14952 17092 14958
rect 17040 14894 17092 14900
rect 16408 14062 16620 14090
rect 16488 14000 16540 14006
rect 16486 13968 16488 13977
rect 16540 13968 16542 13977
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16396 13932 16448 13938
rect 16486 13903 16542 13912
rect 16396 13874 16448 13880
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15764 13326 15792 13806
rect 16028 13728 16080 13734
rect 16028 13670 16080 13676
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 16040 12918 16068 13670
rect 16316 13530 16344 13874
rect 16408 13734 16436 13874
rect 16592 13734 16620 14062
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16396 13728 16448 13734
rect 16396 13670 16448 13676
rect 16580 13728 16632 13734
rect 16580 13670 16632 13676
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16316 13326 16344 13466
rect 16304 13320 16356 13326
rect 16304 13262 16356 13268
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16028 12912 16080 12918
rect 16028 12854 16080 12860
rect 15750 12336 15806 12345
rect 15750 12271 15806 12280
rect 15764 12238 15792 12271
rect 16224 12238 16252 13126
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 16212 12232 16264 12238
rect 16212 12174 16264 12180
rect 15568 11824 15620 11830
rect 15568 11766 15620 11772
rect 15476 11756 15528 11762
rect 15476 11698 15528 11704
rect 15488 11354 15516 11698
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15580 11218 15608 11766
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16028 11688 16080 11694
rect 16028 11630 16080 11636
rect 16040 11354 16068 11630
rect 16132 11558 16160 11698
rect 16396 11688 16448 11694
rect 16396 11630 16448 11636
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 16028 11348 16080 11354
rect 16028 11290 16080 11296
rect 15568 11212 15620 11218
rect 15568 11154 15620 11160
rect 15384 11008 15436 11014
rect 15384 10950 15436 10956
rect 15396 10266 15424 10950
rect 16132 10742 16160 11494
rect 16120 10736 16172 10742
rect 16120 10678 16172 10684
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 16408 10062 16436 11630
rect 16592 11286 16620 12786
rect 16684 11762 16712 14010
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 16856 12776 16908 12782
rect 16960 12764 16988 13262
rect 16908 12736 16988 12764
rect 16856 12718 16908 12724
rect 16868 12442 16896 12718
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 17144 12102 17172 13262
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 16948 12096 17000 12102
rect 16948 12038 17000 12044
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16960 11218 16988 12038
rect 17132 11892 17184 11898
rect 17132 11834 17184 11840
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17052 11354 17080 11698
rect 17040 11348 17092 11354
rect 17040 11290 17092 11296
rect 17144 11234 17172 11834
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 17052 11206 17172 11234
rect 16672 10600 16724 10606
rect 16672 10542 16724 10548
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15396 9518 15424 9930
rect 15672 9654 15700 9998
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 15660 9648 15712 9654
rect 15660 9590 15712 9596
rect 15384 9512 15436 9518
rect 15384 9454 15436 9460
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15292 8900 15344 8906
rect 15292 8842 15344 8848
rect 15396 8838 15424 8978
rect 15672 8974 15700 9590
rect 15948 9586 15976 9862
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 16304 9376 16356 9382
rect 16304 9318 16356 9324
rect 15660 8968 15712 8974
rect 15660 8910 15712 8916
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 14945 8188 15253 8208
rect 14945 8186 14951 8188
rect 15007 8186 15031 8188
rect 15087 8186 15111 8188
rect 15167 8186 15191 8188
rect 15247 8186 15253 8188
rect 15007 8134 15009 8186
rect 15189 8134 15191 8186
rect 14945 8132 14951 8134
rect 15007 8132 15031 8134
rect 15087 8132 15111 8134
rect 15167 8132 15191 8134
rect 15247 8132 15253 8134
rect 14945 8112 15253 8132
rect 15200 7812 15252 7818
rect 15200 7754 15252 7760
rect 15212 7546 15240 7754
rect 15396 7750 15424 8366
rect 15672 7954 15700 8910
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15844 8832 15896 8838
rect 15844 8774 15896 8780
rect 15764 8566 15792 8774
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 15660 7948 15712 7954
rect 15660 7890 15712 7896
rect 15856 7886 15884 8774
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16132 8294 16160 8434
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 15844 7880 15896 7886
rect 15844 7822 15896 7828
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15396 7410 15424 7686
rect 16132 7410 16160 8230
rect 16316 7818 16344 9318
rect 16304 7812 16356 7818
rect 16304 7754 16356 7760
rect 16396 7812 16448 7818
rect 16396 7754 16448 7760
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 14752 7296 14872 7324
rect 16210 7304 16266 7313
rect 14752 6458 14780 7296
rect 16210 7239 16212 7248
rect 16264 7239 16266 7248
rect 16212 7210 16264 7216
rect 14945 7100 15253 7120
rect 14945 7098 14951 7100
rect 15007 7098 15031 7100
rect 15087 7098 15111 7100
rect 15167 7098 15191 7100
rect 15247 7098 15253 7100
rect 15007 7046 15009 7098
rect 15189 7046 15191 7098
rect 14945 7044 14951 7046
rect 15007 7044 15031 7046
rect 15087 7044 15111 7046
rect 15167 7044 15191 7046
rect 15247 7044 15253 7046
rect 14945 7024 15253 7044
rect 16408 6798 16436 7754
rect 16396 6792 16448 6798
rect 16396 6734 16448 6740
rect 14832 6656 14884 6662
rect 14832 6598 14884 6604
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14844 6390 14872 6598
rect 14832 6384 14884 6390
rect 14832 6326 14884 6332
rect 15120 6322 15332 6338
rect 15108 6316 15332 6322
rect 15160 6310 15332 6316
rect 15108 6258 15160 6264
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14200 5222 14412 5250
rect 13634 4720 13690 4729
rect 13634 4655 13690 4664
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14292 4146 14320 4422
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 13832 3738 13860 4082
rect 14004 4072 14056 4078
rect 14004 4014 14056 4020
rect 14096 4072 14148 4078
rect 14096 4014 14148 4020
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 13636 3392 13688 3398
rect 13636 3334 13688 3340
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13648 3097 13676 3334
rect 13634 3088 13690 3097
rect 13634 3023 13690 3032
rect 13542 2952 13598 2961
rect 13542 2887 13598 2896
rect 13740 2854 13768 3334
rect 13832 3126 13860 3674
rect 13924 3194 13952 3878
rect 13912 3188 13964 3194
rect 13912 3130 13964 3136
rect 13820 3120 13872 3126
rect 13820 3062 13872 3068
rect 14016 2922 14044 4014
rect 14108 3126 14136 4014
rect 14188 3460 14240 3466
rect 14188 3402 14240 3408
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 14096 2984 14148 2990
rect 14096 2926 14148 2932
rect 14004 2916 14056 2922
rect 14004 2858 14056 2864
rect 13728 2848 13780 2854
rect 13728 2790 13780 2796
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 14016 2446 14044 2858
rect 14108 2582 14136 2926
rect 14200 2650 14228 3402
rect 14384 2972 14412 5222
rect 14464 5092 14516 5098
rect 14464 5034 14516 5040
rect 14476 3346 14504 5034
rect 14660 4486 14688 6054
rect 14945 6012 15253 6032
rect 14945 6010 14951 6012
rect 15007 6010 15031 6012
rect 15087 6010 15111 6012
rect 15167 6010 15191 6012
rect 15247 6010 15253 6012
rect 15007 5958 15009 6010
rect 15189 5958 15191 6010
rect 14945 5956 14951 5958
rect 15007 5956 15031 5958
rect 15087 5956 15111 5958
rect 15167 5956 15191 5958
rect 15247 5956 15253 5958
rect 14945 5936 15253 5956
rect 15200 5840 15252 5846
rect 15200 5782 15252 5788
rect 15212 5574 15240 5782
rect 15304 5710 15332 6310
rect 16302 6216 16358 6225
rect 16302 6151 16358 6160
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15384 5636 15436 5642
rect 15384 5578 15436 5584
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14648 4480 14700 4486
rect 14648 4422 14700 4428
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14568 3466 14596 3878
rect 14646 3496 14702 3505
rect 14556 3460 14608 3466
rect 14646 3431 14702 3440
rect 14556 3402 14608 3408
rect 14554 3360 14610 3369
rect 14476 3318 14554 3346
rect 14554 3295 14610 3304
rect 14568 3194 14596 3295
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14660 3058 14688 3431
rect 14752 3194 14780 5102
rect 14945 4924 15253 4944
rect 14945 4922 14951 4924
rect 15007 4922 15031 4924
rect 15087 4922 15111 4924
rect 15167 4922 15191 4924
rect 15247 4922 15253 4924
rect 15007 4870 15009 4922
rect 15189 4870 15191 4922
rect 14945 4868 14951 4870
rect 15007 4868 15031 4870
rect 15087 4868 15111 4870
rect 15167 4868 15191 4870
rect 15247 4868 15253 4870
rect 14945 4848 15253 4868
rect 15016 4752 15068 4758
rect 15014 4720 15016 4729
rect 15068 4720 15070 4729
rect 15014 4655 15070 4664
rect 14832 3936 14884 3942
rect 14832 3878 14884 3884
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 14844 3641 14872 3878
rect 14945 3836 15253 3856
rect 14945 3834 14951 3836
rect 15007 3834 15031 3836
rect 15087 3834 15111 3836
rect 15167 3834 15191 3836
rect 15247 3834 15253 3836
rect 15007 3782 15009 3834
rect 15189 3782 15191 3834
rect 14945 3780 14951 3782
rect 15007 3780 15031 3782
rect 15087 3780 15111 3782
rect 15167 3780 15191 3782
rect 15247 3780 15253 3782
rect 14945 3760 15253 3780
rect 15304 3738 15332 3878
rect 15292 3732 15344 3738
rect 15292 3674 15344 3680
rect 14830 3632 14886 3641
rect 14830 3567 14886 3576
rect 14740 3188 14792 3194
rect 14740 3130 14792 3136
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14464 2984 14516 2990
rect 14384 2944 14464 2972
rect 14280 2916 14332 2922
rect 14280 2858 14332 2864
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14096 2576 14148 2582
rect 14096 2518 14148 2524
rect 14292 2514 14320 2858
rect 14384 2854 14412 2944
rect 14464 2926 14516 2932
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 14384 2514 14412 2790
rect 14280 2508 14332 2514
rect 14280 2450 14332 2456
rect 14372 2508 14424 2514
rect 14372 2450 14424 2456
rect 14004 2440 14056 2446
rect 14004 2382 14056 2388
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 12146 2204 12454 2224
rect 12146 2202 12152 2204
rect 12208 2202 12232 2204
rect 12288 2202 12312 2204
rect 12368 2202 12392 2204
rect 12448 2202 12454 2204
rect 12208 2150 12210 2202
rect 12390 2150 12392 2202
rect 12146 2148 12152 2150
rect 12208 2148 12232 2150
rect 12288 2148 12312 2150
rect 12368 2148 12392 2150
rect 12448 2148 12454 2150
rect 12146 2128 12454 2148
rect 14844 1970 14872 3567
rect 14945 2748 15253 2768
rect 14945 2746 14951 2748
rect 15007 2746 15031 2748
rect 15087 2746 15111 2748
rect 15167 2746 15191 2748
rect 15247 2746 15253 2748
rect 15007 2694 15009 2746
rect 15189 2694 15191 2746
rect 14945 2692 14951 2694
rect 15007 2692 15031 2694
rect 15087 2692 15111 2694
rect 15167 2692 15191 2694
rect 15247 2692 15253 2694
rect 14945 2672 15253 2692
rect 15396 2582 15424 5578
rect 16120 5228 16172 5234
rect 16120 5170 16172 5176
rect 16132 5001 16160 5170
rect 16316 5137 16344 6151
rect 16408 5642 16436 6734
rect 16396 5636 16448 5642
rect 16396 5578 16448 5584
rect 16408 5166 16436 5578
rect 16500 5370 16528 9998
rect 16684 8974 16712 10542
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16764 10260 16816 10266
rect 16764 10202 16816 10208
rect 16776 9042 16804 10202
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16868 9110 16896 9454
rect 16856 9104 16908 9110
rect 16856 9046 16908 9052
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 16672 8968 16724 8974
rect 16672 8910 16724 8916
rect 16764 7880 16816 7886
rect 16764 7822 16816 7828
rect 16672 7812 16724 7818
rect 16672 7754 16724 7760
rect 16684 6730 16712 7754
rect 16776 7274 16804 7822
rect 16868 7342 16896 9046
rect 16960 9042 16988 10406
rect 17052 9382 17080 11206
rect 17236 11150 17264 12038
rect 17328 11354 17356 12718
rect 17408 12640 17460 12646
rect 17408 12582 17460 12588
rect 17316 11348 17368 11354
rect 17316 11290 17368 11296
rect 17420 11218 17448 12582
rect 17512 11898 17540 18414
rect 17684 18216 17736 18222
rect 17590 18184 17646 18193
rect 17684 18158 17736 18164
rect 17590 18119 17646 18128
rect 17604 16522 17632 18119
rect 17696 17814 17724 18158
rect 17684 17808 17736 17814
rect 17684 17750 17736 17756
rect 18156 17610 18184 19790
rect 18326 19751 18382 19760
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 18248 18970 18276 19654
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18326 18728 18382 18737
rect 18326 18663 18328 18672
rect 18380 18663 18382 18672
rect 18328 18634 18380 18640
rect 18236 18624 18288 18630
rect 18236 18566 18288 18572
rect 18144 17604 18196 17610
rect 18144 17546 18196 17552
rect 17744 17436 18052 17456
rect 17744 17434 17750 17436
rect 17806 17434 17830 17436
rect 17886 17434 17910 17436
rect 17966 17434 17990 17436
rect 18046 17434 18052 17436
rect 17806 17382 17808 17434
rect 17988 17382 17990 17434
rect 17744 17380 17750 17382
rect 17806 17380 17830 17382
rect 17886 17380 17910 17382
rect 17966 17380 17990 17382
rect 18046 17380 18052 17382
rect 17744 17360 18052 17380
rect 18156 17270 18184 17546
rect 18248 17542 18276 18566
rect 18236 17536 18288 17542
rect 18236 17478 18288 17484
rect 18144 17264 18196 17270
rect 18144 17206 18196 17212
rect 18156 16794 18184 17206
rect 18432 16998 18460 20878
rect 18524 18426 18552 21966
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18708 21622 18736 21830
rect 18696 21616 18748 21622
rect 18696 21558 18748 21564
rect 18880 21004 18932 21010
rect 18880 20946 18932 20952
rect 18604 20800 18656 20806
rect 18604 20742 18656 20748
rect 18616 20602 18644 20742
rect 18604 20596 18656 20602
rect 18604 20538 18656 20544
rect 18616 19922 18644 20538
rect 18604 19916 18656 19922
rect 18604 19858 18656 19864
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18616 19310 18644 19654
rect 18604 19304 18656 19310
rect 18604 19246 18656 19252
rect 18512 18420 18564 18426
rect 18512 18362 18564 18368
rect 18512 18284 18564 18290
rect 18512 18226 18564 18232
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 17592 16516 17644 16522
rect 17592 16458 17644 16464
rect 17744 16348 18052 16368
rect 17744 16346 17750 16348
rect 17806 16346 17830 16348
rect 17886 16346 17910 16348
rect 17966 16346 17990 16348
rect 18046 16346 18052 16348
rect 17806 16294 17808 16346
rect 17988 16294 17990 16346
rect 17744 16292 17750 16294
rect 17806 16292 17830 16294
rect 17886 16292 17910 16294
rect 17966 16292 17990 16294
rect 18046 16292 18052 16294
rect 17744 16272 18052 16292
rect 18156 16096 18184 16730
rect 18236 16108 18288 16114
rect 18156 16068 18236 16096
rect 18236 16050 18288 16056
rect 18524 15910 18552 18226
rect 18616 18086 18644 19246
rect 18696 18760 18748 18766
rect 18696 18702 18748 18708
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18708 17338 18736 18702
rect 18892 17746 18920 20946
rect 18984 19961 19012 23800
rect 19154 22128 19210 22137
rect 19154 22063 19210 22072
rect 19064 21888 19116 21894
rect 19064 21830 19116 21836
rect 19076 21622 19104 21830
rect 19064 21616 19116 21622
rect 19064 21558 19116 21564
rect 19168 21146 19196 22063
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19432 22024 19484 22030
rect 19432 21966 19484 21972
rect 19260 21894 19288 21966
rect 19248 21888 19300 21894
rect 19248 21830 19300 21836
rect 19338 21720 19394 21729
rect 19444 21690 19472 21966
rect 19628 21690 19656 23800
rect 20272 22438 20300 23800
rect 20916 23746 20944 23800
rect 21008 23746 21036 23854
rect 20916 23718 21036 23746
rect 20442 23624 20498 23633
rect 20442 23559 20498 23568
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 19984 22092 20036 22098
rect 19984 22034 20036 22040
rect 19708 21956 19760 21962
rect 19708 21898 19760 21904
rect 19338 21655 19394 21664
rect 19432 21684 19484 21690
rect 19248 21344 19300 21350
rect 19248 21286 19300 21292
rect 19260 21146 19288 21286
rect 19156 21140 19208 21146
rect 19156 21082 19208 21088
rect 19248 21140 19300 21146
rect 19248 21082 19300 21088
rect 19352 20482 19380 21655
rect 19432 21626 19484 21632
rect 19616 21684 19668 21690
rect 19616 21626 19668 21632
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19616 21344 19668 21350
rect 19616 21286 19668 21292
rect 19430 20768 19486 20777
rect 19430 20703 19486 20712
rect 19076 20454 19380 20482
rect 19076 20398 19104 20454
rect 19064 20392 19116 20398
rect 19248 20392 19300 20398
rect 19064 20334 19116 20340
rect 19154 20360 19210 20369
rect 19248 20334 19300 20340
rect 19154 20295 19210 20304
rect 19064 20256 19116 20262
rect 19064 20198 19116 20204
rect 18970 19952 19026 19961
rect 18970 19887 19026 19896
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18984 18630 19012 19790
rect 19076 18766 19104 20198
rect 19168 20058 19196 20295
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19260 19802 19288 20334
rect 19340 19848 19392 19854
rect 19260 19796 19340 19802
rect 19260 19790 19392 19796
rect 19260 19774 19380 19790
rect 19260 19514 19288 19774
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19156 19304 19208 19310
rect 19156 19246 19208 19252
rect 19064 18760 19116 18766
rect 19064 18702 19116 18708
rect 18972 18624 19024 18630
rect 18972 18566 19024 18572
rect 18880 17740 18932 17746
rect 18880 17682 18932 17688
rect 18984 17626 19012 18566
rect 19064 18216 19116 18222
rect 19064 18158 19116 18164
rect 18892 17598 19012 17626
rect 18696 17332 18748 17338
rect 18696 17274 18748 17280
rect 18892 16454 18920 17598
rect 19076 17542 19104 18158
rect 19168 18086 19196 19246
rect 19340 19168 19392 19174
rect 19340 19110 19392 19116
rect 19352 18902 19380 19110
rect 19340 18896 19392 18902
rect 19340 18838 19392 18844
rect 19248 18420 19300 18426
rect 19248 18362 19300 18368
rect 19156 18080 19208 18086
rect 19156 18022 19208 18028
rect 19064 17536 19116 17542
rect 19064 17478 19116 17484
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18696 16040 18748 16046
rect 18696 15982 18748 15988
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 17696 15434 17724 15846
rect 17972 15706 18000 15846
rect 17960 15700 18012 15706
rect 17960 15642 18012 15648
rect 18052 15700 18104 15706
rect 18052 15642 18104 15648
rect 18064 15570 18092 15642
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 18052 15564 18104 15570
rect 18052 15506 18104 15512
rect 18144 15496 18196 15502
rect 18144 15438 18196 15444
rect 17592 15428 17644 15434
rect 17592 15370 17644 15376
rect 17684 15428 17736 15434
rect 17684 15370 17736 15376
rect 17604 14618 17632 15370
rect 17744 15260 18052 15280
rect 17744 15258 17750 15260
rect 17806 15258 17830 15260
rect 17886 15258 17910 15260
rect 17966 15258 17990 15260
rect 18046 15258 18052 15260
rect 17806 15206 17808 15258
rect 17988 15206 17990 15258
rect 17744 15204 17750 15206
rect 17806 15204 17830 15206
rect 17886 15204 17910 15206
rect 17966 15204 17990 15206
rect 18046 15204 18052 15206
rect 17744 15184 18052 15204
rect 18156 15026 18184 15438
rect 18144 15020 18196 15026
rect 18144 14962 18196 14968
rect 17592 14612 17644 14618
rect 17592 14554 17644 14560
rect 17744 14172 18052 14192
rect 17744 14170 17750 14172
rect 17806 14170 17830 14172
rect 17886 14170 17910 14172
rect 17966 14170 17990 14172
rect 18046 14170 18052 14172
rect 17806 14118 17808 14170
rect 17988 14118 17990 14170
rect 17744 14116 17750 14118
rect 17806 14116 17830 14118
rect 17886 14116 17910 14118
rect 17966 14116 17990 14118
rect 18046 14116 18052 14118
rect 17744 14096 18052 14116
rect 18156 13938 18184 14962
rect 18340 14958 18368 15574
rect 18708 15162 18736 15982
rect 18800 15706 18828 16050
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18892 15502 18920 15846
rect 18984 15638 19012 17070
rect 19064 15972 19116 15978
rect 19064 15914 19116 15920
rect 18972 15632 19024 15638
rect 18972 15574 19024 15580
rect 18880 15496 18932 15502
rect 18880 15438 18932 15444
rect 18696 15156 18748 15162
rect 18696 15098 18748 15104
rect 18512 15020 18564 15026
rect 18512 14962 18564 14968
rect 18328 14952 18380 14958
rect 18328 14894 18380 14900
rect 18524 14414 18552 14962
rect 18880 14884 18932 14890
rect 18880 14826 18932 14832
rect 18512 14408 18564 14414
rect 18512 14350 18564 14356
rect 18892 14346 18920 14826
rect 18880 14340 18932 14346
rect 18880 14282 18932 14288
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 17684 13932 17736 13938
rect 17604 13892 17684 13920
rect 17604 11898 17632 13892
rect 17684 13874 17736 13880
rect 18144 13932 18196 13938
rect 18144 13874 18196 13880
rect 17744 13084 18052 13104
rect 17744 13082 17750 13084
rect 17806 13082 17830 13084
rect 17886 13082 17910 13084
rect 17966 13082 17990 13084
rect 18046 13082 18052 13084
rect 17806 13030 17808 13082
rect 17988 13030 17990 13082
rect 17744 13028 17750 13030
rect 17806 13028 17830 13030
rect 17886 13028 17910 13030
rect 17966 13028 17990 13030
rect 18046 13028 18052 13030
rect 17744 13008 18052 13028
rect 18156 12918 18184 13874
rect 18420 13864 18472 13870
rect 18420 13806 18472 13812
rect 18236 13184 18288 13190
rect 18236 13126 18288 13132
rect 18328 13184 18380 13190
rect 18328 13126 18380 13132
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 18156 12442 18184 12854
rect 17868 12436 17920 12442
rect 17868 12378 17920 12384
rect 18144 12436 18196 12442
rect 18144 12378 18196 12384
rect 17880 12209 17908 12378
rect 17866 12200 17922 12209
rect 17866 12135 17922 12144
rect 18144 12164 18196 12170
rect 18248 12152 18276 13126
rect 18196 12124 18276 12152
rect 18144 12106 18196 12112
rect 17744 11996 18052 12016
rect 17744 11994 17750 11996
rect 17806 11994 17830 11996
rect 17886 11994 17910 11996
rect 17966 11994 17990 11996
rect 18046 11994 18052 11996
rect 17806 11942 17808 11994
rect 17988 11942 17990 11994
rect 17744 11940 17750 11942
rect 17806 11940 17830 11942
rect 17886 11940 17910 11942
rect 17966 11940 17990 11942
rect 18046 11940 18052 11942
rect 17744 11920 18052 11940
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17500 11280 17552 11286
rect 17500 11222 17552 11228
rect 17408 11212 17460 11218
rect 17408 11154 17460 11160
rect 17224 11144 17276 11150
rect 17224 11086 17276 11092
rect 17512 10810 17540 11222
rect 17604 11218 17632 11834
rect 18340 11830 18368 13126
rect 18432 11830 18460 13806
rect 18616 12986 18644 14214
rect 19076 13938 19104 15914
rect 19168 14958 19196 18022
rect 19260 17882 19288 18362
rect 19444 18358 19472 20703
rect 19536 20330 19564 21286
rect 19628 21078 19656 21286
rect 19616 21072 19668 21078
rect 19616 21014 19668 21020
rect 19720 20602 19748 21898
rect 19892 21888 19944 21894
rect 19892 21830 19944 21836
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 19708 20596 19760 20602
rect 19708 20538 19760 20544
rect 19812 20505 19840 21286
rect 19904 21049 19932 21830
rect 19996 21418 20024 22034
rect 20456 21894 20484 23559
rect 20543 22332 20851 22352
rect 20543 22330 20549 22332
rect 20605 22330 20629 22332
rect 20685 22330 20709 22332
rect 20765 22330 20789 22332
rect 20845 22330 20851 22332
rect 20605 22278 20607 22330
rect 20787 22278 20789 22330
rect 20543 22276 20549 22278
rect 20605 22276 20629 22278
rect 20685 22276 20709 22278
rect 20765 22276 20789 22278
rect 20845 22276 20851 22278
rect 20543 22256 20851 22276
rect 20628 22024 20680 22030
rect 20548 21984 20628 22012
rect 20444 21888 20496 21894
rect 20166 21856 20222 21865
rect 20444 21830 20496 21836
rect 20166 21791 20222 21800
rect 19984 21412 20036 21418
rect 19984 21354 20036 21360
rect 20180 21146 20208 21791
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20364 21146 20392 21490
rect 20548 21434 20576 21984
rect 20628 21966 20680 21972
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 20916 21865 20944 21966
rect 20902 21856 20958 21865
rect 20902 21791 20958 21800
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 20456 21406 20576 21434
rect 20168 21140 20220 21146
rect 20168 21082 20220 21088
rect 20352 21140 20404 21146
rect 20352 21082 20404 21088
rect 19890 21040 19946 21049
rect 19890 20975 19946 20984
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 19984 20936 20036 20942
rect 19984 20878 20036 20884
rect 19798 20496 19854 20505
rect 19616 20460 19668 20466
rect 19798 20431 19854 20440
rect 19616 20402 19668 20408
rect 19524 20324 19576 20330
rect 19524 20266 19576 20272
rect 19628 20210 19656 20402
rect 19536 20182 19656 20210
rect 19536 19281 19564 20182
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19628 19417 19656 19654
rect 19614 19408 19670 19417
rect 19614 19343 19670 19352
rect 19522 19272 19578 19281
rect 19522 19207 19578 19216
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19536 18698 19564 19110
rect 19524 18692 19576 18698
rect 19524 18634 19576 18640
rect 19616 18692 19668 18698
rect 19616 18634 19668 18640
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19628 18222 19656 18634
rect 19720 18290 19748 19858
rect 19800 19236 19852 19242
rect 19800 19178 19852 19184
rect 19708 18284 19760 18290
rect 19708 18226 19760 18232
rect 19432 18216 19484 18222
rect 19432 18158 19484 18164
rect 19616 18216 19668 18222
rect 19616 18158 19668 18164
rect 19248 17876 19300 17882
rect 19248 17818 19300 17824
rect 19340 17808 19392 17814
rect 19340 17750 19392 17756
rect 19352 17649 19380 17750
rect 19444 17678 19472 18158
rect 19524 18080 19576 18086
rect 19524 18022 19576 18028
rect 19616 18080 19668 18086
rect 19616 18022 19668 18028
rect 19432 17672 19484 17678
rect 19338 17640 19394 17649
rect 19432 17614 19484 17620
rect 19338 17575 19394 17584
rect 19536 17338 19564 18022
rect 19524 17332 19576 17338
rect 19524 17274 19576 17280
rect 19248 17060 19300 17066
rect 19248 17002 19300 17008
rect 19260 16726 19288 17002
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19536 16726 19564 16934
rect 19248 16720 19300 16726
rect 19248 16662 19300 16668
rect 19524 16720 19576 16726
rect 19524 16662 19576 16668
rect 19260 16590 19288 16662
rect 19248 16584 19300 16590
rect 19248 16526 19300 16532
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19260 15570 19288 16050
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19352 15162 19380 16050
rect 19628 15450 19656 18022
rect 19812 17202 19840 19178
rect 19904 18970 19932 20878
rect 19996 20398 20024 20878
rect 20352 20528 20404 20534
rect 20352 20470 20404 20476
rect 19984 20392 20036 20398
rect 19984 20334 20036 20340
rect 20364 20233 20392 20470
rect 20350 20224 20406 20233
rect 20350 20159 20406 20168
rect 20456 19258 20484 21406
rect 20543 21244 20851 21264
rect 20543 21242 20549 21244
rect 20605 21242 20629 21244
rect 20685 21242 20709 21244
rect 20765 21242 20789 21244
rect 20845 21242 20851 21244
rect 20605 21190 20607 21242
rect 20787 21190 20789 21242
rect 20543 21188 20549 21190
rect 20605 21188 20629 21190
rect 20685 21188 20709 21190
rect 20765 21188 20789 21190
rect 20845 21188 20851 21190
rect 20543 21168 20851 21188
rect 20718 20904 20774 20913
rect 20718 20839 20720 20848
rect 20772 20839 20774 20848
rect 20720 20810 20772 20816
rect 20812 20800 20864 20806
rect 20812 20742 20864 20748
rect 20824 20244 20852 20742
rect 20916 20466 20944 21490
rect 20996 21480 21048 21486
rect 20996 21422 21048 21428
rect 21008 20942 21036 21422
rect 20996 20936 21048 20942
rect 21100 20913 21128 21490
rect 20996 20878 21048 20884
rect 21086 20904 21142 20913
rect 21086 20839 21142 20848
rect 21192 20602 21220 23854
rect 21546 23800 21602 24600
rect 22190 23800 22246 24600
rect 22834 23800 22890 24600
rect 23202 24304 23258 24313
rect 23202 24239 23258 24248
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20996 20460 21048 20466
rect 20996 20402 21048 20408
rect 20824 20216 20944 20244
rect 20543 20156 20851 20176
rect 20543 20154 20549 20156
rect 20605 20154 20629 20156
rect 20685 20154 20709 20156
rect 20765 20154 20789 20156
rect 20845 20154 20851 20156
rect 20605 20102 20607 20154
rect 20787 20102 20789 20154
rect 20543 20100 20549 20102
rect 20605 20100 20629 20102
rect 20685 20100 20709 20102
rect 20765 20100 20789 20102
rect 20845 20100 20851 20102
rect 20543 20080 20851 20100
rect 20718 19816 20774 19825
rect 20640 19774 20718 19802
rect 20640 19446 20668 19774
rect 20916 19786 20944 20216
rect 21008 19922 21036 20402
rect 21376 20346 21404 21422
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21100 20318 21404 20346
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 21100 19802 21128 20318
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 21272 20256 21324 20262
rect 21272 20198 21324 20204
rect 21192 19854 21220 20198
rect 20718 19751 20774 19760
rect 20904 19780 20956 19786
rect 20904 19722 20956 19728
rect 21008 19774 21128 19802
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 20628 19440 20680 19446
rect 20628 19382 20680 19388
rect 20640 19281 20668 19382
rect 20904 19372 20956 19378
rect 20904 19314 20956 19320
rect 20180 19230 20484 19258
rect 20626 19272 20682 19281
rect 19892 18964 19944 18970
rect 19892 18906 19944 18912
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 19800 17196 19852 17202
rect 19800 17138 19852 17144
rect 19800 17060 19852 17066
rect 19800 17002 19852 17008
rect 19708 16992 19760 16998
rect 19708 16934 19760 16940
rect 19720 16658 19748 16934
rect 19708 16652 19760 16658
rect 19708 16594 19760 16600
rect 19812 16046 19840 17002
rect 19800 16040 19852 16046
rect 19800 15982 19852 15988
rect 19812 15570 19840 15982
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 19628 15422 19748 15450
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19616 15360 19668 15366
rect 19616 15302 19668 15308
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19156 14952 19208 14958
rect 19156 14894 19208 14900
rect 19168 14482 19196 14894
rect 19156 14476 19208 14482
rect 19156 14418 19208 14424
rect 19156 14340 19208 14346
rect 19156 14282 19208 14288
rect 19168 14074 19196 14282
rect 19352 14074 19380 15098
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19444 14278 19472 14962
rect 19536 14618 19564 15302
rect 19628 15162 19656 15302
rect 19616 15156 19668 15162
rect 19616 15098 19668 15104
rect 19616 14816 19668 14822
rect 19616 14758 19668 14764
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19156 14068 19208 14074
rect 19156 14010 19208 14016
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 18786 13560 18842 13569
rect 19628 13530 19656 14758
rect 18786 13495 18842 13504
rect 19616 13524 19668 13530
rect 18800 13394 18828 13495
rect 19616 13466 19668 13472
rect 19062 13424 19118 13433
rect 18788 13388 18840 13394
rect 19062 13359 19064 13368
rect 18788 13330 18840 13336
rect 19116 13359 19118 13368
rect 19064 13330 19116 13336
rect 19614 13288 19670 13297
rect 19614 13223 19670 13232
rect 18512 12980 18564 12986
rect 18512 12922 18564 12928
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18524 12170 18552 12922
rect 19248 12640 19300 12646
rect 19248 12582 19300 12588
rect 18604 12368 18656 12374
rect 18602 12336 18604 12345
rect 18656 12336 18658 12345
rect 18602 12271 18658 12280
rect 19064 12232 19116 12238
rect 18602 12200 18658 12209
rect 18512 12164 18564 12170
rect 18602 12135 18658 12144
rect 19062 12200 19064 12209
rect 19116 12200 19118 12209
rect 19062 12135 19118 12144
rect 18512 12106 18564 12112
rect 18616 11898 18644 12135
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 18328 11824 18380 11830
rect 18328 11766 18380 11772
rect 18420 11824 18472 11830
rect 18420 11766 18472 11772
rect 18604 11688 18656 11694
rect 18604 11630 18656 11636
rect 17776 11552 17828 11558
rect 17776 11494 17828 11500
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17788 11150 17816 11494
rect 18616 11218 18644 11630
rect 18972 11552 19024 11558
rect 18972 11494 19024 11500
rect 18984 11286 19012 11494
rect 18972 11280 19024 11286
rect 18972 11222 19024 11228
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 18972 11144 19024 11150
rect 18972 11086 19024 11092
rect 18696 11076 18748 11082
rect 18696 11018 18748 11024
rect 17744 10908 18052 10928
rect 17744 10906 17750 10908
rect 17806 10906 17830 10908
rect 17886 10906 17910 10908
rect 17966 10906 17990 10908
rect 18046 10906 18052 10908
rect 17806 10854 17808 10906
rect 17988 10854 17990 10906
rect 17744 10852 17750 10854
rect 17806 10852 17830 10854
rect 17886 10852 17910 10854
rect 17966 10852 17990 10854
rect 18046 10852 18052 10854
rect 17744 10832 18052 10852
rect 17500 10804 17552 10810
rect 17500 10746 17552 10752
rect 17408 10668 17460 10674
rect 17408 10610 17460 10616
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17236 9926 17264 10542
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17040 9376 17092 9382
rect 17040 9318 17092 9324
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 17144 8634 17172 9862
rect 17420 9586 17448 10610
rect 18708 10606 18736 11018
rect 18984 10674 19012 11086
rect 19260 11082 19288 12582
rect 19628 12442 19656 13223
rect 19720 12850 19748 15422
rect 19904 15026 19932 18702
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 19996 15706 20024 16526
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 19904 14618 19932 14962
rect 19892 14612 19944 14618
rect 19892 14554 19944 14560
rect 20076 14408 20128 14414
rect 20076 14350 20128 14356
rect 19984 14272 20036 14278
rect 19984 14214 20036 14220
rect 19996 13326 20024 14214
rect 20088 14074 20116 14350
rect 20180 14278 20208 19230
rect 20626 19207 20682 19216
rect 20260 19168 20312 19174
rect 20260 19110 20312 19116
rect 20272 18358 20300 19110
rect 20543 19068 20851 19088
rect 20543 19066 20549 19068
rect 20605 19066 20629 19068
rect 20685 19066 20709 19068
rect 20765 19066 20789 19068
rect 20845 19066 20851 19068
rect 20605 19014 20607 19066
rect 20787 19014 20789 19066
rect 20543 19012 20549 19014
rect 20605 19012 20629 19014
rect 20685 19012 20709 19014
rect 20765 19012 20789 19014
rect 20845 19012 20851 19014
rect 20543 18992 20851 19012
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20352 18896 20404 18902
rect 20352 18838 20404 18844
rect 20260 18352 20312 18358
rect 20260 18294 20312 18300
rect 20364 18086 20392 18838
rect 20456 18358 20484 18906
rect 20916 18426 20944 19314
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20444 18352 20496 18358
rect 20444 18294 20496 18300
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 20543 17980 20851 18000
rect 20543 17978 20549 17980
rect 20605 17978 20629 17980
rect 20685 17978 20709 17980
rect 20765 17978 20789 17980
rect 20845 17978 20851 17980
rect 20605 17926 20607 17978
rect 20787 17926 20789 17978
rect 20543 17924 20549 17926
rect 20605 17924 20629 17926
rect 20685 17924 20709 17926
rect 20765 17924 20789 17926
rect 20845 17924 20851 17926
rect 20543 17904 20851 17924
rect 20628 17808 20680 17814
rect 20628 17750 20680 17756
rect 20640 17626 20668 17750
rect 20548 17610 20668 17626
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20536 17604 20668 17610
rect 20588 17598 20668 17604
rect 20536 17546 20588 17552
rect 20732 17542 20760 17614
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20260 16992 20312 16998
rect 20260 16934 20312 16940
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20168 14272 20220 14278
rect 20168 14214 20220 14220
rect 20272 14090 20300 16934
rect 20543 16892 20851 16912
rect 20543 16890 20549 16892
rect 20605 16890 20629 16892
rect 20685 16890 20709 16892
rect 20765 16890 20789 16892
rect 20845 16890 20851 16892
rect 20605 16838 20607 16890
rect 20787 16838 20789 16890
rect 20543 16836 20549 16838
rect 20605 16836 20629 16838
rect 20685 16836 20709 16838
rect 20765 16836 20789 16838
rect 20845 16836 20851 16838
rect 20543 16816 20851 16836
rect 20916 16590 20944 16934
rect 20536 16584 20588 16590
rect 20904 16584 20956 16590
rect 20588 16532 20760 16538
rect 20536 16526 20760 16532
rect 20904 16526 20956 16532
rect 20548 16510 20760 16526
rect 20352 16448 20404 16454
rect 20732 16436 20760 16510
rect 20732 16408 20944 16436
rect 20352 16390 20404 16396
rect 20364 15570 20392 16390
rect 20444 15904 20496 15910
rect 20444 15846 20496 15852
rect 20352 15564 20404 15570
rect 20352 15506 20404 15512
rect 20352 14408 20404 14414
rect 20456 14396 20484 15846
rect 20543 15804 20851 15824
rect 20543 15802 20549 15804
rect 20605 15802 20629 15804
rect 20685 15802 20709 15804
rect 20765 15802 20789 15804
rect 20845 15802 20851 15804
rect 20605 15750 20607 15802
rect 20787 15750 20789 15802
rect 20543 15748 20549 15750
rect 20605 15748 20629 15750
rect 20685 15748 20709 15750
rect 20765 15748 20789 15750
rect 20845 15748 20851 15750
rect 20543 15728 20851 15748
rect 20916 15638 20944 16408
rect 21008 16017 21036 19774
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 21100 17066 21128 19654
rect 21192 18766 21220 19790
rect 21284 19514 21312 20198
rect 21468 20058 21496 20742
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21272 19508 21324 19514
rect 21272 19450 21324 19456
rect 21364 19372 21416 19378
rect 21364 19314 21416 19320
rect 21180 18760 21232 18766
rect 21180 18702 21232 18708
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21284 18290 21312 18566
rect 21272 18284 21324 18290
rect 21272 18226 21324 18232
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 21180 17876 21232 17882
rect 21180 17818 21232 17824
rect 21088 17060 21140 17066
rect 21088 17002 21140 17008
rect 21192 16522 21220 17818
rect 21284 17270 21312 18022
rect 21272 17264 21324 17270
rect 21272 17206 21324 17212
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 20994 16008 21050 16017
rect 20994 15943 21050 15952
rect 20904 15632 20956 15638
rect 20904 15574 20956 15580
rect 20996 15564 21048 15570
rect 20996 15506 21048 15512
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20916 15162 20944 15438
rect 20904 15156 20956 15162
rect 20904 15098 20956 15104
rect 21008 14958 21036 15506
rect 21100 15008 21128 16390
rect 21272 15632 21324 15638
rect 21272 15574 21324 15580
rect 21284 15502 21312 15574
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21284 15162 21312 15302
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 21180 15020 21232 15026
rect 21100 14980 21180 15008
rect 21180 14962 21232 14968
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 20543 14716 20851 14736
rect 20543 14714 20549 14716
rect 20605 14714 20629 14716
rect 20685 14714 20709 14716
rect 20765 14714 20789 14716
rect 20845 14714 20851 14716
rect 20605 14662 20607 14714
rect 20787 14662 20789 14714
rect 20543 14660 20549 14662
rect 20605 14660 20629 14662
rect 20685 14660 20709 14662
rect 20765 14660 20789 14662
rect 20845 14660 20851 14662
rect 20543 14640 20851 14660
rect 21008 14482 21036 14894
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 20404 14368 20484 14396
rect 20720 14408 20772 14414
rect 20352 14350 20404 14356
rect 20720 14350 20772 14356
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 20076 14068 20128 14074
rect 20076 14010 20128 14016
rect 20180 14062 20300 14090
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 20088 12986 20116 13874
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 19708 12844 19760 12850
rect 19760 12804 19840 12832
rect 19708 12786 19760 12792
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 19432 12096 19484 12102
rect 19432 12038 19484 12044
rect 19444 11898 19472 12038
rect 19432 11892 19484 11898
rect 19432 11834 19484 11840
rect 19248 11076 19300 11082
rect 19248 11018 19300 11024
rect 19064 11008 19116 11014
rect 19064 10950 19116 10956
rect 18972 10668 19024 10674
rect 18972 10610 19024 10616
rect 18328 10600 18380 10606
rect 18328 10542 18380 10548
rect 18512 10600 18564 10606
rect 18512 10542 18564 10548
rect 18696 10600 18748 10606
rect 18696 10542 18748 10548
rect 18142 10160 18198 10169
rect 18142 10095 18198 10104
rect 18156 10062 18184 10095
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 17744 9820 18052 9840
rect 17744 9818 17750 9820
rect 17806 9818 17830 9820
rect 17886 9818 17910 9820
rect 17966 9818 17990 9820
rect 18046 9818 18052 9820
rect 17806 9766 17808 9818
rect 17988 9766 17990 9818
rect 17744 9764 17750 9766
rect 17806 9764 17830 9766
rect 17886 9764 17910 9766
rect 17966 9764 17990 9766
rect 18046 9764 18052 9766
rect 17744 9744 18052 9764
rect 18340 9722 18368 10542
rect 18524 10470 18552 10542
rect 18512 10464 18564 10470
rect 18512 10406 18564 10412
rect 18420 9988 18472 9994
rect 18420 9930 18472 9936
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 17408 9580 17460 9586
rect 17408 9522 17460 9528
rect 18432 9518 18460 9930
rect 18604 9920 18656 9926
rect 18604 9862 18656 9868
rect 18616 9586 18644 9862
rect 18708 9722 18736 10542
rect 18984 10062 19012 10610
rect 19076 10606 19104 10950
rect 19720 10810 19748 12582
rect 19812 12238 19840 12804
rect 19892 12776 19944 12782
rect 19892 12718 19944 12724
rect 19800 12232 19852 12238
rect 19800 12174 19852 12180
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19064 10600 19116 10606
rect 19064 10542 19116 10548
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18892 9654 18920 9930
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 18984 9586 19012 9998
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 17316 9512 17368 9518
rect 17316 9454 17368 9460
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 17328 9110 17356 9454
rect 17316 9104 17368 9110
rect 17316 9046 17368 9052
rect 18984 9042 19012 9522
rect 18972 9036 19024 9042
rect 18972 8978 19024 8984
rect 17744 8732 18052 8752
rect 17744 8730 17750 8732
rect 17806 8730 17830 8732
rect 17886 8730 17910 8732
rect 17966 8730 17990 8732
rect 18046 8730 18052 8732
rect 17806 8678 17808 8730
rect 17988 8678 17990 8730
rect 17744 8676 17750 8678
rect 17806 8676 17830 8678
rect 17886 8676 17910 8678
rect 17966 8676 17990 8678
rect 18046 8676 18052 8678
rect 17744 8656 18052 8676
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 18984 8498 19012 8978
rect 19076 8498 19104 10406
rect 19720 10062 19748 10746
rect 19904 10266 19932 12718
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 20076 12096 20128 12102
rect 20076 12038 20128 12044
rect 19996 11694 20024 12038
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19996 11558 20024 11630
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 20088 11370 20116 12038
rect 19996 11342 20116 11370
rect 19892 10260 19944 10266
rect 19892 10202 19944 10208
rect 19708 10056 19760 10062
rect 19708 9998 19760 10004
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 19248 8968 19300 8974
rect 19248 8910 19300 8916
rect 19444 8922 19472 9114
rect 19720 9110 19748 9998
rect 19996 9926 20024 11342
rect 20074 11248 20130 11257
rect 20074 11183 20130 11192
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19708 9104 19760 9110
rect 19708 9046 19760 9052
rect 19616 9036 19668 9042
rect 19616 8978 19668 8984
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 19064 8492 19116 8498
rect 19064 8434 19116 8440
rect 17512 7750 17540 8434
rect 17592 8356 17644 8362
rect 17592 8298 17644 8304
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 16856 7336 16908 7342
rect 16856 7278 16908 7284
rect 16764 7268 16816 7274
rect 16764 7210 16816 7216
rect 16672 6724 16724 6730
rect 16672 6666 16724 6672
rect 16776 6662 16804 7210
rect 17512 6866 17540 7686
rect 17604 7478 17632 8298
rect 18984 8090 19196 8106
rect 18984 8084 19208 8090
rect 18984 8078 19156 8084
rect 18984 7954 19012 8078
rect 19156 8026 19208 8032
rect 19260 7970 19288 8910
rect 19444 8906 19564 8922
rect 19444 8900 19576 8906
rect 19444 8894 19524 8900
rect 19338 8664 19394 8673
rect 19338 8599 19340 8608
rect 19392 8599 19394 8608
rect 19340 8570 19392 8576
rect 18604 7948 18656 7954
rect 18604 7890 18656 7896
rect 18972 7948 19024 7954
rect 18972 7890 19024 7896
rect 19168 7942 19288 7970
rect 17744 7644 18052 7664
rect 17744 7642 17750 7644
rect 17806 7642 17830 7644
rect 17886 7642 17910 7644
rect 17966 7642 17990 7644
rect 18046 7642 18052 7644
rect 17806 7590 17808 7642
rect 17988 7590 17990 7642
rect 17744 7588 17750 7590
rect 17806 7588 17830 7590
rect 17886 7588 17910 7590
rect 17966 7588 17990 7590
rect 18046 7588 18052 7590
rect 17744 7568 18052 7588
rect 17592 7472 17644 7478
rect 17592 7414 17644 7420
rect 18236 7336 18288 7342
rect 18236 7278 18288 7284
rect 17500 6860 17552 6866
rect 17500 6802 17552 6808
rect 18248 6798 18276 7278
rect 18616 7206 18644 7890
rect 18878 7848 18934 7857
rect 19168 7818 19196 7942
rect 19340 7880 19392 7886
rect 19306 7828 19340 7834
rect 19306 7822 19392 7828
rect 18878 7783 18934 7792
rect 19156 7812 19208 7818
rect 18604 7200 18656 7206
rect 18604 7142 18656 7148
rect 18616 6934 18644 7142
rect 18604 6928 18656 6934
rect 18604 6870 18656 6876
rect 18786 6896 18842 6905
rect 18420 6860 18472 6866
rect 18786 6831 18842 6840
rect 18420 6802 18472 6808
rect 17316 6792 17368 6798
rect 18236 6792 18288 6798
rect 17316 6734 17368 6740
rect 18142 6760 18198 6769
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16764 6656 16816 6662
rect 16764 6598 16816 6604
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16592 5370 16620 6598
rect 16960 6458 16988 6598
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 16948 6452 17000 6458
rect 16948 6394 17000 6400
rect 16670 5944 16726 5953
rect 16670 5879 16726 5888
rect 16684 5846 16712 5879
rect 16672 5840 16724 5846
rect 16672 5782 16724 5788
rect 16776 5778 16804 6394
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16764 5772 16816 5778
rect 16764 5714 16816 5720
rect 16764 5568 16816 5574
rect 16764 5510 16816 5516
rect 16488 5364 16540 5370
rect 16488 5306 16540 5312
rect 16580 5364 16632 5370
rect 16776 5352 16804 5510
rect 16580 5306 16632 5312
rect 16684 5324 16804 5352
rect 16684 5250 16712 5324
rect 16500 5222 16712 5250
rect 16960 5234 16988 6054
rect 17052 5370 17080 6258
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17040 5364 17092 5370
rect 17040 5306 17092 5312
rect 16948 5228 17000 5234
rect 16396 5160 16448 5166
rect 16302 5128 16358 5137
rect 16396 5102 16448 5108
rect 16302 5063 16358 5072
rect 16118 4992 16174 5001
rect 16118 4927 16174 4936
rect 15658 4720 15714 4729
rect 15476 4684 15528 4690
rect 15658 4655 15714 4664
rect 15476 4626 15528 4632
rect 15488 3738 15516 4626
rect 15566 4176 15622 4185
rect 15566 4111 15622 4120
rect 15580 3913 15608 4111
rect 15566 3904 15622 3913
rect 15566 3839 15622 3848
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15292 2576 15344 2582
rect 15292 2518 15344 2524
rect 15384 2576 15436 2582
rect 15384 2518 15436 2524
rect 14832 1964 14884 1970
rect 14832 1906 14884 1912
rect 15304 1834 15332 2518
rect 15488 2446 15516 3674
rect 15672 3058 15700 4655
rect 16408 4622 16436 5102
rect 16500 4826 16528 5222
rect 16948 5170 17000 5176
rect 16488 4820 16540 4826
rect 16488 4762 16540 4768
rect 16960 4690 16988 5170
rect 17144 4758 17172 6190
rect 17224 5636 17276 5642
rect 17224 5578 17276 5584
rect 17132 4752 17184 4758
rect 17132 4694 17184 4700
rect 16948 4684 17000 4690
rect 16948 4626 17000 4632
rect 17236 4622 17264 5578
rect 17328 5166 17356 6734
rect 18236 6734 18288 6740
rect 18142 6695 18144 6704
rect 18196 6695 18198 6704
rect 18144 6666 18196 6672
rect 17744 6556 18052 6576
rect 17744 6554 17750 6556
rect 17806 6554 17830 6556
rect 17886 6554 17910 6556
rect 17966 6554 17990 6556
rect 18046 6554 18052 6556
rect 17806 6502 17808 6554
rect 17988 6502 17990 6554
rect 17744 6500 17750 6502
rect 17806 6500 17830 6502
rect 17886 6500 17910 6502
rect 17966 6500 17990 6502
rect 18046 6500 18052 6502
rect 17744 6480 18052 6500
rect 18144 6384 18196 6390
rect 18142 6352 18144 6361
rect 18196 6352 18198 6361
rect 17500 6316 17552 6322
rect 18248 6322 18276 6734
rect 18142 6287 18198 6296
rect 18236 6316 18288 6322
rect 17500 6258 17552 6264
rect 18236 6258 18288 6264
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 17408 6112 17460 6118
rect 17408 6054 17460 6060
rect 17420 5710 17448 6054
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 16408 3534 16436 4558
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16856 4480 16908 4486
rect 16856 4422 16908 4428
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16592 4214 16620 4422
rect 16868 4282 16896 4422
rect 16856 4276 16908 4282
rect 16856 4218 16908 4224
rect 16580 4208 16632 4214
rect 16580 4150 16632 4156
rect 16960 3738 16988 4422
rect 17328 4078 17356 5102
rect 17512 5030 17540 6258
rect 18248 5710 18276 6258
rect 18236 5704 18288 5710
rect 18236 5646 18288 5652
rect 18144 5636 18196 5642
rect 18144 5578 18196 5584
rect 17592 5568 17644 5574
rect 17592 5510 17644 5516
rect 17604 5370 17632 5510
rect 17744 5468 18052 5488
rect 17744 5466 17750 5468
rect 17806 5466 17830 5468
rect 17886 5466 17910 5468
rect 17966 5466 17990 5468
rect 18046 5466 18052 5468
rect 17806 5414 17808 5466
rect 17988 5414 17990 5466
rect 17744 5412 17750 5414
rect 17806 5412 17830 5414
rect 17886 5412 17910 5414
rect 17966 5412 17990 5414
rect 18046 5412 18052 5414
rect 17744 5392 18052 5412
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17592 5160 17644 5166
rect 17592 5102 17644 5108
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17604 4690 17632 5102
rect 17592 4684 17644 4690
rect 17592 4626 17644 4632
rect 17696 4570 17724 5170
rect 18050 4992 18106 5001
rect 18050 4927 18106 4936
rect 18064 4826 18092 4927
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18156 4593 18184 5578
rect 18236 4752 18288 4758
rect 18236 4694 18288 4700
rect 17604 4542 17724 4570
rect 18142 4584 18198 4593
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17512 4146 17540 4422
rect 17604 4282 17632 4542
rect 18142 4519 18198 4528
rect 18248 4486 18276 4694
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 17744 4380 18052 4400
rect 17744 4378 17750 4380
rect 17806 4378 17830 4380
rect 17886 4378 17910 4380
rect 17966 4378 17990 4380
rect 18046 4378 18052 4380
rect 17806 4326 17808 4378
rect 17988 4326 17990 4378
rect 17744 4324 17750 4326
rect 17806 4324 17830 4326
rect 17886 4324 17910 4326
rect 17966 4324 17990 4326
rect 18046 4324 18052 4326
rect 17744 4304 18052 4324
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17868 4208 17920 4214
rect 17868 4150 17920 4156
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 17316 4072 17368 4078
rect 17316 4014 17368 4020
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 17696 3602 17724 4014
rect 17880 4010 17908 4150
rect 18340 4146 18368 6258
rect 18432 5574 18460 6802
rect 18604 6656 18656 6662
rect 18604 6598 18656 6604
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18420 5568 18472 5574
rect 18420 5510 18472 5516
rect 18432 4146 18460 5510
rect 18616 5370 18644 6598
rect 18708 5778 18736 6598
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18604 5364 18656 5370
rect 18604 5306 18656 5312
rect 18800 5098 18828 6831
rect 18892 5642 18920 7783
rect 19306 7806 19380 7822
rect 19306 7800 19334 7806
rect 19156 7754 19208 7760
rect 19260 7772 19334 7800
rect 18972 7744 19024 7750
rect 19260 7698 19288 7772
rect 18972 7686 19024 7692
rect 18984 7478 19012 7686
rect 19076 7670 19288 7698
rect 18972 7472 19024 7478
rect 18972 7414 19024 7420
rect 18880 5636 18932 5642
rect 18880 5578 18932 5584
rect 18880 5364 18932 5370
rect 18880 5306 18932 5312
rect 18788 5092 18840 5098
rect 18788 5034 18840 5040
rect 18892 4826 18920 5306
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18880 4820 18932 4826
rect 18880 4762 18932 4768
rect 18984 4758 19012 5170
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 19076 4604 19104 7670
rect 19338 7576 19394 7585
rect 19338 7511 19340 7520
rect 19392 7511 19394 7520
rect 19340 7482 19392 7488
rect 19340 7200 19392 7206
rect 19340 7142 19392 7148
rect 19156 6928 19208 6934
rect 19352 6905 19380 7142
rect 19156 6870 19208 6876
rect 19338 6896 19394 6905
rect 19168 6780 19196 6870
rect 19444 6866 19472 8894
rect 19524 8842 19576 8848
rect 19628 7274 19656 8978
rect 19616 7268 19668 7274
rect 19616 7210 19668 7216
rect 19338 6831 19394 6840
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 19168 6752 19380 6780
rect 19352 6610 19380 6752
rect 19444 6730 19472 6802
rect 19432 6724 19484 6730
rect 19432 6666 19484 6672
rect 19352 6582 19564 6610
rect 19340 6316 19392 6322
rect 19340 6258 19392 6264
rect 19352 5370 19380 6258
rect 19432 6112 19484 6118
rect 19432 6054 19484 6060
rect 19444 5778 19472 6054
rect 19432 5772 19484 5778
rect 19432 5714 19484 5720
rect 19340 5364 19392 5370
rect 19340 5306 19392 5312
rect 19536 5302 19564 6582
rect 19720 6254 19748 9046
rect 19996 7750 20024 9862
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 19812 7274 19840 7346
rect 19800 7268 19852 7274
rect 19800 7210 19852 7216
rect 19996 6458 20024 7686
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19708 6248 19760 6254
rect 19708 6190 19760 6196
rect 19892 5840 19944 5846
rect 19890 5808 19892 5817
rect 19944 5808 19946 5817
rect 19890 5743 19946 5752
rect 19708 5568 19760 5574
rect 19708 5510 19760 5516
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19248 5092 19300 5098
rect 19248 5034 19300 5040
rect 19260 4826 19288 5034
rect 19444 4826 19472 5170
rect 19614 5128 19670 5137
rect 19614 5063 19670 5072
rect 19248 4820 19300 4826
rect 19248 4762 19300 4768
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19524 4820 19576 4826
rect 19524 4762 19576 4768
rect 19444 4622 19472 4762
rect 18984 4576 19104 4604
rect 19432 4616 19484 4622
rect 18984 4146 19012 4576
rect 19432 4558 19484 4564
rect 19536 4486 19564 4762
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19156 4276 19208 4282
rect 19156 4218 19208 4224
rect 19062 4176 19118 4185
rect 18328 4140 18380 4146
rect 18328 4082 18380 4088
rect 18420 4140 18472 4146
rect 18420 4082 18472 4088
rect 18972 4140 19024 4146
rect 19062 4111 19118 4120
rect 18972 4082 19024 4088
rect 19076 4078 19104 4111
rect 19064 4072 19116 4078
rect 18984 4020 19064 4026
rect 18984 4014 19116 4020
rect 17868 4004 17920 4010
rect 17868 3946 17920 3952
rect 18984 3998 19104 4014
rect 17684 3596 17736 3602
rect 17684 3538 17736 3544
rect 16396 3528 16448 3534
rect 16396 3470 16448 3476
rect 16408 3058 16436 3470
rect 17696 3466 17724 3538
rect 18984 3534 19012 3998
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 18972 3528 19024 3534
rect 18972 3470 19024 3476
rect 17684 3460 17736 3466
rect 17684 3402 17736 3408
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 17408 3392 17460 3398
rect 17408 3334 17460 3340
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 16776 3058 16804 3334
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16580 3052 16632 3058
rect 16580 2994 16632 3000
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16224 2774 16252 2994
rect 16224 2746 16344 2774
rect 16210 2544 16266 2553
rect 16210 2479 16266 2488
rect 16224 2446 16252 2479
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16316 1902 16344 2746
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 16408 1970 16436 2518
rect 16592 2514 16620 2994
rect 17420 2854 17448 3334
rect 17744 3292 18052 3312
rect 17744 3290 17750 3292
rect 17806 3290 17830 3292
rect 17886 3290 17910 3292
rect 17966 3290 17990 3292
rect 18046 3290 18052 3292
rect 17806 3238 17808 3290
rect 17988 3238 17990 3290
rect 17744 3236 17750 3238
rect 17806 3236 17830 3238
rect 17886 3236 17910 3238
rect 17966 3236 17990 3238
rect 18046 3236 18052 3238
rect 17744 3216 18052 3236
rect 18156 2922 18184 3334
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 16580 2508 16632 2514
rect 16580 2450 16632 2456
rect 17040 2372 17092 2378
rect 17040 2314 17092 2320
rect 17052 2038 17080 2314
rect 17512 2106 17540 2586
rect 17744 2204 18052 2224
rect 17744 2202 17750 2204
rect 17806 2202 17830 2204
rect 17886 2202 17910 2204
rect 17966 2202 17990 2204
rect 18046 2202 18052 2204
rect 17806 2150 17808 2202
rect 17988 2150 17990 2202
rect 17744 2148 17750 2150
rect 17806 2148 17830 2150
rect 17886 2148 17910 2150
rect 17966 2148 17990 2150
rect 18046 2148 18052 2150
rect 17744 2128 18052 2148
rect 17500 2100 17552 2106
rect 17500 2042 17552 2048
rect 17040 2032 17092 2038
rect 18156 2009 18184 2858
rect 18248 2446 18276 3470
rect 18328 3392 18380 3398
rect 18328 3334 18380 3340
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 18236 2304 18288 2310
rect 18340 2292 18368 3334
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18288 2264 18368 2292
rect 18236 2246 18288 2252
rect 17040 1974 17092 1980
rect 18142 2000 18198 2009
rect 16396 1964 16448 1970
rect 18142 1935 18198 1944
rect 16396 1906 16448 1912
rect 16304 1896 16356 1902
rect 16304 1838 16356 1844
rect 15292 1828 15344 1834
rect 15292 1770 15344 1776
rect 18248 1766 18276 2246
rect 18432 1873 18460 2994
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 18984 2310 19012 2382
rect 18880 2304 18932 2310
rect 18880 2246 18932 2252
rect 18972 2304 19024 2310
rect 18972 2246 19024 2252
rect 18892 1902 18920 2246
rect 18880 1896 18932 1902
rect 18418 1864 18474 1873
rect 18880 1838 18932 1844
rect 18418 1799 18474 1808
rect 18236 1760 18288 1766
rect 18984 1737 19012 2246
rect 18236 1702 18288 1708
rect 18970 1728 19026 1737
rect 18970 1663 19026 1672
rect 2042 0 2098 800
rect 6090 0 6146 800
rect 10230 0 10286 800
rect 14278 0 14334 800
rect 18418 0 18474 800
rect 19076 377 19104 3878
rect 19168 2854 19196 4218
rect 19536 4196 19564 4422
rect 19628 4282 19656 5063
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 19444 4168 19564 4196
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19260 3097 19288 4082
rect 19444 3602 19472 4168
rect 19628 4026 19656 4218
rect 19536 3998 19656 4026
rect 19536 3913 19564 3998
rect 19616 3936 19668 3942
rect 19522 3904 19578 3913
rect 19616 3878 19668 3884
rect 19522 3839 19578 3848
rect 19432 3596 19484 3602
rect 19432 3538 19484 3544
rect 19628 3534 19656 3878
rect 19616 3528 19668 3534
rect 19616 3470 19668 3476
rect 19340 3120 19392 3126
rect 19246 3088 19302 3097
rect 19340 3062 19392 3068
rect 19246 3023 19302 3032
rect 19260 2922 19288 3023
rect 19248 2916 19300 2922
rect 19248 2858 19300 2864
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 19352 2514 19380 3062
rect 19720 2961 19748 5510
rect 19812 5098 20024 5114
rect 19800 5092 20036 5098
rect 19852 5086 19984 5092
rect 19800 5034 19852 5040
rect 19984 5034 20036 5040
rect 19892 5024 19944 5030
rect 19892 4966 19944 4972
rect 19904 4622 19932 4966
rect 19892 4616 19944 4622
rect 19892 4558 19944 4564
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 19812 4282 19840 4422
rect 19982 4312 20038 4321
rect 19800 4276 19852 4282
rect 19982 4247 20038 4256
rect 19800 4218 19852 4224
rect 19996 4010 20024 4247
rect 20088 4146 20116 11183
rect 20180 7954 20208 14062
rect 20732 14006 20760 14350
rect 20720 14000 20772 14006
rect 20720 13942 20772 13948
rect 20442 13832 20498 13841
rect 20442 13767 20498 13776
rect 20456 13433 20484 13767
rect 20543 13628 20851 13648
rect 20543 13626 20549 13628
rect 20605 13626 20629 13628
rect 20685 13626 20709 13628
rect 20765 13626 20789 13628
rect 20845 13626 20851 13628
rect 20605 13574 20607 13626
rect 20787 13574 20789 13626
rect 20543 13572 20549 13574
rect 20605 13572 20629 13574
rect 20685 13572 20709 13574
rect 20765 13572 20789 13574
rect 20845 13572 20851 13574
rect 20543 13552 20851 13572
rect 20442 13424 20498 13433
rect 20442 13359 20498 13368
rect 20456 13190 20484 13359
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20444 13184 20496 13190
rect 20444 13126 20496 13132
rect 20272 12306 20300 13126
rect 20456 12434 20484 13126
rect 20543 12540 20851 12560
rect 20543 12538 20549 12540
rect 20605 12538 20629 12540
rect 20685 12538 20709 12540
rect 20765 12538 20789 12540
rect 20845 12538 20851 12540
rect 20605 12486 20607 12538
rect 20787 12486 20789 12538
rect 20543 12484 20549 12486
rect 20605 12484 20629 12486
rect 20685 12484 20709 12486
rect 20765 12484 20789 12486
rect 20845 12484 20851 12486
rect 20543 12464 20851 12484
rect 20364 12406 20484 12434
rect 20260 12300 20312 12306
rect 20260 12242 20312 12248
rect 20364 11778 20392 12406
rect 20812 12096 20864 12102
rect 20812 12038 20864 12044
rect 20824 11898 20852 12038
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20272 11750 20392 11778
rect 20272 10554 20300 11750
rect 20352 11688 20404 11694
rect 20352 11630 20404 11636
rect 20364 11354 20392 11630
rect 20916 11558 20944 14350
rect 21192 13462 21220 14962
rect 21272 14000 21324 14006
rect 21272 13942 21324 13948
rect 21180 13456 21232 13462
rect 21180 13398 21232 13404
rect 21284 13394 21312 13942
rect 21088 13388 21140 13394
rect 21088 13330 21140 13336
rect 21272 13388 21324 13394
rect 21272 13330 21324 13336
rect 21100 12986 21128 13330
rect 21088 12980 21140 12986
rect 21088 12922 21140 12928
rect 20994 12880 21050 12889
rect 20994 12815 21050 12824
rect 20904 11552 20956 11558
rect 20904 11494 20956 11500
rect 20543 11452 20851 11472
rect 20543 11450 20549 11452
rect 20605 11450 20629 11452
rect 20685 11450 20709 11452
rect 20765 11450 20789 11452
rect 20845 11450 20851 11452
rect 20605 11398 20607 11450
rect 20787 11398 20789 11450
rect 20543 11396 20549 11398
rect 20605 11396 20629 11398
rect 20685 11396 20709 11398
rect 20765 11396 20789 11398
rect 20845 11396 20851 11398
rect 20543 11376 20851 11396
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20444 11280 20496 11286
rect 20916 11257 20944 11494
rect 21008 11354 21036 12815
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20444 11222 20496 11228
rect 20902 11248 20958 11257
rect 20272 10526 20392 10554
rect 20260 10464 20312 10470
rect 20260 10406 20312 10412
rect 20272 10062 20300 10406
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 20272 8634 20300 9998
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20260 8288 20312 8294
rect 20260 8230 20312 8236
rect 20168 7948 20220 7954
rect 20272 7936 20300 8230
rect 20364 8106 20392 10526
rect 20456 9110 20484 11222
rect 20902 11183 20958 11192
rect 21100 10674 21128 12922
rect 21284 12918 21312 13330
rect 21376 13258 21404 19314
rect 21456 19304 21508 19310
rect 21456 19246 21508 19252
rect 21468 18329 21496 19246
rect 21560 18426 21588 23800
rect 22006 22944 22062 22953
rect 22006 22879 22062 22888
rect 21916 22432 21968 22438
rect 21916 22374 21968 22380
rect 21928 22166 21956 22374
rect 21916 22160 21968 22166
rect 21916 22102 21968 22108
rect 21824 22024 21876 22030
rect 21824 21966 21876 21972
rect 21732 21888 21784 21894
rect 21732 21830 21784 21836
rect 21638 21584 21694 21593
rect 21638 21519 21640 21528
rect 21692 21519 21694 21528
rect 21640 21490 21692 21496
rect 21640 21140 21692 21146
rect 21640 21082 21692 21088
rect 21652 20466 21680 21082
rect 21640 20460 21692 20466
rect 21640 20402 21692 20408
rect 21638 20360 21694 20369
rect 21638 20295 21640 20304
rect 21692 20295 21694 20304
rect 21640 20266 21692 20272
rect 21652 19242 21680 20266
rect 21640 19236 21692 19242
rect 21640 19178 21692 19184
rect 21548 18420 21600 18426
rect 21548 18362 21600 18368
rect 21454 18320 21510 18329
rect 21454 18255 21456 18264
rect 21508 18255 21510 18264
rect 21456 18226 21508 18232
rect 21546 17776 21602 17785
rect 21456 17740 21508 17746
rect 21546 17711 21602 17720
rect 21456 17682 21508 17688
rect 21468 16658 21496 17682
rect 21560 17678 21588 17711
rect 21548 17672 21600 17678
rect 21548 17614 21600 17620
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 21744 16522 21772 21830
rect 21836 21486 21864 21966
rect 22020 21690 22048 22879
rect 22204 22250 22232 23800
rect 22204 22222 22324 22250
rect 22192 22092 22244 22098
rect 22192 22034 22244 22040
rect 22100 22024 22152 22030
rect 22100 21966 22152 21972
rect 22008 21684 22060 21690
rect 22008 21626 22060 21632
rect 22112 21593 22140 21966
rect 22098 21584 22154 21593
rect 22098 21519 22154 21528
rect 21824 21480 21876 21486
rect 21824 21422 21876 21428
rect 21824 21344 21876 21350
rect 21824 21286 21876 21292
rect 21836 18698 21864 21286
rect 21916 20868 21968 20874
rect 21916 20810 21968 20816
rect 21928 18970 21956 20810
rect 22006 20632 22062 20641
rect 22006 20567 22062 20576
rect 22020 20262 22048 20567
rect 22100 20392 22152 20398
rect 22100 20334 22152 20340
rect 22008 20256 22060 20262
rect 22008 20198 22060 20204
rect 22112 19718 22140 20334
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 22204 19530 22232 22034
rect 22296 20641 22324 22222
rect 22560 22228 22612 22234
rect 22560 22170 22612 22176
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 22282 20632 22338 20641
rect 22282 20567 22338 20576
rect 22284 20256 22336 20262
rect 22284 20198 22336 20204
rect 22112 19502 22232 19530
rect 22296 19514 22324 20198
rect 22284 19508 22336 19514
rect 21916 18964 21968 18970
rect 21916 18906 21968 18912
rect 21824 18692 21876 18698
rect 21824 18634 21876 18640
rect 22008 18624 22060 18630
rect 22008 18566 22060 18572
rect 21732 16516 21784 16522
rect 21732 16458 21784 16464
rect 21732 16244 21784 16250
rect 21732 16186 21784 16192
rect 21548 16108 21600 16114
rect 21600 16068 21680 16096
rect 21548 16050 21600 16056
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21548 15904 21600 15910
rect 21548 15846 21600 15852
rect 21468 14958 21496 15846
rect 21456 14952 21508 14958
rect 21456 14894 21508 14900
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 21468 13138 21496 13670
rect 21376 13110 21496 13138
rect 21272 12912 21324 12918
rect 21272 12854 21324 12860
rect 21180 11824 21232 11830
rect 21180 11766 21232 11772
rect 21192 11150 21220 11766
rect 21272 11620 21324 11626
rect 21272 11562 21324 11568
rect 21180 11144 21232 11150
rect 21180 11086 21232 11092
rect 21180 10736 21232 10742
rect 21180 10678 21232 10684
rect 21088 10668 21140 10674
rect 21088 10610 21140 10616
rect 20543 10364 20851 10384
rect 20543 10362 20549 10364
rect 20605 10362 20629 10364
rect 20685 10362 20709 10364
rect 20765 10362 20789 10364
rect 20845 10362 20851 10364
rect 20605 10310 20607 10362
rect 20787 10310 20789 10362
rect 20543 10308 20549 10310
rect 20605 10308 20629 10310
rect 20685 10308 20709 10310
rect 20765 10308 20789 10310
rect 20845 10308 20851 10310
rect 20543 10288 20851 10308
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 20543 9276 20851 9296
rect 20543 9274 20549 9276
rect 20605 9274 20629 9276
rect 20685 9274 20709 9276
rect 20765 9274 20789 9276
rect 20845 9274 20851 9276
rect 20605 9222 20607 9274
rect 20787 9222 20789 9274
rect 20543 9220 20549 9222
rect 20605 9220 20629 9222
rect 20685 9220 20709 9222
rect 20765 9220 20789 9222
rect 20845 9220 20851 9222
rect 20543 9200 20851 9220
rect 20444 9104 20496 9110
rect 20444 9046 20496 9052
rect 20456 8430 20484 9046
rect 20916 8514 20944 10202
rect 21192 9654 21220 10678
rect 21284 10538 21312 11562
rect 21272 10532 21324 10538
rect 21272 10474 21324 10480
rect 21180 9648 21232 9654
rect 21180 9590 21232 9596
rect 21376 9568 21404 13110
rect 21454 12880 21510 12889
rect 21560 12850 21588 15846
rect 21652 13938 21680 16068
rect 21744 14278 21772 16186
rect 22020 14414 22048 18566
rect 22112 17882 22140 19502
rect 22284 19450 22336 19456
rect 22282 19408 22338 19417
rect 22192 19372 22244 19378
rect 22282 19343 22338 19352
rect 22192 19314 22244 19320
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 22112 17338 22140 17818
rect 22204 17513 22232 19314
rect 22190 17504 22246 17513
rect 22190 17439 22246 17448
rect 22296 17338 22324 19343
rect 22100 17332 22152 17338
rect 22100 17274 22152 17280
rect 22284 17332 22336 17338
rect 22284 17274 22336 17280
rect 22100 15700 22152 15706
rect 22100 15642 22152 15648
rect 22112 15094 22140 15642
rect 22388 15434 22416 21830
rect 22468 21548 22520 21554
rect 22468 21490 22520 21496
rect 22480 18426 22508 21490
rect 22572 20058 22600 22170
rect 22744 22024 22796 22030
rect 22848 22001 22876 23800
rect 22744 21966 22796 21972
rect 22834 21992 22890 22001
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 22560 20052 22612 20058
rect 22560 19994 22612 20000
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22572 19417 22600 19654
rect 22558 19408 22614 19417
rect 22558 19343 22614 19352
rect 22664 18850 22692 21490
rect 22572 18822 22692 18850
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22572 17921 22600 18822
rect 22652 18760 22704 18766
rect 22652 18702 22704 18708
rect 22558 17912 22614 17921
rect 22558 17847 22614 17856
rect 22468 16108 22520 16114
rect 22468 16050 22520 16056
rect 22560 16108 22612 16114
rect 22560 16050 22612 16056
rect 22376 15428 22428 15434
rect 22376 15370 22428 15376
rect 22192 15360 22244 15366
rect 22192 15302 22244 15308
rect 22204 15162 22232 15302
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 22376 15020 22428 15026
rect 22376 14962 22428 14968
rect 22100 14816 22152 14822
rect 22100 14758 22152 14764
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 21732 14272 21784 14278
rect 21732 14214 21784 14220
rect 22112 14074 22140 14758
rect 22192 14612 22244 14618
rect 22192 14554 22244 14560
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 22204 13938 22232 14554
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22296 13938 22324 14214
rect 21640 13932 21692 13938
rect 21640 13874 21692 13880
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22388 13818 22416 14962
rect 22296 13790 22416 13818
rect 22008 13252 22060 13258
rect 22008 13194 22060 13200
rect 21824 13184 21876 13190
rect 21824 13126 21876 13132
rect 21836 12986 21864 13126
rect 21824 12980 21876 12986
rect 21824 12922 21876 12928
rect 21454 12815 21510 12824
rect 21548 12844 21600 12850
rect 21468 12442 21496 12815
rect 21548 12786 21600 12792
rect 21732 12844 21784 12850
rect 21732 12786 21784 12792
rect 21456 12436 21508 12442
rect 21456 12378 21508 12384
rect 21640 12368 21692 12374
rect 21640 12310 21692 12316
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21560 11762 21588 12242
rect 21548 11756 21600 11762
rect 21548 11698 21600 11704
rect 21652 11626 21680 12310
rect 21744 12306 21772 12786
rect 21824 12776 21876 12782
rect 21824 12718 21876 12724
rect 21732 12300 21784 12306
rect 21732 12242 21784 12248
rect 21836 12238 21864 12718
rect 22020 12434 22048 13194
rect 21928 12406 22048 12434
rect 22100 12436 22152 12442
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 21732 12164 21784 12170
rect 21732 12106 21784 12112
rect 21640 11620 21692 11626
rect 21640 11562 21692 11568
rect 21640 10464 21692 10470
rect 21640 10406 21692 10412
rect 21652 10198 21680 10406
rect 21640 10192 21692 10198
rect 21640 10134 21692 10140
rect 21548 9580 21600 9586
rect 21376 9540 21496 9568
rect 21180 9512 21232 9518
rect 21180 9454 21232 9460
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20824 8486 20944 8514
rect 20824 8430 20852 8486
rect 20444 8424 20496 8430
rect 20444 8366 20496 8372
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 20904 8424 20956 8430
rect 20904 8366 20956 8372
rect 20543 8188 20851 8208
rect 20543 8186 20549 8188
rect 20605 8186 20629 8188
rect 20685 8186 20709 8188
rect 20765 8186 20789 8188
rect 20845 8186 20851 8188
rect 20605 8134 20607 8186
rect 20787 8134 20789 8186
rect 20543 8132 20549 8134
rect 20605 8132 20629 8134
rect 20685 8132 20709 8134
rect 20765 8132 20789 8134
rect 20845 8132 20851 8134
rect 20543 8112 20851 8132
rect 20364 8078 20484 8106
rect 20916 8090 20944 8366
rect 20272 7908 20392 7936
rect 20168 7890 20220 7896
rect 20180 7546 20208 7890
rect 20168 7540 20220 7546
rect 20168 7482 20220 7488
rect 20364 7342 20392 7908
rect 20168 7336 20220 7342
rect 20168 7278 20220 7284
rect 20352 7336 20404 7342
rect 20352 7278 20404 7284
rect 20180 7002 20208 7278
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 20168 6996 20220 7002
rect 20168 6938 20220 6944
rect 20272 6882 20300 7210
rect 20180 6854 20300 6882
rect 20180 6118 20208 6854
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 20260 6112 20312 6118
rect 20260 6054 20312 6060
rect 20076 4140 20128 4146
rect 20076 4082 20128 4088
rect 19984 4004 20036 4010
rect 19984 3946 20036 3952
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19812 3738 19840 3878
rect 19800 3732 19852 3738
rect 19800 3674 19852 3680
rect 19706 2952 19762 2961
rect 19706 2887 19762 2896
rect 20180 2774 20208 6054
rect 20272 5914 20300 6054
rect 20260 5908 20312 5914
rect 20260 5850 20312 5856
rect 20260 5636 20312 5642
rect 20260 5578 20312 5584
rect 20272 5370 20300 5578
rect 20260 5364 20312 5370
rect 20260 5306 20312 5312
rect 20456 4729 20484 8078
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20824 7546 20852 7686
rect 20812 7540 20864 7546
rect 20864 7500 20944 7528
rect 20812 7482 20864 7488
rect 20543 7100 20851 7120
rect 20543 7098 20549 7100
rect 20605 7098 20629 7100
rect 20685 7098 20709 7100
rect 20765 7098 20789 7100
rect 20845 7098 20851 7100
rect 20605 7046 20607 7098
rect 20787 7046 20789 7098
rect 20543 7044 20549 7046
rect 20605 7044 20629 7046
rect 20685 7044 20709 7046
rect 20765 7044 20789 7046
rect 20845 7044 20851 7046
rect 20543 7024 20851 7044
rect 20812 6928 20864 6934
rect 20812 6870 20864 6876
rect 20824 6798 20852 6870
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20916 6322 20944 7500
rect 20904 6316 20956 6322
rect 20904 6258 20956 6264
rect 20543 6012 20851 6032
rect 20543 6010 20549 6012
rect 20605 6010 20629 6012
rect 20685 6010 20709 6012
rect 20765 6010 20789 6012
rect 20845 6010 20851 6012
rect 20605 5958 20607 6010
rect 20787 5958 20789 6010
rect 20543 5956 20549 5958
rect 20605 5956 20629 5958
rect 20685 5956 20709 5958
rect 20765 5956 20789 5958
rect 20845 5956 20851 5958
rect 20543 5936 20851 5956
rect 21008 5794 21036 9318
rect 21088 9104 21140 9110
rect 21088 9046 21140 9052
rect 20732 5766 21036 5794
rect 20732 5710 20760 5766
rect 20720 5704 20772 5710
rect 20720 5646 20772 5652
rect 20543 4924 20851 4944
rect 20543 4922 20549 4924
rect 20605 4922 20629 4924
rect 20685 4922 20709 4924
rect 20765 4922 20789 4924
rect 20845 4922 20851 4924
rect 20605 4870 20607 4922
rect 20787 4870 20789 4922
rect 20543 4868 20549 4870
rect 20605 4868 20629 4870
rect 20685 4868 20709 4870
rect 20765 4868 20789 4870
rect 20845 4868 20851 4870
rect 20543 4848 20851 4868
rect 20442 4720 20498 4729
rect 21100 4690 21128 9046
rect 21192 8634 21220 9454
rect 21364 9444 21416 9450
rect 21364 9386 21416 9392
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21376 8498 21404 9386
rect 21468 9382 21496 9540
rect 21548 9522 21600 9528
rect 21456 9376 21508 9382
rect 21456 9318 21508 9324
rect 21560 9178 21588 9522
rect 21548 9172 21600 9178
rect 21548 9114 21600 9120
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21548 8424 21600 8430
rect 21548 8366 21600 8372
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 21192 7886 21220 8298
rect 21362 8256 21418 8265
rect 21362 8191 21418 8200
rect 21376 8090 21404 8191
rect 21364 8084 21416 8090
rect 21364 8026 21416 8032
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21272 7880 21324 7886
rect 21272 7822 21324 7828
rect 21180 6792 21232 6798
rect 21284 6780 21312 7822
rect 21364 7812 21416 7818
rect 21364 7754 21416 7760
rect 21376 7546 21404 7754
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21560 7478 21588 8366
rect 21548 7472 21600 7478
rect 21548 7414 21600 7420
rect 21546 7304 21602 7313
rect 21546 7239 21602 7248
rect 21232 6752 21312 6780
rect 21454 6760 21510 6769
rect 21180 6734 21232 6740
rect 21192 5710 21220 6734
rect 21560 6730 21588 7239
rect 21454 6695 21456 6704
rect 21508 6695 21510 6704
rect 21548 6724 21600 6730
rect 21456 6666 21508 6672
rect 21548 6666 21600 6672
rect 21456 5908 21508 5914
rect 21456 5850 21508 5856
rect 21180 5704 21232 5710
rect 21180 5646 21232 5652
rect 21192 4690 21220 5646
rect 21270 4720 21326 4729
rect 20442 4655 20498 4664
rect 21088 4684 21140 4690
rect 21088 4626 21140 4632
rect 21180 4684 21232 4690
rect 21468 4706 21496 5850
rect 21548 5704 21600 5710
rect 21548 5646 21600 5652
rect 21560 5137 21588 5646
rect 21652 5234 21680 10134
rect 21744 9602 21772 12106
rect 21836 10266 21864 12174
rect 21928 10577 21956 12406
rect 22100 12378 22152 12384
rect 22112 11898 22140 12378
rect 22296 12238 22324 13790
rect 22376 13728 22428 13734
rect 22376 13670 22428 13676
rect 22388 12850 22416 13670
rect 22480 13530 22508 16050
rect 22572 14006 22600 16050
rect 22664 15706 22692 18702
rect 22756 16454 22784 21966
rect 22834 21927 22890 21936
rect 22928 21956 22980 21962
rect 22928 21898 22980 21904
rect 22836 21344 22888 21350
rect 22836 21286 22888 21292
rect 22848 19378 22876 21286
rect 22836 19372 22888 19378
rect 22836 19314 22888 19320
rect 22940 19258 22968 21898
rect 23020 20460 23072 20466
rect 23020 20402 23072 20408
rect 23032 20369 23060 20402
rect 23018 20360 23074 20369
rect 23018 20295 23074 20304
rect 23020 20256 23072 20262
rect 23020 20198 23072 20204
rect 23110 20224 23166 20233
rect 23032 19825 23060 20198
rect 23110 20159 23166 20168
rect 23018 19816 23074 19825
rect 23018 19751 23074 19760
rect 23020 19712 23072 19718
rect 23020 19654 23072 19660
rect 23032 19553 23060 19654
rect 23018 19544 23074 19553
rect 23018 19479 23074 19488
rect 22940 19230 23060 19258
rect 22928 19168 22980 19174
rect 22928 19110 22980 19116
rect 22834 18864 22890 18873
rect 22834 18799 22890 18808
rect 22848 18766 22876 18799
rect 22836 18760 22888 18766
rect 22836 18702 22888 18708
rect 22940 18426 22968 19110
rect 22928 18420 22980 18426
rect 22928 18362 22980 18368
rect 23032 18306 23060 19230
rect 23124 18970 23152 20159
rect 23216 19514 23244 24239
rect 23478 23800 23534 24600
rect 24122 23800 24178 24600
rect 23492 21604 23520 23800
rect 24136 21622 24164 23800
rect 23400 21576 23520 21604
rect 24124 21616 24176 21622
rect 23400 20534 23428 21576
rect 24124 21558 24176 21564
rect 23480 21480 23532 21486
rect 23480 21422 23532 21428
rect 23388 20528 23440 20534
rect 23388 20470 23440 20476
rect 23296 20460 23348 20466
rect 23296 20402 23348 20408
rect 23204 19508 23256 19514
rect 23204 19450 23256 19456
rect 23112 18964 23164 18970
rect 23112 18906 23164 18912
rect 23308 18578 23336 20402
rect 22848 18278 23060 18306
rect 23124 18550 23336 18578
rect 22848 17377 22876 18278
rect 22928 18216 22980 18222
rect 22928 18158 22980 18164
rect 22940 17542 22968 18158
rect 23020 18080 23072 18086
rect 23020 18022 23072 18028
rect 22928 17536 22980 17542
rect 22928 17478 22980 17484
rect 22834 17368 22890 17377
rect 22834 17303 22890 17312
rect 22836 17264 22888 17270
rect 22834 17232 22836 17241
rect 22888 17232 22890 17241
rect 22834 17167 22890 17176
rect 22940 17134 22968 17478
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22928 16448 22980 16454
rect 22928 16390 22980 16396
rect 22756 16182 22784 16390
rect 22834 16280 22890 16289
rect 22834 16215 22890 16224
rect 22744 16176 22796 16182
rect 22744 16118 22796 16124
rect 22652 15700 22704 15706
rect 22652 15642 22704 15648
rect 22664 14958 22692 15642
rect 22848 15502 22876 16215
rect 22940 16153 22968 16390
rect 23032 16289 23060 18022
rect 23018 16280 23074 16289
rect 23018 16215 23074 16224
rect 22926 16144 22982 16153
rect 22926 16079 22982 16088
rect 23124 15994 23152 18550
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 23204 16992 23256 16998
rect 23204 16934 23256 16940
rect 22940 15966 23152 15994
rect 22744 15496 22796 15502
rect 22744 15438 22796 15444
rect 22836 15496 22888 15502
rect 22836 15438 22888 15444
rect 22940 15450 22968 15966
rect 23112 15904 23164 15910
rect 23112 15846 23164 15852
rect 22652 14952 22704 14958
rect 22652 14894 22704 14900
rect 22652 14272 22704 14278
rect 22652 14214 22704 14220
rect 22664 14074 22692 14214
rect 22652 14068 22704 14074
rect 22652 14010 22704 14016
rect 22560 14000 22612 14006
rect 22560 13942 22612 13948
rect 22560 13864 22612 13870
rect 22560 13806 22612 13812
rect 22572 13569 22600 13806
rect 22756 13734 22784 15438
rect 22940 15422 23060 15450
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22940 13977 22968 15302
rect 22926 13968 22982 13977
rect 22926 13903 22982 13912
rect 22836 13796 22888 13802
rect 22836 13738 22888 13744
rect 22744 13728 22796 13734
rect 22744 13670 22796 13676
rect 22558 13560 22614 13569
rect 22468 13524 22520 13530
rect 22848 13530 22876 13738
rect 22928 13728 22980 13734
rect 22928 13670 22980 13676
rect 22558 13495 22614 13504
rect 22836 13524 22888 13530
rect 22468 13466 22520 13472
rect 22376 12844 22428 12850
rect 22376 12786 22428 12792
rect 22284 12232 22336 12238
rect 22284 12174 22336 12180
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22100 11688 22152 11694
rect 22100 11630 22152 11636
rect 22112 11286 22140 11630
rect 22100 11280 22152 11286
rect 22100 11222 22152 11228
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 21914 10568 21970 10577
rect 21914 10503 21970 10512
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21916 10260 21968 10266
rect 21916 10202 21968 10208
rect 21928 10169 21956 10202
rect 21914 10160 21970 10169
rect 21824 10124 21876 10130
rect 21914 10095 21970 10104
rect 21824 10066 21876 10072
rect 21836 9722 21864 10066
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 22112 9654 22140 9862
rect 22100 9648 22152 9654
rect 21744 9574 21864 9602
rect 22100 9590 22152 9596
rect 21836 9466 21864 9574
rect 21732 9444 21784 9450
rect 21836 9438 22048 9466
rect 21732 9386 21784 9392
rect 21744 9178 21772 9386
rect 21732 9172 21784 9178
rect 21732 9114 21784 9120
rect 21824 8900 21876 8906
rect 21824 8842 21876 8848
rect 21732 8492 21784 8498
rect 21732 8434 21784 8440
rect 21744 8294 21772 8434
rect 21732 8288 21784 8294
rect 21732 8230 21784 8236
rect 21732 7200 21784 7206
rect 21732 7142 21784 7148
rect 21744 5302 21772 7142
rect 21836 5370 21864 8842
rect 21916 6724 21968 6730
rect 21916 6666 21968 6672
rect 21928 6254 21956 6666
rect 21916 6248 21968 6254
rect 21916 6190 21968 6196
rect 22020 6066 22048 9438
rect 22204 7546 22232 11086
rect 22388 10130 22416 12786
rect 22480 12782 22508 13466
rect 22468 12776 22520 12782
rect 22468 12718 22520 12724
rect 22572 12646 22600 13495
rect 22836 13466 22888 13472
rect 22652 13320 22704 13326
rect 22652 13262 22704 13268
rect 22664 12986 22692 13262
rect 22940 13258 22968 13670
rect 22928 13252 22980 13258
rect 22928 13194 22980 13200
rect 22652 12980 22704 12986
rect 22652 12922 22704 12928
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 22560 12640 22612 12646
rect 22560 12582 22612 12588
rect 22848 12345 22876 12786
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 22834 12336 22890 12345
rect 22834 12271 22890 12280
rect 22468 12164 22520 12170
rect 22468 12106 22520 12112
rect 22480 10810 22508 12106
rect 22652 11552 22704 11558
rect 22652 11494 22704 11500
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22376 10124 22428 10130
rect 22376 10066 22428 10072
rect 22572 9722 22600 10542
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22560 8832 22612 8838
rect 22560 8774 22612 8780
rect 22572 8498 22600 8774
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22284 7812 22336 7818
rect 22284 7754 22336 7760
rect 22192 7540 22244 7546
rect 22192 7482 22244 7488
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22100 7268 22152 7274
rect 22100 7210 22152 7216
rect 22112 7002 22140 7210
rect 22204 7002 22232 7346
rect 22100 6996 22152 7002
rect 22100 6938 22152 6944
rect 22192 6996 22244 7002
rect 22192 6938 22244 6944
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 21928 6038 22048 6066
rect 21824 5364 21876 5370
rect 21824 5306 21876 5312
rect 21732 5296 21784 5302
rect 21732 5238 21784 5244
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 21824 5160 21876 5166
rect 21546 5128 21602 5137
rect 21824 5102 21876 5108
rect 21546 5063 21602 5072
rect 21732 5092 21784 5098
rect 21732 5034 21784 5040
rect 21640 5024 21692 5030
rect 21546 4992 21602 5001
rect 21640 4966 21692 4972
rect 21546 4927 21602 4936
rect 21560 4826 21588 4927
rect 21548 4820 21600 4826
rect 21548 4762 21600 4768
rect 21468 4678 21588 4706
rect 21270 4655 21326 4664
rect 21180 4626 21232 4632
rect 20904 4616 20956 4622
rect 20904 4558 20956 4564
rect 20352 4208 20404 4214
rect 20352 4150 20404 4156
rect 20260 4072 20312 4078
rect 20364 4049 20392 4150
rect 20260 4014 20312 4020
rect 20350 4040 20406 4049
rect 20272 3602 20300 4014
rect 20350 3975 20406 3984
rect 20543 3836 20851 3856
rect 20543 3834 20549 3836
rect 20605 3834 20629 3836
rect 20685 3834 20709 3836
rect 20765 3834 20789 3836
rect 20845 3834 20851 3836
rect 20605 3782 20607 3834
rect 20787 3782 20789 3834
rect 20543 3780 20549 3782
rect 20605 3780 20629 3782
rect 20685 3780 20709 3782
rect 20765 3780 20789 3782
rect 20845 3780 20851 3782
rect 20543 3760 20851 3780
rect 20534 3632 20590 3641
rect 20260 3596 20312 3602
rect 20534 3567 20590 3576
rect 20260 3538 20312 3544
rect 20548 3466 20576 3567
rect 20718 3496 20774 3505
rect 20536 3460 20588 3466
rect 20718 3431 20720 3440
rect 20536 3402 20588 3408
rect 20772 3431 20774 3440
rect 20720 3402 20772 3408
rect 20810 3224 20866 3233
rect 20810 3159 20812 3168
rect 20864 3159 20866 3168
rect 20812 3130 20864 3136
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20180 2746 20392 2774
rect 20364 2514 20392 2746
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 20352 2508 20404 2514
rect 20352 2450 20404 2456
rect 20456 2446 20484 2994
rect 20543 2748 20851 2768
rect 20543 2746 20549 2748
rect 20605 2746 20629 2748
rect 20685 2746 20709 2748
rect 20765 2746 20789 2748
rect 20845 2746 20851 2748
rect 20605 2694 20607 2746
rect 20787 2694 20789 2746
rect 20543 2692 20549 2694
rect 20605 2692 20629 2694
rect 20685 2692 20709 2694
rect 20765 2692 20789 2694
rect 20845 2692 20851 2694
rect 20543 2672 20851 2692
rect 20916 2582 20944 4558
rect 21088 4548 21140 4554
rect 21088 4490 21140 4496
rect 20996 4480 21048 4486
rect 20996 4422 21048 4428
rect 21008 4214 21036 4422
rect 20996 4208 21048 4214
rect 20996 4150 21048 4156
rect 21100 2854 21128 4490
rect 21192 3618 21220 4626
rect 21284 4622 21312 4655
rect 21272 4616 21324 4622
rect 21456 4616 21508 4622
rect 21272 4558 21324 4564
rect 21454 4584 21456 4593
rect 21508 4584 21510 4593
rect 21454 4519 21510 4528
rect 21364 4208 21416 4214
rect 21270 4176 21326 4185
rect 21364 4150 21416 4156
rect 21456 4208 21508 4214
rect 21456 4150 21508 4156
rect 21270 4111 21326 4120
rect 21284 4078 21312 4111
rect 21272 4072 21324 4078
rect 21272 4014 21324 4020
rect 21192 3590 21312 3618
rect 21192 3126 21220 3590
rect 21284 3534 21312 3590
rect 21272 3528 21324 3534
rect 21272 3470 21324 3476
rect 21272 3392 21324 3398
rect 21272 3334 21324 3340
rect 21180 3120 21232 3126
rect 21180 3062 21232 3068
rect 21284 3058 21312 3334
rect 21376 3194 21404 4150
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21362 3088 21418 3097
rect 21272 3052 21324 3058
rect 21468 3074 21496 4150
rect 21560 3890 21588 4678
rect 21652 4214 21680 4966
rect 21744 4554 21772 5034
rect 21732 4548 21784 4554
rect 21732 4490 21784 4496
rect 21640 4208 21692 4214
rect 21640 4150 21692 4156
rect 21732 3936 21784 3942
rect 21560 3884 21732 3890
rect 21560 3878 21784 3884
rect 21560 3862 21772 3878
rect 21560 3126 21588 3862
rect 21640 3392 21692 3398
rect 21640 3334 21692 3340
rect 21418 3046 21496 3074
rect 21548 3120 21600 3126
rect 21548 3062 21600 3068
rect 21362 3023 21364 3032
rect 21272 2994 21324 3000
rect 21416 3023 21418 3032
rect 21364 2994 21416 3000
rect 21088 2848 21140 2854
rect 21088 2790 21140 2796
rect 21548 2848 21600 2854
rect 21548 2790 21600 2796
rect 20720 2576 20772 2582
rect 20720 2518 20772 2524
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 20444 2440 20496 2446
rect 19338 2408 19394 2417
rect 20444 2382 20496 2388
rect 20732 2394 20760 2518
rect 19338 2343 19340 2352
rect 19392 2343 19394 2352
rect 20732 2378 20852 2394
rect 20732 2372 20864 2378
rect 20732 2366 20812 2372
rect 19340 2314 19392 2320
rect 20166 2272 20222 2281
rect 20166 2207 20222 2216
rect 20180 1834 20208 2207
rect 20732 2038 20760 2366
rect 20812 2314 20864 2320
rect 20720 2032 20772 2038
rect 20720 1974 20772 1980
rect 20260 1964 20312 1970
rect 20260 1906 20312 1912
rect 20168 1828 20220 1834
rect 20168 1770 20220 1776
rect 20272 1601 20300 1906
rect 20258 1592 20314 1601
rect 20258 1527 20314 1536
rect 21560 921 21588 2790
rect 21652 2310 21680 3334
rect 21836 2310 21864 5102
rect 21928 2446 21956 6038
rect 22100 5636 22152 5642
rect 22100 5578 22152 5584
rect 22008 4004 22060 4010
rect 22008 3946 22060 3952
rect 22020 2514 22048 3946
rect 22112 2990 22140 5578
rect 22204 5370 22232 6734
rect 22296 6390 22324 7754
rect 22376 7336 22428 7342
rect 22376 7278 22428 7284
rect 22388 6458 22416 7278
rect 22376 6452 22428 6458
rect 22376 6394 22428 6400
rect 22284 6384 22336 6390
rect 22284 6326 22336 6332
rect 22296 6225 22324 6326
rect 22282 6216 22338 6225
rect 22282 6151 22338 6160
rect 22282 5808 22338 5817
rect 22282 5743 22338 5752
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22296 5166 22324 5743
rect 22376 5568 22428 5574
rect 22376 5510 22428 5516
rect 22284 5160 22336 5166
rect 22284 5102 22336 5108
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 22388 2582 22416 5510
rect 22468 4208 22520 4214
rect 22468 4150 22520 4156
rect 22480 2990 22508 4150
rect 22572 3210 22600 8434
rect 22664 7449 22692 11494
rect 22848 10198 22876 12271
rect 22836 10192 22888 10198
rect 22836 10134 22888 10140
rect 22836 9580 22888 9586
rect 22836 9522 22888 9528
rect 22744 8560 22796 8566
rect 22744 8502 22796 8508
rect 22756 7750 22784 8502
rect 22848 8090 22876 9522
rect 22940 8945 22968 12582
rect 23032 12209 23060 15422
rect 23124 14414 23152 15846
rect 23216 15026 23244 16934
rect 23204 15020 23256 15026
rect 23204 14962 23256 14968
rect 23216 14929 23244 14962
rect 23202 14920 23258 14929
rect 23202 14855 23258 14864
rect 23112 14408 23164 14414
rect 23112 14350 23164 14356
rect 23124 14249 23152 14350
rect 23110 14240 23166 14249
rect 23110 14175 23166 14184
rect 23112 13320 23164 13326
rect 23110 13288 23112 13297
rect 23164 13288 23166 13297
rect 23110 13223 23166 13232
rect 23018 12200 23074 12209
rect 23018 12135 23074 12144
rect 23020 12096 23072 12102
rect 23020 12038 23072 12044
rect 23032 11694 23060 12038
rect 23112 11756 23164 11762
rect 23112 11698 23164 11704
rect 23020 11688 23072 11694
rect 23124 11665 23152 11698
rect 23020 11630 23072 11636
rect 23110 11656 23166 11665
rect 23110 11591 23166 11600
rect 23124 11354 23152 11591
rect 23112 11348 23164 11354
rect 23112 11290 23164 11296
rect 23204 11280 23256 11286
rect 23204 11222 23256 11228
rect 23112 11144 23164 11150
rect 23112 11086 23164 11092
rect 23020 11008 23072 11014
rect 23124 10985 23152 11086
rect 23020 10950 23072 10956
rect 23110 10976 23166 10985
rect 23032 10305 23060 10950
rect 23110 10911 23166 10920
rect 23018 10296 23074 10305
rect 23018 10231 23074 10240
rect 23032 10062 23060 10231
rect 23020 10056 23072 10062
rect 23020 9998 23072 10004
rect 23124 9654 23152 10911
rect 23112 9648 23164 9654
rect 23112 9590 23164 9596
rect 23112 9512 23164 9518
rect 23112 9454 23164 9460
rect 22926 8936 22982 8945
rect 22926 8871 22982 8880
rect 23124 8838 23152 9454
rect 23112 8832 23164 8838
rect 23112 8774 23164 8780
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22650 7440 22706 7449
rect 22650 7375 22706 7384
rect 22756 7342 22784 7686
rect 22928 7472 22980 7478
rect 22928 7414 22980 7420
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 22652 6792 22704 6798
rect 22652 6734 22704 6740
rect 22664 3738 22692 6734
rect 22756 4214 22784 7142
rect 22940 5778 22968 7414
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 23032 6905 23060 7346
rect 23018 6896 23074 6905
rect 23018 6831 23074 6840
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 23032 6361 23060 6598
rect 23018 6352 23074 6361
rect 23124 6322 23152 8774
rect 23018 6287 23074 6296
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 22928 5772 22980 5778
rect 22928 5714 22980 5720
rect 23032 5681 23060 6054
rect 22834 5672 22890 5681
rect 22834 5607 22890 5616
rect 23018 5672 23074 5681
rect 23018 5607 23074 5616
rect 22848 5234 22876 5607
rect 23216 5302 23244 11222
rect 23308 10810 23336 17614
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23400 15609 23428 16526
rect 23386 15600 23442 15609
rect 23386 15535 23442 15544
rect 23492 15162 23520 21422
rect 23572 19848 23624 19854
rect 23572 19790 23624 19796
rect 23480 15156 23532 15162
rect 23480 15098 23532 15104
rect 23584 11218 23612 19790
rect 23664 19440 23716 19446
rect 23664 19382 23716 19388
rect 23676 14618 23704 19382
rect 23754 18592 23810 18601
rect 23754 18527 23810 18536
rect 23664 14612 23716 14618
rect 23664 14554 23716 14560
rect 23768 13530 23796 18527
rect 23938 16552 23994 16561
rect 23938 16487 23994 16496
rect 23756 13524 23808 13530
rect 23756 13466 23808 13472
rect 23572 11212 23624 11218
rect 23572 11154 23624 11160
rect 23296 10804 23348 10810
rect 23296 10746 23348 10752
rect 23952 10674 23980 16487
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 23294 9616 23350 9625
rect 23294 9551 23350 9560
rect 23308 8673 23336 9551
rect 23386 8936 23442 8945
rect 23386 8871 23442 8880
rect 23294 8664 23350 8673
rect 23294 8599 23350 8608
rect 23308 7886 23336 8599
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 23400 6866 23428 8871
rect 23388 6860 23440 6866
rect 23388 6802 23440 6808
rect 23204 5296 23256 5302
rect 23204 5238 23256 5244
rect 22836 5228 22888 5234
rect 22836 5170 22888 5176
rect 22744 4208 22796 4214
rect 22744 4150 22796 4156
rect 22848 3738 22876 5170
rect 23112 5024 23164 5030
rect 23112 4966 23164 4972
rect 23020 4480 23072 4486
rect 23020 4422 23072 4428
rect 23032 4146 23060 4422
rect 23020 4140 23072 4146
rect 23020 4082 23072 4088
rect 22652 3732 22704 3738
rect 22652 3674 22704 3680
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 22742 3632 22798 3641
rect 22742 3567 22798 3576
rect 22650 3224 22706 3233
rect 22572 3182 22650 3210
rect 22650 3159 22706 3168
rect 22664 3058 22692 3159
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 22468 2984 22520 2990
rect 22468 2926 22520 2932
rect 22756 2582 22784 3567
rect 22836 2984 22888 2990
rect 22836 2926 22888 2932
rect 22848 2650 22876 2926
rect 22836 2644 22888 2650
rect 22836 2586 22888 2592
rect 22376 2576 22428 2582
rect 22376 2518 22428 2524
rect 22744 2576 22796 2582
rect 22744 2518 22796 2524
rect 22008 2508 22060 2514
rect 22008 2450 22060 2456
rect 23124 2446 23152 4966
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 23112 2440 23164 2446
rect 23112 2382 23164 2388
rect 21640 2304 21692 2310
rect 21640 2246 21692 2252
rect 21824 2304 21876 2310
rect 21824 2246 21876 2252
rect 22468 2100 22520 2106
rect 22468 2042 22520 2048
rect 21546 912 21602 921
rect 21546 847 21602 856
rect 22480 800 22508 2042
rect 19062 368 19118 377
rect 19062 303 19118 312
rect 22466 0 22522 800
<< via2 >>
rect 1582 15272 1638 15328
rect 1398 9152 1454 9208
rect 3755 22330 3811 22332
rect 3835 22330 3891 22332
rect 3915 22330 3971 22332
rect 3995 22330 4051 22332
rect 3755 22278 3801 22330
rect 3801 22278 3811 22330
rect 3835 22278 3865 22330
rect 3865 22278 3877 22330
rect 3877 22278 3891 22330
rect 3915 22278 3929 22330
rect 3929 22278 3941 22330
rect 3941 22278 3971 22330
rect 3995 22278 4005 22330
rect 4005 22278 4051 22330
rect 3755 22276 3811 22278
rect 3835 22276 3891 22278
rect 3915 22276 3971 22278
rect 3995 22276 4051 22278
rect 3755 21242 3811 21244
rect 3835 21242 3891 21244
rect 3915 21242 3971 21244
rect 3995 21242 4051 21244
rect 3755 21190 3801 21242
rect 3801 21190 3811 21242
rect 3835 21190 3865 21242
rect 3865 21190 3877 21242
rect 3877 21190 3891 21242
rect 3915 21190 3929 21242
rect 3929 21190 3941 21242
rect 3941 21190 3971 21242
rect 3995 21190 4005 21242
rect 4005 21190 4051 21242
rect 3755 21188 3811 21190
rect 3835 21188 3891 21190
rect 3915 21188 3971 21190
rect 3995 21188 4051 21190
rect 3422 19236 3478 19272
rect 3422 19216 3424 19236
rect 3424 19216 3476 19236
rect 3476 19216 3478 19236
rect 3755 20154 3811 20156
rect 3835 20154 3891 20156
rect 3915 20154 3971 20156
rect 3995 20154 4051 20156
rect 3755 20102 3801 20154
rect 3801 20102 3811 20154
rect 3835 20102 3865 20154
rect 3865 20102 3877 20154
rect 3877 20102 3891 20154
rect 3915 20102 3929 20154
rect 3929 20102 3941 20154
rect 3941 20102 3971 20154
rect 3995 20102 4005 20154
rect 4005 20102 4051 20154
rect 3755 20100 3811 20102
rect 3835 20100 3891 20102
rect 3915 20100 3971 20102
rect 3995 20100 4051 20102
rect 3755 19066 3811 19068
rect 3835 19066 3891 19068
rect 3915 19066 3971 19068
rect 3995 19066 4051 19068
rect 3755 19014 3801 19066
rect 3801 19014 3811 19066
rect 3835 19014 3865 19066
rect 3865 19014 3877 19066
rect 3877 19014 3891 19066
rect 3915 19014 3929 19066
rect 3929 19014 3941 19066
rect 3941 19014 3971 19066
rect 3995 19014 4005 19066
rect 4005 19014 4051 19066
rect 3755 19012 3811 19014
rect 3835 19012 3891 19014
rect 3915 19012 3971 19014
rect 3995 19012 4051 19014
rect 3698 18128 3754 18184
rect 3755 17978 3811 17980
rect 3835 17978 3891 17980
rect 3915 17978 3971 17980
rect 3995 17978 4051 17980
rect 3755 17926 3801 17978
rect 3801 17926 3811 17978
rect 3835 17926 3865 17978
rect 3865 17926 3877 17978
rect 3877 17926 3891 17978
rect 3915 17926 3929 17978
rect 3929 17926 3941 17978
rect 3941 17926 3971 17978
rect 3995 17926 4005 17978
rect 4005 17926 4051 17978
rect 3755 17924 3811 17926
rect 3835 17924 3891 17926
rect 3915 17924 3971 17926
rect 3995 17924 4051 17926
rect 3882 17720 3938 17776
rect 3755 16890 3811 16892
rect 3835 16890 3891 16892
rect 3915 16890 3971 16892
rect 3995 16890 4051 16892
rect 3755 16838 3801 16890
rect 3801 16838 3811 16890
rect 3835 16838 3865 16890
rect 3865 16838 3877 16890
rect 3877 16838 3891 16890
rect 3915 16838 3929 16890
rect 3929 16838 3941 16890
rect 3941 16838 3971 16890
rect 3995 16838 4005 16890
rect 4005 16838 4051 16890
rect 3755 16836 3811 16838
rect 3835 16836 3891 16838
rect 3915 16836 3971 16838
rect 3995 16836 4051 16838
rect 3755 15802 3811 15804
rect 3835 15802 3891 15804
rect 3915 15802 3971 15804
rect 3995 15802 4051 15804
rect 3755 15750 3801 15802
rect 3801 15750 3811 15802
rect 3835 15750 3865 15802
rect 3865 15750 3877 15802
rect 3877 15750 3891 15802
rect 3915 15750 3929 15802
rect 3929 15750 3941 15802
rect 3941 15750 3971 15802
rect 3995 15750 4005 15802
rect 4005 15750 4051 15802
rect 3755 15748 3811 15750
rect 3835 15748 3891 15750
rect 3915 15748 3971 15750
rect 3995 15748 4051 15750
rect 6554 21786 6610 21788
rect 6634 21786 6690 21788
rect 6714 21786 6770 21788
rect 6794 21786 6850 21788
rect 6554 21734 6600 21786
rect 6600 21734 6610 21786
rect 6634 21734 6664 21786
rect 6664 21734 6676 21786
rect 6676 21734 6690 21786
rect 6714 21734 6728 21786
rect 6728 21734 6740 21786
rect 6740 21734 6770 21786
rect 6794 21734 6804 21786
rect 6804 21734 6850 21786
rect 6554 21732 6610 21734
rect 6634 21732 6690 21734
rect 6714 21732 6770 21734
rect 6794 21732 6850 21734
rect 6554 20698 6610 20700
rect 6634 20698 6690 20700
rect 6714 20698 6770 20700
rect 6794 20698 6850 20700
rect 6554 20646 6600 20698
rect 6600 20646 6610 20698
rect 6634 20646 6664 20698
rect 6664 20646 6676 20698
rect 6676 20646 6690 20698
rect 6714 20646 6728 20698
rect 6728 20646 6740 20698
rect 6740 20646 6770 20698
rect 6794 20646 6804 20698
rect 6804 20646 6850 20698
rect 6554 20644 6610 20646
rect 6634 20644 6690 20646
rect 6714 20644 6770 20646
rect 6794 20644 6850 20646
rect 6554 19610 6610 19612
rect 6634 19610 6690 19612
rect 6714 19610 6770 19612
rect 6794 19610 6850 19612
rect 6554 19558 6600 19610
rect 6600 19558 6610 19610
rect 6634 19558 6664 19610
rect 6664 19558 6676 19610
rect 6676 19558 6690 19610
rect 6714 19558 6728 19610
rect 6728 19558 6740 19610
rect 6740 19558 6770 19610
rect 6794 19558 6804 19610
rect 6804 19558 6850 19610
rect 6554 19556 6610 19558
rect 6634 19556 6690 19558
rect 6714 19556 6770 19558
rect 6794 19556 6850 19558
rect 3755 14714 3811 14716
rect 3835 14714 3891 14716
rect 3915 14714 3971 14716
rect 3995 14714 4051 14716
rect 3755 14662 3801 14714
rect 3801 14662 3811 14714
rect 3835 14662 3865 14714
rect 3865 14662 3877 14714
rect 3877 14662 3891 14714
rect 3915 14662 3929 14714
rect 3929 14662 3941 14714
rect 3941 14662 3971 14714
rect 3995 14662 4005 14714
rect 4005 14662 4051 14714
rect 3755 14660 3811 14662
rect 3835 14660 3891 14662
rect 3915 14660 3971 14662
rect 3995 14660 4051 14662
rect 3755 13626 3811 13628
rect 3835 13626 3891 13628
rect 3915 13626 3971 13628
rect 3995 13626 4051 13628
rect 3755 13574 3801 13626
rect 3801 13574 3811 13626
rect 3835 13574 3865 13626
rect 3865 13574 3877 13626
rect 3877 13574 3891 13626
rect 3915 13574 3929 13626
rect 3929 13574 3941 13626
rect 3941 13574 3971 13626
rect 3995 13574 4005 13626
rect 4005 13574 4051 13626
rect 3755 13572 3811 13574
rect 3835 13572 3891 13574
rect 3915 13572 3971 13574
rect 3995 13572 4051 13574
rect 3755 12538 3811 12540
rect 3835 12538 3891 12540
rect 3915 12538 3971 12540
rect 3995 12538 4051 12540
rect 3755 12486 3801 12538
rect 3801 12486 3811 12538
rect 3835 12486 3865 12538
rect 3865 12486 3877 12538
rect 3877 12486 3891 12538
rect 3915 12486 3929 12538
rect 3929 12486 3941 12538
rect 3941 12486 3971 12538
rect 3995 12486 4005 12538
rect 4005 12486 4051 12538
rect 3755 12484 3811 12486
rect 3835 12484 3891 12486
rect 3915 12484 3971 12486
rect 3995 12484 4051 12486
rect 3755 11450 3811 11452
rect 3835 11450 3891 11452
rect 3915 11450 3971 11452
rect 3995 11450 4051 11452
rect 3755 11398 3801 11450
rect 3801 11398 3811 11450
rect 3835 11398 3865 11450
rect 3865 11398 3877 11450
rect 3877 11398 3891 11450
rect 3915 11398 3929 11450
rect 3929 11398 3941 11450
rect 3941 11398 3971 11450
rect 3995 11398 4005 11450
rect 4005 11398 4051 11450
rect 3755 11396 3811 11398
rect 3835 11396 3891 11398
rect 3915 11396 3971 11398
rect 3995 11396 4051 11398
rect 3755 10362 3811 10364
rect 3835 10362 3891 10364
rect 3915 10362 3971 10364
rect 3995 10362 4051 10364
rect 3755 10310 3801 10362
rect 3801 10310 3811 10362
rect 3835 10310 3865 10362
rect 3865 10310 3877 10362
rect 3877 10310 3891 10362
rect 3915 10310 3929 10362
rect 3929 10310 3941 10362
rect 3941 10310 3971 10362
rect 3995 10310 4005 10362
rect 4005 10310 4051 10362
rect 3755 10308 3811 10310
rect 3835 10308 3891 10310
rect 3915 10308 3971 10310
rect 3995 10308 4051 10310
rect 3755 9274 3811 9276
rect 3835 9274 3891 9276
rect 3915 9274 3971 9276
rect 3995 9274 4051 9276
rect 3755 9222 3801 9274
rect 3801 9222 3811 9274
rect 3835 9222 3865 9274
rect 3865 9222 3877 9274
rect 3877 9222 3891 9274
rect 3915 9222 3929 9274
rect 3929 9222 3941 9274
rect 3941 9222 3971 9274
rect 3995 9222 4005 9274
rect 4005 9222 4051 9274
rect 3755 9220 3811 9222
rect 3835 9220 3891 9222
rect 3915 9220 3971 9222
rect 3995 9220 4051 9222
rect 6554 18522 6610 18524
rect 6634 18522 6690 18524
rect 6714 18522 6770 18524
rect 6794 18522 6850 18524
rect 6554 18470 6600 18522
rect 6600 18470 6610 18522
rect 6634 18470 6664 18522
rect 6664 18470 6676 18522
rect 6676 18470 6690 18522
rect 6714 18470 6728 18522
rect 6728 18470 6740 18522
rect 6740 18470 6770 18522
rect 6794 18470 6804 18522
rect 6804 18470 6850 18522
rect 6554 18468 6610 18470
rect 6634 18468 6690 18470
rect 6714 18468 6770 18470
rect 6794 18468 6850 18470
rect 7010 19488 7066 19544
rect 7010 19388 7012 19408
rect 7012 19388 7064 19408
rect 7064 19388 7066 19408
rect 7010 19352 7066 19388
rect 7194 18844 7196 18864
rect 7196 18844 7248 18864
rect 7248 18844 7250 18864
rect 7194 18808 7250 18844
rect 6550 17720 6606 17776
rect 6554 17434 6610 17436
rect 6634 17434 6690 17436
rect 6714 17434 6770 17436
rect 6794 17434 6850 17436
rect 6554 17382 6600 17434
rect 6600 17382 6610 17434
rect 6634 17382 6664 17434
rect 6664 17382 6676 17434
rect 6676 17382 6690 17434
rect 6714 17382 6728 17434
rect 6728 17382 6740 17434
rect 6740 17382 6770 17434
rect 6794 17382 6804 17434
rect 6804 17382 6850 17434
rect 6554 17380 6610 17382
rect 6634 17380 6690 17382
rect 6714 17380 6770 17382
rect 6794 17380 6850 17382
rect 7102 18164 7104 18184
rect 7104 18164 7156 18184
rect 7156 18164 7158 18184
rect 7102 18128 7158 18164
rect 6554 16346 6610 16348
rect 6634 16346 6690 16348
rect 6714 16346 6770 16348
rect 6794 16346 6850 16348
rect 6554 16294 6600 16346
rect 6600 16294 6610 16346
rect 6634 16294 6664 16346
rect 6664 16294 6676 16346
rect 6676 16294 6690 16346
rect 6714 16294 6728 16346
rect 6728 16294 6740 16346
rect 6740 16294 6770 16346
rect 6794 16294 6804 16346
rect 6804 16294 6850 16346
rect 6554 16292 6610 16294
rect 6634 16292 6690 16294
rect 6714 16292 6770 16294
rect 6794 16292 6850 16294
rect 6554 15258 6610 15260
rect 6634 15258 6690 15260
rect 6714 15258 6770 15260
rect 6794 15258 6850 15260
rect 6554 15206 6600 15258
rect 6600 15206 6610 15258
rect 6634 15206 6664 15258
rect 6664 15206 6676 15258
rect 6676 15206 6690 15258
rect 6714 15206 6728 15258
rect 6728 15206 6740 15258
rect 6740 15206 6770 15258
rect 6794 15206 6804 15258
rect 6804 15206 6850 15258
rect 6554 15204 6610 15206
rect 6634 15204 6690 15206
rect 6714 15204 6770 15206
rect 6794 15204 6850 15206
rect 6554 14170 6610 14172
rect 6634 14170 6690 14172
rect 6714 14170 6770 14172
rect 6794 14170 6850 14172
rect 6554 14118 6600 14170
rect 6600 14118 6610 14170
rect 6634 14118 6664 14170
rect 6664 14118 6676 14170
rect 6676 14118 6690 14170
rect 6714 14118 6728 14170
rect 6728 14118 6740 14170
rect 6740 14118 6770 14170
rect 6794 14118 6804 14170
rect 6804 14118 6850 14170
rect 6554 14116 6610 14118
rect 6634 14116 6690 14118
rect 6714 14116 6770 14118
rect 6794 14116 6850 14118
rect 7654 21392 7710 21448
rect 8482 21528 8538 21584
rect 8574 20984 8630 21040
rect 7838 20032 7894 20088
rect 7838 19352 7894 19408
rect 7470 18128 7526 18184
rect 7562 17620 7564 17640
rect 7564 17620 7616 17640
rect 7616 17620 7618 17640
rect 7562 17584 7618 17620
rect 8114 19352 8170 19408
rect 8022 17856 8078 17912
rect 8206 18264 8262 18320
rect 6554 13082 6610 13084
rect 6634 13082 6690 13084
rect 6714 13082 6770 13084
rect 6794 13082 6850 13084
rect 6554 13030 6600 13082
rect 6600 13030 6610 13082
rect 6634 13030 6664 13082
rect 6664 13030 6676 13082
rect 6676 13030 6690 13082
rect 6714 13030 6728 13082
rect 6728 13030 6740 13082
rect 6740 13030 6770 13082
rect 6794 13030 6804 13082
rect 6804 13030 6850 13082
rect 6554 13028 6610 13030
rect 6634 13028 6690 13030
rect 6714 13028 6770 13030
rect 6794 13028 6850 13030
rect 3755 8186 3811 8188
rect 3835 8186 3891 8188
rect 3915 8186 3971 8188
rect 3995 8186 4051 8188
rect 3755 8134 3801 8186
rect 3801 8134 3811 8186
rect 3835 8134 3865 8186
rect 3865 8134 3877 8186
rect 3877 8134 3891 8186
rect 3915 8134 3929 8186
rect 3929 8134 3941 8186
rect 3941 8134 3971 8186
rect 3995 8134 4005 8186
rect 4005 8134 4051 8186
rect 3755 8132 3811 8134
rect 3835 8132 3891 8134
rect 3915 8132 3971 8134
rect 3995 8132 4051 8134
rect 2870 6160 2926 6216
rect 2502 5616 2558 5672
rect 2226 4120 2282 4176
rect 3755 7098 3811 7100
rect 3835 7098 3891 7100
rect 3915 7098 3971 7100
rect 3995 7098 4051 7100
rect 3755 7046 3801 7098
rect 3801 7046 3811 7098
rect 3835 7046 3865 7098
rect 3865 7046 3877 7098
rect 3877 7046 3891 7098
rect 3915 7046 3929 7098
rect 3929 7046 3941 7098
rect 3941 7046 3971 7098
rect 3995 7046 4005 7098
rect 4005 7046 4051 7098
rect 3755 7044 3811 7046
rect 3835 7044 3891 7046
rect 3915 7044 3971 7046
rect 3995 7044 4051 7046
rect 4158 6840 4214 6896
rect 3755 6010 3811 6012
rect 3835 6010 3891 6012
rect 3915 6010 3971 6012
rect 3995 6010 4051 6012
rect 3755 5958 3801 6010
rect 3801 5958 3811 6010
rect 3835 5958 3865 6010
rect 3865 5958 3877 6010
rect 3877 5958 3891 6010
rect 3915 5958 3929 6010
rect 3929 5958 3941 6010
rect 3941 5958 3971 6010
rect 3995 5958 4005 6010
rect 4005 5958 4051 6010
rect 3755 5956 3811 5958
rect 3835 5956 3891 5958
rect 3915 5956 3971 5958
rect 3995 5956 4051 5958
rect 2962 4548 3018 4584
rect 2962 4528 2964 4548
rect 2964 4528 3016 4548
rect 3016 4528 3018 4548
rect 3238 3440 3294 3496
rect 1398 3032 1454 3088
rect 1582 2896 1638 2952
rect 3330 2352 3386 2408
rect 3755 4922 3811 4924
rect 3835 4922 3891 4924
rect 3915 4922 3971 4924
rect 3995 4922 4051 4924
rect 3755 4870 3801 4922
rect 3801 4870 3811 4922
rect 3835 4870 3865 4922
rect 3865 4870 3877 4922
rect 3877 4870 3891 4922
rect 3915 4870 3929 4922
rect 3929 4870 3941 4922
rect 3941 4870 3971 4922
rect 3995 4870 4005 4922
rect 4005 4870 4051 4922
rect 3755 4868 3811 4870
rect 3835 4868 3891 4870
rect 3915 4868 3971 4870
rect 3995 4868 4051 4870
rect 3974 4004 4030 4040
rect 3974 3984 3976 4004
rect 3976 3984 4028 4004
rect 4028 3984 4030 4004
rect 3755 3834 3811 3836
rect 3835 3834 3891 3836
rect 3915 3834 3971 3836
rect 3995 3834 4051 3836
rect 3755 3782 3801 3834
rect 3801 3782 3811 3834
rect 3835 3782 3865 3834
rect 3865 3782 3877 3834
rect 3877 3782 3891 3834
rect 3915 3782 3929 3834
rect 3929 3782 3941 3834
rect 3941 3782 3971 3834
rect 3995 3782 4005 3834
rect 4005 3782 4051 3834
rect 3755 3780 3811 3782
rect 3835 3780 3891 3782
rect 3915 3780 3971 3782
rect 3995 3780 4051 3782
rect 4802 7248 4858 7304
rect 6554 11994 6610 11996
rect 6634 11994 6690 11996
rect 6714 11994 6770 11996
rect 6794 11994 6850 11996
rect 6554 11942 6600 11994
rect 6600 11942 6610 11994
rect 6634 11942 6664 11994
rect 6664 11942 6676 11994
rect 6676 11942 6690 11994
rect 6714 11942 6728 11994
rect 6728 11942 6740 11994
rect 6740 11942 6770 11994
rect 6794 11942 6804 11994
rect 6804 11942 6850 11994
rect 6554 11940 6610 11942
rect 6634 11940 6690 11942
rect 6714 11940 6770 11942
rect 6794 11940 6850 11942
rect 6554 10906 6610 10908
rect 6634 10906 6690 10908
rect 6714 10906 6770 10908
rect 6794 10906 6850 10908
rect 6554 10854 6600 10906
rect 6600 10854 6610 10906
rect 6634 10854 6664 10906
rect 6664 10854 6676 10906
rect 6676 10854 6690 10906
rect 6714 10854 6728 10906
rect 6728 10854 6740 10906
rect 6740 10854 6770 10906
rect 6794 10854 6804 10906
rect 6804 10854 6850 10906
rect 6554 10852 6610 10854
rect 6634 10852 6690 10854
rect 6714 10852 6770 10854
rect 6794 10852 6850 10854
rect 6554 9818 6610 9820
rect 6634 9818 6690 9820
rect 6714 9818 6770 9820
rect 6794 9818 6850 9820
rect 6554 9766 6600 9818
rect 6600 9766 6610 9818
rect 6634 9766 6664 9818
rect 6664 9766 6676 9818
rect 6676 9766 6690 9818
rect 6714 9766 6728 9818
rect 6728 9766 6740 9818
rect 6740 9766 6770 9818
rect 6794 9766 6804 9818
rect 6804 9766 6850 9818
rect 6554 9764 6610 9766
rect 6634 9764 6690 9766
rect 6714 9764 6770 9766
rect 6794 9764 6850 9766
rect 6554 8730 6610 8732
rect 6634 8730 6690 8732
rect 6714 8730 6770 8732
rect 6794 8730 6850 8732
rect 6554 8678 6600 8730
rect 6600 8678 6610 8730
rect 6634 8678 6664 8730
rect 6664 8678 6676 8730
rect 6676 8678 6690 8730
rect 6714 8678 6728 8730
rect 6728 8678 6740 8730
rect 6740 8678 6770 8730
rect 6794 8678 6804 8730
rect 6804 8678 6850 8730
rect 6554 8676 6610 8678
rect 6634 8676 6690 8678
rect 6714 8676 6770 8678
rect 6794 8676 6850 8678
rect 6554 7642 6610 7644
rect 6634 7642 6690 7644
rect 6714 7642 6770 7644
rect 6794 7642 6850 7644
rect 6554 7590 6600 7642
rect 6600 7590 6610 7642
rect 6634 7590 6664 7642
rect 6664 7590 6676 7642
rect 6676 7590 6690 7642
rect 6714 7590 6728 7642
rect 6728 7590 6740 7642
rect 6740 7590 6770 7642
rect 6794 7590 6804 7642
rect 6804 7590 6850 7642
rect 6554 7588 6610 7590
rect 6634 7588 6690 7590
rect 6714 7588 6770 7590
rect 6794 7588 6850 7590
rect 6554 6554 6610 6556
rect 6634 6554 6690 6556
rect 6714 6554 6770 6556
rect 6794 6554 6850 6556
rect 6554 6502 6600 6554
rect 6600 6502 6610 6554
rect 6634 6502 6664 6554
rect 6664 6502 6676 6554
rect 6676 6502 6690 6554
rect 6714 6502 6728 6554
rect 6728 6502 6740 6554
rect 6740 6502 6770 6554
rect 6794 6502 6804 6554
rect 6804 6502 6850 6554
rect 6554 6500 6610 6502
rect 6634 6500 6690 6502
rect 6714 6500 6770 6502
rect 6794 6500 6850 6502
rect 8666 17756 8668 17776
rect 8668 17756 8720 17776
rect 8720 17756 8722 17776
rect 8666 17720 8722 17756
rect 8666 17584 8722 17640
rect 8850 17856 8906 17912
rect 9353 22330 9409 22332
rect 9433 22330 9489 22332
rect 9513 22330 9569 22332
rect 9593 22330 9649 22332
rect 9353 22278 9399 22330
rect 9399 22278 9409 22330
rect 9433 22278 9463 22330
rect 9463 22278 9475 22330
rect 9475 22278 9489 22330
rect 9513 22278 9527 22330
rect 9527 22278 9539 22330
rect 9539 22278 9569 22330
rect 9593 22278 9603 22330
rect 9603 22278 9649 22330
rect 9353 22276 9409 22278
rect 9433 22276 9489 22278
rect 9513 22276 9569 22278
rect 9593 22276 9649 22278
rect 9126 21972 9128 21992
rect 9128 21972 9180 21992
rect 9180 21972 9182 21992
rect 9126 21936 9182 21972
rect 10138 21936 10194 21992
rect 9034 20848 9090 20904
rect 9678 21392 9734 21448
rect 9353 21242 9409 21244
rect 9433 21242 9489 21244
rect 9513 21242 9569 21244
rect 9593 21242 9649 21244
rect 9353 21190 9399 21242
rect 9399 21190 9409 21242
rect 9433 21190 9463 21242
rect 9463 21190 9475 21242
rect 9475 21190 9489 21242
rect 9513 21190 9527 21242
rect 9527 21190 9539 21242
rect 9539 21190 9569 21242
rect 9593 21190 9603 21242
rect 9603 21190 9649 21242
rect 9353 21188 9409 21190
rect 9433 21188 9489 21190
rect 9513 21188 9569 21190
rect 9593 21188 9649 21190
rect 9310 20884 9312 20904
rect 9312 20884 9364 20904
rect 9364 20884 9366 20904
rect 9310 20848 9366 20884
rect 9218 20304 9274 20360
rect 9353 20154 9409 20156
rect 9433 20154 9489 20156
rect 9513 20154 9569 20156
rect 9593 20154 9649 20156
rect 9353 20102 9399 20154
rect 9399 20102 9409 20154
rect 9433 20102 9463 20154
rect 9463 20102 9475 20154
rect 9475 20102 9489 20154
rect 9513 20102 9527 20154
rect 9527 20102 9539 20154
rect 9539 20102 9569 20154
rect 9593 20102 9603 20154
rect 9603 20102 9649 20154
rect 9353 20100 9409 20102
rect 9433 20100 9489 20102
rect 9513 20100 9569 20102
rect 9593 20100 9649 20102
rect 9678 19760 9734 19816
rect 9353 19066 9409 19068
rect 9433 19066 9489 19068
rect 9513 19066 9569 19068
rect 9593 19066 9649 19068
rect 9353 19014 9399 19066
rect 9399 19014 9409 19066
rect 9433 19014 9463 19066
rect 9463 19014 9475 19066
rect 9475 19014 9489 19066
rect 9513 19014 9527 19066
rect 9527 19014 9539 19066
rect 9539 19014 9569 19066
rect 9593 19014 9603 19066
rect 9603 19014 9649 19066
rect 9353 19012 9409 19014
rect 9433 19012 9489 19014
rect 9513 19012 9569 19014
rect 9593 19012 9649 19014
rect 9310 18844 9312 18864
rect 9312 18844 9364 18864
rect 9364 18844 9366 18864
rect 9310 18808 9366 18844
rect 9353 17978 9409 17980
rect 9433 17978 9489 17980
rect 9513 17978 9569 17980
rect 9593 17978 9649 17980
rect 9353 17926 9399 17978
rect 9399 17926 9409 17978
rect 9433 17926 9463 17978
rect 9463 17926 9475 17978
rect 9475 17926 9489 17978
rect 9513 17926 9527 17978
rect 9527 17926 9539 17978
rect 9539 17926 9569 17978
rect 9593 17926 9603 17978
rect 9603 17926 9649 17978
rect 9353 17924 9409 17926
rect 9433 17924 9489 17926
rect 9513 17924 9569 17926
rect 9593 17924 9649 17926
rect 10138 20304 10194 20360
rect 10230 19760 10286 19816
rect 9770 18164 9772 18184
rect 9772 18164 9824 18184
rect 9824 18164 9826 18184
rect 9770 18128 9826 18164
rect 9126 17040 9182 17096
rect 9353 16890 9409 16892
rect 9433 16890 9489 16892
rect 9513 16890 9569 16892
rect 9593 16890 9649 16892
rect 9353 16838 9399 16890
rect 9399 16838 9409 16890
rect 9433 16838 9463 16890
rect 9463 16838 9475 16890
rect 9475 16838 9489 16890
rect 9513 16838 9527 16890
rect 9527 16838 9539 16890
rect 9539 16838 9569 16890
rect 9593 16838 9603 16890
rect 9603 16838 9649 16890
rect 9353 16836 9409 16838
rect 9433 16836 9489 16838
rect 9513 16836 9569 16838
rect 9593 16836 9649 16838
rect 10046 19508 10102 19544
rect 10046 19488 10048 19508
rect 10048 19488 10100 19508
rect 10100 19488 10102 19508
rect 9353 15802 9409 15804
rect 9433 15802 9489 15804
rect 9513 15802 9569 15804
rect 9593 15802 9649 15804
rect 9353 15750 9399 15802
rect 9399 15750 9409 15802
rect 9433 15750 9463 15802
rect 9463 15750 9475 15802
rect 9475 15750 9489 15802
rect 9513 15750 9527 15802
rect 9527 15750 9539 15802
rect 9539 15750 9569 15802
rect 9593 15750 9603 15802
rect 9603 15750 9649 15802
rect 9353 15748 9409 15750
rect 9433 15748 9489 15750
rect 9513 15748 9569 15750
rect 9593 15748 9649 15750
rect 10506 20848 10562 20904
rect 11150 19760 11206 19816
rect 10874 18572 10876 18592
rect 10876 18572 10928 18592
rect 10928 18572 10930 18592
rect 10874 18536 10930 18572
rect 12162 21972 12164 21992
rect 12164 21972 12216 21992
rect 12216 21972 12218 21992
rect 12162 21936 12218 21972
rect 12438 21956 12494 21992
rect 12438 21936 12440 21956
rect 12440 21936 12492 21956
rect 12492 21936 12494 21956
rect 12152 21786 12208 21788
rect 12232 21786 12288 21788
rect 12312 21786 12368 21788
rect 12392 21786 12448 21788
rect 12152 21734 12198 21786
rect 12198 21734 12208 21786
rect 12232 21734 12262 21786
rect 12262 21734 12274 21786
rect 12274 21734 12288 21786
rect 12312 21734 12326 21786
rect 12326 21734 12338 21786
rect 12338 21734 12368 21786
rect 12392 21734 12402 21786
rect 12402 21734 12448 21786
rect 12152 21732 12208 21734
rect 12232 21732 12288 21734
rect 12312 21732 12368 21734
rect 12392 21732 12448 21734
rect 12152 20698 12208 20700
rect 12232 20698 12288 20700
rect 12312 20698 12368 20700
rect 12392 20698 12448 20700
rect 12152 20646 12198 20698
rect 12198 20646 12208 20698
rect 12232 20646 12262 20698
rect 12262 20646 12274 20698
rect 12274 20646 12288 20698
rect 12312 20646 12326 20698
rect 12326 20646 12338 20698
rect 12338 20646 12368 20698
rect 12392 20646 12402 20698
rect 12402 20646 12448 20698
rect 12152 20644 12208 20646
rect 12232 20644 12288 20646
rect 12312 20644 12368 20646
rect 12392 20644 12448 20646
rect 13266 20440 13322 20496
rect 11150 18400 11206 18456
rect 9353 14714 9409 14716
rect 9433 14714 9489 14716
rect 9513 14714 9569 14716
rect 9593 14714 9649 14716
rect 9353 14662 9399 14714
rect 9399 14662 9409 14714
rect 9433 14662 9463 14714
rect 9463 14662 9475 14714
rect 9475 14662 9489 14714
rect 9513 14662 9527 14714
rect 9527 14662 9539 14714
rect 9539 14662 9569 14714
rect 9593 14662 9603 14714
rect 9603 14662 9649 14714
rect 9353 14660 9409 14662
rect 9433 14660 9489 14662
rect 9513 14660 9569 14662
rect 9593 14660 9649 14662
rect 9353 13626 9409 13628
rect 9433 13626 9489 13628
rect 9513 13626 9569 13628
rect 9593 13626 9649 13628
rect 9353 13574 9399 13626
rect 9399 13574 9409 13626
rect 9433 13574 9463 13626
rect 9463 13574 9475 13626
rect 9475 13574 9489 13626
rect 9513 13574 9527 13626
rect 9527 13574 9539 13626
rect 9539 13574 9569 13626
rect 9593 13574 9603 13626
rect 9603 13574 9649 13626
rect 9353 13572 9409 13574
rect 9433 13572 9489 13574
rect 9513 13572 9569 13574
rect 9593 13572 9649 13574
rect 9353 12538 9409 12540
rect 9433 12538 9489 12540
rect 9513 12538 9569 12540
rect 9593 12538 9649 12540
rect 9353 12486 9399 12538
rect 9399 12486 9409 12538
rect 9433 12486 9463 12538
rect 9463 12486 9475 12538
rect 9475 12486 9489 12538
rect 9513 12486 9527 12538
rect 9527 12486 9539 12538
rect 9539 12486 9569 12538
rect 9593 12486 9603 12538
rect 9603 12486 9649 12538
rect 9353 12484 9409 12486
rect 9433 12484 9489 12486
rect 9513 12484 9569 12486
rect 9593 12484 9649 12486
rect 9353 11450 9409 11452
rect 9433 11450 9489 11452
rect 9513 11450 9569 11452
rect 9593 11450 9649 11452
rect 9353 11398 9399 11450
rect 9399 11398 9409 11450
rect 9433 11398 9463 11450
rect 9463 11398 9475 11450
rect 9475 11398 9489 11450
rect 9513 11398 9527 11450
rect 9527 11398 9539 11450
rect 9539 11398 9569 11450
rect 9593 11398 9603 11450
rect 9603 11398 9649 11450
rect 9353 11396 9409 11398
rect 9433 11396 9489 11398
rect 9513 11396 9569 11398
rect 9593 11396 9649 11398
rect 9353 10362 9409 10364
rect 9433 10362 9489 10364
rect 9513 10362 9569 10364
rect 9593 10362 9649 10364
rect 9353 10310 9399 10362
rect 9399 10310 9409 10362
rect 9433 10310 9463 10362
rect 9463 10310 9475 10362
rect 9475 10310 9489 10362
rect 9513 10310 9527 10362
rect 9527 10310 9539 10362
rect 9539 10310 9569 10362
rect 9593 10310 9603 10362
rect 9603 10310 9649 10362
rect 9353 10308 9409 10310
rect 9433 10308 9489 10310
rect 9513 10308 9569 10310
rect 9593 10308 9649 10310
rect 9353 9274 9409 9276
rect 9433 9274 9489 9276
rect 9513 9274 9569 9276
rect 9593 9274 9649 9276
rect 9353 9222 9399 9274
rect 9399 9222 9409 9274
rect 9433 9222 9463 9274
rect 9463 9222 9475 9274
rect 9475 9222 9489 9274
rect 9513 9222 9527 9274
rect 9527 9222 9539 9274
rect 9539 9222 9569 9274
rect 9593 9222 9603 9274
rect 9603 9222 9649 9274
rect 9353 9220 9409 9222
rect 9433 9220 9489 9222
rect 9513 9220 9569 9222
rect 9593 9220 9649 9222
rect 9353 8186 9409 8188
rect 9433 8186 9489 8188
rect 9513 8186 9569 8188
rect 9593 8186 9649 8188
rect 9353 8134 9399 8186
rect 9399 8134 9409 8186
rect 9433 8134 9463 8186
rect 9463 8134 9475 8186
rect 9475 8134 9489 8186
rect 9513 8134 9527 8186
rect 9527 8134 9539 8186
rect 9539 8134 9569 8186
rect 9593 8134 9603 8186
rect 9603 8134 9649 8186
rect 9353 8132 9409 8134
rect 9433 8132 9489 8134
rect 9513 8132 9569 8134
rect 9593 8132 9649 8134
rect 11242 17176 11298 17232
rect 11702 18808 11758 18864
rect 11702 18536 11758 18592
rect 11702 18128 11758 18184
rect 9034 7792 9090 7848
rect 5446 5072 5502 5128
rect 6554 5466 6610 5468
rect 6634 5466 6690 5468
rect 6714 5466 6770 5468
rect 6794 5466 6850 5468
rect 6554 5414 6600 5466
rect 6600 5414 6610 5466
rect 6634 5414 6664 5466
rect 6664 5414 6676 5466
rect 6676 5414 6690 5466
rect 6714 5414 6728 5466
rect 6728 5414 6740 5466
rect 6740 5414 6770 5466
rect 6794 5414 6804 5466
rect 6804 5414 6850 5466
rect 6554 5412 6610 5414
rect 6634 5412 6690 5414
rect 6714 5412 6770 5414
rect 6794 5412 6850 5414
rect 5354 4664 5410 4720
rect 6554 4378 6610 4380
rect 6634 4378 6690 4380
rect 6714 4378 6770 4380
rect 6794 4378 6850 4380
rect 6554 4326 6600 4378
rect 6600 4326 6610 4378
rect 6634 4326 6664 4378
rect 6664 4326 6676 4378
rect 6676 4326 6690 4378
rect 6714 4326 6728 4378
rect 6728 4326 6740 4378
rect 6740 4326 6770 4378
rect 6794 4326 6804 4378
rect 6804 4326 6850 4378
rect 6554 4324 6610 4326
rect 6634 4324 6690 4326
rect 6714 4324 6770 4326
rect 6794 4324 6850 4326
rect 3755 2746 3811 2748
rect 3835 2746 3891 2748
rect 3915 2746 3971 2748
rect 3995 2746 4051 2748
rect 3755 2694 3801 2746
rect 3801 2694 3811 2746
rect 3835 2694 3865 2746
rect 3865 2694 3877 2746
rect 3877 2694 3891 2746
rect 3915 2694 3929 2746
rect 3929 2694 3941 2746
rect 3941 2694 3971 2746
rect 3995 2694 4005 2746
rect 4005 2694 4051 2746
rect 3755 2692 3811 2694
rect 3835 2692 3891 2694
rect 3915 2692 3971 2694
rect 3995 2692 4051 2694
rect 5906 2524 5908 2544
rect 5908 2524 5960 2544
rect 5960 2524 5962 2544
rect 5906 2488 5962 2524
rect 6554 3290 6610 3292
rect 6634 3290 6690 3292
rect 6714 3290 6770 3292
rect 6794 3290 6850 3292
rect 6554 3238 6600 3290
rect 6600 3238 6610 3290
rect 6634 3238 6664 3290
rect 6664 3238 6676 3290
rect 6676 3238 6690 3290
rect 6714 3238 6728 3290
rect 6728 3238 6740 3290
rect 6740 3238 6770 3290
rect 6794 3238 6804 3290
rect 6804 3238 6850 3290
rect 6554 3236 6610 3238
rect 6634 3236 6690 3238
rect 6714 3236 6770 3238
rect 6794 3236 6850 3238
rect 5354 1944 5410 2000
rect 3974 1808 4030 1864
rect 2962 1672 3018 1728
rect 6826 2760 6882 2816
rect 7102 2488 7158 2544
rect 8114 2896 8170 2952
rect 6554 2202 6610 2204
rect 6634 2202 6690 2204
rect 6714 2202 6770 2204
rect 6794 2202 6850 2204
rect 6554 2150 6600 2202
rect 6600 2150 6610 2202
rect 6634 2150 6664 2202
rect 6664 2150 6676 2202
rect 6676 2150 6690 2202
rect 6714 2150 6728 2202
rect 6728 2150 6740 2202
rect 6740 2150 6770 2202
rect 6794 2150 6804 2202
rect 6804 2150 6850 2202
rect 6554 2148 6610 2150
rect 6634 2148 6690 2150
rect 6714 2148 6770 2150
rect 6794 2148 6850 2150
rect 10598 7404 10654 7440
rect 10598 7384 10600 7404
rect 10600 7384 10652 7404
rect 10652 7384 10654 7404
rect 9353 7098 9409 7100
rect 9433 7098 9489 7100
rect 9513 7098 9569 7100
rect 9593 7098 9649 7100
rect 9353 7046 9399 7098
rect 9399 7046 9409 7098
rect 9433 7046 9463 7098
rect 9463 7046 9475 7098
rect 9475 7046 9489 7098
rect 9513 7046 9527 7098
rect 9527 7046 9539 7098
rect 9539 7046 9569 7098
rect 9593 7046 9603 7098
rect 9603 7046 9649 7098
rect 9353 7044 9409 7046
rect 9433 7044 9489 7046
rect 9513 7044 9569 7046
rect 9593 7044 9649 7046
rect 11978 18400 12034 18456
rect 12152 19610 12208 19612
rect 12232 19610 12288 19612
rect 12312 19610 12368 19612
rect 12392 19610 12448 19612
rect 12152 19558 12198 19610
rect 12198 19558 12208 19610
rect 12232 19558 12262 19610
rect 12262 19558 12274 19610
rect 12274 19558 12288 19610
rect 12312 19558 12326 19610
rect 12326 19558 12338 19610
rect 12338 19558 12368 19610
rect 12392 19558 12402 19610
rect 12402 19558 12448 19610
rect 12152 19556 12208 19558
rect 12232 19556 12288 19558
rect 12312 19556 12368 19558
rect 12392 19556 12448 19558
rect 12152 18522 12208 18524
rect 12232 18522 12288 18524
rect 12312 18522 12368 18524
rect 12392 18522 12448 18524
rect 12152 18470 12198 18522
rect 12198 18470 12208 18522
rect 12232 18470 12262 18522
rect 12262 18470 12274 18522
rect 12274 18470 12288 18522
rect 12312 18470 12326 18522
rect 12326 18470 12338 18522
rect 12338 18470 12368 18522
rect 12392 18470 12402 18522
rect 12402 18470 12448 18522
rect 12152 18468 12208 18470
rect 12232 18468 12288 18470
rect 12312 18468 12368 18470
rect 12392 18468 12448 18470
rect 12152 17434 12208 17436
rect 12232 17434 12288 17436
rect 12312 17434 12368 17436
rect 12392 17434 12448 17436
rect 12152 17382 12198 17434
rect 12198 17382 12208 17434
rect 12232 17382 12262 17434
rect 12262 17382 12274 17434
rect 12274 17382 12288 17434
rect 12312 17382 12326 17434
rect 12326 17382 12338 17434
rect 12338 17382 12368 17434
rect 12392 17382 12402 17434
rect 12402 17382 12448 17434
rect 12152 17380 12208 17382
rect 12232 17380 12288 17382
rect 12312 17380 12368 17382
rect 12392 17380 12448 17382
rect 12152 16346 12208 16348
rect 12232 16346 12288 16348
rect 12312 16346 12368 16348
rect 12392 16346 12448 16348
rect 12152 16294 12198 16346
rect 12198 16294 12208 16346
rect 12232 16294 12262 16346
rect 12262 16294 12274 16346
rect 12274 16294 12288 16346
rect 12312 16294 12326 16346
rect 12326 16294 12338 16346
rect 12338 16294 12368 16346
rect 12392 16294 12402 16346
rect 12402 16294 12448 16346
rect 12152 16292 12208 16294
rect 12232 16292 12288 16294
rect 12312 16292 12368 16294
rect 12392 16292 12448 16294
rect 12152 15258 12208 15260
rect 12232 15258 12288 15260
rect 12312 15258 12368 15260
rect 12392 15258 12448 15260
rect 12152 15206 12198 15258
rect 12198 15206 12208 15258
rect 12232 15206 12262 15258
rect 12262 15206 12274 15258
rect 12274 15206 12288 15258
rect 12312 15206 12326 15258
rect 12326 15206 12338 15258
rect 12338 15206 12368 15258
rect 12392 15206 12402 15258
rect 12402 15206 12448 15258
rect 12152 15204 12208 15206
rect 12232 15204 12288 15206
rect 12312 15204 12368 15206
rect 12392 15204 12448 15206
rect 12152 14170 12208 14172
rect 12232 14170 12288 14172
rect 12312 14170 12368 14172
rect 12392 14170 12448 14172
rect 12152 14118 12198 14170
rect 12198 14118 12208 14170
rect 12232 14118 12262 14170
rect 12262 14118 12274 14170
rect 12274 14118 12288 14170
rect 12312 14118 12326 14170
rect 12326 14118 12338 14170
rect 12338 14118 12368 14170
rect 12392 14118 12402 14170
rect 12402 14118 12448 14170
rect 12152 14116 12208 14118
rect 12232 14116 12288 14118
rect 12312 14116 12368 14118
rect 12392 14116 12448 14118
rect 12152 13082 12208 13084
rect 12232 13082 12288 13084
rect 12312 13082 12368 13084
rect 12392 13082 12448 13084
rect 12152 13030 12198 13082
rect 12198 13030 12208 13082
rect 12232 13030 12262 13082
rect 12262 13030 12274 13082
rect 12274 13030 12288 13082
rect 12312 13030 12326 13082
rect 12326 13030 12338 13082
rect 12338 13030 12368 13082
rect 12392 13030 12402 13082
rect 12402 13030 12448 13082
rect 12152 13028 12208 13030
rect 12232 13028 12288 13030
rect 12312 13028 12368 13030
rect 12392 13028 12448 13030
rect 14951 22330 15007 22332
rect 15031 22330 15087 22332
rect 15111 22330 15167 22332
rect 15191 22330 15247 22332
rect 14951 22278 14997 22330
rect 14997 22278 15007 22330
rect 15031 22278 15061 22330
rect 15061 22278 15073 22330
rect 15073 22278 15087 22330
rect 15111 22278 15125 22330
rect 15125 22278 15137 22330
rect 15137 22278 15167 22330
rect 15191 22278 15201 22330
rect 15201 22278 15247 22330
rect 14951 22276 15007 22278
rect 15031 22276 15087 22278
rect 15111 22276 15167 22278
rect 15191 22276 15247 22278
rect 14646 21664 14702 21720
rect 14462 21392 14518 21448
rect 14094 19896 14150 19952
rect 13634 17720 13690 17776
rect 13634 15952 13690 16008
rect 11794 12824 11850 12880
rect 12152 11994 12208 11996
rect 12232 11994 12288 11996
rect 12312 11994 12368 11996
rect 12392 11994 12448 11996
rect 12152 11942 12198 11994
rect 12198 11942 12208 11994
rect 12232 11942 12262 11994
rect 12262 11942 12274 11994
rect 12274 11942 12288 11994
rect 12312 11942 12326 11994
rect 12326 11942 12338 11994
rect 12338 11942 12368 11994
rect 12392 11942 12402 11994
rect 12402 11942 12448 11994
rect 12152 11940 12208 11942
rect 12232 11940 12288 11942
rect 12312 11940 12368 11942
rect 12392 11940 12448 11942
rect 11794 10512 11850 10568
rect 10230 6704 10286 6760
rect 9353 6010 9409 6012
rect 9433 6010 9489 6012
rect 9513 6010 9569 6012
rect 9593 6010 9649 6012
rect 9353 5958 9399 6010
rect 9399 5958 9409 6010
rect 9433 5958 9463 6010
rect 9463 5958 9475 6010
rect 9475 5958 9489 6010
rect 9513 5958 9527 6010
rect 9527 5958 9539 6010
rect 9539 5958 9569 6010
rect 9593 5958 9603 6010
rect 9603 5958 9649 6010
rect 9353 5956 9409 5958
rect 9433 5956 9489 5958
rect 9513 5956 9569 5958
rect 9593 5956 9649 5958
rect 9353 4922 9409 4924
rect 9433 4922 9489 4924
rect 9513 4922 9569 4924
rect 9593 4922 9649 4924
rect 9353 4870 9399 4922
rect 9399 4870 9409 4922
rect 9433 4870 9463 4922
rect 9463 4870 9475 4922
rect 9475 4870 9489 4922
rect 9513 4870 9527 4922
rect 9527 4870 9539 4922
rect 9539 4870 9569 4922
rect 9593 4870 9603 4922
rect 9603 4870 9649 4922
rect 9353 4868 9409 4870
rect 9433 4868 9489 4870
rect 9513 4868 9569 4870
rect 9593 4868 9649 4870
rect 8298 2796 8300 2816
rect 8300 2796 8352 2816
rect 8352 2796 8354 2816
rect 8298 2760 8354 2796
rect 9353 3834 9409 3836
rect 9433 3834 9489 3836
rect 9513 3834 9569 3836
rect 9593 3834 9649 3836
rect 9353 3782 9399 3834
rect 9399 3782 9409 3834
rect 9433 3782 9463 3834
rect 9463 3782 9475 3834
rect 9475 3782 9489 3834
rect 9513 3782 9527 3834
rect 9527 3782 9539 3834
rect 9539 3782 9569 3834
rect 9593 3782 9603 3834
rect 9603 3782 9649 3834
rect 9353 3780 9409 3782
rect 9433 3780 9489 3782
rect 9513 3780 9569 3782
rect 9593 3780 9649 3782
rect 9126 2932 9128 2952
rect 9128 2932 9180 2952
rect 9180 2932 9182 2952
rect 9126 2896 9182 2932
rect 9353 2746 9409 2748
rect 9433 2746 9489 2748
rect 9513 2746 9569 2748
rect 9593 2746 9649 2748
rect 9353 2694 9399 2746
rect 9399 2694 9409 2746
rect 9433 2694 9463 2746
rect 9463 2694 9475 2746
rect 9475 2694 9489 2746
rect 9513 2694 9527 2746
rect 9527 2694 9539 2746
rect 9539 2694 9569 2746
rect 9593 2694 9603 2746
rect 9603 2694 9649 2746
rect 9353 2692 9409 2694
rect 9433 2692 9489 2694
rect 9513 2692 9569 2694
rect 9593 2692 9649 2694
rect 10966 6316 11022 6352
rect 10966 6296 10968 6316
rect 10968 6296 11020 6316
rect 11020 6296 11022 6316
rect 12152 10906 12208 10908
rect 12232 10906 12288 10908
rect 12312 10906 12368 10908
rect 12392 10906 12448 10908
rect 12152 10854 12198 10906
rect 12198 10854 12208 10906
rect 12232 10854 12262 10906
rect 12262 10854 12274 10906
rect 12274 10854 12288 10906
rect 12312 10854 12326 10906
rect 12326 10854 12338 10906
rect 12338 10854 12368 10906
rect 12392 10854 12402 10906
rect 12402 10854 12448 10906
rect 12152 10852 12208 10854
rect 12232 10852 12288 10854
rect 12312 10852 12368 10854
rect 12392 10852 12448 10854
rect 12152 9818 12208 9820
rect 12232 9818 12288 9820
rect 12312 9818 12368 9820
rect 12392 9818 12448 9820
rect 12152 9766 12198 9818
rect 12198 9766 12208 9818
rect 12232 9766 12262 9818
rect 12262 9766 12274 9818
rect 12274 9766 12288 9818
rect 12312 9766 12326 9818
rect 12326 9766 12338 9818
rect 12338 9766 12368 9818
rect 12392 9766 12402 9818
rect 12402 9766 12448 9818
rect 12152 9764 12208 9766
rect 12232 9764 12288 9766
rect 12312 9764 12368 9766
rect 12392 9764 12448 9766
rect 13634 11192 13690 11248
rect 14002 13776 14058 13832
rect 12898 9424 12954 9480
rect 11886 8880 11942 8936
rect 12152 8730 12208 8732
rect 12232 8730 12288 8732
rect 12312 8730 12368 8732
rect 12392 8730 12448 8732
rect 12152 8678 12198 8730
rect 12198 8678 12208 8730
rect 12232 8678 12262 8730
rect 12262 8678 12274 8730
rect 12274 8678 12288 8730
rect 12312 8678 12326 8730
rect 12326 8678 12338 8730
rect 12338 8678 12368 8730
rect 12392 8678 12402 8730
rect 12402 8678 12448 8730
rect 12152 8676 12208 8678
rect 12232 8676 12288 8678
rect 12312 8676 12368 8678
rect 12392 8676 12448 8678
rect 12152 7642 12208 7644
rect 12232 7642 12288 7644
rect 12312 7642 12368 7644
rect 12392 7642 12448 7644
rect 12152 7590 12198 7642
rect 12198 7590 12208 7642
rect 12232 7590 12262 7642
rect 12262 7590 12274 7642
rect 12274 7590 12288 7642
rect 12312 7590 12326 7642
rect 12326 7590 12338 7642
rect 12338 7590 12368 7642
rect 12392 7590 12402 7642
rect 12402 7590 12448 7642
rect 12152 7588 12208 7590
rect 12232 7588 12288 7590
rect 12312 7588 12368 7590
rect 12392 7588 12448 7590
rect 12152 6554 12208 6556
rect 12232 6554 12288 6556
rect 12312 6554 12368 6556
rect 12392 6554 12448 6556
rect 12152 6502 12198 6554
rect 12198 6502 12208 6554
rect 12232 6502 12262 6554
rect 12262 6502 12274 6554
rect 12274 6502 12288 6554
rect 12312 6502 12326 6554
rect 12326 6502 12338 6554
rect 12338 6502 12368 6554
rect 12392 6502 12402 6554
rect 12402 6502 12448 6554
rect 12152 6500 12208 6502
rect 12232 6500 12288 6502
rect 12312 6500 12368 6502
rect 12392 6500 12448 6502
rect 12152 5466 12208 5468
rect 12232 5466 12288 5468
rect 12312 5466 12368 5468
rect 12392 5466 12448 5468
rect 12152 5414 12198 5466
rect 12198 5414 12208 5466
rect 12232 5414 12262 5466
rect 12262 5414 12274 5466
rect 12274 5414 12288 5466
rect 12312 5414 12326 5466
rect 12326 5414 12338 5466
rect 12338 5414 12368 5466
rect 12392 5414 12402 5466
rect 12402 5414 12448 5466
rect 12152 5412 12208 5414
rect 12232 5412 12288 5414
rect 12312 5412 12368 5414
rect 12392 5412 12448 5414
rect 12152 4378 12208 4380
rect 12232 4378 12288 4380
rect 12312 4378 12368 4380
rect 12392 4378 12448 4380
rect 12152 4326 12198 4378
rect 12198 4326 12208 4378
rect 12232 4326 12262 4378
rect 12262 4326 12274 4378
rect 12274 4326 12288 4378
rect 12312 4326 12326 4378
rect 12326 4326 12338 4378
rect 12338 4326 12368 4378
rect 12392 4326 12402 4378
rect 12402 4326 12448 4378
rect 12152 4324 12208 4326
rect 12232 4324 12288 4326
rect 12312 4324 12368 4326
rect 12392 4324 12448 4326
rect 12152 3290 12208 3292
rect 12232 3290 12288 3292
rect 12312 3290 12368 3292
rect 12392 3290 12448 3292
rect 12152 3238 12198 3290
rect 12198 3238 12208 3290
rect 12232 3238 12262 3290
rect 12262 3238 12274 3290
rect 12274 3238 12288 3290
rect 12312 3238 12326 3290
rect 12326 3238 12338 3290
rect 12338 3238 12368 3290
rect 12392 3238 12402 3290
rect 12402 3238 12448 3290
rect 12152 3236 12208 3238
rect 12232 3236 12288 3238
rect 12312 3236 12368 3238
rect 12392 3236 12448 3238
rect 13542 9696 13598 9752
rect 14370 18400 14426 18456
rect 14951 21242 15007 21244
rect 15031 21242 15087 21244
rect 15111 21242 15167 21244
rect 15191 21242 15247 21244
rect 14951 21190 14997 21242
rect 14997 21190 15007 21242
rect 15031 21190 15061 21242
rect 15061 21190 15073 21242
rect 15073 21190 15087 21242
rect 15111 21190 15125 21242
rect 15125 21190 15137 21242
rect 15137 21190 15167 21242
rect 15191 21190 15201 21242
rect 15201 21190 15247 21242
rect 14951 21188 15007 21190
rect 15031 21188 15087 21190
rect 15111 21188 15167 21190
rect 15191 21188 15247 21190
rect 15474 21256 15530 21312
rect 14922 20848 14978 20904
rect 14830 20304 14886 20360
rect 14951 20154 15007 20156
rect 15031 20154 15087 20156
rect 15111 20154 15167 20156
rect 15191 20154 15247 20156
rect 14951 20102 14997 20154
rect 14997 20102 15007 20154
rect 15031 20102 15061 20154
rect 15061 20102 15073 20154
rect 15073 20102 15087 20154
rect 15111 20102 15125 20154
rect 15125 20102 15137 20154
rect 15137 20102 15167 20154
rect 15191 20102 15201 20154
rect 15201 20102 15247 20154
rect 14951 20100 15007 20102
rect 15031 20100 15087 20102
rect 15111 20100 15167 20102
rect 15191 20100 15247 20102
rect 14951 19066 15007 19068
rect 15031 19066 15087 19068
rect 15111 19066 15167 19068
rect 15191 19066 15247 19068
rect 14951 19014 14997 19066
rect 14997 19014 15007 19066
rect 15031 19014 15061 19066
rect 15061 19014 15073 19066
rect 15073 19014 15087 19066
rect 15111 19014 15125 19066
rect 15125 19014 15137 19066
rect 15137 19014 15167 19066
rect 15191 19014 15201 19066
rect 15201 19014 15247 19066
rect 14951 19012 15007 19014
rect 15031 19012 15087 19014
rect 15111 19012 15167 19014
rect 15191 19012 15247 19014
rect 14951 17978 15007 17980
rect 15031 17978 15087 17980
rect 15111 17978 15167 17980
rect 15191 17978 15247 17980
rect 14951 17926 14997 17978
rect 14997 17926 15007 17978
rect 15031 17926 15061 17978
rect 15061 17926 15073 17978
rect 15073 17926 15087 17978
rect 15111 17926 15125 17978
rect 15125 17926 15137 17978
rect 15137 17926 15167 17978
rect 15191 17926 15201 17978
rect 15201 17926 15247 17978
rect 14951 17924 15007 17926
rect 15031 17924 15087 17926
rect 15111 17924 15167 17926
rect 15191 17924 15247 17926
rect 14951 16890 15007 16892
rect 15031 16890 15087 16892
rect 15111 16890 15167 16892
rect 15191 16890 15247 16892
rect 14951 16838 14997 16890
rect 14997 16838 15007 16890
rect 15031 16838 15061 16890
rect 15061 16838 15073 16890
rect 15073 16838 15087 16890
rect 15111 16838 15125 16890
rect 15125 16838 15137 16890
rect 15137 16838 15167 16890
rect 15191 16838 15201 16890
rect 15201 16838 15247 16890
rect 14951 16836 15007 16838
rect 15031 16836 15087 16838
rect 15111 16836 15167 16838
rect 15191 16836 15247 16838
rect 16118 21664 16174 21720
rect 15934 21392 15990 21448
rect 16118 21392 16174 21448
rect 16210 20576 16266 20632
rect 17038 20984 17094 21040
rect 17750 21786 17806 21788
rect 17830 21786 17886 21788
rect 17910 21786 17966 21788
rect 17990 21786 18046 21788
rect 17750 21734 17796 21786
rect 17796 21734 17806 21786
rect 17830 21734 17860 21786
rect 17860 21734 17872 21786
rect 17872 21734 17886 21786
rect 17910 21734 17924 21786
rect 17924 21734 17936 21786
rect 17936 21734 17966 21786
rect 17990 21734 18000 21786
rect 18000 21734 18046 21786
rect 17750 21732 17806 21734
rect 17830 21732 17886 21734
rect 17910 21732 17966 21734
rect 17990 21732 18046 21734
rect 17590 21528 17646 21584
rect 16026 17584 16082 17640
rect 14951 15802 15007 15804
rect 15031 15802 15087 15804
rect 15111 15802 15167 15804
rect 15191 15802 15247 15804
rect 14951 15750 14997 15802
rect 14997 15750 15007 15802
rect 15031 15750 15061 15802
rect 15061 15750 15073 15802
rect 15073 15750 15087 15802
rect 15111 15750 15125 15802
rect 15125 15750 15137 15802
rect 15137 15750 15167 15802
rect 15191 15750 15201 15802
rect 15201 15750 15247 15802
rect 14951 15748 15007 15750
rect 15031 15748 15087 15750
rect 15111 15748 15167 15750
rect 15191 15748 15247 15750
rect 14951 14714 15007 14716
rect 15031 14714 15087 14716
rect 15111 14714 15167 14716
rect 15191 14714 15247 14716
rect 14951 14662 14997 14714
rect 14997 14662 15007 14714
rect 15031 14662 15061 14714
rect 15061 14662 15073 14714
rect 15073 14662 15087 14714
rect 15111 14662 15125 14714
rect 15125 14662 15137 14714
rect 15137 14662 15167 14714
rect 15191 14662 15201 14714
rect 15201 14662 15247 14714
rect 14951 14660 15007 14662
rect 15031 14660 15087 14662
rect 15111 14660 15167 14662
rect 15191 14660 15247 14662
rect 15566 14864 15622 14920
rect 15934 14864 15990 14920
rect 14951 13626 15007 13628
rect 15031 13626 15087 13628
rect 15111 13626 15167 13628
rect 15191 13626 15247 13628
rect 14951 13574 14997 13626
rect 14997 13574 15007 13626
rect 15031 13574 15061 13626
rect 15061 13574 15073 13626
rect 15073 13574 15087 13626
rect 15111 13574 15125 13626
rect 15125 13574 15137 13626
rect 15137 13574 15167 13626
rect 15191 13574 15201 13626
rect 15201 13574 15247 13626
rect 14951 13572 15007 13574
rect 15031 13572 15087 13574
rect 15111 13572 15167 13574
rect 15191 13572 15247 13574
rect 13634 6160 13690 6216
rect 13634 5752 13690 5808
rect 13726 5636 13782 5672
rect 13726 5616 13728 5636
rect 13728 5616 13780 5636
rect 13780 5616 13782 5636
rect 14462 9696 14518 9752
rect 14951 12538 15007 12540
rect 15031 12538 15087 12540
rect 15111 12538 15167 12540
rect 15191 12538 15247 12540
rect 14951 12486 14997 12538
rect 14997 12486 15007 12538
rect 15031 12486 15061 12538
rect 15061 12486 15073 12538
rect 15073 12486 15087 12538
rect 15111 12486 15125 12538
rect 15125 12486 15137 12538
rect 15137 12486 15167 12538
rect 15191 12486 15201 12538
rect 15201 12486 15247 12538
rect 14951 12484 15007 12486
rect 15031 12484 15087 12486
rect 15111 12484 15167 12486
rect 15191 12484 15247 12486
rect 14951 11450 15007 11452
rect 15031 11450 15087 11452
rect 15111 11450 15167 11452
rect 15191 11450 15247 11452
rect 14951 11398 14997 11450
rect 14997 11398 15007 11450
rect 15031 11398 15061 11450
rect 15061 11398 15073 11450
rect 15073 11398 15087 11450
rect 15111 11398 15125 11450
rect 15125 11398 15137 11450
rect 15137 11398 15167 11450
rect 15191 11398 15201 11450
rect 15201 11398 15247 11450
rect 14951 11396 15007 11398
rect 15031 11396 15087 11398
rect 15111 11396 15167 11398
rect 15191 11396 15247 11398
rect 14951 10362 15007 10364
rect 15031 10362 15087 10364
rect 15111 10362 15167 10364
rect 15191 10362 15247 10364
rect 14951 10310 14997 10362
rect 14997 10310 15007 10362
rect 15031 10310 15061 10362
rect 15061 10310 15073 10362
rect 15073 10310 15087 10362
rect 15111 10310 15125 10362
rect 15125 10310 15137 10362
rect 15137 10310 15167 10362
rect 15191 10310 15201 10362
rect 15201 10310 15247 10362
rect 14951 10308 15007 10310
rect 15031 10308 15087 10310
rect 15111 10308 15167 10310
rect 15191 10308 15247 10310
rect 14951 9274 15007 9276
rect 15031 9274 15087 9276
rect 15111 9274 15167 9276
rect 15191 9274 15247 9276
rect 14951 9222 14997 9274
rect 14997 9222 15007 9274
rect 15031 9222 15061 9274
rect 15061 9222 15073 9274
rect 15073 9222 15087 9274
rect 15111 9222 15125 9274
rect 15125 9222 15137 9274
rect 15137 9222 15167 9274
rect 15191 9222 15201 9274
rect 15201 9222 15247 9274
rect 14951 9220 15007 9222
rect 15031 9220 15087 9222
rect 15111 9220 15167 9222
rect 15191 9220 15247 9222
rect 17130 18420 17186 18456
rect 17130 18400 17132 18420
rect 17132 18400 17184 18420
rect 17184 18400 17186 18420
rect 17750 20698 17806 20700
rect 17830 20698 17886 20700
rect 17910 20698 17966 20700
rect 17990 20698 18046 20700
rect 17750 20646 17796 20698
rect 17796 20646 17806 20698
rect 17830 20646 17860 20698
rect 17860 20646 17872 20698
rect 17872 20646 17886 20698
rect 17910 20646 17924 20698
rect 17924 20646 17936 20698
rect 17936 20646 17966 20698
rect 17990 20646 18000 20698
rect 18000 20646 18046 20698
rect 17750 20644 17806 20646
rect 17830 20644 17886 20646
rect 17910 20644 17966 20646
rect 17990 20644 18046 20646
rect 17590 20440 17646 20496
rect 17958 20476 17960 20496
rect 17960 20476 18012 20496
rect 18012 20476 18014 20496
rect 17958 20440 18014 20476
rect 17590 20032 17646 20088
rect 17750 19610 17806 19612
rect 17830 19610 17886 19612
rect 17910 19610 17966 19612
rect 17990 19610 18046 19612
rect 17750 19558 17796 19610
rect 17796 19558 17806 19610
rect 17830 19558 17860 19610
rect 17860 19558 17872 19610
rect 17872 19558 17886 19610
rect 17910 19558 17924 19610
rect 17924 19558 17936 19610
rect 17936 19558 17966 19610
rect 17990 19558 18000 19610
rect 18000 19558 18046 19610
rect 17750 19556 17806 19558
rect 17830 19556 17886 19558
rect 17910 19556 17966 19558
rect 17990 19556 18046 19558
rect 17498 19352 17554 19408
rect 17866 18692 17922 18728
rect 17866 18672 17868 18692
rect 17868 18672 17920 18692
rect 17920 18672 17922 18692
rect 17750 18522 17806 18524
rect 17830 18522 17886 18524
rect 17910 18522 17966 18524
rect 17990 18522 18046 18524
rect 17750 18470 17796 18522
rect 17796 18470 17806 18522
rect 17830 18470 17860 18522
rect 17860 18470 17872 18522
rect 17872 18470 17886 18522
rect 17910 18470 17924 18522
rect 17924 18470 17936 18522
rect 17936 18470 17966 18522
rect 17990 18470 18000 18522
rect 18000 18470 18046 18522
rect 17750 18468 17806 18470
rect 17830 18468 17886 18470
rect 17910 18468 17966 18470
rect 17990 18468 18046 18470
rect 17038 16088 17094 16144
rect 16486 13948 16488 13968
rect 16488 13948 16540 13968
rect 16540 13948 16542 13968
rect 16486 13912 16542 13948
rect 15750 12280 15806 12336
rect 14951 8186 15007 8188
rect 15031 8186 15087 8188
rect 15111 8186 15167 8188
rect 15191 8186 15247 8188
rect 14951 8134 14997 8186
rect 14997 8134 15007 8186
rect 15031 8134 15061 8186
rect 15061 8134 15073 8186
rect 15073 8134 15087 8186
rect 15111 8134 15125 8186
rect 15125 8134 15137 8186
rect 15137 8134 15167 8186
rect 15191 8134 15201 8186
rect 15201 8134 15247 8186
rect 14951 8132 15007 8134
rect 15031 8132 15087 8134
rect 15111 8132 15167 8134
rect 15191 8132 15247 8134
rect 16210 7268 16266 7304
rect 16210 7248 16212 7268
rect 16212 7248 16264 7268
rect 16264 7248 16266 7268
rect 14951 7098 15007 7100
rect 15031 7098 15087 7100
rect 15111 7098 15167 7100
rect 15191 7098 15247 7100
rect 14951 7046 14997 7098
rect 14997 7046 15007 7098
rect 15031 7046 15061 7098
rect 15061 7046 15073 7098
rect 15073 7046 15087 7098
rect 15111 7046 15125 7098
rect 15125 7046 15137 7098
rect 15137 7046 15167 7098
rect 15191 7046 15201 7098
rect 15201 7046 15247 7098
rect 14951 7044 15007 7046
rect 15031 7044 15087 7046
rect 15111 7044 15167 7046
rect 15191 7044 15247 7046
rect 13634 4664 13690 4720
rect 13634 3032 13690 3088
rect 13542 2896 13598 2952
rect 14951 6010 15007 6012
rect 15031 6010 15087 6012
rect 15111 6010 15167 6012
rect 15191 6010 15247 6012
rect 14951 5958 14997 6010
rect 14997 5958 15007 6010
rect 15031 5958 15061 6010
rect 15061 5958 15073 6010
rect 15073 5958 15087 6010
rect 15111 5958 15125 6010
rect 15125 5958 15137 6010
rect 15137 5958 15167 6010
rect 15191 5958 15201 6010
rect 15201 5958 15247 6010
rect 14951 5956 15007 5958
rect 15031 5956 15087 5958
rect 15111 5956 15167 5958
rect 15191 5956 15247 5958
rect 16302 6160 16358 6216
rect 14646 3440 14702 3496
rect 14554 3304 14610 3360
rect 14951 4922 15007 4924
rect 15031 4922 15087 4924
rect 15111 4922 15167 4924
rect 15191 4922 15247 4924
rect 14951 4870 14997 4922
rect 14997 4870 15007 4922
rect 15031 4870 15061 4922
rect 15061 4870 15073 4922
rect 15073 4870 15087 4922
rect 15111 4870 15125 4922
rect 15125 4870 15137 4922
rect 15137 4870 15167 4922
rect 15191 4870 15201 4922
rect 15201 4870 15247 4922
rect 14951 4868 15007 4870
rect 15031 4868 15087 4870
rect 15111 4868 15167 4870
rect 15191 4868 15247 4870
rect 15014 4700 15016 4720
rect 15016 4700 15068 4720
rect 15068 4700 15070 4720
rect 15014 4664 15070 4700
rect 14951 3834 15007 3836
rect 15031 3834 15087 3836
rect 15111 3834 15167 3836
rect 15191 3834 15247 3836
rect 14951 3782 14997 3834
rect 14997 3782 15007 3834
rect 15031 3782 15061 3834
rect 15061 3782 15073 3834
rect 15073 3782 15087 3834
rect 15111 3782 15125 3834
rect 15125 3782 15137 3834
rect 15137 3782 15167 3834
rect 15191 3782 15201 3834
rect 15201 3782 15247 3834
rect 14951 3780 15007 3782
rect 15031 3780 15087 3782
rect 15111 3780 15167 3782
rect 15191 3780 15247 3782
rect 14830 3576 14886 3632
rect 12152 2202 12208 2204
rect 12232 2202 12288 2204
rect 12312 2202 12368 2204
rect 12392 2202 12448 2204
rect 12152 2150 12198 2202
rect 12198 2150 12208 2202
rect 12232 2150 12262 2202
rect 12262 2150 12274 2202
rect 12274 2150 12288 2202
rect 12312 2150 12326 2202
rect 12326 2150 12338 2202
rect 12338 2150 12368 2202
rect 12392 2150 12402 2202
rect 12402 2150 12448 2202
rect 12152 2148 12208 2150
rect 12232 2148 12288 2150
rect 12312 2148 12368 2150
rect 12392 2148 12448 2150
rect 14951 2746 15007 2748
rect 15031 2746 15087 2748
rect 15111 2746 15167 2748
rect 15191 2746 15247 2748
rect 14951 2694 14997 2746
rect 14997 2694 15007 2746
rect 15031 2694 15061 2746
rect 15061 2694 15073 2746
rect 15073 2694 15087 2746
rect 15111 2694 15125 2746
rect 15125 2694 15137 2746
rect 15137 2694 15167 2746
rect 15191 2694 15201 2746
rect 15201 2694 15247 2746
rect 14951 2692 15007 2694
rect 15031 2692 15087 2694
rect 15111 2692 15167 2694
rect 15191 2692 15247 2694
rect 17590 18128 17646 18184
rect 18326 19760 18382 19816
rect 18326 18692 18382 18728
rect 18326 18672 18328 18692
rect 18328 18672 18380 18692
rect 18380 18672 18382 18692
rect 17750 17434 17806 17436
rect 17830 17434 17886 17436
rect 17910 17434 17966 17436
rect 17990 17434 18046 17436
rect 17750 17382 17796 17434
rect 17796 17382 17806 17434
rect 17830 17382 17860 17434
rect 17860 17382 17872 17434
rect 17872 17382 17886 17434
rect 17910 17382 17924 17434
rect 17924 17382 17936 17434
rect 17936 17382 17966 17434
rect 17990 17382 18000 17434
rect 18000 17382 18046 17434
rect 17750 17380 17806 17382
rect 17830 17380 17886 17382
rect 17910 17380 17966 17382
rect 17990 17380 18046 17382
rect 17750 16346 17806 16348
rect 17830 16346 17886 16348
rect 17910 16346 17966 16348
rect 17990 16346 18046 16348
rect 17750 16294 17796 16346
rect 17796 16294 17806 16346
rect 17830 16294 17860 16346
rect 17860 16294 17872 16346
rect 17872 16294 17886 16346
rect 17910 16294 17924 16346
rect 17924 16294 17936 16346
rect 17936 16294 17966 16346
rect 17990 16294 18000 16346
rect 18000 16294 18046 16346
rect 17750 16292 17806 16294
rect 17830 16292 17886 16294
rect 17910 16292 17966 16294
rect 17990 16292 18046 16294
rect 19154 22072 19210 22128
rect 19338 21664 19394 21720
rect 20442 23568 20498 23624
rect 19430 20712 19486 20768
rect 19154 20304 19210 20360
rect 18970 19896 19026 19952
rect 17750 15258 17806 15260
rect 17830 15258 17886 15260
rect 17910 15258 17966 15260
rect 17990 15258 18046 15260
rect 17750 15206 17796 15258
rect 17796 15206 17806 15258
rect 17830 15206 17860 15258
rect 17860 15206 17872 15258
rect 17872 15206 17886 15258
rect 17910 15206 17924 15258
rect 17924 15206 17936 15258
rect 17936 15206 17966 15258
rect 17990 15206 18000 15258
rect 18000 15206 18046 15258
rect 17750 15204 17806 15206
rect 17830 15204 17886 15206
rect 17910 15204 17966 15206
rect 17990 15204 18046 15206
rect 17750 14170 17806 14172
rect 17830 14170 17886 14172
rect 17910 14170 17966 14172
rect 17990 14170 18046 14172
rect 17750 14118 17796 14170
rect 17796 14118 17806 14170
rect 17830 14118 17860 14170
rect 17860 14118 17872 14170
rect 17872 14118 17886 14170
rect 17910 14118 17924 14170
rect 17924 14118 17936 14170
rect 17936 14118 17966 14170
rect 17990 14118 18000 14170
rect 18000 14118 18046 14170
rect 17750 14116 17806 14118
rect 17830 14116 17886 14118
rect 17910 14116 17966 14118
rect 17990 14116 18046 14118
rect 17750 13082 17806 13084
rect 17830 13082 17886 13084
rect 17910 13082 17966 13084
rect 17990 13082 18046 13084
rect 17750 13030 17796 13082
rect 17796 13030 17806 13082
rect 17830 13030 17860 13082
rect 17860 13030 17872 13082
rect 17872 13030 17886 13082
rect 17910 13030 17924 13082
rect 17924 13030 17936 13082
rect 17936 13030 17966 13082
rect 17990 13030 18000 13082
rect 18000 13030 18046 13082
rect 17750 13028 17806 13030
rect 17830 13028 17886 13030
rect 17910 13028 17966 13030
rect 17990 13028 18046 13030
rect 17866 12144 17922 12200
rect 17750 11994 17806 11996
rect 17830 11994 17886 11996
rect 17910 11994 17966 11996
rect 17990 11994 18046 11996
rect 17750 11942 17796 11994
rect 17796 11942 17806 11994
rect 17830 11942 17860 11994
rect 17860 11942 17872 11994
rect 17872 11942 17886 11994
rect 17910 11942 17924 11994
rect 17924 11942 17936 11994
rect 17936 11942 17966 11994
rect 17990 11942 18000 11994
rect 18000 11942 18046 11994
rect 17750 11940 17806 11942
rect 17830 11940 17886 11942
rect 17910 11940 17966 11942
rect 17990 11940 18046 11942
rect 20549 22330 20605 22332
rect 20629 22330 20685 22332
rect 20709 22330 20765 22332
rect 20789 22330 20845 22332
rect 20549 22278 20595 22330
rect 20595 22278 20605 22330
rect 20629 22278 20659 22330
rect 20659 22278 20671 22330
rect 20671 22278 20685 22330
rect 20709 22278 20723 22330
rect 20723 22278 20735 22330
rect 20735 22278 20765 22330
rect 20789 22278 20799 22330
rect 20799 22278 20845 22330
rect 20549 22276 20605 22278
rect 20629 22276 20685 22278
rect 20709 22276 20765 22278
rect 20789 22276 20845 22278
rect 20166 21800 20222 21856
rect 20902 21800 20958 21856
rect 19890 20984 19946 21040
rect 19798 20440 19854 20496
rect 19614 19352 19670 19408
rect 19522 19216 19578 19272
rect 19338 17584 19394 17640
rect 20350 20168 20406 20224
rect 20549 21242 20605 21244
rect 20629 21242 20685 21244
rect 20709 21242 20765 21244
rect 20789 21242 20845 21244
rect 20549 21190 20595 21242
rect 20595 21190 20605 21242
rect 20629 21190 20659 21242
rect 20659 21190 20671 21242
rect 20671 21190 20685 21242
rect 20709 21190 20723 21242
rect 20723 21190 20735 21242
rect 20735 21190 20765 21242
rect 20789 21190 20799 21242
rect 20799 21190 20845 21242
rect 20549 21188 20605 21190
rect 20629 21188 20685 21190
rect 20709 21188 20765 21190
rect 20789 21188 20845 21190
rect 20718 20868 20774 20904
rect 20718 20848 20720 20868
rect 20720 20848 20772 20868
rect 20772 20848 20774 20868
rect 21086 20848 21142 20904
rect 23202 24248 23258 24304
rect 20549 20154 20605 20156
rect 20629 20154 20685 20156
rect 20709 20154 20765 20156
rect 20789 20154 20845 20156
rect 20549 20102 20595 20154
rect 20595 20102 20605 20154
rect 20629 20102 20659 20154
rect 20659 20102 20671 20154
rect 20671 20102 20685 20154
rect 20709 20102 20723 20154
rect 20723 20102 20735 20154
rect 20735 20102 20765 20154
rect 20789 20102 20799 20154
rect 20799 20102 20845 20154
rect 20549 20100 20605 20102
rect 20629 20100 20685 20102
rect 20709 20100 20765 20102
rect 20789 20100 20845 20102
rect 20718 19760 20774 19816
rect 18786 13504 18842 13560
rect 19062 13388 19118 13424
rect 19062 13368 19064 13388
rect 19064 13368 19116 13388
rect 19116 13368 19118 13388
rect 19614 13232 19670 13288
rect 18602 12316 18604 12336
rect 18604 12316 18656 12336
rect 18656 12316 18658 12336
rect 18602 12280 18658 12316
rect 18602 12144 18658 12200
rect 19062 12180 19064 12200
rect 19064 12180 19116 12200
rect 19116 12180 19118 12200
rect 19062 12144 19118 12180
rect 17750 10906 17806 10908
rect 17830 10906 17886 10908
rect 17910 10906 17966 10908
rect 17990 10906 18046 10908
rect 17750 10854 17796 10906
rect 17796 10854 17806 10906
rect 17830 10854 17860 10906
rect 17860 10854 17872 10906
rect 17872 10854 17886 10906
rect 17910 10854 17924 10906
rect 17924 10854 17936 10906
rect 17936 10854 17966 10906
rect 17990 10854 18000 10906
rect 18000 10854 18046 10906
rect 17750 10852 17806 10854
rect 17830 10852 17886 10854
rect 17910 10852 17966 10854
rect 17990 10852 18046 10854
rect 20626 19216 20682 19272
rect 20549 19066 20605 19068
rect 20629 19066 20685 19068
rect 20709 19066 20765 19068
rect 20789 19066 20845 19068
rect 20549 19014 20595 19066
rect 20595 19014 20605 19066
rect 20629 19014 20659 19066
rect 20659 19014 20671 19066
rect 20671 19014 20685 19066
rect 20709 19014 20723 19066
rect 20723 19014 20735 19066
rect 20735 19014 20765 19066
rect 20789 19014 20799 19066
rect 20799 19014 20845 19066
rect 20549 19012 20605 19014
rect 20629 19012 20685 19014
rect 20709 19012 20765 19014
rect 20789 19012 20845 19014
rect 20549 17978 20605 17980
rect 20629 17978 20685 17980
rect 20709 17978 20765 17980
rect 20789 17978 20845 17980
rect 20549 17926 20595 17978
rect 20595 17926 20605 17978
rect 20629 17926 20659 17978
rect 20659 17926 20671 17978
rect 20671 17926 20685 17978
rect 20709 17926 20723 17978
rect 20723 17926 20735 17978
rect 20735 17926 20765 17978
rect 20789 17926 20799 17978
rect 20799 17926 20845 17978
rect 20549 17924 20605 17926
rect 20629 17924 20685 17926
rect 20709 17924 20765 17926
rect 20789 17924 20845 17926
rect 20549 16890 20605 16892
rect 20629 16890 20685 16892
rect 20709 16890 20765 16892
rect 20789 16890 20845 16892
rect 20549 16838 20595 16890
rect 20595 16838 20605 16890
rect 20629 16838 20659 16890
rect 20659 16838 20671 16890
rect 20671 16838 20685 16890
rect 20709 16838 20723 16890
rect 20723 16838 20735 16890
rect 20735 16838 20765 16890
rect 20789 16838 20799 16890
rect 20799 16838 20845 16890
rect 20549 16836 20605 16838
rect 20629 16836 20685 16838
rect 20709 16836 20765 16838
rect 20789 16836 20845 16838
rect 20549 15802 20605 15804
rect 20629 15802 20685 15804
rect 20709 15802 20765 15804
rect 20789 15802 20845 15804
rect 20549 15750 20595 15802
rect 20595 15750 20605 15802
rect 20629 15750 20659 15802
rect 20659 15750 20671 15802
rect 20671 15750 20685 15802
rect 20709 15750 20723 15802
rect 20723 15750 20735 15802
rect 20735 15750 20765 15802
rect 20789 15750 20799 15802
rect 20799 15750 20845 15802
rect 20549 15748 20605 15750
rect 20629 15748 20685 15750
rect 20709 15748 20765 15750
rect 20789 15748 20845 15750
rect 20994 15952 21050 16008
rect 20549 14714 20605 14716
rect 20629 14714 20685 14716
rect 20709 14714 20765 14716
rect 20789 14714 20845 14716
rect 20549 14662 20595 14714
rect 20595 14662 20605 14714
rect 20629 14662 20659 14714
rect 20659 14662 20671 14714
rect 20671 14662 20685 14714
rect 20709 14662 20723 14714
rect 20723 14662 20735 14714
rect 20735 14662 20765 14714
rect 20789 14662 20799 14714
rect 20799 14662 20845 14714
rect 20549 14660 20605 14662
rect 20629 14660 20685 14662
rect 20709 14660 20765 14662
rect 20789 14660 20845 14662
rect 18142 10104 18198 10160
rect 17750 9818 17806 9820
rect 17830 9818 17886 9820
rect 17910 9818 17966 9820
rect 17990 9818 18046 9820
rect 17750 9766 17796 9818
rect 17796 9766 17806 9818
rect 17830 9766 17860 9818
rect 17860 9766 17872 9818
rect 17872 9766 17886 9818
rect 17910 9766 17924 9818
rect 17924 9766 17936 9818
rect 17936 9766 17966 9818
rect 17990 9766 18000 9818
rect 18000 9766 18046 9818
rect 17750 9764 17806 9766
rect 17830 9764 17886 9766
rect 17910 9764 17966 9766
rect 17990 9764 18046 9766
rect 17750 8730 17806 8732
rect 17830 8730 17886 8732
rect 17910 8730 17966 8732
rect 17990 8730 18046 8732
rect 17750 8678 17796 8730
rect 17796 8678 17806 8730
rect 17830 8678 17860 8730
rect 17860 8678 17872 8730
rect 17872 8678 17886 8730
rect 17910 8678 17924 8730
rect 17924 8678 17936 8730
rect 17936 8678 17966 8730
rect 17990 8678 18000 8730
rect 18000 8678 18046 8730
rect 17750 8676 17806 8678
rect 17830 8676 17886 8678
rect 17910 8676 17966 8678
rect 17990 8676 18046 8678
rect 20074 11192 20130 11248
rect 19338 8628 19394 8664
rect 19338 8608 19340 8628
rect 19340 8608 19392 8628
rect 19392 8608 19394 8628
rect 17750 7642 17806 7644
rect 17830 7642 17886 7644
rect 17910 7642 17966 7644
rect 17990 7642 18046 7644
rect 17750 7590 17796 7642
rect 17796 7590 17806 7642
rect 17830 7590 17860 7642
rect 17860 7590 17872 7642
rect 17872 7590 17886 7642
rect 17910 7590 17924 7642
rect 17924 7590 17936 7642
rect 17936 7590 17966 7642
rect 17990 7590 18000 7642
rect 18000 7590 18046 7642
rect 17750 7588 17806 7590
rect 17830 7588 17886 7590
rect 17910 7588 17966 7590
rect 17990 7588 18046 7590
rect 18878 7792 18934 7848
rect 18786 6840 18842 6896
rect 16670 5888 16726 5944
rect 16302 5072 16358 5128
rect 16118 4936 16174 4992
rect 15658 4664 15714 4720
rect 15566 4120 15622 4176
rect 15566 3848 15622 3904
rect 18142 6724 18198 6760
rect 18142 6704 18144 6724
rect 18144 6704 18196 6724
rect 18196 6704 18198 6724
rect 17750 6554 17806 6556
rect 17830 6554 17886 6556
rect 17910 6554 17966 6556
rect 17990 6554 18046 6556
rect 17750 6502 17796 6554
rect 17796 6502 17806 6554
rect 17830 6502 17860 6554
rect 17860 6502 17872 6554
rect 17872 6502 17886 6554
rect 17910 6502 17924 6554
rect 17924 6502 17936 6554
rect 17936 6502 17966 6554
rect 17990 6502 18000 6554
rect 18000 6502 18046 6554
rect 17750 6500 17806 6502
rect 17830 6500 17886 6502
rect 17910 6500 17966 6502
rect 17990 6500 18046 6502
rect 18142 6332 18144 6352
rect 18144 6332 18196 6352
rect 18196 6332 18198 6352
rect 18142 6296 18198 6332
rect 17750 5466 17806 5468
rect 17830 5466 17886 5468
rect 17910 5466 17966 5468
rect 17990 5466 18046 5468
rect 17750 5414 17796 5466
rect 17796 5414 17806 5466
rect 17830 5414 17860 5466
rect 17860 5414 17872 5466
rect 17872 5414 17886 5466
rect 17910 5414 17924 5466
rect 17924 5414 17936 5466
rect 17936 5414 17966 5466
rect 17990 5414 18000 5466
rect 18000 5414 18046 5466
rect 17750 5412 17806 5414
rect 17830 5412 17886 5414
rect 17910 5412 17966 5414
rect 17990 5412 18046 5414
rect 18050 4936 18106 4992
rect 18142 4528 18198 4584
rect 17750 4378 17806 4380
rect 17830 4378 17886 4380
rect 17910 4378 17966 4380
rect 17990 4378 18046 4380
rect 17750 4326 17796 4378
rect 17796 4326 17806 4378
rect 17830 4326 17860 4378
rect 17860 4326 17872 4378
rect 17872 4326 17886 4378
rect 17910 4326 17924 4378
rect 17924 4326 17936 4378
rect 17936 4326 17966 4378
rect 17990 4326 18000 4378
rect 18000 4326 18046 4378
rect 17750 4324 17806 4326
rect 17830 4324 17886 4326
rect 17910 4324 17966 4326
rect 17990 4324 18046 4326
rect 19338 7540 19394 7576
rect 19338 7520 19340 7540
rect 19340 7520 19392 7540
rect 19392 7520 19394 7540
rect 19338 6840 19394 6896
rect 19890 5788 19892 5808
rect 19892 5788 19944 5808
rect 19944 5788 19946 5808
rect 19890 5752 19946 5788
rect 19614 5072 19670 5128
rect 19062 4120 19118 4176
rect 16210 2488 16266 2544
rect 17750 3290 17806 3292
rect 17830 3290 17886 3292
rect 17910 3290 17966 3292
rect 17990 3290 18046 3292
rect 17750 3238 17796 3290
rect 17796 3238 17806 3290
rect 17830 3238 17860 3290
rect 17860 3238 17872 3290
rect 17872 3238 17886 3290
rect 17910 3238 17924 3290
rect 17924 3238 17936 3290
rect 17936 3238 17966 3290
rect 17990 3238 18000 3290
rect 18000 3238 18046 3290
rect 17750 3236 17806 3238
rect 17830 3236 17886 3238
rect 17910 3236 17966 3238
rect 17990 3236 18046 3238
rect 17750 2202 17806 2204
rect 17830 2202 17886 2204
rect 17910 2202 17966 2204
rect 17990 2202 18046 2204
rect 17750 2150 17796 2202
rect 17796 2150 17806 2202
rect 17830 2150 17860 2202
rect 17860 2150 17872 2202
rect 17872 2150 17886 2202
rect 17910 2150 17924 2202
rect 17924 2150 17936 2202
rect 17936 2150 17966 2202
rect 17990 2150 18000 2202
rect 18000 2150 18046 2202
rect 17750 2148 17806 2150
rect 17830 2148 17886 2150
rect 17910 2148 17966 2150
rect 17990 2148 18046 2150
rect 18142 1944 18198 2000
rect 18418 1808 18474 1864
rect 18970 1672 19026 1728
rect 19522 3848 19578 3904
rect 19246 3032 19302 3088
rect 19982 4256 20038 4312
rect 20442 13776 20498 13832
rect 20549 13626 20605 13628
rect 20629 13626 20685 13628
rect 20709 13626 20765 13628
rect 20789 13626 20845 13628
rect 20549 13574 20595 13626
rect 20595 13574 20605 13626
rect 20629 13574 20659 13626
rect 20659 13574 20671 13626
rect 20671 13574 20685 13626
rect 20709 13574 20723 13626
rect 20723 13574 20735 13626
rect 20735 13574 20765 13626
rect 20789 13574 20799 13626
rect 20799 13574 20845 13626
rect 20549 13572 20605 13574
rect 20629 13572 20685 13574
rect 20709 13572 20765 13574
rect 20789 13572 20845 13574
rect 20442 13368 20498 13424
rect 20549 12538 20605 12540
rect 20629 12538 20685 12540
rect 20709 12538 20765 12540
rect 20789 12538 20845 12540
rect 20549 12486 20595 12538
rect 20595 12486 20605 12538
rect 20629 12486 20659 12538
rect 20659 12486 20671 12538
rect 20671 12486 20685 12538
rect 20709 12486 20723 12538
rect 20723 12486 20735 12538
rect 20735 12486 20765 12538
rect 20789 12486 20799 12538
rect 20799 12486 20845 12538
rect 20549 12484 20605 12486
rect 20629 12484 20685 12486
rect 20709 12484 20765 12486
rect 20789 12484 20845 12486
rect 20994 12824 21050 12880
rect 20549 11450 20605 11452
rect 20629 11450 20685 11452
rect 20709 11450 20765 11452
rect 20789 11450 20845 11452
rect 20549 11398 20595 11450
rect 20595 11398 20605 11450
rect 20629 11398 20659 11450
rect 20659 11398 20671 11450
rect 20671 11398 20685 11450
rect 20709 11398 20723 11450
rect 20723 11398 20735 11450
rect 20735 11398 20765 11450
rect 20789 11398 20799 11450
rect 20799 11398 20845 11450
rect 20549 11396 20605 11398
rect 20629 11396 20685 11398
rect 20709 11396 20765 11398
rect 20789 11396 20845 11398
rect 20902 11192 20958 11248
rect 22006 22888 22062 22944
rect 21638 21548 21694 21584
rect 21638 21528 21640 21548
rect 21640 21528 21692 21548
rect 21692 21528 21694 21548
rect 21638 20324 21694 20360
rect 21638 20304 21640 20324
rect 21640 20304 21692 20324
rect 21692 20304 21694 20324
rect 21454 18284 21510 18320
rect 21454 18264 21456 18284
rect 21456 18264 21508 18284
rect 21508 18264 21510 18284
rect 21546 17720 21602 17776
rect 22098 21528 22154 21584
rect 22006 20576 22062 20632
rect 22282 20576 22338 20632
rect 20549 10362 20605 10364
rect 20629 10362 20685 10364
rect 20709 10362 20765 10364
rect 20789 10362 20845 10364
rect 20549 10310 20595 10362
rect 20595 10310 20605 10362
rect 20629 10310 20659 10362
rect 20659 10310 20671 10362
rect 20671 10310 20685 10362
rect 20709 10310 20723 10362
rect 20723 10310 20735 10362
rect 20735 10310 20765 10362
rect 20789 10310 20799 10362
rect 20799 10310 20845 10362
rect 20549 10308 20605 10310
rect 20629 10308 20685 10310
rect 20709 10308 20765 10310
rect 20789 10308 20845 10310
rect 20549 9274 20605 9276
rect 20629 9274 20685 9276
rect 20709 9274 20765 9276
rect 20789 9274 20845 9276
rect 20549 9222 20595 9274
rect 20595 9222 20605 9274
rect 20629 9222 20659 9274
rect 20659 9222 20671 9274
rect 20671 9222 20685 9274
rect 20709 9222 20723 9274
rect 20723 9222 20735 9274
rect 20735 9222 20765 9274
rect 20789 9222 20799 9274
rect 20799 9222 20845 9274
rect 20549 9220 20605 9222
rect 20629 9220 20685 9222
rect 20709 9220 20765 9222
rect 20789 9220 20845 9222
rect 21454 12824 21510 12880
rect 22282 19352 22338 19408
rect 22190 17448 22246 17504
rect 22558 19352 22614 19408
rect 22558 17856 22614 17912
rect 20549 8186 20605 8188
rect 20629 8186 20685 8188
rect 20709 8186 20765 8188
rect 20789 8186 20845 8188
rect 20549 8134 20595 8186
rect 20595 8134 20605 8186
rect 20629 8134 20659 8186
rect 20659 8134 20671 8186
rect 20671 8134 20685 8186
rect 20709 8134 20723 8186
rect 20723 8134 20735 8186
rect 20735 8134 20765 8186
rect 20789 8134 20799 8186
rect 20799 8134 20845 8186
rect 20549 8132 20605 8134
rect 20629 8132 20685 8134
rect 20709 8132 20765 8134
rect 20789 8132 20845 8134
rect 19706 2896 19762 2952
rect 20549 7098 20605 7100
rect 20629 7098 20685 7100
rect 20709 7098 20765 7100
rect 20789 7098 20845 7100
rect 20549 7046 20595 7098
rect 20595 7046 20605 7098
rect 20629 7046 20659 7098
rect 20659 7046 20671 7098
rect 20671 7046 20685 7098
rect 20709 7046 20723 7098
rect 20723 7046 20735 7098
rect 20735 7046 20765 7098
rect 20789 7046 20799 7098
rect 20799 7046 20845 7098
rect 20549 7044 20605 7046
rect 20629 7044 20685 7046
rect 20709 7044 20765 7046
rect 20789 7044 20845 7046
rect 20549 6010 20605 6012
rect 20629 6010 20685 6012
rect 20709 6010 20765 6012
rect 20789 6010 20845 6012
rect 20549 5958 20595 6010
rect 20595 5958 20605 6010
rect 20629 5958 20659 6010
rect 20659 5958 20671 6010
rect 20671 5958 20685 6010
rect 20709 5958 20723 6010
rect 20723 5958 20735 6010
rect 20735 5958 20765 6010
rect 20789 5958 20799 6010
rect 20799 5958 20845 6010
rect 20549 5956 20605 5958
rect 20629 5956 20685 5958
rect 20709 5956 20765 5958
rect 20789 5956 20845 5958
rect 20549 4922 20605 4924
rect 20629 4922 20685 4924
rect 20709 4922 20765 4924
rect 20789 4922 20845 4924
rect 20549 4870 20595 4922
rect 20595 4870 20605 4922
rect 20629 4870 20659 4922
rect 20659 4870 20671 4922
rect 20671 4870 20685 4922
rect 20709 4870 20723 4922
rect 20723 4870 20735 4922
rect 20735 4870 20765 4922
rect 20789 4870 20799 4922
rect 20799 4870 20845 4922
rect 20549 4868 20605 4870
rect 20629 4868 20685 4870
rect 20709 4868 20765 4870
rect 20789 4868 20845 4870
rect 20442 4664 20498 4720
rect 21362 8200 21418 8256
rect 21546 7248 21602 7304
rect 21454 6724 21510 6760
rect 21454 6704 21456 6724
rect 21456 6704 21508 6724
rect 21508 6704 21510 6724
rect 21270 4664 21326 4720
rect 22834 21936 22890 21992
rect 23018 20304 23074 20360
rect 23110 20168 23166 20224
rect 23018 19760 23074 19816
rect 23018 19488 23074 19544
rect 22834 18808 22890 18864
rect 22834 17312 22890 17368
rect 22834 17212 22836 17232
rect 22836 17212 22888 17232
rect 22888 17212 22890 17232
rect 22834 17176 22890 17212
rect 22834 16224 22890 16280
rect 23018 16224 23074 16280
rect 22926 16088 22982 16144
rect 22926 13912 22982 13968
rect 22558 13504 22614 13560
rect 21914 10512 21970 10568
rect 21914 10104 21970 10160
rect 22834 12280 22890 12336
rect 21546 5072 21602 5128
rect 21546 4936 21602 4992
rect 20350 3984 20406 4040
rect 20549 3834 20605 3836
rect 20629 3834 20685 3836
rect 20709 3834 20765 3836
rect 20789 3834 20845 3836
rect 20549 3782 20595 3834
rect 20595 3782 20605 3834
rect 20629 3782 20659 3834
rect 20659 3782 20671 3834
rect 20671 3782 20685 3834
rect 20709 3782 20723 3834
rect 20723 3782 20735 3834
rect 20735 3782 20765 3834
rect 20789 3782 20799 3834
rect 20799 3782 20845 3834
rect 20549 3780 20605 3782
rect 20629 3780 20685 3782
rect 20709 3780 20765 3782
rect 20789 3780 20845 3782
rect 20534 3576 20590 3632
rect 20718 3460 20774 3496
rect 20718 3440 20720 3460
rect 20720 3440 20772 3460
rect 20772 3440 20774 3460
rect 20810 3188 20866 3224
rect 20810 3168 20812 3188
rect 20812 3168 20864 3188
rect 20864 3168 20866 3188
rect 20549 2746 20605 2748
rect 20629 2746 20685 2748
rect 20709 2746 20765 2748
rect 20789 2746 20845 2748
rect 20549 2694 20595 2746
rect 20595 2694 20605 2746
rect 20629 2694 20659 2746
rect 20659 2694 20671 2746
rect 20671 2694 20685 2746
rect 20709 2694 20723 2746
rect 20723 2694 20735 2746
rect 20735 2694 20765 2746
rect 20789 2694 20799 2746
rect 20799 2694 20845 2746
rect 20549 2692 20605 2694
rect 20629 2692 20685 2694
rect 20709 2692 20765 2694
rect 20789 2692 20845 2694
rect 21454 4564 21456 4584
rect 21456 4564 21508 4584
rect 21508 4564 21510 4584
rect 21454 4528 21510 4564
rect 21270 4120 21326 4176
rect 21362 3052 21418 3088
rect 21362 3032 21364 3052
rect 21364 3032 21416 3052
rect 21416 3032 21418 3052
rect 19338 2372 19394 2408
rect 19338 2352 19340 2372
rect 19340 2352 19392 2372
rect 19392 2352 19394 2372
rect 20166 2216 20222 2272
rect 20258 1536 20314 1592
rect 22282 6160 22338 6216
rect 22282 5752 22338 5808
rect 23202 14864 23258 14920
rect 23110 14184 23166 14240
rect 23110 13268 23112 13288
rect 23112 13268 23164 13288
rect 23164 13268 23166 13288
rect 23110 13232 23166 13268
rect 23018 12144 23074 12200
rect 23110 11600 23166 11656
rect 23110 10920 23166 10976
rect 23018 10240 23074 10296
rect 22926 8880 22982 8936
rect 22650 7384 22706 7440
rect 23018 6840 23074 6896
rect 23018 6296 23074 6352
rect 22834 5616 22890 5672
rect 23018 5616 23074 5672
rect 23386 15544 23442 15600
rect 23754 18536 23810 18592
rect 23938 16496 23994 16552
rect 23294 9560 23350 9616
rect 23386 8880 23442 8936
rect 23294 8608 23350 8664
rect 22742 3576 22798 3632
rect 22650 3168 22706 3224
rect 21546 856 21602 912
rect 19062 312 19118 368
<< metal3 >>
rect 23197 24306 23263 24309
rect 23800 24306 24600 24336
rect 23197 24304 24600 24306
rect 23197 24248 23202 24304
rect 23258 24248 24600 24304
rect 23197 24246 24600 24248
rect 23197 24243 23263 24246
rect 23800 24216 24600 24246
rect 20437 23626 20503 23629
rect 23800 23626 24600 23656
rect 20437 23624 24600 23626
rect 20437 23568 20442 23624
rect 20498 23568 24600 23624
rect 20437 23566 24600 23568
rect 20437 23563 20503 23566
rect 23800 23536 24600 23566
rect 22001 22946 22067 22949
rect 23800 22946 24600 22976
rect 22001 22944 24600 22946
rect 22001 22888 22006 22944
rect 22062 22888 24600 22944
rect 22001 22886 24600 22888
rect 22001 22883 22067 22886
rect 23800 22856 24600 22886
rect 3743 22336 4063 22337
rect 3743 22272 3751 22336
rect 3815 22272 3831 22336
rect 3895 22272 3911 22336
rect 3975 22272 3991 22336
rect 4055 22272 4063 22336
rect 3743 22271 4063 22272
rect 9341 22336 9661 22337
rect 9341 22272 9349 22336
rect 9413 22272 9429 22336
rect 9493 22272 9509 22336
rect 9573 22272 9589 22336
rect 9653 22272 9661 22336
rect 9341 22271 9661 22272
rect 14939 22336 15259 22337
rect 14939 22272 14947 22336
rect 15011 22272 15027 22336
rect 15091 22272 15107 22336
rect 15171 22272 15187 22336
rect 15251 22272 15259 22336
rect 14939 22271 15259 22272
rect 20537 22336 20857 22337
rect 20537 22272 20545 22336
rect 20609 22272 20625 22336
rect 20689 22272 20705 22336
rect 20769 22272 20785 22336
rect 20849 22272 20857 22336
rect 20537 22271 20857 22272
rect 23800 22266 24600 22296
rect 22050 22206 24600 22266
rect 19149 22130 19215 22133
rect 22050 22130 22110 22206
rect 23800 22176 24600 22206
rect 19149 22128 22110 22130
rect 19149 22072 19154 22128
rect 19210 22072 22110 22128
rect 19149 22070 22110 22072
rect 19149 22067 19215 22070
rect 9121 21996 9187 21997
rect 9070 21932 9076 21996
rect 9140 21994 9187 21996
rect 10133 21994 10199 21997
rect 12157 21994 12223 21997
rect 9140 21992 9232 21994
rect 9182 21936 9232 21992
rect 9140 21934 9232 21936
rect 10133 21992 12223 21994
rect 10133 21936 10138 21992
rect 10194 21936 12162 21992
rect 12218 21936 12223 21992
rect 10133 21934 12223 21936
rect 9140 21932 9187 21934
rect 9121 21931 9187 21932
rect 10133 21931 10199 21934
rect 12157 21931 12223 21934
rect 12433 21994 12499 21997
rect 22829 21994 22895 21997
rect 12433 21992 22895 21994
rect 12433 21936 12438 21992
rect 12494 21936 22834 21992
rect 22890 21936 22895 21992
rect 12433 21934 22895 21936
rect 12433 21931 12499 21934
rect 22829 21931 22895 21934
rect 20161 21858 20227 21861
rect 20897 21858 20963 21861
rect 20161 21856 20963 21858
rect 20161 21800 20166 21856
rect 20222 21800 20902 21856
rect 20958 21800 20963 21856
rect 20161 21798 20963 21800
rect 20161 21795 20227 21798
rect 20897 21795 20963 21798
rect 6542 21792 6862 21793
rect 6542 21728 6550 21792
rect 6614 21728 6630 21792
rect 6694 21728 6710 21792
rect 6774 21728 6790 21792
rect 6854 21728 6862 21792
rect 6542 21727 6862 21728
rect 12140 21792 12460 21793
rect 12140 21728 12148 21792
rect 12212 21728 12228 21792
rect 12292 21728 12308 21792
rect 12372 21728 12388 21792
rect 12452 21728 12460 21792
rect 12140 21727 12460 21728
rect 17738 21792 18058 21793
rect 17738 21728 17746 21792
rect 17810 21728 17826 21792
rect 17890 21728 17906 21792
rect 17970 21728 17986 21792
rect 18050 21728 18058 21792
rect 17738 21727 18058 21728
rect 14641 21722 14707 21725
rect 16113 21722 16179 21725
rect 14641 21720 16179 21722
rect 14641 21664 14646 21720
rect 14702 21664 16118 21720
rect 16174 21664 16179 21720
rect 14641 21662 16179 21664
rect 14641 21659 14707 21662
rect 16113 21659 16179 21662
rect 19333 21722 19399 21725
rect 19333 21720 22386 21722
rect 19333 21664 19338 21720
rect 19394 21664 22386 21720
rect 19333 21662 22386 21664
rect 19333 21659 19399 21662
rect 8477 21586 8543 21589
rect 17585 21586 17651 21589
rect 21633 21586 21699 21589
rect 22093 21586 22159 21589
rect 8477 21584 17651 21586
rect 8477 21528 8482 21584
rect 8538 21528 17590 21584
rect 17646 21528 17651 21584
rect 8477 21526 17651 21528
rect 8477 21523 8543 21526
rect 17585 21523 17651 21526
rect 17726 21584 21699 21586
rect 17726 21528 21638 21584
rect 21694 21528 21699 21584
rect 17726 21526 21699 21528
rect 0 21360 800 21480
rect 7649 21450 7715 21453
rect 9673 21450 9739 21453
rect 7649 21448 9739 21450
rect 7649 21392 7654 21448
rect 7710 21392 9678 21448
rect 9734 21392 9739 21448
rect 7649 21390 9739 21392
rect 7649 21387 7715 21390
rect 9673 21387 9739 21390
rect 14457 21450 14523 21453
rect 15929 21450 15995 21453
rect 14457 21448 15995 21450
rect 14457 21392 14462 21448
rect 14518 21392 15934 21448
rect 15990 21392 15995 21448
rect 14457 21390 15995 21392
rect 14457 21387 14523 21390
rect 15929 21387 15995 21390
rect 16113 21450 16179 21453
rect 17726 21450 17786 21526
rect 21633 21523 21699 21526
rect 22050 21584 22159 21586
rect 22050 21528 22098 21584
rect 22154 21528 22159 21584
rect 22050 21523 22159 21528
rect 22326 21586 22386 21662
rect 23800 21586 24600 21616
rect 22326 21526 24600 21586
rect 22050 21450 22110 21523
rect 23800 21496 24600 21526
rect 16113 21448 17786 21450
rect 16113 21392 16118 21448
rect 16174 21392 17786 21448
rect 16113 21390 17786 21392
rect 20302 21390 22110 21450
rect 16113 21387 16179 21390
rect 15469 21314 15535 21317
rect 20302 21314 20362 21390
rect 15469 21312 20362 21314
rect 15469 21256 15474 21312
rect 15530 21256 20362 21312
rect 15469 21254 20362 21256
rect 15469 21251 15535 21254
rect 3743 21248 4063 21249
rect 3743 21184 3751 21248
rect 3815 21184 3831 21248
rect 3895 21184 3911 21248
rect 3975 21184 3991 21248
rect 4055 21184 4063 21248
rect 3743 21183 4063 21184
rect 9341 21248 9661 21249
rect 9341 21184 9349 21248
rect 9413 21184 9429 21248
rect 9493 21184 9509 21248
rect 9573 21184 9589 21248
rect 9653 21184 9661 21248
rect 9341 21183 9661 21184
rect 14939 21248 15259 21249
rect 14939 21184 14947 21248
rect 15011 21184 15027 21248
rect 15091 21184 15107 21248
rect 15171 21184 15187 21248
rect 15251 21184 15259 21248
rect 14939 21183 15259 21184
rect 20537 21248 20857 21249
rect 20537 21184 20545 21248
rect 20609 21184 20625 21248
rect 20689 21184 20705 21248
rect 20769 21184 20785 21248
rect 20849 21184 20857 21248
rect 20537 21183 20857 21184
rect 8569 21042 8635 21045
rect 17033 21042 17099 21045
rect 8569 21040 17099 21042
rect 8569 20984 8574 21040
rect 8630 20984 17038 21040
rect 17094 20984 17099 21040
rect 8569 20982 17099 20984
rect 8569 20979 8635 20982
rect 17033 20979 17099 20982
rect 19374 20980 19380 21044
rect 19444 21042 19450 21044
rect 19885 21042 19951 21045
rect 19444 21040 19951 21042
rect 19444 20984 19890 21040
rect 19946 20984 19951 21040
rect 19444 20982 19951 20984
rect 19444 20980 19450 20982
rect 19885 20979 19951 20982
rect 9029 20906 9095 20909
rect 9305 20906 9371 20909
rect 9029 20904 9371 20906
rect 9029 20848 9034 20904
rect 9090 20848 9310 20904
rect 9366 20848 9371 20904
rect 9029 20846 9371 20848
rect 9029 20843 9095 20846
rect 9305 20843 9371 20846
rect 10501 20906 10567 20909
rect 14917 20906 14983 20909
rect 20713 20906 20779 20909
rect 10501 20904 14842 20906
rect 10501 20848 10506 20904
rect 10562 20848 14842 20904
rect 10501 20846 14842 20848
rect 10501 20843 10567 20846
rect 14782 20770 14842 20846
rect 14917 20904 20779 20906
rect 14917 20848 14922 20904
rect 14978 20848 20718 20904
rect 20774 20848 20779 20904
rect 14917 20846 20779 20848
rect 14917 20843 14983 20846
rect 20713 20843 20779 20846
rect 21081 20906 21147 20909
rect 21214 20906 21220 20908
rect 21081 20904 21220 20906
rect 21081 20848 21086 20904
rect 21142 20848 21220 20904
rect 21081 20846 21220 20848
rect 21081 20843 21147 20846
rect 21214 20844 21220 20846
rect 21284 20844 21290 20908
rect 23800 20906 24600 20936
rect 22050 20846 24600 20906
rect 19425 20770 19491 20773
rect 22050 20770 22110 20846
rect 23800 20816 24600 20846
rect 14782 20710 16130 20770
rect 6542 20704 6862 20705
rect 6542 20640 6550 20704
rect 6614 20640 6630 20704
rect 6694 20640 6710 20704
rect 6774 20640 6790 20704
rect 6854 20640 6862 20704
rect 6542 20639 6862 20640
rect 12140 20704 12460 20705
rect 12140 20640 12148 20704
rect 12212 20640 12228 20704
rect 12292 20640 12308 20704
rect 12372 20640 12388 20704
rect 12452 20640 12460 20704
rect 12140 20639 12460 20640
rect 16070 20634 16130 20710
rect 19425 20768 22110 20770
rect 19425 20712 19430 20768
rect 19486 20712 22110 20768
rect 19425 20710 22110 20712
rect 19425 20707 19491 20710
rect 17738 20704 18058 20705
rect 17738 20640 17746 20704
rect 17810 20640 17826 20704
rect 17890 20640 17906 20704
rect 17970 20640 17986 20704
rect 18050 20640 18058 20704
rect 17738 20639 18058 20640
rect 16205 20634 16271 20637
rect 16070 20632 16271 20634
rect 16070 20576 16210 20632
rect 16266 20576 16271 20632
rect 16070 20574 16271 20576
rect 16205 20571 16271 20574
rect 22001 20634 22067 20637
rect 22277 20634 22343 20637
rect 22001 20632 22343 20634
rect 22001 20576 22006 20632
rect 22062 20576 22282 20632
rect 22338 20576 22343 20632
rect 22001 20574 22343 20576
rect 22001 20571 22067 20574
rect 22277 20571 22343 20574
rect 13261 20498 13327 20501
rect 17585 20498 17651 20501
rect 13261 20496 17651 20498
rect 13261 20440 13266 20496
rect 13322 20440 17590 20496
rect 17646 20440 17651 20496
rect 13261 20438 17651 20440
rect 13261 20435 13327 20438
rect 17585 20435 17651 20438
rect 17953 20498 18019 20501
rect 19793 20498 19859 20501
rect 17953 20496 19859 20498
rect 17953 20440 17958 20496
rect 18014 20440 19798 20496
rect 19854 20440 19859 20496
rect 17953 20438 19859 20440
rect 17953 20435 18019 20438
rect 19793 20435 19859 20438
rect 9213 20362 9279 20365
rect 10133 20362 10199 20365
rect 9213 20360 10199 20362
rect 9213 20304 9218 20360
rect 9274 20304 10138 20360
rect 10194 20304 10199 20360
rect 9213 20302 10199 20304
rect 9213 20299 9279 20302
rect 10133 20299 10199 20302
rect 14825 20362 14891 20365
rect 19149 20362 19215 20365
rect 21633 20362 21699 20365
rect 14825 20360 19074 20362
rect 14825 20304 14830 20360
rect 14886 20304 19074 20360
rect 14825 20302 19074 20304
rect 14825 20299 14891 20302
rect 19014 20226 19074 20302
rect 19149 20360 21699 20362
rect 19149 20304 19154 20360
rect 19210 20304 21638 20360
rect 21694 20304 21699 20360
rect 19149 20302 21699 20304
rect 19149 20299 19215 20302
rect 21633 20299 21699 20302
rect 22870 20300 22876 20364
rect 22940 20362 22946 20364
rect 23013 20362 23079 20365
rect 22940 20360 23079 20362
rect 22940 20304 23018 20360
rect 23074 20304 23079 20360
rect 22940 20302 23079 20304
rect 22940 20300 22946 20302
rect 23013 20299 23079 20302
rect 20345 20226 20411 20229
rect 19014 20224 20411 20226
rect 19014 20168 20350 20224
rect 20406 20168 20411 20224
rect 19014 20166 20411 20168
rect 20345 20163 20411 20166
rect 23105 20226 23171 20229
rect 23800 20226 24600 20256
rect 23105 20224 24600 20226
rect 23105 20168 23110 20224
rect 23166 20168 24600 20224
rect 23105 20166 24600 20168
rect 23105 20163 23171 20166
rect 3743 20160 4063 20161
rect 3743 20096 3751 20160
rect 3815 20096 3831 20160
rect 3895 20096 3911 20160
rect 3975 20096 3991 20160
rect 4055 20096 4063 20160
rect 3743 20095 4063 20096
rect 9341 20160 9661 20161
rect 9341 20096 9349 20160
rect 9413 20096 9429 20160
rect 9493 20096 9509 20160
rect 9573 20096 9589 20160
rect 9653 20096 9661 20160
rect 9341 20095 9661 20096
rect 14939 20160 15259 20161
rect 14939 20096 14947 20160
rect 15011 20096 15027 20160
rect 15091 20096 15107 20160
rect 15171 20096 15187 20160
rect 15251 20096 15259 20160
rect 14939 20095 15259 20096
rect 20537 20160 20857 20161
rect 20537 20096 20545 20160
rect 20609 20096 20625 20160
rect 20689 20096 20705 20160
rect 20769 20096 20785 20160
rect 20849 20096 20857 20160
rect 23800 20136 24600 20166
rect 20537 20095 20857 20096
rect 7833 20090 7899 20093
rect 7966 20090 7972 20092
rect 7833 20088 7972 20090
rect 7833 20032 7838 20088
rect 7894 20032 7972 20088
rect 7833 20030 7972 20032
rect 7833 20027 7899 20030
rect 7966 20028 7972 20030
rect 8036 20028 8042 20092
rect 17585 20090 17651 20093
rect 17585 20088 20362 20090
rect 17585 20032 17590 20088
rect 17646 20032 20362 20088
rect 17585 20030 20362 20032
rect 17585 20027 17651 20030
rect 14089 19954 14155 19957
rect 18965 19954 19031 19957
rect 14089 19952 19031 19954
rect 14089 19896 14094 19952
rect 14150 19896 18970 19952
rect 19026 19896 19031 19952
rect 14089 19894 19031 19896
rect 14089 19891 14155 19894
rect 18965 19891 19031 19894
rect 9673 19818 9739 19821
rect 10225 19818 10291 19821
rect 9673 19816 10291 19818
rect 9673 19760 9678 19816
rect 9734 19760 10230 19816
rect 10286 19760 10291 19816
rect 9673 19758 10291 19760
rect 9673 19755 9739 19758
rect 10225 19755 10291 19758
rect 11145 19818 11211 19821
rect 18321 19818 18387 19821
rect 11145 19816 18387 19818
rect 11145 19760 11150 19816
rect 11206 19760 18326 19816
rect 18382 19760 18387 19816
rect 11145 19758 18387 19760
rect 11145 19755 11211 19758
rect 18321 19755 18387 19758
rect 6542 19616 6862 19617
rect 6542 19552 6550 19616
rect 6614 19552 6630 19616
rect 6694 19552 6710 19616
rect 6774 19552 6790 19616
rect 6854 19552 6862 19616
rect 6542 19551 6862 19552
rect 12140 19616 12460 19617
rect 12140 19552 12148 19616
rect 12212 19552 12228 19616
rect 12292 19552 12308 19616
rect 12372 19552 12388 19616
rect 12452 19552 12460 19616
rect 12140 19551 12460 19552
rect 17738 19616 18058 19617
rect 17738 19552 17746 19616
rect 17810 19552 17826 19616
rect 17890 19552 17906 19616
rect 17970 19552 17986 19616
rect 18050 19552 18058 19616
rect 17738 19551 18058 19552
rect 7005 19546 7071 19549
rect 10041 19546 10107 19549
rect 7005 19544 10107 19546
rect 7005 19488 7010 19544
rect 7066 19488 10046 19544
rect 10102 19488 10107 19544
rect 7005 19486 10107 19488
rect 20302 19546 20362 20030
rect 20713 19818 20779 19821
rect 23013 19818 23079 19821
rect 20713 19816 23079 19818
rect 20713 19760 20718 19816
rect 20774 19760 23018 19816
rect 23074 19760 23079 19816
rect 20713 19758 23079 19760
rect 20713 19755 20779 19758
rect 23013 19755 23079 19758
rect 23013 19546 23079 19549
rect 23800 19546 24600 19576
rect 20302 19486 22110 19546
rect 7005 19483 7071 19486
rect 10041 19483 10107 19486
rect 7005 19410 7071 19413
rect 7833 19410 7899 19413
rect 8109 19410 8175 19413
rect 7005 19408 8175 19410
rect 7005 19352 7010 19408
rect 7066 19352 7838 19408
rect 7894 19352 8114 19408
rect 8170 19352 8175 19408
rect 7005 19350 8175 19352
rect 7005 19347 7071 19350
rect 7833 19347 7899 19350
rect 8109 19347 8175 19350
rect 17493 19410 17559 19413
rect 19609 19410 19675 19413
rect 17493 19408 19675 19410
rect 17493 19352 17498 19408
rect 17554 19352 19614 19408
rect 19670 19352 19675 19408
rect 17493 19350 19675 19352
rect 22050 19410 22110 19486
rect 23013 19544 24600 19546
rect 23013 19488 23018 19544
rect 23074 19488 24600 19544
rect 23013 19486 24600 19488
rect 23013 19483 23079 19486
rect 23800 19456 24600 19486
rect 22277 19410 22343 19413
rect 22553 19410 22619 19413
rect 22050 19408 22619 19410
rect 22050 19352 22282 19408
rect 22338 19352 22558 19408
rect 22614 19352 22619 19408
rect 22050 19350 22619 19352
rect 17493 19347 17559 19350
rect 19609 19347 19675 19350
rect 22277 19347 22343 19350
rect 22553 19347 22619 19350
rect 3417 19274 3483 19277
rect 19517 19274 19583 19277
rect 20621 19274 20687 19277
rect 3417 19272 20687 19274
rect 3417 19216 3422 19272
rect 3478 19216 19522 19272
rect 19578 19216 20626 19272
rect 20682 19216 20687 19272
rect 3417 19214 20687 19216
rect 3417 19211 3483 19214
rect 19517 19211 19583 19214
rect 20621 19211 20687 19214
rect 3743 19072 4063 19073
rect 3743 19008 3751 19072
rect 3815 19008 3831 19072
rect 3895 19008 3911 19072
rect 3975 19008 3991 19072
rect 4055 19008 4063 19072
rect 3743 19007 4063 19008
rect 9341 19072 9661 19073
rect 9341 19008 9349 19072
rect 9413 19008 9429 19072
rect 9493 19008 9509 19072
rect 9573 19008 9589 19072
rect 9653 19008 9661 19072
rect 9341 19007 9661 19008
rect 14939 19072 15259 19073
rect 14939 19008 14947 19072
rect 15011 19008 15027 19072
rect 15091 19008 15107 19072
rect 15171 19008 15187 19072
rect 15251 19008 15259 19072
rect 14939 19007 15259 19008
rect 20537 19072 20857 19073
rect 20537 19008 20545 19072
rect 20609 19008 20625 19072
rect 20689 19008 20705 19072
rect 20769 19008 20785 19072
rect 20849 19008 20857 19072
rect 20537 19007 20857 19008
rect 7189 18866 7255 18869
rect 9305 18866 9371 18869
rect 7189 18864 9371 18866
rect 7189 18808 7194 18864
rect 7250 18808 9310 18864
rect 9366 18808 9371 18864
rect 7189 18806 9371 18808
rect 7189 18803 7255 18806
rect 9305 18803 9371 18806
rect 11697 18866 11763 18869
rect 22829 18866 22895 18869
rect 23800 18866 24600 18896
rect 11697 18864 22895 18866
rect 11697 18808 11702 18864
rect 11758 18808 22834 18864
rect 22890 18808 22895 18864
rect 11697 18806 22895 18808
rect 11697 18803 11763 18806
rect 22829 18803 22895 18806
rect 23614 18806 24600 18866
rect 17861 18730 17927 18733
rect 18321 18730 18387 18733
rect 17861 18728 18387 18730
rect 17861 18672 17866 18728
rect 17922 18672 18326 18728
rect 18382 18672 18387 18728
rect 17861 18670 18387 18672
rect 17861 18667 17927 18670
rect 18321 18667 18387 18670
rect 10869 18594 10935 18597
rect 11697 18594 11763 18597
rect 10869 18592 11763 18594
rect 10869 18536 10874 18592
rect 10930 18536 11702 18592
rect 11758 18536 11763 18592
rect 10869 18534 11763 18536
rect 23614 18594 23674 18806
rect 23800 18776 24600 18806
rect 23749 18594 23815 18597
rect 23614 18592 23815 18594
rect 23614 18536 23754 18592
rect 23810 18536 23815 18592
rect 23614 18534 23815 18536
rect 10869 18531 10935 18534
rect 11697 18531 11763 18534
rect 23749 18531 23815 18534
rect 6542 18528 6862 18529
rect 6542 18464 6550 18528
rect 6614 18464 6630 18528
rect 6694 18464 6710 18528
rect 6774 18464 6790 18528
rect 6854 18464 6862 18528
rect 6542 18463 6862 18464
rect 12140 18528 12460 18529
rect 12140 18464 12148 18528
rect 12212 18464 12228 18528
rect 12292 18464 12308 18528
rect 12372 18464 12388 18528
rect 12452 18464 12460 18528
rect 12140 18463 12460 18464
rect 17738 18528 18058 18529
rect 17738 18464 17746 18528
rect 17810 18464 17826 18528
rect 17890 18464 17906 18528
rect 17970 18464 17986 18528
rect 18050 18464 18058 18528
rect 17738 18463 18058 18464
rect 11145 18458 11211 18461
rect 11973 18458 12039 18461
rect 11145 18456 12039 18458
rect 11145 18400 11150 18456
rect 11206 18400 11978 18456
rect 12034 18400 12039 18456
rect 11145 18398 12039 18400
rect 11145 18395 11211 18398
rect 11973 18395 12039 18398
rect 14365 18458 14431 18461
rect 17125 18458 17191 18461
rect 14365 18456 17191 18458
rect 14365 18400 14370 18456
rect 14426 18400 17130 18456
rect 17186 18400 17191 18456
rect 14365 18398 17191 18400
rect 14365 18395 14431 18398
rect 17125 18395 17191 18398
rect 8201 18322 8267 18325
rect 21449 18322 21515 18325
rect 23800 18322 24600 18352
rect 8201 18320 21515 18322
rect 8201 18264 8206 18320
rect 8262 18264 21454 18320
rect 21510 18264 21515 18320
rect 8201 18262 21515 18264
rect 8201 18259 8267 18262
rect 21449 18259 21515 18262
rect 22050 18262 24600 18322
rect 3693 18186 3759 18189
rect 3558 18184 3759 18186
rect 3558 18128 3698 18184
rect 3754 18128 3759 18184
rect 3558 18126 3759 18128
rect 3558 17778 3618 18126
rect 3693 18123 3759 18126
rect 7097 18186 7163 18189
rect 7465 18186 7531 18189
rect 7097 18184 7531 18186
rect 7097 18128 7102 18184
rect 7158 18128 7470 18184
rect 7526 18128 7531 18184
rect 7097 18126 7531 18128
rect 7097 18123 7163 18126
rect 7465 18123 7531 18126
rect 9765 18186 9831 18189
rect 11697 18186 11763 18189
rect 9765 18184 11763 18186
rect 9765 18128 9770 18184
rect 9826 18128 11702 18184
rect 11758 18128 11763 18184
rect 9765 18126 11763 18128
rect 9765 18123 9831 18126
rect 11697 18123 11763 18126
rect 17585 18186 17651 18189
rect 22050 18186 22110 18262
rect 23800 18232 24600 18262
rect 17585 18184 22110 18186
rect 17585 18128 17590 18184
rect 17646 18128 22110 18184
rect 17585 18126 22110 18128
rect 17585 18123 17651 18126
rect 3743 17984 4063 17985
rect 3743 17920 3751 17984
rect 3815 17920 3831 17984
rect 3895 17920 3911 17984
rect 3975 17920 3991 17984
rect 4055 17920 4063 17984
rect 3743 17919 4063 17920
rect 9341 17984 9661 17985
rect 9341 17920 9349 17984
rect 9413 17920 9429 17984
rect 9493 17920 9509 17984
rect 9573 17920 9589 17984
rect 9653 17920 9661 17984
rect 9341 17919 9661 17920
rect 14939 17984 15259 17985
rect 14939 17920 14947 17984
rect 15011 17920 15027 17984
rect 15091 17920 15107 17984
rect 15171 17920 15187 17984
rect 15251 17920 15259 17984
rect 14939 17919 15259 17920
rect 20537 17984 20857 17985
rect 20537 17920 20545 17984
rect 20609 17920 20625 17984
rect 20689 17920 20705 17984
rect 20769 17920 20785 17984
rect 20849 17920 20857 17984
rect 20537 17919 20857 17920
rect 8017 17914 8083 17917
rect 8845 17914 8911 17917
rect 8017 17912 8911 17914
rect 8017 17856 8022 17912
rect 8078 17856 8850 17912
rect 8906 17856 8911 17912
rect 8017 17854 8911 17856
rect 8017 17851 8083 17854
rect 8845 17851 8911 17854
rect 21030 17852 21036 17916
rect 21100 17914 21106 17916
rect 22553 17914 22619 17917
rect 21100 17912 22619 17914
rect 21100 17856 22558 17912
rect 22614 17856 22619 17912
rect 21100 17854 22619 17856
rect 21100 17852 21106 17854
rect 22553 17851 22619 17854
rect 3877 17778 3943 17781
rect 3558 17776 3943 17778
rect 3558 17720 3882 17776
rect 3938 17720 3943 17776
rect 3558 17718 3943 17720
rect 3877 17715 3943 17718
rect 6545 17778 6611 17781
rect 8661 17778 8727 17781
rect 6545 17776 8727 17778
rect 6545 17720 6550 17776
rect 6606 17720 8666 17776
rect 8722 17720 8727 17776
rect 6545 17718 8727 17720
rect 6545 17715 6611 17718
rect 8661 17715 8727 17718
rect 13629 17778 13695 17781
rect 21541 17778 21607 17781
rect 13629 17776 21607 17778
rect 13629 17720 13634 17776
rect 13690 17720 21546 17776
rect 21602 17720 21607 17776
rect 13629 17718 21607 17720
rect 13629 17715 13695 17718
rect 21541 17715 21607 17718
rect 7557 17642 7623 17645
rect 8661 17642 8727 17645
rect 7557 17640 8727 17642
rect 7557 17584 7562 17640
rect 7618 17584 8666 17640
rect 8722 17584 8727 17640
rect 7557 17582 8727 17584
rect 7557 17579 7623 17582
rect 8661 17579 8727 17582
rect 16021 17642 16087 17645
rect 19333 17642 19399 17645
rect 23800 17642 24600 17672
rect 16021 17640 18338 17642
rect 16021 17584 16026 17640
rect 16082 17584 18338 17640
rect 16021 17582 18338 17584
rect 16021 17579 16087 17582
rect 6542 17440 6862 17441
rect 6542 17376 6550 17440
rect 6614 17376 6630 17440
rect 6694 17376 6710 17440
rect 6774 17376 6790 17440
rect 6854 17376 6862 17440
rect 6542 17375 6862 17376
rect 12140 17440 12460 17441
rect 12140 17376 12148 17440
rect 12212 17376 12228 17440
rect 12292 17376 12308 17440
rect 12372 17376 12388 17440
rect 12452 17376 12460 17440
rect 12140 17375 12460 17376
rect 17738 17440 18058 17441
rect 17738 17376 17746 17440
rect 17810 17376 17826 17440
rect 17890 17376 17906 17440
rect 17970 17376 17986 17440
rect 18050 17376 18058 17440
rect 17738 17375 18058 17376
rect 18278 17370 18338 17582
rect 19333 17640 24600 17642
rect 19333 17584 19338 17640
rect 19394 17584 24600 17640
rect 19333 17582 24600 17584
rect 19333 17579 19399 17582
rect 23800 17552 24600 17582
rect 20294 17444 20300 17508
rect 20364 17506 20370 17508
rect 22185 17506 22251 17509
rect 20364 17504 22251 17506
rect 20364 17448 22190 17504
rect 22246 17448 22251 17504
rect 20364 17446 22251 17448
rect 20364 17444 20370 17446
rect 22185 17443 22251 17446
rect 22829 17370 22895 17373
rect 18278 17368 22895 17370
rect 18278 17312 22834 17368
rect 22890 17312 22895 17368
rect 18278 17310 22895 17312
rect 22829 17307 22895 17310
rect 11237 17234 11303 17237
rect 22829 17234 22895 17237
rect 11237 17232 22895 17234
rect 11237 17176 11242 17232
rect 11298 17176 22834 17232
rect 22890 17176 22895 17232
rect 11237 17174 22895 17176
rect 11237 17171 11303 17174
rect 22829 17171 22895 17174
rect 9121 17100 9187 17101
rect 9070 17098 9076 17100
rect 9030 17038 9076 17098
rect 9140 17096 9187 17100
rect 9182 17040 9187 17096
rect 9070 17036 9076 17038
rect 9140 17036 9187 17040
rect 9121 17035 9187 17036
rect 23800 16962 24600 16992
rect 23614 16902 24600 16962
rect 3743 16896 4063 16897
rect 3743 16832 3751 16896
rect 3815 16832 3831 16896
rect 3895 16832 3911 16896
rect 3975 16832 3991 16896
rect 4055 16832 4063 16896
rect 3743 16831 4063 16832
rect 9341 16896 9661 16897
rect 9341 16832 9349 16896
rect 9413 16832 9429 16896
rect 9493 16832 9509 16896
rect 9573 16832 9589 16896
rect 9653 16832 9661 16896
rect 9341 16831 9661 16832
rect 14939 16896 15259 16897
rect 14939 16832 14947 16896
rect 15011 16832 15027 16896
rect 15091 16832 15107 16896
rect 15171 16832 15187 16896
rect 15251 16832 15259 16896
rect 14939 16831 15259 16832
rect 20537 16896 20857 16897
rect 20537 16832 20545 16896
rect 20609 16832 20625 16896
rect 20689 16832 20705 16896
rect 20769 16832 20785 16896
rect 20849 16832 20857 16896
rect 20537 16831 20857 16832
rect 23614 16690 23674 16902
rect 23800 16872 24600 16902
rect 23614 16630 24042 16690
rect 23982 16557 24042 16630
rect 23933 16552 24042 16557
rect 23933 16496 23938 16552
rect 23994 16496 24042 16552
rect 23933 16494 24042 16496
rect 23933 16491 23999 16494
rect 6542 16352 6862 16353
rect 6542 16288 6550 16352
rect 6614 16288 6630 16352
rect 6694 16288 6710 16352
rect 6774 16288 6790 16352
rect 6854 16288 6862 16352
rect 6542 16287 6862 16288
rect 12140 16352 12460 16353
rect 12140 16288 12148 16352
rect 12212 16288 12228 16352
rect 12292 16288 12308 16352
rect 12372 16288 12388 16352
rect 12452 16288 12460 16352
rect 12140 16287 12460 16288
rect 17738 16352 18058 16353
rect 17738 16288 17746 16352
rect 17810 16288 17826 16352
rect 17890 16288 17906 16352
rect 17970 16288 17986 16352
rect 18050 16288 18058 16352
rect 17738 16287 18058 16288
rect 22829 16282 22895 16285
rect 23013 16282 23079 16285
rect 23800 16282 24600 16312
rect 22829 16280 24600 16282
rect 22829 16224 22834 16280
rect 22890 16224 23018 16280
rect 23074 16224 24600 16280
rect 22829 16222 24600 16224
rect 22829 16219 22895 16222
rect 23013 16219 23079 16222
rect 23800 16192 24600 16222
rect 17033 16146 17099 16149
rect 22921 16146 22987 16149
rect 17033 16144 22987 16146
rect 17033 16088 17038 16144
rect 17094 16088 22926 16144
rect 22982 16088 22987 16144
rect 17033 16086 22987 16088
rect 17033 16083 17099 16086
rect 22921 16083 22987 16086
rect 13629 16010 13695 16013
rect 20989 16010 21055 16013
rect 13629 16008 21055 16010
rect 13629 15952 13634 16008
rect 13690 15952 20994 16008
rect 21050 15952 21055 16008
rect 13629 15950 21055 15952
rect 13629 15947 13695 15950
rect 20989 15947 21055 15950
rect 3743 15808 4063 15809
rect 3743 15744 3751 15808
rect 3815 15744 3831 15808
rect 3895 15744 3911 15808
rect 3975 15744 3991 15808
rect 4055 15744 4063 15808
rect 3743 15743 4063 15744
rect 9341 15808 9661 15809
rect 9341 15744 9349 15808
rect 9413 15744 9429 15808
rect 9493 15744 9509 15808
rect 9573 15744 9589 15808
rect 9653 15744 9661 15808
rect 9341 15743 9661 15744
rect 14939 15808 15259 15809
rect 14939 15744 14947 15808
rect 15011 15744 15027 15808
rect 15091 15744 15107 15808
rect 15171 15744 15187 15808
rect 15251 15744 15259 15808
rect 14939 15743 15259 15744
rect 20537 15808 20857 15809
rect 20537 15744 20545 15808
rect 20609 15744 20625 15808
rect 20689 15744 20705 15808
rect 20769 15744 20785 15808
rect 20849 15744 20857 15808
rect 20537 15743 20857 15744
rect 23381 15602 23447 15605
rect 23800 15602 24600 15632
rect 23381 15600 24600 15602
rect 23381 15544 23386 15600
rect 23442 15544 24600 15600
rect 23381 15542 24600 15544
rect 23381 15539 23447 15542
rect 23800 15512 24600 15542
rect 0 15330 800 15360
rect 1577 15330 1643 15333
rect 0 15328 1643 15330
rect 0 15272 1582 15328
rect 1638 15272 1643 15328
rect 0 15270 1643 15272
rect 0 15240 800 15270
rect 1577 15267 1643 15270
rect 6542 15264 6862 15265
rect 6542 15200 6550 15264
rect 6614 15200 6630 15264
rect 6694 15200 6710 15264
rect 6774 15200 6790 15264
rect 6854 15200 6862 15264
rect 6542 15199 6862 15200
rect 12140 15264 12460 15265
rect 12140 15200 12148 15264
rect 12212 15200 12228 15264
rect 12292 15200 12308 15264
rect 12372 15200 12388 15264
rect 12452 15200 12460 15264
rect 12140 15199 12460 15200
rect 17738 15264 18058 15265
rect 17738 15200 17746 15264
rect 17810 15200 17826 15264
rect 17890 15200 17906 15264
rect 17970 15200 17986 15264
rect 18050 15200 18058 15264
rect 17738 15199 18058 15200
rect 15561 14922 15627 14925
rect 15929 14922 15995 14925
rect 21214 14922 21220 14924
rect 15561 14920 21220 14922
rect 15561 14864 15566 14920
rect 15622 14864 15934 14920
rect 15990 14864 21220 14920
rect 15561 14862 21220 14864
rect 15561 14859 15627 14862
rect 15929 14859 15995 14862
rect 21214 14860 21220 14862
rect 21284 14860 21290 14924
rect 23197 14922 23263 14925
rect 23800 14922 24600 14952
rect 23197 14920 24600 14922
rect 23197 14864 23202 14920
rect 23258 14864 24600 14920
rect 23197 14862 24600 14864
rect 23197 14859 23263 14862
rect 23800 14832 24600 14862
rect 3743 14720 4063 14721
rect 3743 14656 3751 14720
rect 3815 14656 3831 14720
rect 3895 14656 3911 14720
rect 3975 14656 3991 14720
rect 4055 14656 4063 14720
rect 3743 14655 4063 14656
rect 9341 14720 9661 14721
rect 9341 14656 9349 14720
rect 9413 14656 9429 14720
rect 9493 14656 9509 14720
rect 9573 14656 9589 14720
rect 9653 14656 9661 14720
rect 9341 14655 9661 14656
rect 14939 14720 15259 14721
rect 14939 14656 14947 14720
rect 15011 14656 15027 14720
rect 15091 14656 15107 14720
rect 15171 14656 15187 14720
rect 15251 14656 15259 14720
rect 14939 14655 15259 14656
rect 20537 14720 20857 14721
rect 20537 14656 20545 14720
rect 20609 14656 20625 14720
rect 20689 14656 20705 14720
rect 20769 14656 20785 14720
rect 20849 14656 20857 14720
rect 20537 14655 20857 14656
rect 23105 14242 23171 14245
rect 23800 14242 24600 14272
rect 23105 14240 24600 14242
rect 23105 14184 23110 14240
rect 23166 14184 24600 14240
rect 23105 14182 24600 14184
rect 23105 14179 23171 14182
rect 6542 14176 6862 14177
rect 6542 14112 6550 14176
rect 6614 14112 6630 14176
rect 6694 14112 6710 14176
rect 6774 14112 6790 14176
rect 6854 14112 6862 14176
rect 6542 14111 6862 14112
rect 12140 14176 12460 14177
rect 12140 14112 12148 14176
rect 12212 14112 12228 14176
rect 12292 14112 12308 14176
rect 12372 14112 12388 14176
rect 12452 14112 12460 14176
rect 12140 14111 12460 14112
rect 17738 14176 18058 14177
rect 17738 14112 17746 14176
rect 17810 14112 17826 14176
rect 17890 14112 17906 14176
rect 17970 14112 17986 14176
rect 18050 14112 18058 14176
rect 23800 14152 24600 14182
rect 17738 14111 18058 14112
rect 16481 13970 16547 13973
rect 22921 13970 22987 13973
rect 16481 13968 22987 13970
rect 16481 13912 16486 13968
rect 16542 13912 22926 13968
rect 22982 13912 22987 13968
rect 16481 13910 22987 13912
rect 16481 13907 16547 13910
rect 22921 13907 22987 13910
rect 13997 13834 14063 13837
rect 20437 13834 20503 13837
rect 13997 13832 20503 13834
rect 13997 13776 14002 13832
rect 14058 13776 20442 13832
rect 20498 13776 20503 13832
rect 13997 13774 20503 13776
rect 13997 13771 14063 13774
rect 20437 13771 20503 13774
rect 3743 13632 4063 13633
rect 3743 13568 3751 13632
rect 3815 13568 3831 13632
rect 3895 13568 3911 13632
rect 3975 13568 3991 13632
rect 4055 13568 4063 13632
rect 3743 13567 4063 13568
rect 9341 13632 9661 13633
rect 9341 13568 9349 13632
rect 9413 13568 9429 13632
rect 9493 13568 9509 13632
rect 9573 13568 9589 13632
rect 9653 13568 9661 13632
rect 9341 13567 9661 13568
rect 14939 13632 15259 13633
rect 14939 13568 14947 13632
rect 15011 13568 15027 13632
rect 15091 13568 15107 13632
rect 15171 13568 15187 13632
rect 15251 13568 15259 13632
rect 14939 13567 15259 13568
rect 20537 13632 20857 13633
rect 20537 13568 20545 13632
rect 20609 13568 20625 13632
rect 20689 13568 20705 13632
rect 20769 13568 20785 13632
rect 20849 13568 20857 13632
rect 20537 13567 20857 13568
rect 18781 13562 18847 13565
rect 20294 13562 20300 13564
rect 18781 13560 20300 13562
rect 18781 13504 18786 13560
rect 18842 13504 20300 13560
rect 18781 13502 20300 13504
rect 18781 13499 18847 13502
rect 20294 13500 20300 13502
rect 20364 13500 20370 13564
rect 22553 13562 22619 13565
rect 23800 13562 24600 13592
rect 22553 13560 24600 13562
rect 22553 13504 22558 13560
rect 22614 13504 24600 13560
rect 22553 13502 24600 13504
rect 22553 13499 22619 13502
rect 23800 13472 24600 13502
rect 19057 13426 19123 13429
rect 19374 13426 19380 13428
rect 19057 13424 19380 13426
rect 19057 13368 19062 13424
rect 19118 13368 19380 13424
rect 19057 13366 19380 13368
rect 19057 13363 19123 13366
rect 19374 13364 19380 13366
rect 19444 13364 19450 13428
rect 20437 13426 20503 13429
rect 21030 13426 21036 13428
rect 20437 13424 21036 13426
rect 20437 13368 20442 13424
rect 20498 13368 21036 13424
rect 20437 13366 21036 13368
rect 20437 13363 20503 13366
rect 21030 13364 21036 13366
rect 21100 13364 21106 13428
rect 19609 13290 19675 13293
rect 23105 13290 23171 13293
rect 19609 13288 23306 13290
rect 19609 13232 19614 13288
rect 19670 13232 23110 13288
rect 23166 13232 23306 13288
rect 19609 13230 23306 13232
rect 19609 13227 19675 13230
rect 23105 13227 23171 13230
rect 6542 13088 6862 13089
rect 6542 13024 6550 13088
rect 6614 13024 6630 13088
rect 6694 13024 6710 13088
rect 6774 13024 6790 13088
rect 6854 13024 6862 13088
rect 6542 13023 6862 13024
rect 12140 13088 12460 13089
rect 12140 13024 12148 13088
rect 12212 13024 12228 13088
rect 12292 13024 12308 13088
rect 12372 13024 12388 13088
rect 12452 13024 12460 13088
rect 12140 13023 12460 13024
rect 17738 13088 18058 13089
rect 17738 13024 17746 13088
rect 17810 13024 17826 13088
rect 17890 13024 17906 13088
rect 17970 13024 17986 13088
rect 18050 13024 18058 13088
rect 17738 13023 18058 13024
rect 11789 12882 11855 12885
rect 16798 12882 16804 12884
rect 11789 12880 16804 12882
rect 11789 12824 11794 12880
rect 11850 12824 16804 12880
rect 11789 12822 16804 12824
rect 11789 12819 11855 12822
rect 16798 12820 16804 12822
rect 16868 12882 16874 12884
rect 20989 12882 21055 12885
rect 21449 12882 21515 12885
rect 16868 12880 21515 12882
rect 16868 12824 20994 12880
rect 21050 12824 21454 12880
rect 21510 12824 21515 12880
rect 16868 12822 21515 12824
rect 23246 12882 23306 13230
rect 23800 12882 24600 12912
rect 23246 12822 24600 12882
rect 16868 12820 16874 12822
rect 20989 12819 21055 12822
rect 21449 12819 21515 12822
rect 23800 12792 24600 12822
rect 3743 12544 4063 12545
rect 3743 12480 3751 12544
rect 3815 12480 3831 12544
rect 3895 12480 3911 12544
rect 3975 12480 3991 12544
rect 4055 12480 4063 12544
rect 3743 12479 4063 12480
rect 9341 12544 9661 12545
rect 9341 12480 9349 12544
rect 9413 12480 9429 12544
rect 9493 12480 9509 12544
rect 9573 12480 9589 12544
rect 9653 12480 9661 12544
rect 9341 12479 9661 12480
rect 14939 12544 15259 12545
rect 14939 12480 14947 12544
rect 15011 12480 15027 12544
rect 15091 12480 15107 12544
rect 15171 12480 15187 12544
rect 15251 12480 15259 12544
rect 14939 12479 15259 12480
rect 20537 12544 20857 12545
rect 20537 12480 20545 12544
rect 20609 12480 20625 12544
rect 20689 12480 20705 12544
rect 20769 12480 20785 12544
rect 20849 12480 20857 12544
rect 20537 12479 20857 12480
rect 15745 12338 15811 12341
rect 18597 12338 18663 12341
rect 15745 12336 18663 12338
rect 15745 12280 15750 12336
rect 15806 12280 18602 12336
rect 18658 12280 18663 12336
rect 15745 12278 18663 12280
rect 15745 12275 15811 12278
rect 18597 12275 18663 12278
rect 22829 12338 22895 12341
rect 23800 12338 24600 12368
rect 22829 12336 24600 12338
rect 22829 12280 22834 12336
rect 22890 12280 24600 12336
rect 22829 12278 24600 12280
rect 22829 12275 22895 12278
rect 23800 12248 24600 12278
rect 17861 12202 17927 12205
rect 18597 12202 18663 12205
rect 17861 12200 18663 12202
rect 17861 12144 17866 12200
rect 17922 12144 18602 12200
rect 18658 12144 18663 12200
rect 17861 12142 18663 12144
rect 17861 12139 17927 12142
rect 18597 12139 18663 12142
rect 19057 12202 19123 12205
rect 23013 12202 23079 12205
rect 19057 12200 23079 12202
rect 19057 12144 19062 12200
rect 19118 12144 23018 12200
rect 23074 12144 23079 12200
rect 19057 12142 23079 12144
rect 19057 12139 19123 12142
rect 23013 12139 23079 12142
rect 6542 12000 6862 12001
rect 6542 11936 6550 12000
rect 6614 11936 6630 12000
rect 6694 11936 6710 12000
rect 6774 11936 6790 12000
rect 6854 11936 6862 12000
rect 6542 11935 6862 11936
rect 12140 12000 12460 12001
rect 12140 11936 12148 12000
rect 12212 11936 12228 12000
rect 12292 11936 12308 12000
rect 12372 11936 12388 12000
rect 12452 11936 12460 12000
rect 12140 11935 12460 11936
rect 17738 12000 18058 12001
rect 17738 11936 17746 12000
rect 17810 11936 17826 12000
rect 17890 11936 17906 12000
rect 17970 11936 17986 12000
rect 18050 11936 18058 12000
rect 17738 11935 18058 11936
rect 23105 11658 23171 11661
rect 23800 11658 24600 11688
rect 23105 11656 24600 11658
rect 23105 11600 23110 11656
rect 23166 11600 24600 11656
rect 23105 11598 24600 11600
rect 23105 11595 23171 11598
rect 23800 11568 24600 11598
rect 3743 11456 4063 11457
rect 3743 11392 3751 11456
rect 3815 11392 3831 11456
rect 3895 11392 3911 11456
rect 3975 11392 3991 11456
rect 4055 11392 4063 11456
rect 3743 11391 4063 11392
rect 9341 11456 9661 11457
rect 9341 11392 9349 11456
rect 9413 11392 9429 11456
rect 9493 11392 9509 11456
rect 9573 11392 9589 11456
rect 9653 11392 9661 11456
rect 9341 11391 9661 11392
rect 14939 11456 15259 11457
rect 14939 11392 14947 11456
rect 15011 11392 15027 11456
rect 15091 11392 15107 11456
rect 15171 11392 15187 11456
rect 15251 11392 15259 11456
rect 14939 11391 15259 11392
rect 20537 11456 20857 11457
rect 20537 11392 20545 11456
rect 20609 11392 20625 11456
rect 20689 11392 20705 11456
rect 20769 11392 20785 11456
rect 20849 11392 20857 11456
rect 20537 11391 20857 11392
rect 13629 11250 13695 11253
rect 16614 11250 16620 11252
rect 13629 11248 16620 11250
rect 13629 11192 13634 11248
rect 13690 11192 16620 11248
rect 13629 11190 16620 11192
rect 13629 11187 13695 11190
rect 16614 11188 16620 11190
rect 16684 11188 16690 11252
rect 20069 11250 20135 11253
rect 20897 11250 20963 11253
rect 20069 11248 20963 11250
rect 20069 11192 20074 11248
rect 20130 11192 20902 11248
rect 20958 11192 20963 11248
rect 20069 11190 20963 11192
rect 20069 11187 20135 11190
rect 20897 11187 20963 11190
rect 23105 10978 23171 10981
rect 23800 10978 24600 11008
rect 23105 10976 24600 10978
rect 23105 10920 23110 10976
rect 23166 10920 24600 10976
rect 23105 10918 24600 10920
rect 23105 10915 23171 10918
rect 6542 10912 6862 10913
rect 6542 10848 6550 10912
rect 6614 10848 6630 10912
rect 6694 10848 6710 10912
rect 6774 10848 6790 10912
rect 6854 10848 6862 10912
rect 6542 10847 6862 10848
rect 12140 10912 12460 10913
rect 12140 10848 12148 10912
rect 12212 10848 12228 10912
rect 12292 10848 12308 10912
rect 12372 10848 12388 10912
rect 12452 10848 12460 10912
rect 12140 10847 12460 10848
rect 17738 10912 18058 10913
rect 17738 10848 17746 10912
rect 17810 10848 17826 10912
rect 17890 10848 17906 10912
rect 17970 10848 17986 10912
rect 18050 10848 18058 10912
rect 23800 10888 24600 10918
rect 17738 10847 18058 10848
rect 11789 10570 11855 10573
rect 21909 10570 21975 10573
rect 11789 10568 21975 10570
rect 11789 10512 11794 10568
rect 11850 10512 21914 10568
rect 21970 10512 21975 10568
rect 11789 10510 21975 10512
rect 11789 10507 11855 10510
rect 21909 10507 21975 10510
rect 3743 10368 4063 10369
rect 3743 10304 3751 10368
rect 3815 10304 3831 10368
rect 3895 10304 3911 10368
rect 3975 10304 3991 10368
rect 4055 10304 4063 10368
rect 3743 10303 4063 10304
rect 9341 10368 9661 10369
rect 9341 10304 9349 10368
rect 9413 10304 9429 10368
rect 9493 10304 9509 10368
rect 9573 10304 9589 10368
rect 9653 10304 9661 10368
rect 9341 10303 9661 10304
rect 14939 10368 15259 10369
rect 14939 10304 14947 10368
rect 15011 10304 15027 10368
rect 15091 10304 15107 10368
rect 15171 10304 15187 10368
rect 15251 10304 15259 10368
rect 14939 10303 15259 10304
rect 20537 10368 20857 10369
rect 20537 10304 20545 10368
rect 20609 10304 20625 10368
rect 20689 10304 20705 10368
rect 20769 10304 20785 10368
rect 20849 10304 20857 10368
rect 20537 10303 20857 10304
rect 23013 10298 23079 10301
rect 23800 10298 24600 10328
rect 23013 10296 24600 10298
rect 23013 10240 23018 10296
rect 23074 10240 24600 10296
rect 23013 10238 24600 10240
rect 23013 10235 23079 10238
rect 23800 10208 24600 10238
rect 18137 10162 18203 10165
rect 21909 10162 21975 10165
rect 18137 10160 21975 10162
rect 18137 10104 18142 10160
rect 18198 10104 21914 10160
rect 21970 10104 21975 10160
rect 18137 10102 21975 10104
rect 18137 10099 18203 10102
rect 21909 10099 21975 10102
rect 6542 9824 6862 9825
rect 6542 9760 6550 9824
rect 6614 9760 6630 9824
rect 6694 9760 6710 9824
rect 6774 9760 6790 9824
rect 6854 9760 6862 9824
rect 6542 9759 6862 9760
rect 12140 9824 12460 9825
rect 12140 9760 12148 9824
rect 12212 9760 12228 9824
rect 12292 9760 12308 9824
rect 12372 9760 12388 9824
rect 12452 9760 12460 9824
rect 12140 9759 12460 9760
rect 17738 9824 18058 9825
rect 17738 9760 17746 9824
rect 17810 9760 17826 9824
rect 17890 9760 17906 9824
rect 17970 9760 17986 9824
rect 18050 9760 18058 9824
rect 17738 9759 18058 9760
rect 13537 9754 13603 9757
rect 14457 9754 14523 9757
rect 13537 9752 14523 9754
rect 13537 9696 13542 9752
rect 13598 9696 14462 9752
rect 14518 9696 14523 9752
rect 13537 9694 14523 9696
rect 13537 9691 13603 9694
rect 14457 9691 14523 9694
rect 23289 9618 23355 9621
rect 23800 9618 24600 9648
rect 23289 9616 24600 9618
rect 23289 9560 23294 9616
rect 23350 9560 24600 9616
rect 23289 9558 24600 9560
rect 23289 9555 23355 9558
rect 23800 9528 24600 9558
rect 12893 9482 12959 9485
rect 16798 9482 16804 9484
rect 12893 9480 16804 9482
rect 12893 9424 12898 9480
rect 12954 9424 16804 9480
rect 12893 9422 16804 9424
rect 12893 9419 12959 9422
rect 16798 9420 16804 9422
rect 16868 9420 16874 9484
rect 3743 9280 4063 9281
rect 0 9210 800 9240
rect 3743 9216 3751 9280
rect 3815 9216 3831 9280
rect 3895 9216 3911 9280
rect 3975 9216 3991 9280
rect 4055 9216 4063 9280
rect 3743 9215 4063 9216
rect 9341 9280 9661 9281
rect 9341 9216 9349 9280
rect 9413 9216 9429 9280
rect 9493 9216 9509 9280
rect 9573 9216 9589 9280
rect 9653 9216 9661 9280
rect 9341 9215 9661 9216
rect 14939 9280 15259 9281
rect 14939 9216 14947 9280
rect 15011 9216 15027 9280
rect 15091 9216 15107 9280
rect 15171 9216 15187 9280
rect 15251 9216 15259 9280
rect 14939 9215 15259 9216
rect 20537 9280 20857 9281
rect 20537 9216 20545 9280
rect 20609 9216 20625 9280
rect 20689 9216 20705 9280
rect 20769 9216 20785 9280
rect 20849 9216 20857 9280
rect 20537 9215 20857 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 11881 8938 11947 8941
rect 22921 8938 22987 8941
rect 11881 8936 22987 8938
rect 11881 8880 11886 8936
rect 11942 8880 22926 8936
rect 22982 8880 22987 8936
rect 11881 8878 22987 8880
rect 11881 8875 11947 8878
rect 22921 8875 22987 8878
rect 23381 8938 23447 8941
rect 23800 8938 24600 8968
rect 23381 8936 24600 8938
rect 23381 8880 23386 8936
rect 23442 8880 24600 8936
rect 23381 8878 24600 8880
rect 23381 8875 23447 8878
rect 23800 8848 24600 8878
rect 6542 8736 6862 8737
rect 6542 8672 6550 8736
rect 6614 8672 6630 8736
rect 6694 8672 6710 8736
rect 6774 8672 6790 8736
rect 6854 8672 6862 8736
rect 6542 8671 6862 8672
rect 12140 8736 12460 8737
rect 12140 8672 12148 8736
rect 12212 8672 12228 8736
rect 12292 8672 12308 8736
rect 12372 8672 12388 8736
rect 12452 8672 12460 8736
rect 12140 8671 12460 8672
rect 17738 8736 18058 8737
rect 17738 8672 17746 8736
rect 17810 8672 17826 8736
rect 17890 8672 17906 8736
rect 17970 8672 17986 8736
rect 18050 8672 18058 8736
rect 17738 8671 18058 8672
rect 19333 8666 19399 8669
rect 23289 8666 23355 8669
rect 19333 8664 23355 8666
rect 19333 8608 19338 8664
rect 19394 8608 23294 8664
rect 23350 8608 23355 8664
rect 19333 8606 23355 8608
rect 19333 8603 19399 8606
rect 23289 8603 23355 8606
rect 21357 8258 21423 8261
rect 23800 8258 24600 8288
rect 21357 8256 24600 8258
rect 21357 8200 21362 8256
rect 21418 8200 24600 8256
rect 21357 8198 24600 8200
rect 21357 8195 21423 8198
rect 3743 8192 4063 8193
rect 3743 8128 3751 8192
rect 3815 8128 3831 8192
rect 3895 8128 3911 8192
rect 3975 8128 3991 8192
rect 4055 8128 4063 8192
rect 3743 8127 4063 8128
rect 9341 8192 9661 8193
rect 9341 8128 9349 8192
rect 9413 8128 9429 8192
rect 9493 8128 9509 8192
rect 9573 8128 9589 8192
rect 9653 8128 9661 8192
rect 9341 8127 9661 8128
rect 14939 8192 15259 8193
rect 14939 8128 14947 8192
rect 15011 8128 15027 8192
rect 15091 8128 15107 8192
rect 15171 8128 15187 8192
rect 15251 8128 15259 8192
rect 14939 8127 15259 8128
rect 20537 8192 20857 8193
rect 20537 8128 20545 8192
rect 20609 8128 20625 8192
rect 20689 8128 20705 8192
rect 20769 8128 20785 8192
rect 20849 8128 20857 8192
rect 23800 8168 24600 8198
rect 20537 8127 20857 8128
rect 9029 7850 9095 7853
rect 18873 7850 18939 7853
rect 9029 7848 18939 7850
rect 9029 7792 9034 7848
rect 9090 7792 18878 7848
rect 18934 7792 18939 7848
rect 9029 7790 18939 7792
rect 9029 7787 9095 7790
rect 18873 7787 18939 7790
rect 6542 7648 6862 7649
rect 6542 7584 6550 7648
rect 6614 7584 6630 7648
rect 6694 7584 6710 7648
rect 6774 7584 6790 7648
rect 6854 7584 6862 7648
rect 6542 7583 6862 7584
rect 12140 7648 12460 7649
rect 12140 7584 12148 7648
rect 12212 7584 12228 7648
rect 12292 7584 12308 7648
rect 12372 7584 12388 7648
rect 12452 7584 12460 7648
rect 12140 7583 12460 7584
rect 17738 7648 18058 7649
rect 17738 7584 17746 7648
rect 17810 7584 17826 7648
rect 17890 7584 17906 7648
rect 17970 7584 17986 7648
rect 18050 7584 18058 7648
rect 17738 7583 18058 7584
rect 19333 7578 19399 7581
rect 23800 7578 24600 7608
rect 19333 7576 24600 7578
rect 19333 7520 19338 7576
rect 19394 7520 24600 7576
rect 19333 7518 24600 7520
rect 19333 7515 19399 7518
rect 23800 7488 24600 7518
rect 10593 7442 10659 7445
rect 22645 7442 22711 7445
rect 10593 7440 22711 7442
rect 10593 7384 10598 7440
rect 10654 7384 22650 7440
rect 22706 7384 22711 7440
rect 10593 7382 22711 7384
rect 10593 7379 10659 7382
rect 22645 7379 22711 7382
rect 4797 7306 4863 7309
rect 16205 7306 16271 7309
rect 21541 7306 21607 7309
rect 4797 7304 21607 7306
rect 4797 7248 4802 7304
rect 4858 7248 16210 7304
rect 16266 7248 21546 7304
rect 21602 7248 21607 7304
rect 4797 7246 21607 7248
rect 4797 7243 4863 7246
rect 16205 7243 16271 7246
rect 21541 7243 21607 7246
rect 3743 7104 4063 7105
rect 3743 7040 3751 7104
rect 3815 7040 3831 7104
rect 3895 7040 3911 7104
rect 3975 7040 3991 7104
rect 4055 7040 4063 7104
rect 3743 7039 4063 7040
rect 9341 7104 9661 7105
rect 9341 7040 9349 7104
rect 9413 7040 9429 7104
rect 9493 7040 9509 7104
rect 9573 7040 9589 7104
rect 9653 7040 9661 7104
rect 9341 7039 9661 7040
rect 14939 7104 15259 7105
rect 14939 7040 14947 7104
rect 15011 7040 15027 7104
rect 15091 7040 15107 7104
rect 15171 7040 15187 7104
rect 15251 7040 15259 7104
rect 14939 7039 15259 7040
rect 20537 7104 20857 7105
rect 20537 7040 20545 7104
rect 20609 7040 20625 7104
rect 20689 7040 20705 7104
rect 20769 7040 20785 7104
rect 20849 7040 20857 7104
rect 20537 7039 20857 7040
rect 4153 6898 4219 6901
rect 18781 6898 18847 6901
rect 4153 6896 18847 6898
rect 4153 6840 4158 6896
rect 4214 6840 18786 6896
rect 18842 6840 18847 6896
rect 4153 6838 18847 6840
rect 4153 6835 4219 6838
rect 18781 6835 18847 6838
rect 19333 6898 19399 6901
rect 23013 6898 23079 6901
rect 23800 6898 24600 6928
rect 19333 6896 24600 6898
rect 19333 6840 19338 6896
rect 19394 6840 23018 6896
rect 23074 6840 24600 6896
rect 19333 6838 24600 6840
rect 19333 6835 19399 6838
rect 23013 6835 23079 6838
rect 23800 6808 24600 6838
rect 10225 6762 10291 6765
rect 18137 6762 18203 6765
rect 21449 6762 21515 6765
rect 10225 6760 21515 6762
rect 10225 6704 10230 6760
rect 10286 6704 18142 6760
rect 18198 6704 21454 6760
rect 21510 6704 21515 6760
rect 10225 6702 21515 6704
rect 10225 6699 10291 6702
rect 18137 6699 18203 6702
rect 21449 6699 21515 6702
rect 6542 6560 6862 6561
rect 6542 6496 6550 6560
rect 6614 6496 6630 6560
rect 6694 6496 6710 6560
rect 6774 6496 6790 6560
rect 6854 6496 6862 6560
rect 6542 6495 6862 6496
rect 12140 6560 12460 6561
rect 12140 6496 12148 6560
rect 12212 6496 12228 6560
rect 12292 6496 12308 6560
rect 12372 6496 12388 6560
rect 12452 6496 12460 6560
rect 12140 6495 12460 6496
rect 17738 6560 18058 6561
rect 17738 6496 17746 6560
rect 17810 6496 17826 6560
rect 17890 6496 17906 6560
rect 17970 6496 17986 6560
rect 18050 6496 18058 6560
rect 17738 6495 18058 6496
rect 10961 6354 11027 6357
rect 18137 6354 18203 6357
rect 10961 6352 18203 6354
rect 10961 6296 10966 6352
rect 11022 6296 18142 6352
rect 18198 6296 18203 6352
rect 10961 6294 18203 6296
rect 10961 6291 11027 6294
rect 18137 6291 18203 6294
rect 23013 6354 23079 6357
rect 23800 6354 24600 6384
rect 23013 6352 24600 6354
rect 23013 6296 23018 6352
rect 23074 6296 24600 6352
rect 23013 6294 24600 6296
rect 23013 6291 23079 6294
rect 23800 6264 24600 6294
rect 2865 6218 2931 6221
rect 13629 6218 13695 6221
rect 2865 6216 13695 6218
rect 2865 6160 2870 6216
rect 2926 6160 13634 6216
rect 13690 6160 13695 6216
rect 2865 6158 13695 6160
rect 2865 6155 2931 6158
rect 13629 6155 13695 6158
rect 16297 6218 16363 6221
rect 22277 6218 22343 6221
rect 16297 6216 22343 6218
rect 16297 6160 16302 6216
rect 16358 6160 22282 6216
rect 22338 6160 22343 6216
rect 16297 6158 22343 6160
rect 16297 6155 16363 6158
rect 22277 6155 22343 6158
rect 3743 6016 4063 6017
rect 3743 5952 3751 6016
rect 3815 5952 3831 6016
rect 3895 5952 3911 6016
rect 3975 5952 3991 6016
rect 4055 5952 4063 6016
rect 3743 5951 4063 5952
rect 9341 6016 9661 6017
rect 9341 5952 9349 6016
rect 9413 5952 9429 6016
rect 9493 5952 9509 6016
rect 9573 5952 9589 6016
rect 9653 5952 9661 6016
rect 9341 5951 9661 5952
rect 14939 6016 15259 6017
rect 14939 5952 14947 6016
rect 15011 5952 15027 6016
rect 15091 5952 15107 6016
rect 15171 5952 15187 6016
rect 15251 5952 15259 6016
rect 14939 5951 15259 5952
rect 20537 6016 20857 6017
rect 20537 5952 20545 6016
rect 20609 5952 20625 6016
rect 20689 5952 20705 6016
rect 20769 5952 20785 6016
rect 20849 5952 20857 6016
rect 20537 5951 20857 5952
rect 16665 5948 16731 5949
rect 16614 5884 16620 5948
rect 16684 5946 16731 5948
rect 16684 5944 16776 5946
rect 16726 5888 16776 5944
rect 16684 5886 16776 5888
rect 16684 5884 16731 5886
rect 16665 5883 16731 5884
rect 13629 5810 13695 5813
rect 19885 5810 19951 5813
rect 22277 5810 22343 5813
rect 13629 5808 22343 5810
rect 13629 5752 13634 5808
rect 13690 5752 19890 5808
rect 19946 5752 22282 5808
rect 22338 5752 22343 5808
rect 13629 5750 22343 5752
rect 13629 5747 13695 5750
rect 19885 5747 19951 5750
rect 22277 5747 22343 5750
rect 2497 5674 2563 5677
rect 13721 5674 13787 5677
rect 22829 5674 22895 5677
rect 2497 5672 22895 5674
rect 2497 5616 2502 5672
rect 2558 5616 13726 5672
rect 13782 5616 22834 5672
rect 22890 5616 22895 5672
rect 2497 5614 22895 5616
rect 2497 5611 2563 5614
rect 13721 5611 13787 5614
rect 22829 5611 22895 5614
rect 23013 5674 23079 5677
rect 23800 5674 24600 5704
rect 23013 5672 24600 5674
rect 23013 5616 23018 5672
rect 23074 5616 24600 5672
rect 23013 5614 24600 5616
rect 23013 5611 23079 5614
rect 23800 5584 24600 5614
rect 6542 5472 6862 5473
rect 6542 5408 6550 5472
rect 6614 5408 6630 5472
rect 6694 5408 6710 5472
rect 6774 5408 6790 5472
rect 6854 5408 6862 5472
rect 6542 5407 6862 5408
rect 12140 5472 12460 5473
rect 12140 5408 12148 5472
rect 12212 5408 12228 5472
rect 12292 5408 12308 5472
rect 12372 5408 12388 5472
rect 12452 5408 12460 5472
rect 12140 5407 12460 5408
rect 17738 5472 18058 5473
rect 17738 5408 17746 5472
rect 17810 5408 17826 5472
rect 17890 5408 17906 5472
rect 17970 5408 17986 5472
rect 18050 5408 18058 5472
rect 17738 5407 18058 5408
rect 5441 5130 5507 5133
rect 16297 5130 16363 5133
rect 5441 5128 16363 5130
rect 5441 5072 5446 5128
rect 5502 5072 16302 5128
rect 16358 5072 16363 5128
rect 5441 5070 16363 5072
rect 5441 5067 5507 5070
rect 16297 5067 16363 5070
rect 19609 5130 19675 5133
rect 21541 5130 21607 5133
rect 19609 5128 21607 5130
rect 19609 5072 19614 5128
rect 19670 5072 21546 5128
rect 21602 5072 21607 5128
rect 19609 5070 21607 5072
rect 19609 5067 19675 5070
rect 21541 5067 21607 5070
rect 16113 4994 16179 4997
rect 18045 4994 18111 4997
rect 16113 4992 18111 4994
rect 16113 4936 16118 4992
rect 16174 4936 18050 4992
rect 18106 4936 18111 4992
rect 16113 4934 18111 4936
rect 16113 4931 16179 4934
rect 18045 4931 18111 4934
rect 21541 4994 21607 4997
rect 23800 4994 24600 5024
rect 21541 4992 24600 4994
rect 21541 4936 21546 4992
rect 21602 4936 24600 4992
rect 21541 4934 24600 4936
rect 21541 4931 21607 4934
rect 3743 4928 4063 4929
rect 3743 4864 3751 4928
rect 3815 4864 3831 4928
rect 3895 4864 3911 4928
rect 3975 4864 3991 4928
rect 4055 4864 4063 4928
rect 3743 4863 4063 4864
rect 9341 4928 9661 4929
rect 9341 4864 9349 4928
rect 9413 4864 9429 4928
rect 9493 4864 9509 4928
rect 9573 4864 9589 4928
rect 9653 4864 9661 4928
rect 9341 4863 9661 4864
rect 14939 4928 15259 4929
rect 14939 4864 14947 4928
rect 15011 4864 15027 4928
rect 15091 4864 15107 4928
rect 15171 4864 15187 4928
rect 15251 4864 15259 4928
rect 14939 4863 15259 4864
rect 20537 4928 20857 4929
rect 20537 4864 20545 4928
rect 20609 4864 20625 4928
rect 20689 4864 20705 4928
rect 20769 4864 20785 4928
rect 20849 4864 20857 4928
rect 23800 4904 24600 4934
rect 20537 4863 20857 4864
rect 15518 4798 18522 4858
rect 5349 4722 5415 4725
rect 13629 4722 13695 4725
rect 5349 4720 13695 4722
rect 5349 4664 5354 4720
rect 5410 4664 13634 4720
rect 13690 4664 13695 4720
rect 5349 4662 13695 4664
rect 5349 4659 5415 4662
rect 13629 4659 13695 4662
rect 15009 4722 15075 4725
rect 15518 4722 15578 4798
rect 15009 4720 15578 4722
rect 15009 4664 15014 4720
rect 15070 4664 15578 4720
rect 15009 4662 15578 4664
rect 15653 4722 15719 4725
rect 18462 4722 18522 4798
rect 20437 4722 20503 4725
rect 21265 4722 21331 4725
rect 15653 4720 18338 4722
rect 15653 4664 15658 4720
rect 15714 4664 18338 4720
rect 15653 4662 18338 4664
rect 18462 4720 21331 4722
rect 18462 4664 20442 4720
rect 20498 4664 21270 4720
rect 21326 4664 21331 4720
rect 18462 4662 21331 4664
rect 15009 4659 15075 4662
rect 15653 4659 15719 4662
rect 2957 4586 3023 4589
rect 18137 4586 18203 4589
rect 2957 4584 18203 4586
rect 2957 4528 2962 4584
rect 3018 4528 18142 4584
rect 18198 4528 18203 4584
rect 2957 4526 18203 4528
rect 18278 4586 18338 4662
rect 20437 4659 20503 4662
rect 21265 4659 21331 4662
rect 21449 4586 21515 4589
rect 18278 4584 21515 4586
rect 18278 4528 21454 4584
rect 21510 4528 21515 4584
rect 18278 4526 21515 4528
rect 2957 4523 3023 4526
rect 18137 4523 18203 4526
rect 21449 4523 21515 4526
rect 6542 4384 6862 4385
rect 6542 4320 6550 4384
rect 6614 4320 6630 4384
rect 6694 4320 6710 4384
rect 6774 4320 6790 4384
rect 6854 4320 6862 4384
rect 6542 4319 6862 4320
rect 12140 4384 12460 4385
rect 12140 4320 12148 4384
rect 12212 4320 12228 4384
rect 12292 4320 12308 4384
rect 12372 4320 12388 4384
rect 12452 4320 12460 4384
rect 12140 4319 12460 4320
rect 17738 4384 18058 4385
rect 17738 4320 17746 4384
rect 17810 4320 17826 4384
rect 17890 4320 17906 4384
rect 17970 4320 17986 4384
rect 18050 4320 18058 4384
rect 17738 4319 18058 4320
rect 19977 4314 20043 4317
rect 23800 4314 24600 4344
rect 19977 4312 24600 4314
rect 19977 4256 19982 4312
rect 20038 4256 24600 4312
rect 19977 4254 24600 4256
rect 19977 4251 20043 4254
rect 23800 4224 24600 4254
rect 2221 4178 2287 4181
rect 15561 4178 15627 4181
rect 2221 4176 15627 4178
rect 2221 4120 2226 4176
rect 2282 4120 15566 4176
rect 15622 4120 15627 4176
rect 2221 4118 15627 4120
rect 2221 4115 2287 4118
rect 15561 4115 15627 4118
rect 19057 4178 19123 4181
rect 21265 4178 21331 4181
rect 19057 4176 21331 4178
rect 19057 4120 19062 4176
rect 19118 4120 21270 4176
rect 21326 4120 21331 4176
rect 19057 4118 21331 4120
rect 19057 4115 19123 4118
rect 21265 4115 21331 4118
rect 3969 4042 4035 4045
rect 20345 4042 20411 4045
rect 3969 4040 20411 4042
rect 3969 3984 3974 4040
rect 4030 3984 20350 4040
rect 20406 3984 20411 4040
rect 3969 3982 20411 3984
rect 3969 3979 4035 3982
rect 20345 3979 20411 3982
rect 15561 3906 15627 3909
rect 19517 3906 19583 3909
rect 15561 3904 19583 3906
rect 15561 3848 15566 3904
rect 15622 3848 19522 3904
rect 19578 3848 19583 3904
rect 15561 3846 19583 3848
rect 15561 3843 15627 3846
rect 19517 3843 19583 3846
rect 3743 3840 4063 3841
rect 3743 3776 3751 3840
rect 3815 3776 3831 3840
rect 3895 3776 3911 3840
rect 3975 3776 3991 3840
rect 4055 3776 4063 3840
rect 3743 3775 4063 3776
rect 9341 3840 9661 3841
rect 9341 3776 9349 3840
rect 9413 3776 9429 3840
rect 9493 3776 9509 3840
rect 9573 3776 9589 3840
rect 9653 3776 9661 3840
rect 9341 3775 9661 3776
rect 14939 3840 15259 3841
rect 14939 3776 14947 3840
rect 15011 3776 15027 3840
rect 15091 3776 15107 3840
rect 15171 3776 15187 3840
rect 15251 3776 15259 3840
rect 14939 3775 15259 3776
rect 20537 3840 20857 3841
rect 20537 3776 20545 3840
rect 20609 3776 20625 3840
rect 20689 3776 20705 3840
rect 20769 3776 20785 3840
rect 20849 3776 20857 3840
rect 20537 3775 20857 3776
rect 14825 3634 14891 3637
rect 20529 3634 20595 3637
rect 14825 3632 20595 3634
rect 14825 3576 14830 3632
rect 14886 3576 20534 3632
rect 20590 3576 20595 3632
rect 14825 3574 20595 3576
rect 14825 3571 14891 3574
rect 20529 3571 20595 3574
rect 22737 3634 22803 3637
rect 23800 3634 24600 3664
rect 22737 3632 24600 3634
rect 22737 3576 22742 3632
rect 22798 3576 24600 3632
rect 22737 3574 24600 3576
rect 22737 3571 22803 3574
rect 23800 3544 24600 3574
rect 3233 3498 3299 3501
rect 14641 3498 14707 3501
rect 20713 3498 20779 3501
rect 3233 3496 14707 3498
rect 3233 3440 3238 3496
rect 3294 3440 14646 3496
rect 14702 3440 14707 3496
rect 3233 3438 14707 3440
rect 3233 3435 3299 3438
rect 14641 3435 14707 3438
rect 14782 3496 20779 3498
rect 14782 3440 20718 3496
rect 20774 3440 20779 3496
rect 14782 3438 20779 3440
rect 14549 3362 14615 3365
rect 14782 3362 14842 3438
rect 20713 3435 20779 3438
rect 14549 3360 14842 3362
rect 14549 3304 14554 3360
rect 14610 3304 14842 3360
rect 14549 3302 14842 3304
rect 14549 3299 14615 3302
rect 6542 3296 6862 3297
rect 6542 3232 6550 3296
rect 6614 3232 6630 3296
rect 6694 3232 6710 3296
rect 6774 3232 6790 3296
rect 6854 3232 6862 3296
rect 6542 3231 6862 3232
rect 12140 3296 12460 3297
rect 12140 3232 12148 3296
rect 12212 3232 12228 3296
rect 12292 3232 12308 3296
rect 12372 3232 12388 3296
rect 12452 3232 12460 3296
rect 12140 3231 12460 3232
rect 17738 3296 18058 3297
rect 17738 3232 17746 3296
rect 17810 3232 17826 3296
rect 17890 3232 17906 3296
rect 17970 3232 17986 3296
rect 18050 3232 18058 3296
rect 17738 3231 18058 3232
rect 20805 3226 20871 3229
rect 22645 3226 22711 3229
rect 20805 3224 22711 3226
rect 20805 3168 20810 3224
rect 20866 3168 22650 3224
rect 22706 3168 22711 3224
rect 20805 3166 22711 3168
rect 20805 3163 20871 3166
rect 22645 3163 22711 3166
rect 0 3090 800 3120
rect 1393 3090 1459 3093
rect 0 3088 1459 3090
rect 0 3032 1398 3088
rect 1454 3032 1459 3088
rect 0 3030 1459 3032
rect 0 3000 800 3030
rect 1393 3027 1459 3030
rect 13629 3090 13695 3093
rect 19241 3090 19307 3093
rect 21357 3090 21423 3093
rect 13629 3088 19307 3090
rect 13629 3032 13634 3088
rect 13690 3032 19246 3088
rect 19302 3032 19307 3088
rect 13629 3030 19307 3032
rect 13629 3027 13695 3030
rect 19241 3027 19307 3030
rect 19566 3088 21423 3090
rect 19566 3032 21362 3088
rect 21418 3032 21423 3088
rect 19566 3030 21423 3032
rect 1577 2954 1643 2957
rect 8109 2954 8175 2957
rect 1577 2952 8175 2954
rect 1577 2896 1582 2952
rect 1638 2896 8114 2952
rect 8170 2896 8175 2952
rect 1577 2894 8175 2896
rect 1577 2891 1643 2894
rect 8109 2891 8175 2894
rect 9121 2954 9187 2957
rect 13537 2954 13603 2957
rect 19566 2954 19626 3030
rect 21357 3027 21423 3030
rect 9121 2952 19626 2954
rect 9121 2896 9126 2952
rect 9182 2896 13542 2952
rect 13598 2896 19626 2952
rect 9121 2894 19626 2896
rect 19701 2954 19767 2957
rect 23800 2954 24600 2984
rect 19701 2952 24600 2954
rect 19701 2896 19706 2952
rect 19762 2896 24600 2952
rect 19701 2894 24600 2896
rect 9121 2891 9187 2894
rect 13537 2891 13603 2894
rect 19701 2891 19767 2894
rect 23800 2864 24600 2894
rect 6821 2818 6887 2821
rect 8293 2818 8359 2821
rect 6821 2816 8359 2818
rect 6821 2760 6826 2816
rect 6882 2760 8298 2816
rect 8354 2760 8359 2816
rect 6821 2758 8359 2760
rect 6821 2755 6887 2758
rect 8293 2755 8359 2758
rect 3743 2752 4063 2753
rect 3743 2688 3751 2752
rect 3815 2688 3831 2752
rect 3895 2688 3911 2752
rect 3975 2688 3991 2752
rect 4055 2688 4063 2752
rect 3743 2687 4063 2688
rect 9341 2752 9661 2753
rect 9341 2688 9349 2752
rect 9413 2688 9429 2752
rect 9493 2688 9509 2752
rect 9573 2688 9589 2752
rect 9653 2688 9661 2752
rect 9341 2687 9661 2688
rect 14939 2752 15259 2753
rect 14939 2688 14947 2752
rect 15011 2688 15027 2752
rect 15091 2688 15107 2752
rect 15171 2688 15187 2752
rect 15251 2688 15259 2752
rect 14939 2687 15259 2688
rect 20537 2752 20857 2753
rect 20537 2688 20545 2752
rect 20609 2688 20625 2752
rect 20689 2688 20705 2752
rect 20769 2688 20785 2752
rect 20849 2688 20857 2752
rect 20537 2687 20857 2688
rect 5901 2546 5967 2549
rect 7097 2546 7163 2549
rect 5901 2544 7163 2546
rect 5901 2488 5906 2544
rect 5962 2488 7102 2544
rect 7158 2488 7163 2544
rect 5901 2486 7163 2488
rect 5901 2483 5967 2486
rect 7097 2483 7163 2486
rect 16205 2546 16271 2549
rect 16614 2546 16620 2548
rect 16205 2544 16620 2546
rect 16205 2488 16210 2544
rect 16266 2488 16620 2544
rect 16205 2486 16620 2488
rect 16205 2483 16271 2486
rect 16614 2484 16620 2486
rect 16684 2484 16690 2548
rect 3325 2410 3391 2413
rect 19333 2410 19399 2413
rect 3325 2408 19399 2410
rect 3325 2352 3330 2408
rect 3386 2352 19338 2408
rect 19394 2352 19399 2408
rect 3325 2350 19399 2352
rect 3325 2347 3391 2350
rect 19333 2347 19399 2350
rect 20161 2274 20227 2277
rect 23800 2274 24600 2304
rect 20161 2272 24600 2274
rect 20161 2216 20166 2272
rect 20222 2216 24600 2272
rect 20161 2214 24600 2216
rect 20161 2211 20227 2214
rect 6542 2208 6862 2209
rect 6542 2144 6550 2208
rect 6614 2144 6630 2208
rect 6694 2144 6710 2208
rect 6774 2144 6790 2208
rect 6854 2144 6862 2208
rect 6542 2143 6862 2144
rect 12140 2208 12460 2209
rect 12140 2144 12148 2208
rect 12212 2144 12228 2208
rect 12292 2144 12308 2208
rect 12372 2144 12388 2208
rect 12452 2144 12460 2208
rect 12140 2143 12460 2144
rect 17738 2208 18058 2209
rect 17738 2144 17746 2208
rect 17810 2144 17826 2208
rect 17890 2144 17906 2208
rect 17970 2144 17986 2208
rect 18050 2144 18058 2208
rect 23800 2184 24600 2214
rect 17738 2143 18058 2144
rect 5349 2002 5415 2005
rect 18137 2002 18203 2005
rect 5349 2000 18203 2002
rect 5349 1944 5354 2000
rect 5410 1944 18142 2000
rect 18198 1944 18203 2000
rect 5349 1942 18203 1944
rect 5349 1939 5415 1942
rect 18137 1939 18203 1942
rect 3969 1866 4035 1869
rect 18413 1866 18479 1869
rect 3969 1864 18479 1866
rect 3969 1808 3974 1864
rect 4030 1808 18418 1864
rect 18474 1808 18479 1864
rect 3969 1806 18479 1808
rect 3969 1803 4035 1806
rect 18413 1803 18479 1806
rect 2957 1730 3023 1733
rect 18965 1730 19031 1733
rect 2957 1728 19031 1730
rect 2957 1672 2962 1728
rect 3018 1672 18970 1728
rect 19026 1672 19031 1728
rect 2957 1670 19031 1672
rect 2957 1667 3023 1670
rect 18965 1667 19031 1670
rect 20253 1594 20319 1597
rect 23800 1594 24600 1624
rect 20253 1592 24600 1594
rect 20253 1536 20258 1592
rect 20314 1536 24600 1592
rect 20253 1534 24600 1536
rect 20253 1531 20319 1534
rect 23800 1504 24600 1534
rect 21541 914 21607 917
rect 23800 914 24600 944
rect 21541 912 24600 914
rect 21541 856 21546 912
rect 21602 856 24600 912
rect 21541 854 24600 856
rect 21541 851 21607 854
rect 23800 824 24600 854
rect 19057 370 19123 373
rect 23800 370 24600 400
rect 19057 368 24600 370
rect 19057 312 19062 368
rect 19118 312 24600 368
rect 19057 310 24600 312
rect 19057 307 19123 310
rect 23800 280 24600 310
<< via3 >>
rect 3751 22332 3815 22336
rect 3751 22276 3755 22332
rect 3755 22276 3811 22332
rect 3811 22276 3815 22332
rect 3751 22272 3815 22276
rect 3831 22332 3895 22336
rect 3831 22276 3835 22332
rect 3835 22276 3891 22332
rect 3891 22276 3895 22332
rect 3831 22272 3895 22276
rect 3911 22332 3975 22336
rect 3911 22276 3915 22332
rect 3915 22276 3971 22332
rect 3971 22276 3975 22332
rect 3911 22272 3975 22276
rect 3991 22332 4055 22336
rect 3991 22276 3995 22332
rect 3995 22276 4051 22332
rect 4051 22276 4055 22332
rect 3991 22272 4055 22276
rect 9349 22332 9413 22336
rect 9349 22276 9353 22332
rect 9353 22276 9409 22332
rect 9409 22276 9413 22332
rect 9349 22272 9413 22276
rect 9429 22332 9493 22336
rect 9429 22276 9433 22332
rect 9433 22276 9489 22332
rect 9489 22276 9493 22332
rect 9429 22272 9493 22276
rect 9509 22332 9573 22336
rect 9509 22276 9513 22332
rect 9513 22276 9569 22332
rect 9569 22276 9573 22332
rect 9509 22272 9573 22276
rect 9589 22332 9653 22336
rect 9589 22276 9593 22332
rect 9593 22276 9649 22332
rect 9649 22276 9653 22332
rect 9589 22272 9653 22276
rect 14947 22332 15011 22336
rect 14947 22276 14951 22332
rect 14951 22276 15007 22332
rect 15007 22276 15011 22332
rect 14947 22272 15011 22276
rect 15027 22332 15091 22336
rect 15027 22276 15031 22332
rect 15031 22276 15087 22332
rect 15087 22276 15091 22332
rect 15027 22272 15091 22276
rect 15107 22332 15171 22336
rect 15107 22276 15111 22332
rect 15111 22276 15167 22332
rect 15167 22276 15171 22332
rect 15107 22272 15171 22276
rect 15187 22332 15251 22336
rect 15187 22276 15191 22332
rect 15191 22276 15247 22332
rect 15247 22276 15251 22332
rect 15187 22272 15251 22276
rect 20545 22332 20609 22336
rect 20545 22276 20549 22332
rect 20549 22276 20605 22332
rect 20605 22276 20609 22332
rect 20545 22272 20609 22276
rect 20625 22332 20689 22336
rect 20625 22276 20629 22332
rect 20629 22276 20685 22332
rect 20685 22276 20689 22332
rect 20625 22272 20689 22276
rect 20705 22332 20769 22336
rect 20705 22276 20709 22332
rect 20709 22276 20765 22332
rect 20765 22276 20769 22332
rect 20705 22272 20769 22276
rect 20785 22332 20849 22336
rect 20785 22276 20789 22332
rect 20789 22276 20845 22332
rect 20845 22276 20849 22332
rect 20785 22272 20849 22276
rect 9076 21992 9140 21996
rect 9076 21936 9126 21992
rect 9126 21936 9140 21992
rect 9076 21932 9140 21936
rect 6550 21788 6614 21792
rect 6550 21732 6554 21788
rect 6554 21732 6610 21788
rect 6610 21732 6614 21788
rect 6550 21728 6614 21732
rect 6630 21788 6694 21792
rect 6630 21732 6634 21788
rect 6634 21732 6690 21788
rect 6690 21732 6694 21788
rect 6630 21728 6694 21732
rect 6710 21788 6774 21792
rect 6710 21732 6714 21788
rect 6714 21732 6770 21788
rect 6770 21732 6774 21788
rect 6710 21728 6774 21732
rect 6790 21788 6854 21792
rect 6790 21732 6794 21788
rect 6794 21732 6850 21788
rect 6850 21732 6854 21788
rect 6790 21728 6854 21732
rect 12148 21788 12212 21792
rect 12148 21732 12152 21788
rect 12152 21732 12208 21788
rect 12208 21732 12212 21788
rect 12148 21728 12212 21732
rect 12228 21788 12292 21792
rect 12228 21732 12232 21788
rect 12232 21732 12288 21788
rect 12288 21732 12292 21788
rect 12228 21728 12292 21732
rect 12308 21788 12372 21792
rect 12308 21732 12312 21788
rect 12312 21732 12368 21788
rect 12368 21732 12372 21788
rect 12308 21728 12372 21732
rect 12388 21788 12452 21792
rect 12388 21732 12392 21788
rect 12392 21732 12448 21788
rect 12448 21732 12452 21788
rect 12388 21728 12452 21732
rect 17746 21788 17810 21792
rect 17746 21732 17750 21788
rect 17750 21732 17806 21788
rect 17806 21732 17810 21788
rect 17746 21728 17810 21732
rect 17826 21788 17890 21792
rect 17826 21732 17830 21788
rect 17830 21732 17886 21788
rect 17886 21732 17890 21788
rect 17826 21728 17890 21732
rect 17906 21788 17970 21792
rect 17906 21732 17910 21788
rect 17910 21732 17966 21788
rect 17966 21732 17970 21788
rect 17906 21728 17970 21732
rect 17986 21788 18050 21792
rect 17986 21732 17990 21788
rect 17990 21732 18046 21788
rect 18046 21732 18050 21788
rect 17986 21728 18050 21732
rect 3751 21244 3815 21248
rect 3751 21188 3755 21244
rect 3755 21188 3811 21244
rect 3811 21188 3815 21244
rect 3751 21184 3815 21188
rect 3831 21244 3895 21248
rect 3831 21188 3835 21244
rect 3835 21188 3891 21244
rect 3891 21188 3895 21244
rect 3831 21184 3895 21188
rect 3911 21244 3975 21248
rect 3911 21188 3915 21244
rect 3915 21188 3971 21244
rect 3971 21188 3975 21244
rect 3911 21184 3975 21188
rect 3991 21244 4055 21248
rect 3991 21188 3995 21244
rect 3995 21188 4051 21244
rect 4051 21188 4055 21244
rect 3991 21184 4055 21188
rect 9349 21244 9413 21248
rect 9349 21188 9353 21244
rect 9353 21188 9409 21244
rect 9409 21188 9413 21244
rect 9349 21184 9413 21188
rect 9429 21244 9493 21248
rect 9429 21188 9433 21244
rect 9433 21188 9489 21244
rect 9489 21188 9493 21244
rect 9429 21184 9493 21188
rect 9509 21244 9573 21248
rect 9509 21188 9513 21244
rect 9513 21188 9569 21244
rect 9569 21188 9573 21244
rect 9509 21184 9573 21188
rect 9589 21244 9653 21248
rect 9589 21188 9593 21244
rect 9593 21188 9649 21244
rect 9649 21188 9653 21244
rect 9589 21184 9653 21188
rect 14947 21244 15011 21248
rect 14947 21188 14951 21244
rect 14951 21188 15007 21244
rect 15007 21188 15011 21244
rect 14947 21184 15011 21188
rect 15027 21244 15091 21248
rect 15027 21188 15031 21244
rect 15031 21188 15087 21244
rect 15087 21188 15091 21244
rect 15027 21184 15091 21188
rect 15107 21244 15171 21248
rect 15107 21188 15111 21244
rect 15111 21188 15167 21244
rect 15167 21188 15171 21244
rect 15107 21184 15171 21188
rect 15187 21244 15251 21248
rect 15187 21188 15191 21244
rect 15191 21188 15247 21244
rect 15247 21188 15251 21244
rect 15187 21184 15251 21188
rect 20545 21244 20609 21248
rect 20545 21188 20549 21244
rect 20549 21188 20605 21244
rect 20605 21188 20609 21244
rect 20545 21184 20609 21188
rect 20625 21244 20689 21248
rect 20625 21188 20629 21244
rect 20629 21188 20685 21244
rect 20685 21188 20689 21244
rect 20625 21184 20689 21188
rect 20705 21244 20769 21248
rect 20705 21188 20709 21244
rect 20709 21188 20765 21244
rect 20765 21188 20769 21244
rect 20705 21184 20769 21188
rect 20785 21244 20849 21248
rect 20785 21188 20789 21244
rect 20789 21188 20845 21244
rect 20845 21188 20849 21244
rect 20785 21184 20849 21188
rect 19380 20980 19444 21044
rect 21220 20844 21284 20908
rect 6550 20700 6614 20704
rect 6550 20644 6554 20700
rect 6554 20644 6610 20700
rect 6610 20644 6614 20700
rect 6550 20640 6614 20644
rect 6630 20700 6694 20704
rect 6630 20644 6634 20700
rect 6634 20644 6690 20700
rect 6690 20644 6694 20700
rect 6630 20640 6694 20644
rect 6710 20700 6774 20704
rect 6710 20644 6714 20700
rect 6714 20644 6770 20700
rect 6770 20644 6774 20700
rect 6710 20640 6774 20644
rect 6790 20700 6854 20704
rect 6790 20644 6794 20700
rect 6794 20644 6850 20700
rect 6850 20644 6854 20700
rect 6790 20640 6854 20644
rect 12148 20700 12212 20704
rect 12148 20644 12152 20700
rect 12152 20644 12208 20700
rect 12208 20644 12212 20700
rect 12148 20640 12212 20644
rect 12228 20700 12292 20704
rect 12228 20644 12232 20700
rect 12232 20644 12288 20700
rect 12288 20644 12292 20700
rect 12228 20640 12292 20644
rect 12308 20700 12372 20704
rect 12308 20644 12312 20700
rect 12312 20644 12368 20700
rect 12368 20644 12372 20700
rect 12308 20640 12372 20644
rect 12388 20700 12452 20704
rect 12388 20644 12392 20700
rect 12392 20644 12448 20700
rect 12448 20644 12452 20700
rect 12388 20640 12452 20644
rect 17746 20700 17810 20704
rect 17746 20644 17750 20700
rect 17750 20644 17806 20700
rect 17806 20644 17810 20700
rect 17746 20640 17810 20644
rect 17826 20700 17890 20704
rect 17826 20644 17830 20700
rect 17830 20644 17886 20700
rect 17886 20644 17890 20700
rect 17826 20640 17890 20644
rect 17906 20700 17970 20704
rect 17906 20644 17910 20700
rect 17910 20644 17966 20700
rect 17966 20644 17970 20700
rect 17906 20640 17970 20644
rect 17986 20700 18050 20704
rect 17986 20644 17990 20700
rect 17990 20644 18046 20700
rect 18046 20644 18050 20700
rect 17986 20640 18050 20644
rect 22876 20300 22940 20364
rect 3751 20156 3815 20160
rect 3751 20100 3755 20156
rect 3755 20100 3811 20156
rect 3811 20100 3815 20156
rect 3751 20096 3815 20100
rect 3831 20156 3895 20160
rect 3831 20100 3835 20156
rect 3835 20100 3891 20156
rect 3891 20100 3895 20156
rect 3831 20096 3895 20100
rect 3911 20156 3975 20160
rect 3911 20100 3915 20156
rect 3915 20100 3971 20156
rect 3971 20100 3975 20156
rect 3911 20096 3975 20100
rect 3991 20156 4055 20160
rect 3991 20100 3995 20156
rect 3995 20100 4051 20156
rect 4051 20100 4055 20156
rect 3991 20096 4055 20100
rect 9349 20156 9413 20160
rect 9349 20100 9353 20156
rect 9353 20100 9409 20156
rect 9409 20100 9413 20156
rect 9349 20096 9413 20100
rect 9429 20156 9493 20160
rect 9429 20100 9433 20156
rect 9433 20100 9489 20156
rect 9489 20100 9493 20156
rect 9429 20096 9493 20100
rect 9509 20156 9573 20160
rect 9509 20100 9513 20156
rect 9513 20100 9569 20156
rect 9569 20100 9573 20156
rect 9509 20096 9573 20100
rect 9589 20156 9653 20160
rect 9589 20100 9593 20156
rect 9593 20100 9649 20156
rect 9649 20100 9653 20156
rect 9589 20096 9653 20100
rect 14947 20156 15011 20160
rect 14947 20100 14951 20156
rect 14951 20100 15007 20156
rect 15007 20100 15011 20156
rect 14947 20096 15011 20100
rect 15027 20156 15091 20160
rect 15027 20100 15031 20156
rect 15031 20100 15087 20156
rect 15087 20100 15091 20156
rect 15027 20096 15091 20100
rect 15107 20156 15171 20160
rect 15107 20100 15111 20156
rect 15111 20100 15167 20156
rect 15167 20100 15171 20156
rect 15107 20096 15171 20100
rect 15187 20156 15251 20160
rect 15187 20100 15191 20156
rect 15191 20100 15247 20156
rect 15247 20100 15251 20156
rect 15187 20096 15251 20100
rect 20545 20156 20609 20160
rect 20545 20100 20549 20156
rect 20549 20100 20605 20156
rect 20605 20100 20609 20156
rect 20545 20096 20609 20100
rect 20625 20156 20689 20160
rect 20625 20100 20629 20156
rect 20629 20100 20685 20156
rect 20685 20100 20689 20156
rect 20625 20096 20689 20100
rect 20705 20156 20769 20160
rect 20705 20100 20709 20156
rect 20709 20100 20765 20156
rect 20765 20100 20769 20156
rect 20705 20096 20769 20100
rect 20785 20156 20849 20160
rect 20785 20100 20789 20156
rect 20789 20100 20845 20156
rect 20845 20100 20849 20156
rect 20785 20096 20849 20100
rect 7972 20028 8036 20092
rect 6550 19612 6614 19616
rect 6550 19556 6554 19612
rect 6554 19556 6610 19612
rect 6610 19556 6614 19612
rect 6550 19552 6614 19556
rect 6630 19612 6694 19616
rect 6630 19556 6634 19612
rect 6634 19556 6690 19612
rect 6690 19556 6694 19612
rect 6630 19552 6694 19556
rect 6710 19612 6774 19616
rect 6710 19556 6714 19612
rect 6714 19556 6770 19612
rect 6770 19556 6774 19612
rect 6710 19552 6774 19556
rect 6790 19612 6854 19616
rect 6790 19556 6794 19612
rect 6794 19556 6850 19612
rect 6850 19556 6854 19612
rect 6790 19552 6854 19556
rect 12148 19612 12212 19616
rect 12148 19556 12152 19612
rect 12152 19556 12208 19612
rect 12208 19556 12212 19612
rect 12148 19552 12212 19556
rect 12228 19612 12292 19616
rect 12228 19556 12232 19612
rect 12232 19556 12288 19612
rect 12288 19556 12292 19612
rect 12228 19552 12292 19556
rect 12308 19612 12372 19616
rect 12308 19556 12312 19612
rect 12312 19556 12368 19612
rect 12368 19556 12372 19612
rect 12308 19552 12372 19556
rect 12388 19612 12452 19616
rect 12388 19556 12392 19612
rect 12392 19556 12448 19612
rect 12448 19556 12452 19612
rect 12388 19552 12452 19556
rect 17746 19612 17810 19616
rect 17746 19556 17750 19612
rect 17750 19556 17806 19612
rect 17806 19556 17810 19612
rect 17746 19552 17810 19556
rect 17826 19612 17890 19616
rect 17826 19556 17830 19612
rect 17830 19556 17886 19612
rect 17886 19556 17890 19612
rect 17826 19552 17890 19556
rect 17906 19612 17970 19616
rect 17906 19556 17910 19612
rect 17910 19556 17966 19612
rect 17966 19556 17970 19612
rect 17906 19552 17970 19556
rect 17986 19612 18050 19616
rect 17986 19556 17990 19612
rect 17990 19556 18046 19612
rect 18046 19556 18050 19612
rect 17986 19552 18050 19556
rect 3751 19068 3815 19072
rect 3751 19012 3755 19068
rect 3755 19012 3811 19068
rect 3811 19012 3815 19068
rect 3751 19008 3815 19012
rect 3831 19068 3895 19072
rect 3831 19012 3835 19068
rect 3835 19012 3891 19068
rect 3891 19012 3895 19068
rect 3831 19008 3895 19012
rect 3911 19068 3975 19072
rect 3911 19012 3915 19068
rect 3915 19012 3971 19068
rect 3971 19012 3975 19068
rect 3911 19008 3975 19012
rect 3991 19068 4055 19072
rect 3991 19012 3995 19068
rect 3995 19012 4051 19068
rect 4051 19012 4055 19068
rect 3991 19008 4055 19012
rect 9349 19068 9413 19072
rect 9349 19012 9353 19068
rect 9353 19012 9409 19068
rect 9409 19012 9413 19068
rect 9349 19008 9413 19012
rect 9429 19068 9493 19072
rect 9429 19012 9433 19068
rect 9433 19012 9489 19068
rect 9489 19012 9493 19068
rect 9429 19008 9493 19012
rect 9509 19068 9573 19072
rect 9509 19012 9513 19068
rect 9513 19012 9569 19068
rect 9569 19012 9573 19068
rect 9509 19008 9573 19012
rect 9589 19068 9653 19072
rect 9589 19012 9593 19068
rect 9593 19012 9649 19068
rect 9649 19012 9653 19068
rect 9589 19008 9653 19012
rect 14947 19068 15011 19072
rect 14947 19012 14951 19068
rect 14951 19012 15007 19068
rect 15007 19012 15011 19068
rect 14947 19008 15011 19012
rect 15027 19068 15091 19072
rect 15027 19012 15031 19068
rect 15031 19012 15087 19068
rect 15087 19012 15091 19068
rect 15027 19008 15091 19012
rect 15107 19068 15171 19072
rect 15107 19012 15111 19068
rect 15111 19012 15167 19068
rect 15167 19012 15171 19068
rect 15107 19008 15171 19012
rect 15187 19068 15251 19072
rect 15187 19012 15191 19068
rect 15191 19012 15247 19068
rect 15247 19012 15251 19068
rect 15187 19008 15251 19012
rect 20545 19068 20609 19072
rect 20545 19012 20549 19068
rect 20549 19012 20605 19068
rect 20605 19012 20609 19068
rect 20545 19008 20609 19012
rect 20625 19068 20689 19072
rect 20625 19012 20629 19068
rect 20629 19012 20685 19068
rect 20685 19012 20689 19068
rect 20625 19008 20689 19012
rect 20705 19068 20769 19072
rect 20705 19012 20709 19068
rect 20709 19012 20765 19068
rect 20765 19012 20769 19068
rect 20705 19008 20769 19012
rect 20785 19068 20849 19072
rect 20785 19012 20789 19068
rect 20789 19012 20845 19068
rect 20845 19012 20849 19068
rect 20785 19008 20849 19012
rect 6550 18524 6614 18528
rect 6550 18468 6554 18524
rect 6554 18468 6610 18524
rect 6610 18468 6614 18524
rect 6550 18464 6614 18468
rect 6630 18524 6694 18528
rect 6630 18468 6634 18524
rect 6634 18468 6690 18524
rect 6690 18468 6694 18524
rect 6630 18464 6694 18468
rect 6710 18524 6774 18528
rect 6710 18468 6714 18524
rect 6714 18468 6770 18524
rect 6770 18468 6774 18524
rect 6710 18464 6774 18468
rect 6790 18524 6854 18528
rect 6790 18468 6794 18524
rect 6794 18468 6850 18524
rect 6850 18468 6854 18524
rect 6790 18464 6854 18468
rect 12148 18524 12212 18528
rect 12148 18468 12152 18524
rect 12152 18468 12208 18524
rect 12208 18468 12212 18524
rect 12148 18464 12212 18468
rect 12228 18524 12292 18528
rect 12228 18468 12232 18524
rect 12232 18468 12288 18524
rect 12288 18468 12292 18524
rect 12228 18464 12292 18468
rect 12308 18524 12372 18528
rect 12308 18468 12312 18524
rect 12312 18468 12368 18524
rect 12368 18468 12372 18524
rect 12308 18464 12372 18468
rect 12388 18524 12452 18528
rect 12388 18468 12392 18524
rect 12392 18468 12448 18524
rect 12448 18468 12452 18524
rect 12388 18464 12452 18468
rect 17746 18524 17810 18528
rect 17746 18468 17750 18524
rect 17750 18468 17806 18524
rect 17806 18468 17810 18524
rect 17746 18464 17810 18468
rect 17826 18524 17890 18528
rect 17826 18468 17830 18524
rect 17830 18468 17886 18524
rect 17886 18468 17890 18524
rect 17826 18464 17890 18468
rect 17906 18524 17970 18528
rect 17906 18468 17910 18524
rect 17910 18468 17966 18524
rect 17966 18468 17970 18524
rect 17906 18464 17970 18468
rect 17986 18524 18050 18528
rect 17986 18468 17990 18524
rect 17990 18468 18046 18524
rect 18046 18468 18050 18524
rect 17986 18464 18050 18468
rect 3751 17980 3815 17984
rect 3751 17924 3755 17980
rect 3755 17924 3811 17980
rect 3811 17924 3815 17980
rect 3751 17920 3815 17924
rect 3831 17980 3895 17984
rect 3831 17924 3835 17980
rect 3835 17924 3891 17980
rect 3891 17924 3895 17980
rect 3831 17920 3895 17924
rect 3911 17980 3975 17984
rect 3911 17924 3915 17980
rect 3915 17924 3971 17980
rect 3971 17924 3975 17980
rect 3911 17920 3975 17924
rect 3991 17980 4055 17984
rect 3991 17924 3995 17980
rect 3995 17924 4051 17980
rect 4051 17924 4055 17980
rect 3991 17920 4055 17924
rect 9349 17980 9413 17984
rect 9349 17924 9353 17980
rect 9353 17924 9409 17980
rect 9409 17924 9413 17980
rect 9349 17920 9413 17924
rect 9429 17980 9493 17984
rect 9429 17924 9433 17980
rect 9433 17924 9489 17980
rect 9489 17924 9493 17980
rect 9429 17920 9493 17924
rect 9509 17980 9573 17984
rect 9509 17924 9513 17980
rect 9513 17924 9569 17980
rect 9569 17924 9573 17980
rect 9509 17920 9573 17924
rect 9589 17980 9653 17984
rect 9589 17924 9593 17980
rect 9593 17924 9649 17980
rect 9649 17924 9653 17980
rect 9589 17920 9653 17924
rect 14947 17980 15011 17984
rect 14947 17924 14951 17980
rect 14951 17924 15007 17980
rect 15007 17924 15011 17980
rect 14947 17920 15011 17924
rect 15027 17980 15091 17984
rect 15027 17924 15031 17980
rect 15031 17924 15087 17980
rect 15087 17924 15091 17980
rect 15027 17920 15091 17924
rect 15107 17980 15171 17984
rect 15107 17924 15111 17980
rect 15111 17924 15167 17980
rect 15167 17924 15171 17980
rect 15107 17920 15171 17924
rect 15187 17980 15251 17984
rect 15187 17924 15191 17980
rect 15191 17924 15247 17980
rect 15247 17924 15251 17980
rect 15187 17920 15251 17924
rect 20545 17980 20609 17984
rect 20545 17924 20549 17980
rect 20549 17924 20605 17980
rect 20605 17924 20609 17980
rect 20545 17920 20609 17924
rect 20625 17980 20689 17984
rect 20625 17924 20629 17980
rect 20629 17924 20685 17980
rect 20685 17924 20689 17980
rect 20625 17920 20689 17924
rect 20705 17980 20769 17984
rect 20705 17924 20709 17980
rect 20709 17924 20765 17980
rect 20765 17924 20769 17980
rect 20705 17920 20769 17924
rect 20785 17980 20849 17984
rect 20785 17924 20789 17980
rect 20789 17924 20845 17980
rect 20845 17924 20849 17980
rect 20785 17920 20849 17924
rect 21036 17852 21100 17916
rect 6550 17436 6614 17440
rect 6550 17380 6554 17436
rect 6554 17380 6610 17436
rect 6610 17380 6614 17436
rect 6550 17376 6614 17380
rect 6630 17436 6694 17440
rect 6630 17380 6634 17436
rect 6634 17380 6690 17436
rect 6690 17380 6694 17436
rect 6630 17376 6694 17380
rect 6710 17436 6774 17440
rect 6710 17380 6714 17436
rect 6714 17380 6770 17436
rect 6770 17380 6774 17436
rect 6710 17376 6774 17380
rect 6790 17436 6854 17440
rect 6790 17380 6794 17436
rect 6794 17380 6850 17436
rect 6850 17380 6854 17436
rect 6790 17376 6854 17380
rect 12148 17436 12212 17440
rect 12148 17380 12152 17436
rect 12152 17380 12208 17436
rect 12208 17380 12212 17436
rect 12148 17376 12212 17380
rect 12228 17436 12292 17440
rect 12228 17380 12232 17436
rect 12232 17380 12288 17436
rect 12288 17380 12292 17436
rect 12228 17376 12292 17380
rect 12308 17436 12372 17440
rect 12308 17380 12312 17436
rect 12312 17380 12368 17436
rect 12368 17380 12372 17436
rect 12308 17376 12372 17380
rect 12388 17436 12452 17440
rect 12388 17380 12392 17436
rect 12392 17380 12448 17436
rect 12448 17380 12452 17436
rect 12388 17376 12452 17380
rect 17746 17436 17810 17440
rect 17746 17380 17750 17436
rect 17750 17380 17806 17436
rect 17806 17380 17810 17436
rect 17746 17376 17810 17380
rect 17826 17436 17890 17440
rect 17826 17380 17830 17436
rect 17830 17380 17886 17436
rect 17886 17380 17890 17436
rect 17826 17376 17890 17380
rect 17906 17436 17970 17440
rect 17906 17380 17910 17436
rect 17910 17380 17966 17436
rect 17966 17380 17970 17436
rect 17906 17376 17970 17380
rect 17986 17436 18050 17440
rect 17986 17380 17990 17436
rect 17990 17380 18046 17436
rect 18046 17380 18050 17436
rect 17986 17376 18050 17380
rect 20300 17444 20364 17508
rect 9076 17096 9140 17100
rect 9076 17040 9126 17096
rect 9126 17040 9140 17096
rect 9076 17036 9140 17040
rect 3751 16892 3815 16896
rect 3751 16836 3755 16892
rect 3755 16836 3811 16892
rect 3811 16836 3815 16892
rect 3751 16832 3815 16836
rect 3831 16892 3895 16896
rect 3831 16836 3835 16892
rect 3835 16836 3891 16892
rect 3891 16836 3895 16892
rect 3831 16832 3895 16836
rect 3911 16892 3975 16896
rect 3911 16836 3915 16892
rect 3915 16836 3971 16892
rect 3971 16836 3975 16892
rect 3911 16832 3975 16836
rect 3991 16892 4055 16896
rect 3991 16836 3995 16892
rect 3995 16836 4051 16892
rect 4051 16836 4055 16892
rect 3991 16832 4055 16836
rect 9349 16892 9413 16896
rect 9349 16836 9353 16892
rect 9353 16836 9409 16892
rect 9409 16836 9413 16892
rect 9349 16832 9413 16836
rect 9429 16892 9493 16896
rect 9429 16836 9433 16892
rect 9433 16836 9489 16892
rect 9489 16836 9493 16892
rect 9429 16832 9493 16836
rect 9509 16892 9573 16896
rect 9509 16836 9513 16892
rect 9513 16836 9569 16892
rect 9569 16836 9573 16892
rect 9509 16832 9573 16836
rect 9589 16892 9653 16896
rect 9589 16836 9593 16892
rect 9593 16836 9649 16892
rect 9649 16836 9653 16892
rect 9589 16832 9653 16836
rect 14947 16892 15011 16896
rect 14947 16836 14951 16892
rect 14951 16836 15007 16892
rect 15007 16836 15011 16892
rect 14947 16832 15011 16836
rect 15027 16892 15091 16896
rect 15027 16836 15031 16892
rect 15031 16836 15087 16892
rect 15087 16836 15091 16892
rect 15027 16832 15091 16836
rect 15107 16892 15171 16896
rect 15107 16836 15111 16892
rect 15111 16836 15167 16892
rect 15167 16836 15171 16892
rect 15107 16832 15171 16836
rect 15187 16892 15251 16896
rect 15187 16836 15191 16892
rect 15191 16836 15247 16892
rect 15247 16836 15251 16892
rect 15187 16832 15251 16836
rect 20545 16892 20609 16896
rect 20545 16836 20549 16892
rect 20549 16836 20605 16892
rect 20605 16836 20609 16892
rect 20545 16832 20609 16836
rect 20625 16892 20689 16896
rect 20625 16836 20629 16892
rect 20629 16836 20685 16892
rect 20685 16836 20689 16892
rect 20625 16832 20689 16836
rect 20705 16892 20769 16896
rect 20705 16836 20709 16892
rect 20709 16836 20765 16892
rect 20765 16836 20769 16892
rect 20705 16832 20769 16836
rect 20785 16892 20849 16896
rect 20785 16836 20789 16892
rect 20789 16836 20845 16892
rect 20845 16836 20849 16892
rect 20785 16832 20849 16836
rect 6550 16348 6614 16352
rect 6550 16292 6554 16348
rect 6554 16292 6610 16348
rect 6610 16292 6614 16348
rect 6550 16288 6614 16292
rect 6630 16348 6694 16352
rect 6630 16292 6634 16348
rect 6634 16292 6690 16348
rect 6690 16292 6694 16348
rect 6630 16288 6694 16292
rect 6710 16348 6774 16352
rect 6710 16292 6714 16348
rect 6714 16292 6770 16348
rect 6770 16292 6774 16348
rect 6710 16288 6774 16292
rect 6790 16348 6854 16352
rect 6790 16292 6794 16348
rect 6794 16292 6850 16348
rect 6850 16292 6854 16348
rect 6790 16288 6854 16292
rect 12148 16348 12212 16352
rect 12148 16292 12152 16348
rect 12152 16292 12208 16348
rect 12208 16292 12212 16348
rect 12148 16288 12212 16292
rect 12228 16348 12292 16352
rect 12228 16292 12232 16348
rect 12232 16292 12288 16348
rect 12288 16292 12292 16348
rect 12228 16288 12292 16292
rect 12308 16348 12372 16352
rect 12308 16292 12312 16348
rect 12312 16292 12368 16348
rect 12368 16292 12372 16348
rect 12308 16288 12372 16292
rect 12388 16348 12452 16352
rect 12388 16292 12392 16348
rect 12392 16292 12448 16348
rect 12448 16292 12452 16348
rect 12388 16288 12452 16292
rect 17746 16348 17810 16352
rect 17746 16292 17750 16348
rect 17750 16292 17806 16348
rect 17806 16292 17810 16348
rect 17746 16288 17810 16292
rect 17826 16348 17890 16352
rect 17826 16292 17830 16348
rect 17830 16292 17886 16348
rect 17886 16292 17890 16348
rect 17826 16288 17890 16292
rect 17906 16348 17970 16352
rect 17906 16292 17910 16348
rect 17910 16292 17966 16348
rect 17966 16292 17970 16348
rect 17906 16288 17970 16292
rect 17986 16348 18050 16352
rect 17986 16292 17990 16348
rect 17990 16292 18046 16348
rect 18046 16292 18050 16348
rect 17986 16288 18050 16292
rect 3751 15804 3815 15808
rect 3751 15748 3755 15804
rect 3755 15748 3811 15804
rect 3811 15748 3815 15804
rect 3751 15744 3815 15748
rect 3831 15804 3895 15808
rect 3831 15748 3835 15804
rect 3835 15748 3891 15804
rect 3891 15748 3895 15804
rect 3831 15744 3895 15748
rect 3911 15804 3975 15808
rect 3911 15748 3915 15804
rect 3915 15748 3971 15804
rect 3971 15748 3975 15804
rect 3911 15744 3975 15748
rect 3991 15804 4055 15808
rect 3991 15748 3995 15804
rect 3995 15748 4051 15804
rect 4051 15748 4055 15804
rect 3991 15744 4055 15748
rect 9349 15804 9413 15808
rect 9349 15748 9353 15804
rect 9353 15748 9409 15804
rect 9409 15748 9413 15804
rect 9349 15744 9413 15748
rect 9429 15804 9493 15808
rect 9429 15748 9433 15804
rect 9433 15748 9489 15804
rect 9489 15748 9493 15804
rect 9429 15744 9493 15748
rect 9509 15804 9573 15808
rect 9509 15748 9513 15804
rect 9513 15748 9569 15804
rect 9569 15748 9573 15804
rect 9509 15744 9573 15748
rect 9589 15804 9653 15808
rect 9589 15748 9593 15804
rect 9593 15748 9649 15804
rect 9649 15748 9653 15804
rect 9589 15744 9653 15748
rect 14947 15804 15011 15808
rect 14947 15748 14951 15804
rect 14951 15748 15007 15804
rect 15007 15748 15011 15804
rect 14947 15744 15011 15748
rect 15027 15804 15091 15808
rect 15027 15748 15031 15804
rect 15031 15748 15087 15804
rect 15087 15748 15091 15804
rect 15027 15744 15091 15748
rect 15107 15804 15171 15808
rect 15107 15748 15111 15804
rect 15111 15748 15167 15804
rect 15167 15748 15171 15804
rect 15107 15744 15171 15748
rect 15187 15804 15251 15808
rect 15187 15748 15191 15804
rect 15191 15748 15247 15804
rect 15247 15748 15251 15804
rect 15187 15744 15251 15748
rect 20545 15804 20609 15808
rect 20545 15748 20549 15804
rect 20549 15748 20605 15804
rect 20605 15748 20609 15804
rect 20545 15744 20609 15748
rect 20625 15804 20689 15808
rect 20625 15748 20629 15804
rect 20629 15748 20685 15804
rect 20685 15748 20689 15804
rect 20625 15744 20689 15748
rect 20705 15804 20769 15808
rect 20705 15748 20709 15804
rect 20709 15748 20765 15804
rect 20765 15748 20769 15804
rect 20705 15744 20769 15748
rect 20785 15804 20849 15808
rect 20785 15748 20789 15804
rect 20789 15748 20845 15804
rect 20845 15748 20849 15804
rect 20785 15744 20849 15748
rect 6550 15260 6614 15264
rect 6550 15204 6554 15260
rect 6554 15204 6610 15260
rect 6610 15204 6614 15260
rect 6550 15200 6614 15204
rect 6630 15260 6694 15264
rect 6630 15204 6634 15260
rect 6634 15204 6690 15260
rect 6690 15204 6694 15260
rect 6630 15200 6694 15204
rect 6710 15260 6774 15264
rect 6710 15204 6714 15260
rect 6714 15204 6770 15260
rect 6770 15204 6774 15260
rect 6710 15200 6774 15204
rect 6790 15260 6854 15264
rect 6790 15204 6794 15260
rect 6794 15204 6850 15260
rect 6850 15204 6854 15260
rect 6790 15200 6854 15204
rect 12148 15260 12212 15264
rect 12148 15204 12152 15260
rect 12152 15204 12208 15260
rect 12208 15204 12212 15260
rect 12148 15200 12212 15204
rect 12228 15260 12292 15264
rect 12228 15204 12232 15260
rect 12232 15204 12288 15260
rect 12288 15204 12292 15260
rect 12228 15200 12292 15204
rect 12308 15260 12372 15264
rect 12308 15204 12312 15260
rect 12312 15204 12368 15260
rect 12368 15204 12372 15260
rect 12308 15200 12372 15204
rect 12388 15260 12452 15264
rect 12388 15204 12392 15260
rect 12392 15204 12448 15260
rect 12448 15204 12452 15260
rect 12388 15200 12452 15204
rect 17746 15260 17810 15264
rect 17746 15204 17750 15260
rect 17750 15204 17806 15260
rect 17806 15204 17810 15260
rect 17746 15200 17810 15204
rect 17826 15260 17890 15264
rect 17826 15204 17830 15260
rect 17830 15204 17886 15260
rect 17886 15204 17890 15260
rect 17826 15200 17890 15204
rect 17906 15260 17970 15264
rect 17906 15204 17910 15260
rect 17910 15204 17966 15260
rect 17966 15204 17970 15260
rect 17906 15200 17970 15204
rect 17986 15260 18050 15264
rect 17986 15204 17990 15260
rect 17990 15204 18046 15260
rect 18046 15204 18050 15260
rect 17986 15200 18050 15204
rect 21220 14860 21284 14924
rect 3751 14716 3815 14720
rect 3751 14660 3755 14716
rect 3755 14660 3811 14716
rect 3811 14660 3815 14716
rect 3751 14656 3815 14660
rect 3831 14716 3895 14720
rect 3831 14660 3835 14716
rect 3835 14660 3891 14716
rect 3891 14660 3895 14716
rect 3831 14656 3895 14660
rect 3911 14716 3975 14720
rect 3911 14660 3915 14716
rect 3915 14660 3971 14716
rect 3971 14660 3975 14716
rect 3911 14656 3975 14660
rect 3991 14716 4055 14720
rect 3991 14660 3995 14716
rect 3995 14660 4051 14716
rect 4051 14660 4055 14716
rect 3991 14656 4055 14660
rect 9349 14716 9413 14720
rect 9349 14660 9353 14716
rect 9353 14660 9409 14716
rect 9409 14660 9413 14716
rect 9349 14656 9413 14660
rect 9429 14716 9493 14720
rect 9429 14660 9433 14716
rect 9433 14660 9489 14716
rect 9489 14660 9493 14716
rect 9429 14656 9493 14660
rect 9509 14716 9573 14720
rect 9509 14660 9513 14716
rect 9513 14660 9569 14716
rect 9569 14660 9573 14716
rect 9509 14656 9573 14660
rect 9589 14716 9653 14720
rect 9589 14660 9593 14716
rect 9593 14660 9649 14716
rect 9649 14660 9653 14716
rect 9589 14656 9653 14660
rect 14947 14716 15011 14720
rect 14947 14660 14951 14716
rect 14951 14660 15007 14716
rect 15007 14660 15011 14716
rect 14947 14656 15011 14660
rect 15027 14716 15091 14720
rect 15027 14660 15031 14716
rect 15031 14660 15087 14716
rect 15087 14660 15091 14716
rect 15027 14656 15091 14660
rect 15107 14716 15171 14720
rect 15107 14660 15111 14716
rect 15111 14660 15167 14716
rect 15167 14660 15171 14716
rect 15107 14656 15171 14660
rect 15187 14716 15251 14720
rect 15187 14660 15191 14716
rect 15191 14660 15247 14716
rect 15247 14660 15251 14716
rect 15187 14656 15251 14660
rect 20545 14716 20609 14720
rect 20545 14660 20549 14716
rect 20549 14660 20605 14716
rect 20605 14660 20609 14716
rect 20545 14656 20609 14660
rect 20625 14716 20689 14720
rect 20625 14660 20629 14716
rect 20629 14660 20685 14716
rect 20685 14660 20689 14716
rect 20625 14656 20689 14660
rect 20705 14716 20769 14720
rect 20705 14660 20709 14716
rect 20709 14660 20765 14716
rect 20765 14660 20769 14716
rect 20705 14656 20769 14660
rect 20785 14716 20849 14720
rect 20785 14660 20789 14716
rect 20789 14660 20845 14716
rect 20845 14660 20849 14716
rect 20785 14656 20849 14660
rect 6550 14172 6614 14176
rect 6550 14116 6554 14172
rect 6554 14116 6610 14172
rect 6610 14116 6614 14172
rect 6550 14112 6614 14116
rect 6630 14172 6694 14176
rect 6630 14116 6634 14172
rect 6634 14116 6690 14172
rect 6690 14116 6694 14172
rect 6630 14112 6694 14116
rect 6710 14172 6774 14176
rect 6710 14116 6714 14172
rect 6714 14116 6770 14172
rect 6770 14116 6774 14172
rect 6710 14112 6774 14116
rect 6790 14172 6854 14176
rect 6790 14116 6794 14172
rect 6794 14116 6850 14172
rect 6850 14116 6854 14172
rect 6790 14112 6854 14116
rect 12148 14172 12212 14176
rect 12148 14116 12152 14172
rect 12152 14116 12208 14172
rect 12208 14116 12212 14172
rect 12148 14112 12212 14116
rect 12228 14172 12292 14176
rect 12228 14116 12232 14172
rect 12232 14116 12288 14172
rect 12288 14116 12292 14172
rect 12228 14112 12292 14116
rect 12308 14172 12372 14176
rect 12308 14116 12312 14172
rect 12312 14116 12368 14172
rect 12368 14116 12372 14172
rect 12308 14112 12372 14116
rect 12388 14172 12452 14176
rect 12388 14116 12392 14172
rect 12392 14116 12448 14172
rect 12448 14116 12452 14172
rect 12388 14112 12452 14116
rect 17746 14172 17810 14176
rect 17746 14116 17750 14172
rect 17750 14116 17806 14172
rect 17806 14116 17810 14172
rect 17746 14112 17810 14116
rect 17826 14172 17890 14176
rect 17826 14116 17830 14172
rect 17830 14116 17886 14172
rect 17886 14116 17890 14172
rect 17826 14112 17890 14116
rect 17906 14172 17970 14176
rect 17906 14116 17910 14172
rect 17910 14116 17966 14172
rect 17966 14116 17970 14172
rect 17906 14112 17970 14116
rect 17986 14172 18050 14176
rect 17986 14116 17990 14172
rect 17990 14116 18046 14172
rect 18046 14116 18050 14172
rect 17986 14112 18050 14116
rect 3751 13628 3815 13632
rect 3751 13572 3755 13628
rect 3755 13572 3811 13628
rect 3811 13572 3815 13628
rect 3751 13568 3815 13572
rect 3831 13628 3895 13632
rect 3831 13572 3835 13628
rect 3835 13572 3891 13628
rect 3891 13572 3895 13628
rect 3831 13568 3895 13572
rect 3911 13628 3975 13632
rect 3911 13572 3915 13628
rect 3915 13572 3971 13628
rect 3971 13572 3975 13628
rect 3911 13568 3975 13572
rect 3991 13628 4055 13632
rect 3991 13572 3995 13628
rect 3995 13572 4051 13628
rect 4051 13572 4055 13628
rect 3991 13568 4055 13572
rect 9349 13628 9413 13632
rect 9349 13572 9353 13628
rect 9353 13572 9409 13628
rect 9409 13572 9413 13628
rect 9349 13568 9413 13572
rect 9429 13628 9493 13632
rect 9429 13572 9433 13628
rect 9433 13572 9489 13628
rect 9489 13572 9493 13628
rect 9429 13568 9493 13572
rect 9509 13628 9573 13632
rect 9509 13572 9513 13628
rect 9513 13572 9569 13628
rect 9569 13572 9573 13628
rect 9509 13568 9573 13572
rect 9589 13628 9653 13632
rect 9589 13572 9593 13628
rect 9593 13572 9649 13628
rect 9649 13572 9653 13628
rect 9589 13568 9653 13572
rect 14947 13628 15011 13632
rect 14947 13572 14951 13628
rect 14951 13572 15007 13628
rect 15007 13572 15011 13628
rect 14947 13568 15011 13572
rect 15027 13628 15091 13632
rect 15027 13572 15031 13628
rect 15031 13572 15087 13628
rect 15087 13572 15091 13628
rect 15027 13568 15091 13572
rect 15107 13628 15171 13632
rect 15107 13572 15111 13628
rect 15111 13572 15167 13628
rect 15167 13572 15171 13628
rect 15107 13568 15171 13572
rect 15187 13628 15251 13632
rect 15187 13572 15191 13628
rect 15191 13572 15247 13628
rect 15247 13572 15251 13628
rect 15187 13568 15251 13572
rect 20545 13628 20609 13632
rect 20545 13572 20549 13628
rect 20549 13572 20605 13628
rect 20605 13572 20609 13628
rect 20545 13568 20609 13572
rect 20625 13628 20689 13632
rect 20625 13572 20629 13628
rect 20629 13572 20685 13628
rect 20685 13572 20689 13628
rect 20625 13568 20689 13572
rect 20705 13628 20769 13632
rect 20705 13572 20709 13628
rect 20709 13572 20765 13628
rect 20765 13572 20769 13628
rect 20705 13568 20769 13572
rect 20785 13628 20849 13632
rect 20785 13572 20789 13628
rect 20789 13572 20845 13628
rect 20845 13572 20849 13628
rect 20785 13568 20849 13572
rect 20300 13500 20364 13564
rect 19380 13364 19444 13428
rect 21036 13364 21100 13428
rect 6550 13084 6614 13088
rect 6550 13028 6554 13084
rect 6554 13028 6610 13084
rect 6610 13028 6614 13084
rect 6550 13024 6614 13028
rect 6630 13084 6694 13088
rect 6630 13028 6634 13084
rect 6634 13028 6690 13084
rect 6690 13028 6694 13084
rect 6630 13024 6694 13028
rect 6710 13084 6774 13088
rect 6710 13028 6714 13084
rect 6714 13028 6770 13084
rect 6770 13028 6774 13084
rect 6710 13024 6774 13028
rect 6790 13084 6854 13088
rect 6790 13028 6794 13084
rect 6794 13028 6850 13084
rect 6850 13028 6854 13084
rect 6790 13024 6854 13028
rect 12148 13084 12212 13088
rect 12148 13028 12152 13084
rect 12152 13028 12208 13084
rect 12208 13028 12212 13084
rect 12148 13024 12212 13028
rect 12228 13084 12292 13088
rect 12228 13028 12232 13084
rect 12232 13028 12288 13084
rect 12288 13028 12292 13084
rect 12228 13024 12292 13028
rect 12308 13084 12372 13088
rect 12308 13028 12312 13084
rect 12312 13028 12368 13084
rect 12368 13028 12372 13084
rect 12308 13024 12372 13028
rect 12388 13084 12452 13088
rect 12388 13028 12392 13084
rect 12392 13028 12448 13084
rect 12448 13028 12452 13084
rect 12388 13024 12452 13028
rect 17746 13084 17810 13088
rect 17746 13028 17750 13084
rect 17750 13028 17806 13084
rect 17806 13028 17810 13084
rect 17746 13024 17810 13028
rect 17826 13084 17890 13088
rect 17826 13028 17830 13084
rect 17830 13028 17886 13084
rect 17886 13028 17890 13084
rect 17826 13024 17890 13028
rect 17906 13084 17970 13088
rect 17906 13028 17910 13084
rect 17910 13028 17966 13084
rect 17966 13028 17970 13084
rect 17906 13024 17970 13028
rect 17986 13084 18050 13088
rect 17986 13028 17990 13084
rect 17990 13028 18046 13084
rect 18046 13028 18050 13084
rect 17986 13024 18050 13028
rect 16804 12820 16868 12884
rect 3751 12540 3815 12544
rect 3751 12484 3755 12540
rect 3755 12484 3811 12540
rect 3811 12484 3815 12540
rect 3751 12480 3815 12484
rect 3831 12540 3895 12544
rect 3831 12484 3835 12540
rect 3835 12484 3891 12540
rect 3891 12484 3895 12540
rect 3831 12480 3895 12484
rect 3911 12540 3975 12544
rect 3911 12484 3915 12540
rect 3915 12484 3971 12540
rect 3971 12484 3975 12540
rect 3911 12480 3975 12484
rect 3991 12540 4055 12544
rect 3991 12484 3995 12540
rect 3995 12484 4051 12540
rect 4051 12484 4055 12540
rect 3991 12480 4055 12484
rect 9349 12540 9413 12544
rect 9349 12484 9353 12540
rect 9353 12484 9409 12540
rect 9409 12484 9413 12540
rect 9349 12480 9413 12484
rect 9429 12540 9493 12544
rect 9429 12484 9433 12540
rect 9433 12484 9489 12540
rect 9489 12484 9493 12540
rect 9429 12480 9493 12484
rect 9509 12540 9573 12544
rect 9509 12484 9513 12540
rect 9513 12484 9569 12540
rect 9569 12484 9573 12540
rect 9509 12480 9573 12484
rect 9589 12540 9653 12544
rect 9589 12484 9593 12540
rect 9593 12484 9649 12540
rect 9649 12484 9653 12540
rect 9589 12480 9653 12484
rect 14947 12540 15011 12544
rect 14947 12484 14951 12540
rect 14951 12484 15007 12540
rect 15007 12484 15011 12540
rect 14947 12480 15011 12484
rect 15027 12540 15091 12544
rect 15027 12484 15031 12540
rect 15031 12484 15087 12540
rect 15087 12484 15091 12540
rect 15027 12480 15091 12484
rect 15107 12540 15171 12544
rect 15107 12484 15111 12540
rect 15111 12484 15167 12540
rect 15167 12484 15171 12540
rect 15107 12480 15171 12484
rect 15187 12540 15251 12544
rect 15187 12484 15191 12540
rect 15191 12484 15247 12540
rect 15247 12484 15251 12540
rect 15187 12480 15251 12484
rect 20545 12540 20609 12544
rect 20545 12484 20549 12540
rect 20549 12484 20605 12540
rect 20605 12484 20609 12540
rect 20545 12480 20609 12484
rect 20625 12540 20689 12544
rect 20625 12484 20629 12540
rect 20629 12484 20685 12540
rect 20685 12484 20689 12540
rect 20625 12480 20689 12484
rect 20705 12540 20769 12544
rect 20705 12484 20709 12540
rect 20709 12484 20765 12540
rect 20765 12484 20769 12540
rect 20705 12480 20769 12484
rect 20785 12540 20849 12544
rect 20785 12484 20789 12540
rect 20789 12484 20845 12540
rect 20845 12484 20849 12540
rect 20785 12480 20849 12484
rect 6550 11996 6614 12000
rect 6550 11940 6554 11996
rect 6554 11940 6610 11996
rect 6610 11940 6614 11996
rect 6550 11936 6614 11940
rect 6630 11996 6694 12000
rect 6630 11940 6634 11996
rect 6634 11940 6690 11996
rect 6690 11940 6694 11996
rect 6630 11936 6694 11940
rect 6710 11996 6774 12000
rect 6710 11940 6714 11996
rect 6714 11940 6770 11996
rect 6770 11940 6774 11996
rect 6710 11936 6774 11940
rect 6790 11996 6854 12000
rect 6790 11940 6794 11996
rect 6794 11940 6850 11996
rect 6850 11940 6854 11996
rect 6790 11936 6854 11940
rect 12148 11996 12212 12000
rect 12148 11940 12152 11996
rect 12152 11940 12208 11996
rect 12208 11940 12212 11996
rect 12148 11936 12212 11940
rect 12228 11996 12292 12000
rect 12228 11940 12232 11996
rect 12232 11940 12288 11996
rect 12288 11940 12292 11996
rect 12228 11936 12292 11940
rect 12308 11996 12372 12000
rect 12308 11940 12312 11996
rect 12312 11940 12368 11996
rect 12368 11940 12372 11996
rect 12308 11936 12372 11940
rect 12388 11996 12452 12000
rect 12388 11940 12392 11996
rect 12392 11940 12448 11996
rect 12448 11940 12452 11996
rect 12388 11936 12452 11940
rect 17746 11996 17810 12000
rect 17746 11940 17750 11996
rect 17750 11940 17806 11996
rect 17806 11940 17810 11996
rect 17746 11936 17810 11940
rect 17826 11996 17890 12000
rect 17826 11940 17830 11996
rect 17830 11940 17886 11996
rect 17886 11940 17890 11996
rect 17826 11936 17890 11940
rect 17906 11996 17970 12000
rect 17906 11940 17910 11996
rect 17910 11940 17966 11996
rect 17966 11940 17970 11996
rect 17906 11936 17970 11940
rect 17986 11996 18050 12000
rect 17986 11940 17990 11996
rect 17990 11940 18046 11996
rect 18046 11940 18050 11996
rect 17986 11936 18050 11940
rect 3751 11452 3815 11456
rect 3751 11396 3755 11452
rect 3755 11396 3811 11452
rect 3811 11396 3815 11452
rect 3751 11392 3815 11396
rect 3831 11452 3895 11456
rect 3831 11396 3835 11452
rect 3835 11396 3891 11452
rect 3891 11396 3895 11452
rect 3831 11392 3895 11396
rect 3911 11452 3975 11456
rect 3911 11396 3915 11452
rect 3915 11396 3971 11452
rect 3971 11396 3975 11452
rect 3911 11392 3975 11396
rect 3991 11452 4055 11456
rect 3991 11396 3995 11452
rect 3995 11396 4051 11452
rect 4051 11396 4055 11452
rect 3991 11392 4055 11396
rect 9349 11452 9413 11456
rect 9349 11396 9353 11452
rect 9353 11396 9409 11452
rect 9409 11396 9413 11452
rect 9349 11392 9413 11396
rect 9429 11452 9493 11456
rect 9429 11396 9433 11452
rect 9433 11396 9489 11452
rect 9489 11396 9493 11452
rect 9429 11392 9493 11396
rect 9509 11452 9573 11456
rect 9509 11396 9513 11452
rect 9513 11396 9569 11452
rect 9569 11396 9573 11452
rect 9509 11392 9573 11396
rect 9589 11452 9653 11456
rect 9589 11396 9593 11452
rect 9593 11396 9649 11452
rect 9649 11396 9653 11452
rect 9589 11392 9653 11396
rect 14947 11452 15011 11456
rect 14947 11396 14951 11452
rect 14951 11396 15007 11452
rect 15007 11396 15011 11452
rect 14947 11392 15011 11396
rect 15027 11452 15091 11456
rect 15027 11396 15031 11452
rect 15031 11396 15087 11452
rect 15087 11396 15091 11452
rect 15027 11392 15091 11396
rect 15107 11452 15171 11456
rect 15107 11396 15111 11452
rect 15111 11396 15167 11452
rect 15167 11396 15171 11452
rect 15107 11392 15171 11396
rect 15187 11452 15251 11456
rect 15187 11396 15191 11452
rect 15191 11396 15247 11452
rect 15247 11396 15251 11452
rect 15187 11392 15251 11396
rect 20545 11452 20609 11456
rect 20545 11396 20549 11452
rect 20549 11396 20605 11452
rect 20605 11396 20609 11452
rect 20545 11392 20609 11396
rect 20625 11452 20689 11456
rect 20625 11396 20629 11452
rect 20629 11396 20685 11452
rect 20685 11396 20689 11452
rect 20625 11392 20689 11396
rect 20705 11452 20769 11456
rect 20705 11396 20709 11452
rect 20709 11396 20765 11452
rect 20765 11396 20769 11452
rect 20705 11392 20769 11396
rect 20785 11452 20849 11456
rect 20785 11396 20789 11452
rect 20789 11396 20845 11452
rect 20845 11396 20849 11452
rect 20785 11392 20849 11396
rect 16620 11188 16684 11252
rect 6550 10908 6614 10912
rect 6550 10852 6554 10908
rect 6554 10852 6610 10908
rect 6610 10852 6614 10908
rect 6550 10848 6614 10852
rect 6630 10908 6694 10912
rect 6630 10852 6634 10908
rect 6634 10852 6690 10908
rect 6690 10852 6694 10908
rect 6630 10848 6694 10852
rect 6710 10908 6774 10912
rect 6710 10852 6714 10908
rect 6714 10852 6770 10908
rect 6770 10852 6774 10908
rect 6710 10848 6774 10852
rect 6790 10908 6854 10912
rect 6790 10852 6794 10908
rect 6794 10852 6850 10908
rect 6850 10852 6854 10908
rect 6790 10848 6854 10852
rect 12148 10908 12212 10912
rect 12148 10852 12152 10908
rect 12152 10852 12208 10908
rect 12208 10852 12212 10908
rect 12148 10848 12212 10852
rect 12228 10908 12292 10912
rect 12228 10852 12232 10908
rect 12232 10852 12288 10908
rect 12288 10852 12292 10908
rect 12228 10848 12292 10852
rect 12308 10908 12372 10912
rect 12308 10852 12312 10908
rect 12312 10852 12368 10908
rect 12368 10852 12372 10908
rect 12308 10848 12372 10852
rect 12388 10908 12452 10912
rect 12388 10852 12392 10908
rect 12392 10852 12448 10908
rect 12448 10852 12452 10908
rect 12388 10848 12452 10852
rect 17746 10908 17810 10912
rect 17746 10852 17750 10908
rect 17750 10852 17806 10908
rect 17806 10852 17810 10908
rect 17746 10848 17810 10852
rect 17826 10908 17890 10912
rect 17826 10852 17830 10908
rect 17830 10852 17886 10908
rect 17886 10852 17890 10908
rect 17826 10848 17890 10852
rect 17906 10908 17970 10912
rect 17906 10852 17910 10908
rect 17910 10852 17966 10908
rect 17966 10852 17970 10908
rect 17906 10848 17970 10852
rect 17986 10908 18050 10912
rect 17986 10852 17990 10908
rect 17990 10852 18046 10908
rect 18046 10852 18050 10908
rect 17986 10848 18050 10852
rect 3751 10364 3815 10368
rect 3751 10308 3755 10364
rect 3755 10308 3811 10364
rect 3811 10308 3815 10364
rect 3751 10304 3815 10308
rect 3831 10364 3895 10368
rect 3831 10308 3835 10364
rect 3835 10308 3891 10364
rect 3891 10308 3895 10364
rect 3831 10304 3895 10308
rect 3911 10364 3975 10368
rect 3911 10308 3915 10364
rect 3915 10308 3971 10364
rect 3971 10308 3975 10364
rect 3911 10304 3975 10308
rect 3991 10364 4055 10368
rect 3991 10308 3995 10364
rect 3995 10308 4051 10364
rect 4051 10308 4055 10364
rect 3991 10304 4055 10308
rect 9349 10364 9413 10368
rect 9349 10308 9353 10364
rect 9353 10308 9409 10364
rect 9409 10308 9413 10364
rect 9349 10304 9413 10308
rect 9429 10364 9493 10368
rect 9429 10308 9433 10364
rect 9433 10308 9489 10364
rect 9489 10308 9493 10364
rect 9429 10304 9493 10308
rect 9509 10364 9573 10368
rect 9509 10308 9513 10364
rect 9513 10308 9569 10364
rect 9569 10308 9573 10364
rect 9509 10304 9573 10308
rect 9589 10364 9653 10368
rect 9589 10308 9593 10364
rect 9593 10308 9649 10364
rect 9649 10308 9653 10364
rect 9589 10304 9653 10308
rect 14947 10364 15011 10368
rect 14947 10308 14951 10364
rect 14951 10308 15007 10364
rect 15007 10308 15011 10364
rect 14947 10304 15011 10308
rect 15027 10364 15091 10368
rect 15027 10308 15031 10364
rect 15031 10308 15087 10364
rect 15087 10308 15091 10364
rect 15027 10304 15091 10308
rect 15107 10364 15171 10368
rect 15107 10308 15111 10364
rect 15111 10308 15167 10364
rect 15167 10308 15171 10364
rect 15107 10304 15171 10308
rect 15187 10364 15251 10368
rect 15187 10308 15191 10364
rect 15191 10308 15247 10364
rect 15247 10308 15251 10364
rect 15187 10304 15251 10308
rect 20545 10364 20609 10368
rect 20545 10308 20549 10364
rect 20549 10308 20605 10364
rect 20605 10308 20609 10364
rect 20545 10304 20609 10308
rect 20625 10364 20689 10368
rect 20625 10308 20629 10364
rect 20629 10308 20685 10364
rect 20685 10308 20689 10364
rect 20625 10304 20689 10308
rect 20705 10364 20769 10368
rect 20705 10308 20709 10364
rect 20709 10308 20765 10364
rect 20765 10308 20769 10364
rect 20705 10304 20769 10308
rect 20785 10364 20849 10368
rect 20785 10308 20789 10364
rect 20789 10308 20845 10364
rect 20845 10308 20849 10364
rect 20785 10304 20849 10308
rect 6550 9820 6614 9824
rect 6550 9764 6554 9820
rect 6554 9764 6610 9820
rect 6610 9764 6614 9820
rect 6550 9760 6614 9764
rect 6630 9820 6694 9824
rect 6630 9764 6634 9820
rect 6634 9764 6690 9820
rect 6690 9764 6694 9820
rect 6630 9760 6694 9764
rect 6710 9820 6774 9824
rect 6710 9764 6714 9820
rect 6714 9764 6770 9820
rect 6770 9764 6774 9820
rect 6710 9760 6774 9764
rect 6790 9820 6854 9824
rect 6790 9764 6794 9820
rect 6794 9764 6850 9820
rect 6850 9764 6854 9820
rect 6790 9760 6854 9764
rect 12148 9820 12212 9824
rect 12148 9764 12152 9820
rect 12152 9764 12208 9820
rect 12208 9764 12212 9820
rect 12148 9760 12212 9764
rect 12228 9820 12292 9824
rect 12228 9764 12232 9820
rect 12232 9764 12288 9820
rect 12288 9764 12292 9820
rect 12228 9760 12292 9764
rect 12308 9820 12372 9824
rect 12308 9764 12312 9820
rect 12312 9764 12368 9820
rect 12368 9764 12372 9820
rect 12308 9760 12372 9764
rect 12388 9820 12452 9824
rect 12388 9764 12392 9820
rect 12392 9764 12448 9820
rect 12448 9764 12452 9820
rect 12388 9760 12452 9764
rect 17746 9820 17810 9824
rect 17746 9764 17750 9820
rect 17750 9764 17806 9820
rect 17806 9764 17810 9820
rect 17746 9760 17810 9764
rect 17826 9820 17890 9824
rect 17826 9764 17830 9820
rect 17830 9764 17886 9820
rect 17886 9764 17890 9820
rect 17826 9760 17890 9764
rect 17906 9820 17970 9824
rect 17906 9764 17910 9820
rect 17910 9764 17966 9820
rect 17966 9764 17970 9820
rect 17906 9760 17970 9764
rect 17986 9820 18050 9824
rect 17986 9764 17990 9820
rect 17990 9764 18046 9820
rect 18046 9764 18050 9820
rect 17986 9760 18050 9764
rect 16804 9420 16868 9484
rect 3751 9276 3815 9280
rect 3751 9220 3755 9276
rect 3755 9220 3811 9276
rect 3811 9220 3815 9276
rect 3751 9216 3815 9220
rect 3831 9276 3895 9280
rect 3831 9220 3835 9276
rect 3835 9220 3891 9276
rect 3891 9220 3895 9276
rect 3831 9216 3895 9220
rect 3911 9276 3975 9280
rect 3911 9220 3915 9276
rect 3915 9220 3971 9276
rect 3971 9220 3975 9276
rect 3911 9216 3975 9220
rect 3991 9276 4055 9280
rect 3991 9220 3995 9276
rect 3995 9220 4051 9276
rect 4051 9220 4055 9276
rect 3991 9216 4055 9220
rect 9349 9276 9413 9280
rect 9349 9220 9353 9276
rect 9353 9220 9409 9276
rect 9409 9220 9413 9276
rect 9349 9216 9413 9220
rect 9429 9276 9493 9280
rect 9429 9220 9433 9276
rect 9433 9220 9489 9276
rect 9489 9220 9493 9276
rect 9429 9216 9493 9220
rect 9509 9276 9573 9280
rect 9509 9220 9513 9276
rect 9513 9220 9569 9276
rect 9569 9220 9573 9276
rect 9509 9216 9573 9220
rect 9589 9276 9653 9280
rect 9589 9220 9593 9276
rect 9593 9220 9649 9276
rect 9649 9220 9653 9276
rect 9589 9216 9653 9220
rect 14947 9276 15011 9280
rect 14947 9220 14951 9276
rect 14951 9220 15007 9276
rect 15007 9220 15011 9276
rect 14947 9216 15011 9220
rect 15027 9276 15091 9280
rect 15027 9220 15031 9276
rect 15031 9220 15087 9276
rect 15087 9220 15091 9276
rect 15027 9216 15091 9220
rect 15107 9276 15171 9280
rect 15107 9220 15111 9276
rect 15111 9220 15167 9276
rect 15167 9220 15171 9276
rect 15107 9216 15171 9220
rect 15187 9276 15251 9280
rect 15187 9220 15191 9276
rect 15191 9220 15247 9276
rect 15247 9220 15251 9276
rect 15187 9216 15251 9220
rect 20545 9276 20609 9280
rect 20545 9220 20549 9276
rect 20549 9220 20605 9276
rect 20605 9220 20609 9276
rect 20545 9216 20609 9220
rect 20625 9276 20689 9280
rect 20625 9220 20629 9276
rect 20629 9220 20685 9276
rect 20685 9220 20689 9276
rect 20625 9216 20689 9220
rect 20705 9276 20769 9280
rect 20705 9220 20709 9276
rect 20709 9220 20765 9276
rect 20765 9220 20769 9276
rect 20705 9216 20769 9220
rect 20785 9276 20849 9280
rect 20785 9220 20789 9276
rect 20789 9220 20845 9276
rect 20845 9220 20849 9276
rect 20785 9216 20849 9220
rect 6550 8732 6614 8736
rect 6550 8676 6554 8732
rect 6554 8676 6610 8732
rect 6610 8676 6614 8732
rect 6550 8672 6614 8676
rect 6630 8732 6694 8736
rect 6630 8676 6634 8732
rect 6634 8676 6690 8732
rect 6690 8676 6694 8732
rect 6630 8672 6694 8676
rect 6710 8732 6774 8736
rect 6710 8676 6714 8732
rect 6714 8676 6770 8732
rect 6770 8676 6774 8732
rect 6710 8672 6774 8676
rect 6790 8732 6854 8736
rect 6790 8676 6794 8732
rect 6794 8676 6850 8732
rect 6850 8676 6854 8732
rect 6790 8672 6854 8676
rect 12148 8732 12212 8736
rect 12148 8676 12152 8732
rect 12152 8676 12208 8732
rect 12208 8676 12212 8732
rect 12148 8672 12212 8676
rect 12228 8732 12292 8736
rect 12228 8676 12232 8732
rect 12232 8676 12288 8732
rect 12288 8676 12292 8732
rect 12228 8672 12292 8676
rect 12308 8732 12372 8736
rect 12308 8676 12312 8732
rect 12312 8676 12368 8732
rect 12368 8676 12372 8732
rect 12308 8672 12372 8676
rect 12388 8732 12452 8736
rect 12388 8676 12392 8732
rect 12392 8676 12448 8732
rect 12448 8676 12452 8732
rect 12388 8672 12452 8676
rect 17746 8732 17810 8736
rect 17746 8676 17750 8732
rect 17750 8676 17806 8732
rect 17806 8676 17810 8732
rect 17746 8672 17810 8676
rect 17826 8732 17890 8736
rect 17826 8676 17830 8732
rect 17830 8676 17886 8732
rect 17886 8676 17890 8732
rect 17826 8672 17890 8676
rect 17906 8732 17970 8736
rect 17906 8676 17910 8732
rect 17910 8676 17966 8732
rect 17966 8676 17970 8732
rect 17906 8672 17970 8676
rect 17986 8732 18050 8736
rect 17986 8676 17990 8732
rect 17990 8676 18046 8732
rect 18046 8676 18050 8732
rect 17986 8672 18050 8676
rect 3751 8188 3815 8192
rect 3751 8132 3755 8188
rect 3755 8132 3811 8188
rect 3811 8132 3815 8188
rect 3751 8128 3815 8132
rect 3831 8188 3895 8192
rect 3831 8132 3835 8188
rect 3835 8132 3891 8188
rect 3891 8132 3895 8188
rect 3831 8128 3895 8132
rect 3911 8188 3975 8192
rect 3911 8132 3915 8188
rect 3915 8132 3971 8188
rect 3971 8132 3975 8188
rect 3911 8128 3975 8132
rect 3991 8188 4055 8192
rect 3991 8132 3995 8188
rect 3995 8132 4051 8188
rect 4051 8132 4055 8188
rect 3991 8128 4055 8132
rect 9349 8188 9413 8192
rect 9349 8132 9353 8188
rect 9353 8132 9409 8188
rect 9409 8132 9413 8188
rect 9349 8128 9413 8132
rect 9429 8188 9493 8192
rect 9429 8132 9433 8188
rect 9433 8132 9489 8188
rect 9489 8132 9493 8188
rect 9429 8128 9493 8132
rect 9509 8188 9573 8192
rect 9509 8132 9513 8188
rect 9513 8132 9569 8188
rect 9569 8132 9573 8188
rect 9509 8128 9573 8132
rect 9589 8188 9653 8192
rect 9589 8132 9593 8188
rect 9593 8132 9649 8188
rect 9649 8132 9653 8188
rect 9589 8128 9653 8132
rect 14947 8188 15011 8192
rect 14947 8132 14951 8188
rect 14951 8132 15007 8188
rect 15007 8132 15011 8188
rect 14947 8128 15011 8132
rect 15027 8188 15091 8192
rect 15027 8132 15031 8188
rect 15031 8132 15087 8188
rect 15087 8132 15091 8188
rect 15027 8128 15091 8132
rect 15107 8188 15171 8192
rect 15107 8132 15111 8188
rect 15111 8132 15167 8188
rect 15167 8132 15171 8188
rect 15107 8128 15171 8132
rect 15187 8188 15251 8192
rect 15187 8132 15191 8188
rect 15191 8132 15247 8188
rect 15247 8132 15251 8188
rect 15187 8128 15251 8132
rect 20545 8188 20609 8192
rect 20545 8132 20549 8188
rect 20549 8132 20605 8188
rect 20605 8132 20609 8188
rect 20545 8128 20609 8132
rect 20625 8188 20689 8192
rect 20625 8132 20629 8188
rect 20629 8132 20685 8188
rect 20685 8132 20689 8188
rect 20625 8128 20689 8132
rect 20705 8188 20769 8192
rect 20705 8132 20709 8188
rect 20709 8132 20765 8188
rect 20765 8132 20769 8188
rect 20705 8128 20769 8132
rect 20785 8188 20849 8192
rect 20785 8132 20789 8188
rect 20789 8132 20845 8188
rect 20845 8132 20849 8188
rect 20785 8128 20849 8132
rect 6550 7644 6614 7648
rect 6550 7588 6554 7644
rect 6554 7588 6610 7644
rect 6610 7588 6614 7644
rect 6550 7584 6614 7588
rect 6630 7644 6694 7648
rect 6630 7588 6634 7644
rect 6634 7588 6690 7644
rect 6690 7588 6694 7644
rect 6630 7584 6694 7588
rect 6710 7644 6774 7648
rect 6710 7588 6714 7644
rect 6714 7588 6770 7644
rect 6770 7588 6774 7644
rect 6710 7584 6774 7588
rect 6790 7644 6854 7648
rect 6790 7588 6794 7644
rect 6794 7588 6850 7644
rect 6850 7588 6854 7644
rect 6790 7584 6854 7588
rect 12148 7644 12212 7648
rect 12148 7588 12152 7644
rect 12152 7588 12208 7644
rect 12208 7588 12212 7644
rect 12148 7584 12212 7588
rect 12228 7644 12292 7648
rect 12228 7588 12232 7644
rect 12232 7588 12288 7644
rect 12288 7588 12292 7644
rect 12228 7584 12292 7588
rect 12308 7644 12372 7648
rect 12308 7588 12312 7644
rect 12312 7588 12368 7644
rect 12368 7588 12372 7644
rect 12308 7584 12372 7588
rect 12388 7644 12452 7648
rect 12388 7588 12392 7644
rect 12392 7588 12448 7644
rect 12448 7588 12452 7644
rect 12388 7584 12452 7588
rect 17746 7644 17810 7648
rect 17746 7588 17750 7644
rect 17750 7588 17806 7644
rect 17806 7588 17810 7644
rect 17746 7584 17810 7588
rect 17826 7644 17890 7648
rect 17826 7588 17830 7644
rect 17830 7588 17886 7644
rect 17886 7588 17890 7644
rect 17826 7584 17890 7588
rect 17906 7644 17970 7648
rect 17906 7588 17910 7644
rect 17910 7588 17966 7644
rect 17966 7588 17970 7644
rect 17906 7584 17970 7588
rect 17986 7644 18050 7648
rect 17986 7588 17990 7644
rect 17990 7588 18046 7644
rect 18046 7588 18050 7644
rect 17986 7584 18050 7588
rect 3751 7100 3815 7104
rect 3751 7044 3755 7100
rect 3755 7044 3811 7100
rect 3811 7044 3815 7100
rect 3751 7040 3815 7044
rect 3831 7100 3895 7104
rect 3831 7044 3835 7100
rect 3835 7044 3891 7100
rect 3891 7044 3895 7100
rect 3831 7040 3895 7044
rect 3911 7100 3975 7104
rect 3911 7044 3915 7100
rect 3915 7044 3971 7100
rect 3971 7044 3975 7100
rect 3911 7040 3975 7044
rect 3991 7100 4055 7104
rect 3991 7044 3995 7100
rect 3995 7044 4051 7100
rect 4051 7044 4055 7100
rect 3991 7040 4055 7044
rect 9349 7100 9413 7104
rect 9349 7044 9353 7100
rect 9353 7044 9409 7100
rect 9409 7044 9413 7100
rect 9349 7040 9413 7044
rect 9429 7100 9493 7104
rect 9429 7044 9433 7100
rect 9433 7044 9489 7100
rect 9489 7044 9493 7100
rect 9429 7040 9493 7044
rect 9509 7100 9573 7104
rect 9509 7044 9513 7100
rect 9513 7044 9569 7100
rect 9569 7044 9573 7100
rect 9509 7040 9573 7044
rect 9589 7100 9653 7104
rect 9589 7044 9593 7100
rect 9593 7044 9649 7100
rect 9649 7044 9653 7100
rect 9589 7040 9653 7044
rect 14947 7100 15011 7104
rect 14947 7044 14951 7100
rect 14951 7044 15007 7100
rect 15007 7044 15011 7100
rect 14947 7040 15011 7044
rect 15027 7100 15091 7104
rect 15027 7044 15031 7100
rect 15031 7044 15087 7100
rect 15087 7044 15091 7100
rect 15027 7040 15091 7044
rect 15107 7100 15171 7104
rect 15107 7044 15111 7100
rect 15111 7044 15167 7100
rect 15167 7044 15171 7100
rect 15107 7040 15171 7044
rect 15187 7100 15251 7104
rect 15187 7044 15191 7100
rect 15191 7044 15247 7100
rect 15247 7044 15251 7100
rect 15187 7040 15251 7044
rect 20545 7100 20609 7104
rect 20545 7044 20549 7100
rect 20549 7044 20605 7100
rect 20605 7044 20609 7100
rect 20545 7040 20609 7044
rect 20625 7100 20689 7104
rect 20625 7044 20629 7100
rect 20629 7044 20685 7100
rect 20685 7044 20689 7100
rect 20625 7040 20689 7044
rect 20705 7100 20769 7104
rect 20705 7044 20709 7100
rect 20709 7044 20765 7100
rect 20765 7044 20769 7100
rect 20705 7040 20769 7044
rect 20785 7100 20849 7104
rect 20785 7044 20789 7100
rect 20789 7044 20845 7100
rect 20845 7044 20849 7100
rect 20785 7040 20849 7044
rect 6550 6556 6614 6560
rect 6550 6500 6554 6556
rect 6554 6500 6610 6556
rect 6610 6500 6614 6556
rect 6550 6496 6614 6500
rect 6630 6556 6694 6560
rect 6630 6500 6634 6556
rect 6634 6500 6690 6556
rect 6690 6500 6694 6556
rect 6630 6496 6694 6500
rect 6710 6556 6774 6560
rect 6710 6500 6714 6556
rect 6714 6500 6770 6556
rect 6770 6500 6774 6556
rect 6710 6496 6774 6500
rect 6790 6556 6854 6560
rect 6790 6500 6794 6556
rect 6794 6500 6850 6556
rect 6850 6500 6854 6556
rect 6790 6496 6854 6500
rect 12148 6556 12212 6560
rect 12148 6500 12152 6556
rect 12152 6500 12208 6556
rect 12208 6500 12212 6556
rect 12148 6496 12212 6500
rect 12228 6556 12292 6560
rect 12228 6500 12232 6556
rect 12232 6500 12288 6556
rect 12288 6500 12292 6556
rect 12228 6496 12292 6500
rect 12308 6556 12372 6560
rect 12308 6500 12312 6556
rect 12312 6500 12368 6556
rect 12368 6500 12372 6556
rect 12308 6496 12372 6500
rect 12388 6556 12452 6560
rect 12388 6500 12392 6556
rect 12392 6500 12448 6556
rect 12448 6500 12452 6556
rect 12388 6496 12452 6500
rect 17746 6556 17810 6560
rect 17746 6500 17750 6556
rect 17750 6500 17806 6556
rect 17806 6500 17810 6556
rect 17746 6496 17810 6500
rect 17826 6556 17890 6560
rect 17826 6500 17830 6556
rect 17830 6500 17886 6556
rect 17886 6500 17890 6556
rect 17826 6496 17890 6500
rect 17906 6556 17970 6560
rect 17906 6500 17910 6556
rect 17910 6500 17966 6556
rect 17966 6500 17970 6556
rect 17906 6496 17970 6500
rect 17986 6556 18050 6560
rect 17986 6500 17990 6556
rect 17990 6500 18046 6556
rect 18046 6500 18050 6556
rect 17986 6496 18050 6500
rect 3751 6012 3815 6016
rect 3751 5956 3755 6012
rect 3755 5956 3811 6012
rect 3811 5956 3815 6012
rect 3751 5952 3815 5956
rect 3831 6012 3895 6016
rect 3831 5956 3835 6012
rect 3835 5956 3891 6012
rect 3891 5956 3895 6012
rect 3831 5952 3895 5956
rect 3911 6012 3975 6016
rect 3911 5956 3915 6012
rect 3915 5956 3971 6012
rect 3971 5956 3975 6012
rect 3911 5952 3975 5956
rect 3991 6012 4055 6016
rect 3991 5956 3995 6012
rect 3995 5956 4051 6012
rect 4051 5956 4055 6012
rect 3991 5952 4055 5956
rect 9349 6012 9413 6016
rect 9349 5956 9353 6012
rect 9353 5956 9409 6012
rect 9409 5956 9413 6012
rect 9349 5952 9413 5956
rect 9429 6012 9493 6016
rect 9429 5956 9433 6012
rect 9433 5956 9489 6012
rect 9489 5956 9493 6012
rect 9429 5952 9493 5956
rect 9509 6012 9573 6016
rect 9509 5956 9513 6012
rect 9513 5956 9569 6012
rect 9569 5956 9573 6012
rect 9509 5952 9573 5956
rect 9589 6012 9653 6016
rect 9589 5956 9593 6012
rect 9593 5956 9649 6012
rect 9649 5956 9653 6012
rect 9589 5952 9653 5956
rect 14947 6012 15011 6016
rect 14947 5956 14951 6012
rect 14951 5956 15007 6012
rect 15007 5956 15011 6012
rect 14947 5952 15011 5956
rect 15027 6012 15091 6016
rect 15027 5956 15031 6012
rect 15031 5956 15087 6012
rect 15087 5956 15091 6012
rect 15027 5952 15091 5956
rect 15107 6012 15171 6016
rect 15107 5956 15111 6012
rect 15111 5956 15167 6012
rect 15167 5956 15171 6012
rect 15107 5952 15171 5956
rect 15187 6012 15251 6016
rect 15187 5956 15191 6012
rect 15191 5956 15247 6012
rect 15247 5956 15251 6012
rect 15187 5952 15251 5956
rect 20545 6012 20609 6016
rect 20545 5956 20549 6012
rect 20549 5956 20605 6012
rect 20605 5956 20609 6012
rect 20545 5952 20609 5956
rect 20625 6012 20689 6016
rect 20625 5956 20629 6012
rect 20629 5956 20685 6012
rect 20685 5956 20689 6012
rect 20625 5952 20689 5956
rect 20705 6012 20769 6016
rect 20705 5956 20709 6012
rect 20709 5956 20765 6012
rect 20765 5956 20769 6012
rect 20705 5952 20769 5956
rect 20785 6012 20849 6016
rect 20785 5956 20789 6012
rect 20789 5956 20845 6012
rect 20845 5956 20849 6012
rect 20785 5952 20849 5956
rect 16620 5944 16684 5948
rect 16620 5888 16670 5944
rect 16670 5888 16684 5944
rect 16620 5884 16684 5888
rect 6550 5468 6614 5472
rect 6550 5412 6554 5468
rect 6554 5412 6610 5468
rect 6610 5412 6614 5468
rect 6550 5408 6614 5412
rect 6630 5468 6694 5472
rect 6630 5412 6634 5468
rect 6634 5412 6690 5468
rect 6690 5412 6694 5468
rect 6630 5408 6694 5412
rect 6710 5468 6774 5472
rect 6710 5412 6714 5468
rect 6714 5412 6770 5468
rect 6770 5412 6774 5468
rect 6710 5408 6774 5412
rect 6790 5468 6854 5472
rect 6790 5412 6794 5468
rect 6794 5412 6850 5468
rect 6850 5412 6854 5468
rect 6790 5408 6854 5412
rect 12148 5468 12212 5472
rect 12148 5412 12152 5468
rect 12152 5412 12208 5468
rect 12208 5412 12212 5468
rect 12148 5408 12212 5412
rect 12228 5468 12292 5472
rect 12228 5412 12232 5468
rect 12232 5412 12288 5468
rect 12288 5412 12292 5468
rect 12228 5408 12292 5412
rect 12308 5468 12372 5472
rect 12308 5412 12312 5468
rect 12312 5412 12368 5468
rect 12368 5412 12372 5468
rect 12308 5408 12372 5412
rect 12388 5468 12452 5472
rect 12388 5412 12392 5468
rect 12392 5412 12448 5468
rect 12448 5412 12452 5468
rect 12388 5408 12452 5412
rect 17746 5468 17810 5472
rect 17746 5412 17750 5468
rect 17750 5412 17806 5468
rect 17806 5412 17810 5468
rect 17746 5408 17810 5412
rect 17826 5468 17890 5472
rect 17826 5412 17830 5468
rect 17830 5412 17886 5468
rect 17886 5412 17890 5468
rect 17826 5408 17890 5412
rect 17906 5468 17970 5472
rect 17906 5412 17910 5468
rect 17910 5412 17966 5468
rect 17966 5412 17970 5468
rect 17906 5408 17970 5412
rect 17986 5468 18050 5472
rect 17986 5412 17990 5468
rect 17990 5412 18046 5468
rect 18046 5412 18050 5468
rect 17986 5408 18050 5412
rect 3751 4924 3815 4928
rect 3751 4868 3755 4924
rect 3755 4868 3811 4924
rect 3811 4868 3815 4924
rect 3751 4864 3815 4868
rect 3831 4924 3895 4928
rect 3831 4868 3835 4924
rect 3835 4868 3891 4924
rect 3891 4868 3895 4924
rect 3831 4864 3895 4868
rect 3911 4924 3975 4928
rect 3911 4868 3915 4924
rect 3915 4868 3971 4924
rect 3971 4868 3975 4924
rect 3911 4864 3975 4868
rect 3991 4924 4055 4928
rect 3991 4868 3995 4924
rect 3995 4868 4051 4924
rect 4051 4868 4055 4924
rect 3991 4864 4055 4868
rect 9349 4924 9413 4928
rect 9349 4868 9353 4924
rect 9353 4868 9409 4924
rect 9409 4868 9413 4924
rect 9349 4864 9413 4868
rect 9429 4924 9493 4928
rect 9429 4868 9433 4924
rect 9433 4868 9489 4924
rect 9489 4868 9493 4924
rect 9429 4864 9493 4868
rect 9509 4924 9573 4928
rect 9509 4868 9513 4924
rect 9513 4868 9569 4924
rect 9569 4868 9573 4924
rect 9509 4864 9573 4868
rect 9589 4924 9653 4928
rect 9589 4868 9593 4924
rect 9593 4868 9649 4924
rect 9649 4868 9653 4924
rect 9589 4864 9653 4868
rect 14947 4924 15011 4928
rect 14947 4868 14951 4924
rect 14951 4868 15007 4924
rect 15007 4868 15011 4924
rect 14947 4864 15011 4868
rect 15027 4924 15091 4928
rect 15027 4868 15031 4924
rect 15031 4868 15087 4924
rect 15087 4868 15091 4924
rect 15027 4864 15091 4868
rect 15107 4924 15171 4928
rect 15107 4868 15111 4924
rect 15111 4868 15167 4924
rect 15167 4868 15171 4924
rect 15107 4864 15171 4868
rect 15187 4924 15251 4928
rect 15187 4868 15191 4924
rect 15191 4868 15247 4924
rect 15247 4868 15251 4924
rect 15187 4864 15251 4868
rect 20545 4924 20609 4928
rect 20545 4868 20549 4924
rect 20549 4868 20605 4924
rect 20605 4868 20609 4924
rect 20545 4864 20609 4868
rect 20625 4924 20689 4928
rect 20625 4868 20629 4924
rect 20629 4868 20685 4924
rect 20685 4868 20689 4924
rect 20625 4864 20689 4868
rect 20705 4924 20769 4928
rect 20705 4868 20709 4924
rect 20709 4868 20765 4924
rect 20765 4868 20769 4924
rect 20705 4864 20769 4868
rect 20785 4924 20849 4928
rect 20785 4868 20789 4924
rect 20789 4868 20845 4924
rect 20845 4868 20849 4924
rect 20785 4864 20849 4868
rect 6550 4380 6614 4384
rect 6550 4324 6554 4380
rect 6554 4324 6610 4380
rect 6610 4324 6614 4380
rect 6550 4320 6614 4324
rect 6630 4380 6694 4384
rect 6630 4324 6634 4380
rect 6634 4324 6690 4380
rect 6690 4324 6694 4380
rect 6630 4320 6694 4324
rect 6710 4380 6774 4384
rect 6710 4324 6714 4380
rect 6714 4324 6770 4380
rect 6770 4324 6774 4380
rect 6710 4320 6774 4324
rect 6790 4380 6854 4384
rect 6790 4324 6794 4380
rect 6794 4324 6850 4380
rect 6850 4324 6854 4380
rect 6790 4320 6854 4324
rect 12148 4380 12212 4384
rect 12148 4324 12152 4380
rect 12152 4324 12208 4380
rect 12208 4324 12212 4380
rect 12148 4320 12212 4324
rect 12228 4380 12292 4384
rect 12228 4324 12232 4380
rect 12232 4324 12288 4380
rect 12288 4324 12292 4380
rect 12228 4320 12292 4324
rect 12308 4380 12372 4384
rect 12308 4324 12312 4380
rect 12312 4324 12368 4380
rect 12368 4324 12372 4380
rect 12308 4320 12372 4324
rect 12388 4380 12452 4384
rect 12388 4324 12392 4380
rect 12392 4324 12448 4380
rect 12448 4324 12452 4380
rect 12388 4320 12452 4324
rect 17746 4380 17810 4384
rect 17746 4324 17750 4380
rect 17750 4324 17806 4380
rect 17806 4324 17810 4380
rect 17746 4320 17810 4324
rect 17826 4380 17890 4384
rect 17826 4324 17830 4380
rect 17830 4324 17886 4380
rect 17886 4324 17890 4380
rect 17826 4320 17890 4324
rect 17906 4380 17970 4384
rect 17906 4324 17910 4380
rect 17910 4324 17966 4380
rect 17966 4324 17970 4380
rect 17906 4320 17970 4324
rect 17986 4380 18050 4384
rect 17986 4324 17990 4380
rect 17990 4324 18046 4380
rect 18046 4324 18050 4380
rect 17986 4320 18050 4324
rect 3751 3836 3815 3840
rect 3751 3780 3755 3836
rect 3755 3780 3811 3836
rect 3811 3780 3815 3836
rect 3751 3776 3815 3780
rect 3831 3836 3895 3840
rect 3831 3780 3835 3836
rect 3835 3780 3891 3836
rect 3891 3780 3895 3836
rect 3831 3776 3895 3780
rect 3911 3836 3975 3840
rect 3911 3780 3915 3836
rect 3915 3780 3971 3836
rect 3971 3780 3975 3836
rect 3911 3776 3975 3780
rect 3991 3836 4055 3840
rect 3991 3780 3995 3836
rect 3995 3780 4051 3836
rect 4051 3780 4055 3836
rect 3991 3776 4055 3780
rect 9349 3836 9413 3840
rect 9349 3780 9353 3836
rect 9353 3780 9409 3836
rect 9409 3780 9413 3836
rect 9349 3776 9413 3780
rect 9429 3836 9493 3840
rect 9429 3780 9433 3836
rect 9433 3780 9489 3836
rect 9489 3780 9493 3836
rect 9429 3776 9493 3780
rect 9509 3836 9573 3840
rect 9509 3780 9513 3836
rect 9513 3780 9569 3836
rect 9569 3780 9573 3836
rect 9509 3776 9573 3780
rect 9589 3836 9653 3840
rect 9589 3780 9593 3836
rect 9593 3780 9649 3836
rect 9649 3780 9653 3836
rect 9589 3776 9653 3780
rect 14947 3836 15011 3840
rect 14947 3780 14951 3836
rect 14951 3780 15007 3836
rect 15007 3780 15011 3836
rect 14947 3776 15011 3780
rect 15027 3836 15091 3840
rect 15027 3780 15031 3836
rect 15031 3780 15087 3836
rect 15087 3780 15091 3836
rect 15027 3776 15091 3780
rect 15107 3836 15171 3840
rect 15107 3780 15111 3836
rect 15111 3780 15167 3836
rect 15167 3780 15171 3836
rect 15107 3776 15171 3780
rect 15187 3836 15251 3840
rect 15187 3780 15191 3836
rect 15191 3780 15247 3836
rect 15247 3780 15251 3836
rect 15187 3776 15251 3780
rect 20545 3836 20609 3840
rect 20545 3780 20549 3836
rect 20549 3780 20605 3836
rect 20605 3780 20609 3836
rect 20545 3776 20609 3780
rect 20625 3836 20689 3840
rect 20625 3780 20629 3836
rect 20629 3780 20685 3836
rect 20685 3780 20689 3836
rect 20625 3776 20689 3780
rect 20705 3836 20769 3840
rect 20705 3780 20709 3836
rect 20709 3780 20765 3836
rect 20765 3780 20769 3836
rect 20705 3776 20769 3780
rect 20785 3836 20849 3840
rect 20785 3780 20789 3836
rect 20789 3780 20845 3836
rect 20845 3780 20849 3836
rect 20785 3776 20849 3780
rect 6550 3292 6614 3296
rect 6550 3236 6554 3292
rect 6554 3236 6610 3292
rect 6610 3236 6614 3292
rect 6550 3232 6614 3236
rect 6630 3292 6694 3296
rect 6630 3236 6634 3292
rect 6634 3236 6690 3292
rect 6690 3236 6694 3292
rect 6630 3232 6694 3236
rect 6710 3292 6774 3296
rect 6710 3236 6714 3292
rect 6714 3236 6770 3292
rect 6770 3236 6774 3292
rect 6710 3232 6774 3236
rect 6790 3292 6854 3296
rect 6790 3236 6794 3292
rect 6794 3236 6850 3292
rect 6850 3236 6854 3292
rect 6790 3232 6854 3236
rect 12148 3292 12212 3296
rect 12148 3236 12152 3292
rect 12152 3236 12208 3292
rect 12208 3236 12212 3292
rect 12148 3232 12212 3236
rect 12228 3292 12292 3296
rect 12228 3236 12232 3292
rect 12232 3236 12288 3292
rect 12288 3236 12292 3292
rect 12228 3232 12292 3236
rect 12308 3292 12372 3296
rect 12308 3236 12312 3292
rect 12312 3236 12368 3292
rect 12368 3236 12372 3292
rect 12308 3232 12372 3236
rect 12388 3292 12452 3296
rect 12388 3236 12392 3292
rect 12392 3236 12448 3292
rect 12448 3236 12452 3292
rect 12388 3232 12452 3236
rect 17746 3292 17810 3296
rect 17746 3236 17750 3292
rect 17750 3236 17806 3292
rect 17806 3236 17810 3292
rect 17746 3232 17810 3236
rect 17826 3292 17890 3296
rect 17826 3236 17830 3292
rect 17830 3236 17886 3292
rect 17886 3236 17890 3292
rect 17826 3232 17890 3236
rect 17906 3292 17970 3296
rect 17906 3236 17910 3292
rect 17910 3236 17966 3292
rect 17966 3236 17970 3292
rect 17906 3232 17970 3236
rect 17986 3292 18050 3296
rect 17986 3236 17990 3292
rect 17990 3236 18046 3292
rect 18046 3236 18050 3292
rect 17986 3232 18050 3236
rect 3751 2748 3815 2752
rect 3751 2692 3755 2748
rect 3755 2692 3811 2748
rect 3811 2692 3815 2748
rect 3751 2688 3815 2692
rect 3831 2748 3895 2752
rect 3831 2692 3835 2748
rect 3835 2692 3891 2748
rect 3891 2692 3895 2748
rect 3831 2688 3895 2692
rect 3911 2748 3975 2752
rect 3911 2692 3915 2748
rect 3915 2692 3971 2748
rect 3971 2692 3975 2748
rect 3911 2688 3975 2692
rect 3991 2748 4055 2752
rect 3991 2692 3995 2748
rect 3995 2692 4051 2748
rect 4051 2692 4055 2748
rect 3991 2688 4055 2692
rect 9349 2748 9413 2752
rect 9349 2692 9353 2748
rect 9353 2692 9409 2748
rect 9409 2692 9413 2748
rect 9349 2688 9413 2692
rect 9429 2748 9493 2752
rect 9429 2692 9433 2748
rect 9433 2692 9489 2748
rect 9489 2692 9493 2748
rect 9429 2688 9493 2692
rect 9509 2748 9573 2752
rect 9509 2692 9513 2748
rect 9513 2692 9569 2748
rect 9569 2692 9573 2748
rect 9509 2688 9573 2692
rect 9589 2748 9653 2752
rect 9589 2692 9593 2748
rect 9593 2692 9649 2748
rect 9649 2692 9653 2748
rect 9589 2688 9653 2692
rect 14947 2748 15011 2752
rect 14947 2692 14951 2748
rect 14951 2692 15007 2748
rect 15007 2692 15011 2748
rect 14947 2688 15011 2692
rect 15027 2748 15091 2752
rect 15027 2692 15031 2748
rect 15031 2692 15087 2748
rect 15087 2692 15091 2748
rect 15027 2688 15091 2692
rect 15107 2748 15171 2752
rect 15107 2692 15111 2748
rect 15111 2692 15167 2748
rect 15167 2692 15171 2748
rect 15107 2688 15171 2692
rect 15187 2748 15251 2752
rect 15187 2692 15191 2748
rect 15191 2692 15247 2748
rect 15247 2692 15251 2748
rect 15187 2688 15251 2692
rect 20545 2748 20609 2752
rect 20545 2692 20549 2748
rect 20549 2692 20605 2748
rect 20605 2692 20609 2748
rect 20545 2688 20609 2692
rect 20625 2748 20689 2752
rect 20625 2692 20629 2748
rect 20629 2692 20685 2748
rect 20685 2692 20689 2748
rect 20625 2688 20689 2692
rect 20705 2748 20769 2752
rect 20705 2692 20709 2748
rect 20709 2692 20765 2748
rect 20765 2692 20769 2748
rect 20705 2688 20769 2692
rect 20785 2748 20849 2752
rect 20785 2692 20789 2748
rect 20789 2692 20845 2748
rect 20845 2692 20849 2748
rect 20785 2688 20849 2692
rect 16620 2484 16684 2548
rect 6550 2204 6614 2208
rect 6550 2148 6554 2204
rect 6554 2148 6610 2204
rect 6610 2148 6614 2204
rect 6550 2144 6614 2148
rect 6630 2204 6694 2208
rect 6630 2148 6634 2204
rect 6634 2148 6690 2204
rect 6690 2148 6694 2204
rect 6630 2144 6694 2148
rect 6710 2204 6774 2208
rect 6710 2148 6714 2204
rect 6714 2148 6770 2204
rect 6770 2148 6774 2204
rect 6710 2144 6774 2148
rect 6790 2204 6854 2208
rect 6790 2148 6794 2204
rect 6794 2148 6850 2204
rect 6850 2148 6854 2204
rect 6790 2144 6854 2148
rect 12148 2204 12212 2208
rect 12148 2148 12152 2204
rect 12152 2148 12208 2204
rect 12208 2148 12212 2204
rect 12148 2144 12212 2148
rect 12228 2204 12292 2208
rect 12228 2148 12232 2204
rect 12232 2148 12288 2204
rect 12288 2148 12292 2204
rect 12228 2144 12292 2148
rect 12308 2204 12372 2208
rect 12308 2148 12312 2204
rect 12312 2148 12368 2204
rect 12368 2148 12372 2204
rect 12308 2144 12372 2148
rect 12388 2204 12452 2208
rect 12388 2148 12392 2204
rect 12392 2148 12448 2204
rect 12448 2148 12452 2204
rect 12388 2144 12452 2148
rect 17746 2204 17810 2208
rect 17746 2148 17750 2204
rect 17750 2148 17806 2204
rect 17806 2148 17810 2204
rect 17746 2144 17810 2148
rect 17826 2204 17890 2208
rect 17826 2148 17830 2204
rect 17830 2148 17886 2204
rect 17886 2148 17890 2204
rect 17826 2144 17890 2148
rect 17906 2204 17970 2208
rect 17906 2148 17910 2204
rect 17910 2148 17966 2204
rect 17966 2148 17970 2204
rect 17906 2144 17970 2148
rect 17986 2204 18050 2208
rect 17986 2148 17990 2204
rect 17990 2148 18046 2204
rect 18046 2148 18050 2204
rect 17986 2144 18050 2148
<< metal4 >>
rect 3743 22336 4063 22352
rect 3743 22272 3751 22336
rect 3815 22272 3831 22336
rect 3895 22272 3911 22336
rect 3975 22272 3991 22336
rect 4055 22272 4063 22336
rect 3743 21248 4063 22272
rect 3743 21184 3751 21248
rect 3815 21184 3831 21248
rect 3895 21184 3911 21248
rect 3975 21184 3991 21248
rect 4055 21184 4063 21248
rect 3743 20160 4063 21184
rect 3743 20096 3751 20160
rect 3815 20096 3831 20160
rect 3895 20096 3911 20160
rect 3975 20096 3991 20160
rect 4055 20096 4063 20160
rect 3743 19072 4063 20096
rect 3743 19008 3751 19072
rect 3815 19008 3831 19072
rect 3895 19008 3911 19072
rect 3975 19008 3991 19072
rect 4055 19008 4063 19072
rect 3743 17984 4063 19008
rect 3743 17920 3751 17984
rect 3815 17920 3831 17984
rect 3895 17920 3911 17984
rect 3975 17920 3991 17984
rect 4055 17920 4063 17984
rect 3743 16896 4063 17920
rect 3743 16832 3751 16896
rect 3815 16832 3831 16896
rect 3895 16832 3911 16896
rect 3975 16832 3991 16896
rect 4055 16832 4063 16896
rect 3743 15808 4063 16832
rect 3743 15744 3751 15808
rect 3815 15744 3831 15808
rect 3895 15744 3911 15808
rect 3975 15744 3991 15808
rect 4055 15744 4063 15808
rect 3743 14720 4063 15744
rect 3743 14656 3751 14720
rect 3815 14656 3831 14720
rect 3895 14656 3911 14720
rect 3975 14656 3991 14720
rect 4055 14656 4063 14720
rect 3743 13632 4063 14656
rect 3743 13568 3751 13632
rect 3815 13568 3831 13632
rect 3895 13568 3911 13632
rect 3975 13568 3991 13632
rect 4055 13568 4063 13632
rect 3743 12544 4063 13568
rect 3743 12480 3751 12544
rect 3815 12480 3831 12544
rect 3895 12480 3911 12544
rect 3975 12480 3991 12544
rect 4055 12480 4063 12544
rect 3743 11456 4063 12480
rect 3743 11392 3751 11456
rect 3815 11392 3831 11456
rect 3895 11392 3911 11456
rect 3975 11392 3991 11456
rect 4055 11392 4063 11456
rect 3743 10368 4063 11392
rect 3743 10304 3751 10368
rect 3815 10304 3831 10368
rect 3895 10304 3911 10368
rect 3975 10304 3991 10368
rect 4055 10304 4063 10368
rect 3743 9280 4063 10304
rect 3743 9216 3751 9280
rect 3815 9216 3831 9280
rect 3895 9216 3911 9280
rect 3975 9216 3991 9280
rect 4055 9216 4063 9280
rect 3743 8192 4063 9216
rect 3743 8128 3751 8192
rect 3815 8128 3831 8192
rect 3895 8128 3911 8192
rect 3975 8128 3991 8192
rect 4055 8128 4063 8192
rect 3743 7104 4063 8128
rect 3743 7040 3751 7104
rect 3815 7040 3831 7104
rect 3895 7040 3911 7104
rect 3975 7040 3991 7104
rect 4055 7040 4063 7104
rect 3743 6016 4063 7040
rect 3743 5952 3751 6016
rect 3815 5952 3831 6016
rect 3895 5952 3911 6016
rect 3975 5952 3991 6016
rect 4055 5952 4063 6016
rect 3743 4928 4063 5952
rect 3743 4864 3751 4928
rect 3815 4864 3831 4928
rect 3895 4864 3911 4928
rect 3975 4864 3991 4928
rect 4055 4864 4063 4928
rect 3743 3840 4063 4864
rect 3743 3776 3751 3840
rect 3815 3776 3831 3840
rect 3895 3776 3911 3840
rect 3975 3776 3991 3840
rect 4055 3776 4063 3840
rect 3743 2752 4063 3776
rect 3743 2688 3751 2752
rect 3815 2688 3831 2752
rect 3895 2688 3911 2752
rect 3975 2688 3991 2752
rect 4055 2688 4063 2752
rect 3743 2128 4063 2688
rect 6542 21792 6862 22352
rect 9341 22336 9661 22352
rect 9341 22272 9349 22336
rect 9413 22272 9429 22336
rect 9493 22272 9509 22336
rect 9573 22272 9589 22336
rect 9653 22272 9661 22336
rect 9075 21996 9141 21997
rect 9075 21932 9076 21996
rect 9140 21932 9141 21996
rect 9075 21931 9141 21932
rect 6542 21728 6550 21792
rect 6614 21728 6630 21792
rect 6694 21728 6710 21792
rect 6774 21728 6790 21792
rect 6854 21728 6862 21792
rect 6542 20704 6862 21728
rect 6542 20640 6550 20704
rect 6614 20640 6630 20704
rect 6694 20640 6710 20704
rect 6774 20640 6790 20704
rect 6854 20640 6862 20704
rect 6542 19616 6862 20640
rect 6542 19552 6550 19616
rect 6614 19552 6630 19616
rect 6694 19552 6710 19616
rect 6774 19552 6790 19616
rect 6854 19552 6862 19616
rect 6542 18528 6862 19552
rect 6542 18464 6550 18528
rect 6614 18464 6630 18528
rect 6694 18464 6710 18528
rect 6774 18464 6790 18528
rect 6854 18464 6862 18528
rect 6542 17440 6862 18464
rect 6542 17376 6550 17440
rect 6614 17376 6630 17440
rect 6694 17376 6710 17440
rect 6774 17376 6790 17440
rect 6854 17376 6862 17440
rect 6542 16352 6862 17376
rect 9078 17101 9138 21931
rect 9341 21248 9661 22272
rect 9341 21184 9349 21248
rect 9413 21184 9429 21248
rect 9493 21184 9509 21248
rect 9573 21184 9589 21248
rect 9653 21184 9661 21248
rect 9341 20160 9661 21184
rect 9341 20096 9349 20160
rect 9413 20096 9429 20160
rect 9493 20096 9509 20160
rect 9573 20096 9589 20160
rect 9653 20096 9661 20160
rect 9341 19072 9661 20096
rect 9341 19008 9349 19072
rect 9413 19008 9429 19072
rect 9493 19008 9509 19072
rect 9573 19008 9589 19072
rect 9653 19008 9661 19072
rect 9341 17984 9661 19008
rect 9341 17920 9349 17984
rect 9413 17920 9429 17984
rect 9493 17920 9509 17984
rect 9573 17920 9589 17984
rect 9653 17920 9661 17984
rect 9075 17100 9141 17101
rect 9075 17036 9076 17100
rect 9140 17036 9141 17100
rect 9075 17035 9141 17036
rect 6542 16288 6550 16352
rect 6614 16288 6630 16352
rect 6694 16288 6710 16352
rect 6774 16288 6790 16352
rect 6854 16288 6862 16352
rect 6542 15264 6862 16288
rect 6542 15200 6550 15264
rect 6614 15200 6630 15264
rect 6694 15200 6710 15264
rect 6774 15200 6790 15264
rect 6854 15200 6862 15264
rect 6542 14176 6862 15200
rect 6542 14112 6550 14176
rect 6614 14112 6630 14176
rect 6694 14112 6710 14176
rect 6774 14112 6790 14176
rect 6854 14112 6862 14176
rect 6542 13088 6862 14112
rect 6542 13024 6550 13088
rect 6614 13024 6630 13088
rect 6694 13024 6710 13088
rect 6774 13024 6790 13088
rect 6854 13024 6862 13088
rect 6542 12000 6862 13024
rect 6542 11936 6550 12000
rect 6614 11936 6630 12000
rect 6694 11936 6710 12000
rect 6774 11936 6790 12000
rect 6854 11936 6862 12000
rect 6542 10912 6862 11936
rect 6542 10848 6550 10912
rect 6614 10848 6630 10912
rect 6694 10848 6710 10912
rect 6774 10848 6790 10912
rect 6854 10848 6862 10912
rect 6542 9824 6862 10848
rect 6542 9760 6550 9824
rect 6614 9760 6630 9824
rect 6694 9760 6710 9824
rect 6774 9760 6790 9824
rect 6854 9760 6862 9824
rect 6542 8736 6862 9760
rect 6542 8672 6550 8736
rect 6614 8672 6630 8736
rect 6694 8672 6710 8736
rect 6774 8672 6790 8736
rect 6854 8672 6862 8736
rect 6542 7648 6862 8672
rect 6542 7584 6550 7648
rect 6614 7584 6630 7648
rect 6694 7584 6710 7648
rect 6774 7584 6790 7648
rect 6854 7584 6862 7648
rect 6542 6560 6862 7584
rect 6542 6496 6550 6560
rect 6614 6496 6630 6560
rect 6694 6496 6710 6560
rect 6774 6496 6790 6560
rect 6854 6496 6862 6560
rect 6542 5472 6862 6496
rect 6542 5408 6550 5472
rect 6614 5408 6630 5472
rect 6694 5408 6710 5472
rect 6774 5408 6790 5472
rect 6854 5408 6862 5472
rect 6542 4384 6862 5408
rect 6542 4320 6550 4384
rect 6614 4320 6630 4384
rect 6694 4320 6710 4384
rect 6774 4320 6790 4384
rect 6854 4320 6862 4384
rect 6542 3296 6862 4320
rect 6542 3232 6550 3296
rect 6614 3232 6630 3296
rect 6694 3232 6710 3296
rect 6774 3232 6790 3296
rect 6854 3232 6862 3296
rect 6542 2208 6862 3232
rect 6542 2144 6550 2208
rect 6614 2144 6630 2208
rect 6694 2144 6710 2208
rect 6774 2144 6790 2208
rect 6854 2144 6862 2208
rect 6542 2128 6862 2144
rect 9341 16896 9661 17920
rect 9341 16832 9349 16896
rect 9413 16832 9429 16896
rect 9493 16832 9509 16896
rect 9573 16832 9589 16896
rect 9653 16832 9661 16896
rect 9341 15808 9661 16832
rect 9341 15744 9349 15808
rect 9413 15744 9429 15808
rect 9493 15744 9509 15808
rect 9573 15744 9589 15808
rect 9653 15744 9661 15808
rect 9341 14720 9661 15744
rect 9341 14656 9349 14720
rect 9413 14656 9429 14720
rect 9493 14656 9509 14720
rect 9573 14656 9589 14720
rect 9653 14656 9661 14720
rect 9341 13632 9661 14656
rect 9341 13568 9349 13632
rect 9413 13568 9429 13632
rect 9493 13568 9509 13632
rect 9573 13568 9589 13632
rect 9653 13568 9661 13632
rect 9341 12544 9661 13568
rect 9341 12480 9349 12544
rect 9413 12480 9429 12544
rect 9493 12480 9509 12544
rect 9573 12480 9589 12544
rect 9653 12480 9661 12544
rect 9341 11456 9661 12480
rect 9341 11392 9349 11456
rect 9413 11392 9429 11456
rect 9493 11392 9509 11456
rect 9573 11392 9589 11456
rect 9653 11392 9661 11456
rect 9341 10368 9661 11392
rect 9341 10304 9349 10368
rect 9413 10304 9429 10368
rect 9493 10304 9509 10368
rect 9573 10304 9589 10368
rect 9653 10304 9661 10368
rect 9341 9280 9661 10304
rect 9341 9216 9349 9280
rect 9413 9216 9429 9280
rect 9493 9216 9509 9280
rect 9573 9216 9589 9280
rect 9653 9216 9661 9280
rect 9341 8192 9661 9216
rect 9341 8128 9349 8192
rect 9413 8128 9429 8192
rect 9493 8128 9509 8192
rect 9573 8128 9589 8192
rect 9653 8128 9661 8192
rect 9341 7104 9661 8128
rect 9341 7040 9349 7104
rect 9413 7040 9429 7104
rect 9493 7040 9509 7104
rect 9573 7040 9589 7104
rect 9653 7040 9661 7104
rect 9341 6016 9661 7040
rect 9341 5952 9349 6016
rect 9413 5952 9429 6016
rect 9493 5952 9509 6016
rect 9573 5952 9589 6016
rect 9653 5952 9661 6016
rect 9341 4928 9661 5952
rect 9341 4864 9349 4928
rect 9413 4864 9429 4928
rect 9493 4864 9509 4928
rect 9573 4864 9589 4928
rect 9653 4864 9661 4928
rect 9341 3840 9661 4864
rect 9341 3776 9349 3840
rect 9413 3776 9429 3840
rect 9493 3776 9509 3840
rect 9573 3776 9589 3840
rect 9653 3776 9661 3840
rect 9341 2752 9661 3776
rect 9341 2688 9349 2752
rect 9413 2688 9429 2752
rect 9493 2688 9509 2752
rect 9573 2688 9589 2752
rect 9653 2688 9661 2752
rect 9341 2128 9661 2688
rect 12140 21792 12460 22352
rect 12140 21728 12148 21792
rect 12212 21728 12228 21792
rect 12292 21728 12308 21792
rect 12372 21728 12388 21792
rect 12452 21728 12460 21792
rect 12140 20704 12460 21728
rect 12140 20640 12148 20704
rect 12212 20640 12228 20704
rect 12292 20640 12308 20704
rect 12372 20640 12388 20704
rect 12452 20640 12460 20704
rect 12140 19616 12460 20640
rect 12140 19552 12148 19616
rect 12212 19552 12228 19616
rect 12292 19552 12308 19616
rect 12372 19552 12388 19616
rect 12452 19552 12460 19616
rect 12140 18528 12460 19552
rect 12140 18464 12148 18528
rect 12212 18464 12228 18528
rect 12292 18464 12308 18528
rect 12372 18464 12388 18528
rect 12452 18464 12460 18528
rect 12140 17440 12460 18464
rect 12140 17376 12148 17440
rect 12212 17376 12228 17440
rect 12292 17376 12308 17440
rect 12372 17376 12388 17440
rect 12452 17376 12460 17440
rect 12140 16352 12460 17376
rect 12140 16288 12148 16352
rect 12212 16288 12228 16352
rect 12292 16288 12308 16352
rect 12372 16288 12388 16352
rect 12452 16288 12460 16352
rect 12140 15264 12460 16288
rect 12140 15200 12148 15264
rect 12212 15200 12228 15264
rect 12292 15200 12308 15264
rect 12372 15200 12388 15264
rect 12452 15200 12460 15264
rect 12140 14176 12460 15200
rect 12140 14112 12148 14176
rect 12212 14112 12228 14176
rect 12292 14112 12308 14176
rect 12372 14112 12388 14176
rect 12452 14112 12460 14176
rect 12140 13088 12460 14112
rect 12140 13024 12148 13088
rect 12212 13024 12228 13088
rect 12292 13024 12308 13088
rect 12372 13024 12388 13088
rect 12452 13024 12460 13088
rect 12140 12000 12460 13024
rect 12140 11936 12148 12000
rect 12212 11936 12228 12000
rect 12292 11936 12308 12000
rect 12372 11936 12388 12000
rect 12452 11936 12460 12000
rect 12140 10912 12460 11936
rect 12140 10848 12148 10912
rect 12212 10848 12228 10912
rect 12292 10848 12308 10912
rect 12372 10848 12388 10912
rect 12452 10848 12460 10912
rect 12140 9824 12460 10848
rect 12140 9760 12148 9824
rect 12212 9760 12228 9824
rect 12292 9760 12308 9824
rect 12372 9760 12388 9824
rect 12452 9760 12460 9824
rect 12140 8736 12460 9760
rect 12140 8672 12148 8736
rect 12212 8672 12228 8736
rect 12292 8672 12308 8736
rect 12372 8672 12388 8736
rect 12452 8672 12460 8736
rect 12140 7648 12460 8672
rect 12140 7584 12148 7648
rect 12212 7584 12228 7648
rect 12292 7584 12308 7648
rect 12372 7584 12388 7648
rect 12452 7584 12460 7648
rect 12140 6560 12460 7584
rect 12140 6496 12148 6560
rect 12212 6496 12228 6560
rect 12292 6496 12308 6560
rect 12372 6496 12388 6560
rect 12452 6496 12460 6560
rect 12140 5472 12460 6496
rect 12140 5408 12148 5472
rect 12212 5408 12228 5472
rect 12292 5408 12308 5472
rect 12372 5408 12388 5472
rect 12452 5408 12460 5472
rect 12140 4384 12460 5408
rect 12140 4320 12148 4384
rect 12212 4320 12228 4384
rect 12292 4320 12308 4384
rect 12372 4320 12388 4384
rect 12452 4320 12460 4384
rect 12140 3296 12460 4320
rect 12140 3232 12148 3296
rect 12212 3232 12228 3296
rect 12292 3232 12308 3296
rect 12372 3232 12388 3296
rect 12452 3232 12460 3296
rect 12140 2208 12460 3232
rect 12140 2144 12148 2208
rect 12212 2144 12228 2208
rect 12292 2144 12308 2208
rect 12372 2144 12388 2208
rect 12452 2144 12460 2208
rect 12140 2128 12460 2144
rect 14939 22336 15259 22352
rect 14939 22272 14947 22336
rect 15011 22272 15027 22336
rect 15091 22272 15107 22336
rect 15171 22272 15187 22336
rect 15251 22272 15259 22336
rect 14939 21248 15259 22272
rect 14939 21184 14947 21248
rect 15011 21184 15027 21248
rect 15091 21184 15107 21248
rect 15171 21184 15187 21248
rect 15251 21184 15259 21248
rect 14939 20160 15259 21184
rect 14939 20096 14947 20160
rect 15011 20096 15027 20160
rect 15091 20096 15107 20160
rect 15171 20096 15187 20160
rect 15251 20096 15259 20160
rect 14939 19072 15259 20096
rect 14939 19008 14947 19072
rect 15011 19008 15027 19072
rect 15091 19008 15107 19072
rect 15171 19008 15187 19072
rect 15251 19008 15259 19072
rect 14939 17984 15259 19008
rect 14939 17920 14947 17984
rect 15011 17920 15027 17984
rect 15091 17920 15107 17984
rect 15171 17920 15187 17984
rect 15251 17920 15259 17984
rect 14939 16896 15259 17920
rect 14939 16832 14947 16896
rect 15011 16832 15027 16896
rect 15091 16832 15107 16896
rect 15171 16832 15187 16896
rect 15251 16832 15259 16896
rect 14939 15808 15259 16832
rect 14939 15744 14947 15808
rect 15011 15744 15027 15808
rect 15091 15744 15107 15808
rect 15171 15744 15187 15808
rect 15251 15744 15259 15808
rect 14939 14720 15259 15744
rect 14939 14656 14947 14720
rect 15011 14656 15027 14720
rect 15091 14656 15107 14720
rect 15171 14656 15187 14720
rect 15251 14656 15259 14720
rect 14939 13632 15259 14656
rect 14939 13568 14947 13632
rect 15011 13568 15027 13632
rect 15091 13568 15107 13632
rect 15171 13568 15187 13632
rect 15251 13568 15259 13632
rect 14939 12544 15259 13568
rect 17738 21792 18058 22352
rect 17738 21728 17746 21792
rect 17810 21728 17826 21792
rect 17890 21728 17906 21792
rect 17970 21728 17986 21792
rect 18050 21728 18058 21792
rect 17738 20704 18058 21728
rect 20537 22336 20857 22352
rect 20537 22272 20545 22336
rect 20609 22272 20625 22336
rect 20689 22272 20705 22336
rect 20769 22272 20785 22336
rect 20849 22272 20857 22336
rect 20537 21248 20857 22272
rect 20537 21184 20545 21248
rect 20609 21184 20625 21248
rect 20689 21184 20705 21248
rect 20769 21184 20785 21248
rect 20849 21184 20857 21248
rect 19379 21044 19445 21045
rect 19379 20980 19380 21044
rect 19444 20980 19445 21044
rect 19379 20979 19445 20980
rect 17738 20640 17746 20704
rect 17810 20640 17826 20704
rect 17890 20640 17906 20704
rect 17970 20640 17986 20704
rect 18050 20640 18058 20704
rect 17738 19616 18058 20640
rect 17738 19552 17746 19616
rect 17810 19552 17826 19616
rect 17890 19552 17906 19616
rect 17970 19552 17986 19616
rect 18050 19552 18058 19616
rect 17738 18528 18058 19552
rect 17738 18464 17746 18528
rect 17810 18464 17826 18528
rect 17890 18464 17906 18528
rect 17970 18464 17986 18528
rect 18050 18464 18058 18528
rect 17738 17440 18058 18464
rect 17738 17376 17746 17440
rect 17810 17376 17826 17440
rect 17890 17376 17906 17440
rect 17970 17376 17986 17440
rect 18050 17376 18058 17440
rect 17738 16352 18058 17376
rect 17738 16288 17746 16352
rect 17810 16288 17826 16352
rect 17890 16288 17906 16352
rect 17970 16288 17986 16352
rect 18050 16288 18058 16352
rect 17738 15264 18058 16288
rect 17738 15200 17746 15264
rect 17810 15200 17826 15264
rect 17890 15200 17906 15264
rect 17970 15200 17986 15264
rect 18050 15200 18058 15264
rect 17738 14176 18058 15200
rect 17738 14112 17746 14176
rect 17810 14112 17826 14176
rect 17890 14112 17906 14176
rect 17970 14112 17986 14176
rect 18050 14112 18058 14176
rect 17738 13088 18058 14112
rect 19382 13429 19442 20979
rect 20537 20160 20857 21184
rect 21219 20908 21285 20909
rect 21219 20844 21220 20908
rect 21284 20844 21285 20908
rect 21219 20843 21285 20844
rect 20537 20096 20545 20160
rect 20609 20096 20625 20160
rect 20689 20096 20705 20160
rect 20769 20096 20785 20160
rect 20849 20096 20857 20160
rect 20537 19072 20857 20096
rect 20537 19008 20545 19072
rect 20609 19008 20625 19072
rect 20689 19008 20705 19072
rect 20769 19008 20785 19072
rect 20849 19008 20857 19072
rect 20537 17984 20857 19008
rect 20537 17920 20545 17984
rect 20609 17920 20625 17984
rect 20689 17920 20705 17984
rect 20769 17920 20785 17984
rect 20849 17920 20857 17984
rect 20299 17508 20365 17509
rect 20299 17444 20300 17508
rect 20364 17444 20365 17508
rect 20299 17443 20365 17444
rect 20302 13565 20362 17443
rect 20537 16896 20857 17920
rect 21035 17916 21101 17917
rect 21035 17852 21036 17916
rect 21100 17852 21101 17916
rect 21035 17851 21101 17852
rect 20537 16832 20545 16896
rect 20609 16832 20625 16896
rect 20689 16832 20705 16896
rect 20769 16832 20785 16896
rect 20849 16832 20857 16896
rect 20537 15808 20857 16832
rect 20537 15744 20545 15808
rect 20609 15744 20625 15808
rect 20689 15744 20705 15808
rect 20769 15744 20785 15808
rect 20849 15744 20857 15808
rect 20537 14720 20857 15744
rect 20537 14656 20545 14720
rect 20609 14656 20625 14720
rect 20689 14656 20705 14720
rect 20769 14656 20785 14720
rect 20849 14656 20857 14720
rect 20537 13632 20857 14656
rect 20537 13568 20545 13632
rect 20609 13568 20625 13632
rect 20689 13568 20705 13632
rect 20769 13568 20785 13632
rect 20849 13568 20857 13632
rect 20299 13564 20365 13565
rect 20299 13500 20300 13564
rect 20364 13500 20365 13564
rect 20299 13499 20365 13500
rect 19379 13428 19445 13429
rect 19379 13364 19380 13428
rect 19444 13364 19445 13428
rect 19379 13363 19445 13364
rect 17738 13024 17746 13088
rect 17810 13024 17826 13088
rect 17890 13024 17906 13088
rect 17970 13024 17986 13088
rect 18050 13024 18058 13088
rect 16803 12884 16869 12885
rect 16803 12820 16804 12884
rect 16868 12820 16869 12884
rect 16803 12819 16869 12820
rect 14939 12480 14947 12544
rect 15011 12480 15027 12544
rect 15091 12480 15107 12544
rect 15171 12480 15187 12544
rect 15251 12480 15259 12544
rect 14939 11456 15259 12480
rect 14939 11392 14947 11456
rect 15011 11392 15027 11456
rect 15091 11392 15107 11456
rect 15171 11392 15187 11456
rect 15251 11392 15259 11456
rect 14939 10368 15259 11392
rect 16619 11252 16685 11253
rect 16619 11188 16620 11252
rect 16684 11188 16685 11252
rect 16619 11187 16685 11188
rect 14939 10304 14947 10368
rect 15011 10304 15027 10368
rect 15091 10304 15107 10368
rect 15171 10304 15187 10368
rect 15251 10304 15259 10368
rect 14939 9280 15259 10304
rect 14939 9216 14947 9280
rect 15011 9216 15027 9280
rect 15091 9216 15107 9280
rect 15171 9216 15187 9280
rect 15251 9216 15259 9280
rect 14939 8192 15259 9216
rect 14939 8128 14947 8192
rect 15011 8128 15027 8192
rect 15091 8128 15107 8192
rect 15171 8128 15187 8192
rect 15251 8128 15259 8192
rect 14939 7104 15259 8128
rect 14939 7040 14947 7104
rect 15011 7040 15027 7104
rect 15091 7040 15107 7104
rect 15171 7040 15187 7104
rect 15251 7040 15259 7104
rect 14939 6016 15259 7040
rect 14939 5952 14947 6016
rect 15011 5952 15027 6016
rect 15091 5952 15107 6016
rect 15171 5952 15187 6016
rect 15251 5952 15259 6016
rect 14939 4928 15259 5952
rect 16622 5949 16682 11187
rect 16806 9485 16866 12819
rect 17738 12000 18058 13024
rect 17738 11936 17746 12000
rect 17810 11936 17826 12000
rect 17890 11936 17906 12000
rect 17970 11936 17986 12000
rect 18050 11936 18058 12000
rect 17738 10912 18058 11936
rect 17738 10848 17746 10912
rect 17810 10848 17826 10912
rect 17890 10848 17906 10912
rect 17970 10848 17986 10912
rect 18050 10848 18058 10912
rect 17738 9824 18058 10848
rect 17738 9760 17746 9824
rect 17810 9760 17826 9824
rect 17890 9760 17906 9824
rect 17970 9760 17986 9824
rect 18050 9760 18058 9824
rect 16803 9484 16869 9485
rect 16803 9420 16804 9484
rect 16868 9420 16869 9484
rect 16803 9419 16869 9420
rect 17738 8736 18058 9760
rect 17738 8672 17746 8736
rect 17810 8672 17826 8736
rect 17890 8672 17906 8736
rect 17970 8672 17986 8736
rect 18050 8672 18058 8736
rect 17738 7648 18058 8672
rect 17738 7584 17746 7648
rect 17810 7584 17826 7648
rect 17890 7584 17906 7648
rect 17970 7584 17986 7648
rect 18050 7584 18058 7648
rect 17738 6560 18058 7584
rect 17738 6496 17746 6560
rect 17810 6496 17826 6560
rect 17890 6496 17906 6560
rect 17970 6496 17986 6560
rect 18050 6496 18058 6560
rect 16619 5948 16685 5949
rect 16619 5884 16620 5948
rect 16684 5884 16685 5948
rect 16619 5883 16685 5884
rect 14939 4864 14947 4928
rect 15011 4864 15027 4928
rect 15091 4864 15107 4928
rect 15171 4864 15187 4928
rect 15251 4864 15259 4928
rect 14939 3840 15259 4864
rect 14939 3776 14947 3840
rect 15011 3776 15027 3840
rect 15091 3776 15107 3840
rect 15171 3776 15187 3840
rect 15251 3776 15259 3840
rect 14939 2752 15259 3776
rect 14939 2688 14947 2752
rect 15011 2688 15027 2752
rect 15091 2688 15107 2752
rect 15171 2688 15187 2752
rect 15251 2688 15259 2752
rect 14939 2128 15259 2688
rect 16622 2549 16682 5883
rect 17738 5472 18058 6496
rect 17738 5408 17746 5472
rect 17810 5408 17826 5472
rect 17890 5408 17906 5472
rect 17970 5408 17986 5472
rect 18050 5408 18058 5472
rect 17738 4384 18058 5408
rect 17738 4320 17746 4384
rect 17810 4320 17826 4384
rect 17890 4320 17906 4384
rect 17970 4320 17986 4384
rect 18050 4320 18058 4384
rect 17738 3296 18058 4320
rect 17738 3232 17746 3296
rect 17810 3232 17826 3296
rect 17890 3232 17906 3296
rect 17970 3232 17986 3296
rect 18050 3232 18058 3296
rect 16619 2548 16685 2549
rect 16619 2484 16620 2548
rect 16684 2484 16685 2548
rect 16619 2483 16685 2484
rect 17738 2208 18058 3232
rect 17738 2144 17746 2208
rect 17810 2144 17826 2208
rect 17890 2144 17906 2208
rect 17970 2144 17986 2208
rect 18050 2144 18058 2208
rect 17738 2128 18058 2144
rect 20537 12544 20857 13568
rect 21038 13429 21098 17851
rect 21222 14925 21282 20843
rect 22875 20364 22941 20365
rect 22875 20300 22876 20364
rect 22940 20300 22941 20364
rect 22875 20299 22941 20300
rect 22878 20178 22938 20299
rect 21219 14924 21285 14925
rect 21219 14860 21220 14924
rect 21284 14860 21285 14924
rect 21219 14859 21285 14860
rect 21035 13428 21101 13429
rect 21035 13364 21036 13428
rect 21100 13364 21101 13428
rect 21035 13363 21101 13364
rect 20537 12480 20545 12544
rect 20609 12480 20625 12544
rect 20689 12480 20705 12544
rect 20769 12480 20785 12544
rect 20849 12480 20857 12544
rect 20537 11456 20857 12480
rect 20537 11392 20545 11456
rect 20609 11392 20625 11456
rect 20689 11392 20705 11456
rect 20769 11392 20785 11456
rect 20849 11392 20857 11456
rect 20537 10368 20857 11392
rect 20537 10304 20545 10368
rect 20609 10304 20625 10368
rect 20689 10304 20705 10368
rect 20769 10304 20785 10368
rect 20849 10304 20857 10368
rect 20537 9280 20857 10304
rect 20537 9216 20545 9280
rect 20609 9216 20625 9280
rect 20689 9216 20705 9280
rect 20769 9216 20785 9280
rect 20849 9216 20857 9280
rect 20537 8192 20857 9216
rect 20537 8128 20545 8192
rect 20609 8128 20625 8192
rect 20689 8128 20705 8192
rect 20769 8128 20785 8192
rect 20849 8128 20857 8192
rect 20537 7104 20857 8128
rect 20537 7040 20545 7104
rect 20609 7040 20625 7104
rect 20689 7040 20705 7104
rect 20769 7040 20785 7104
rect 20849 7040 20857 7104
rect 20537 6016 20857 7040
rect 20537 5952 20545 6016
rect 20609 5952 20625 6016
rect 20689 5952 20705 6016
rect 20769 5952 20785 6016
rect 20849 5952 20857 6016
rect 20537 4928 20857 5952
rect 20537 4864 20545 4928
rect 20609 4864 20625 4928
rect 20689 4864 20705 4928
rect 20769 4864 20785 4928
rect 20849 4864 20857 4928
rect 20537 3840 20857 4864
rect 20537 3776 20545 3840
rect 20609 3776 20625 3840
rect 20689 3776 20705 3840
rect 20769 3776 20785 3840
rect 20849 3776 20857 3840
rect 20537 2752 20857 3776
rect 20537 2688 20545 2752
rect 20609 2688 20625 2752
rect 20689 2688 20705 2752
rect 20769 2688 20785 2752
rect 20849 2688 20857 2752
rect 20537 2128 20857 2688
<< via4 >>
rect 7886 20092 8122 20178
rect 7886 20028 7972 20092
rect 7972 20028 8036 20092
rect 8036 20028 8122 20092
rect 7886 19942 8122 20028
rect 22790 19942 23026 20178
<< metal5 >>
rect 7844 20178 23068 20220
rect 7844 19942 7886 20178
rect 8122 19942 22790 20178
rect 23026 19942 23068 20178
rect 7844 19900 23068 19942
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_E_FTB01_A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17940 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_FTB00_A
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_Test_en_W_FTB01_A
timestamp 1649977179
transform 1 0 1656 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform 1 0 8648 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform -1 0 1564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform -1 0 13984 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform -1 0 11684 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform -1 0 13984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__75__A
timestamp 1649977179
transform 1 0 2300 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__76__A
timestamp 1649977179
transform -1 0 2668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__77__A
timestamp 1649977179
transform 1 0 2668 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__78__A
timestamp 1649977179
transform 1 0 3220 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__79__A
timestamp 1649977179
transform 1 0 4048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__81__A
timestamp 1649977179
transform 1 0 3128 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__82__A
timestamp 1649977179
transform 1 0 4600 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_0_N_in_A
timestamp 1649977179
transform -1 0 16192 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 6440 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 5336 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 6532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 10948 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 14168 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 13984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform -1 0 21160 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk_A
timestamp 1649977179
transform -1 0 19412 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold71_A
timestamp 1649977179
transform -1 0 2576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold105_A
timestamp 1649977179
transform -1 0 3956 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold118_A
timestamp 1649977179
transform -1 0 3312 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold139_A
timestamp 1649977179
transform -1 0 3312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold150_A
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold178_A
timestamp 1649977179
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hold194_A
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 2300 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 16560 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 1840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 9108 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 20240 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 18400 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 23184 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 20884 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 22908 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 19688 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 20240 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 23184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 23184 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 18860 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 23184 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 19136 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform 1 0 12328 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform 1 0 17020 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 22908 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 6532 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 13800 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 11408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 14260 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 22816 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 14260 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 11408 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 7084 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 4784 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 8924 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform 1 0 8648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 16560 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 6256 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 7268 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 4324 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9752 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A0
timestamp 1649977179
transform 1 0 9016 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6__A1
timestamp 1649977179
transform -1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A0
timestamp 1649977179
transform -1 0 9016 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7__A1
timestamp 1649977179
transform -1 0 13616 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__A
timestamp 1649977179
transform -1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11__D
timestamp 1649977179
transform -1 0 19136 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13__D
timestamp 1649977179
transform -1 0 15088 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15__D
timestamp 1649977179
transform -1 0 19872 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16__D
timestamp 1649977179
transform -1 0 14720 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 14904 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0__S
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0__D
timestamp 1649977179
transform -1 0 18308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1__D
timestamp 1649977179
transform -1 0 22816 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0__S
timestamp 1649977179
transform -1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1__A
timestamp 1649977179
transform 1 0 11684 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2__A
timestamp 1649977179
transform 1 0 10488 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0__B
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 20884 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output38_A
timestamp 1649977179
transform 1 0 13064 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output45_A
timestamp 1649977179
transform 1 0 12420 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output50_A
timestamp 1649977179
transform -1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output54_A
timestamp 1649977179
transform 1 0 14904 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output62_A
timestamp 1649977179
transform 1 0 14904 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output64_A
timestamp 1649977179
transform 1 0 15916 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output66_A
timestamp 1649977179
transform 1 0 13524 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output68_A
timestamp 1649977179
transform -1 0 19136 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output70_A
timestamp 1649977179
transform -1 0 22816 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1649977179
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1649977179
transform -1 0 23184 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output78_A
timestamp 1649977179
transform -1 0 18400 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1649977179
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_6 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1656 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_47
timestamp 1649977179
transform 1 0 5428 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_64
timestamp 1649977179
transform 1 0 6992 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_19
timestamp 1649977179
transform 1 0 2852 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_68
timestamp 1649977179
transform 1 0 7360 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_129
timestamp 1649977179
transform 1 0 12972 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_11
timestamp 1649977179
transform 1 0 2116 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_131
timestamp 1649977179
transform 1 0 13156 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_21
timestamp 1649977179
transform 1 0 3036 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_75
timestamp 1649977179
transform 1 0 8004 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_128
timestamp 1649977179
transform 1 0 12880 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_239
timestamp 1649977179
transform 1 0 23092 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_19
timestamp 1649977179
transform 1 0 2852 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_79
timestamp 1649977179
transform 1 0 8372 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1649977179
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_220
timestamp 1649977179
transform 1 0 21344 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_7_15 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_26
timestamp 1649977179
transform 1 0 3496 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_65
timestamp 1649977179
transform 1 0 7084 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_95
timestamp 1649977179
transform 1 0 9844 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_126
timestamp 1649977179
transform 1 0 12696 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_151
timestamp 1649977179
transform 1 0 14996 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_16
timestamp 1649977179
transform 1 0 2576 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_58
timestamp 1649977179
transform 1 0 6440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_182
timestamp 1649977179
transform 1 0 17848 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_213
timestamp 1649977179
transform 1 0 20700 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_22
timestamp 1649977179
transform 1 0 3128 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_71
timestamp 1649977179
transform 1 0 7636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_185
timestamp 1649977179
transform 1 0 18124 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_220
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_235
timestamp 1649977179
transform 1 0 22724 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_71
timestamp 1649977179
transform 1 0 7636 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_75
timestamp 1649977179
transform 1 0 8004 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_157
timestamp 1649977179
transform 1 0 15548 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_161
timestamp 1649977179
transform 1 0 15916 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_186
timestamp 1649977179
transform 1 0 18216 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_9
timestamp 1649977179
transform 1 0 1932 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_44
timestamp 1649977179
transform 1 0 5152 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_65
timestamp 1649977179
transform 1 0 7084 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_103
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_117
timestamp 1649977179
transform 1 0 11868 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_185
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_239
timestamp 1649977179
transform 1 0 23092 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_64
timestamp 1649977179
transform 1 0 6992 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_12_103
timestamp 1649977179
transform 1 0 10580 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_135
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_168
timestamp 1649977179
transform 1 0 16560 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_178
timestamp 1649977179
transform 1 0 17480 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_203
timestamp 1649977179
transform 1 0 19780 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_223
timestamp 1649977179
transform 1 0 21620 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_8
timestamp 1649977179
transform 1 0 1840 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_127
timestamp 1649977179
transform 1 0 12788 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_131
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_23
timestamp 1649977179
transform 1 0 3220 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_38
timestamp 1649977179
transform 1 0 4600 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_64
timestamp 1649977179
transform 1 0 6992 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_94
timestamp 1649977179
transform 1 0 9752 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_111
timestamp 1649977179
transform 1 0 11316 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_117
timestamp 1649977179
transform 1 0 11868 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_137
timestamp 1649977179
transform 1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_115
timestamp 1649977179
transform 1 0 11684 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_119
timestamp 1649977179
transform 1 0 12052 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_178
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_182
timestamp 1649977179
transform 1 0 17848 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_207
timestamp 1649977179
transform 1 0 20148 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_236
timestamp 1649977179
transform 1 0 22816 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_23
timestamp 1649977179
transform 1 0 3220 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1649977179
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_120
timestamp 1649977179
transform 1 0 12144 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_182
timestamp 1649977179
transform 1 0 17848 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_236
timestamp 1649977179
transform 1 0 22816 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_94
timestamp 1649977179
transform 1 0 9752 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_123
timestamp 1649977179
transform 1 0 12420 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_142
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1649977179
transform 1 0 16928 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_9
timestamp 1649977179
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1649977179
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_45
timestamp 1649977179
transform 1 0 5244 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_51
timestamp 1649977179
transform 1 0 5796 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_88
timestamp 1649977179
transform 1 0 9200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_114
timestamp 1649977179
transform 1 0 11592 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_193
timestamp 1649977179
transform 1 0 18860 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_7
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_24
timestamp 1649977179
transform 1 0 3312 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_34
timestamp 1649977179
transform 1 0 4232 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_45
timestamp 1649977179
transform 1 0 5244 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_63
timestamp 1649977179
transform 1 0 6900 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_122
timestamp 1649977179
transform 1 0 12328 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_158
timestamp 1649977179
transform 1 0 15640 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_202
timestamp 1649977179
transform 1 0 19688 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_47
timestamp 1649977179
transform 1 0 5428 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_123
timestamp 1649977179
transform 1 0 12420 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_147
timestamp 1649977179
transform 1 0 14628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_172
timestamp 1649977179
transform 1 0 16928 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_206
timestamp 1649977179
transform 1 0 20056 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_97
timestamp 1649977179
transform 1 0 10028 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_129
timestamp 1649977179
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_180
timestamp 1649977179
transform 1 0 17664 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_32
timestamp 1649977179
transform 1 0 4048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1649977179
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_111
timestamp 1649977179
transform 1 0 11316 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_73
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_130
timestamp 1649977179
transform 1 0 13064 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_194
timestamp 1649977179
transform 1 0 18952 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_56
timestamp 1649977179
transform 1 0 6256 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1649977179
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_114
timestamp 1649977179
transform 1 0 11592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_123
timestamp 1649977179
transform 1 0 12420 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_131
timestamp 1649977179
transform 1 0 13156 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_192
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_94
timestamp 1649977179
transform 1 0 9752 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_24
timestamp 1649977179
transform 1 0 3312 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_110
timestamp 1649977179
transform 1 0 11224 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_208
timestamp 1649977179
transform 1 0 20240 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_109
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_96
timestamp 1649977179
transform 1 0 9936 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_65
timestamp 1649977179
transform 1 0 7084 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_141
timestamp 1649977179
transform 1 0 14076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_151
timestamp 1649977179
transform 1 0 14996 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_136
timestamp 1649977179
transform 1 0 13616 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_210
timestamp 1649977179
transform 1 0 20424 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_235
timestamp 1649977179
transform 1 0 22724 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_50
timestamp 1649977179
transform 1 0 5704 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1649977179
transform 1 0 6624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_135
timestamp 1649977179
transform 1 0 13524 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_207
timestamp 1649977179
transform 1 0 20148 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_37
timestamp 1649977179
transform 1 0 4508 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_128
timestamp 1649977179
transform 1 0 12880 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_116
timestamp 1649977179
transform 1 0 11776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_174
timestamp 1649977179
transform 1 0 17112 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_185
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_207
timestamp 1649977179
transform 1 0 20148 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_51
timestamp 1649977179
transform 1 0 5796 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_96
timestamp 1649977179
transform 1 0 9936 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_191
timestamp 1649977179
transform 1 0 18676 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_24
timestamp 1649977179
transform 1 0 3312 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_41
timestamp 1649977179
transform 1 0 4876 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_47
timestamp 1649977179
transform 1 0 5428 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_83
timestamp 1649977179
transform 1 0 8740 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_61
timestamp 1649977179
transform 1 0 6716 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_113
timestamp 1649977179
transform 1 0 11500 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_36_149
timestamp 1649977179
transform 1 0 14812 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 23460 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 23460 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 23460 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 23460 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 23460 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 23460 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 23460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 23460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 23460 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 23460 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 23460 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 23460 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 23460 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 23460 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 23460 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 23460 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 23460 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 23460 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 23460 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 23460 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 23460 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 23460 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 23460 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 23460 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 23460 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 23460 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 23460 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 23460 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 23460 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 23460 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 23460 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 23460 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 23460 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 6256 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 11408 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 16560 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 21712 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_E_FTB01 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21068 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  Test_en_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6624 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_W_FTB01
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform -1 0 8556 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform -1 0 1840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform -1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform -1 0 11776 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform -1 0 13984 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform -1 0 11960 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform -1 0 16560 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform 1 0 22632 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform 1 0 20700 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1649977179
transform 1 0 2024 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1649977179
transform 1 0 2668 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp 1649977179
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1649977179
transform -1 0 2024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_0_FTB00
timestamp 1649977179
transform -1 0 16928 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12144 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk_0_N_in
timestamp 1649977179
transform -1 0 14536 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk_0_N_in
timestamp 1649977179
transform -1 0 11408 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk_0_N_in
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_0_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5428 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_1_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform -1 0 4784 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_2_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 9384 0 -1 7616
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_3_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 9568 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_4_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 4324 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_5_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 4048 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_6_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 9936 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_7_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_8_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform -1 0 16560 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_9_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_10_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 19688 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_11_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 19872 0 1 8704
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_12_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 14536 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_13_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 15272 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_14_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 19872 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  clkbuf_4_15_0_ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 19412 0 1 18496
box -38 -48 1050 592
use sky130_fd_sc_hd__conb_1  grid_clb_105 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8832 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1649977179
transform -1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1649977179
transform -1 0 6348 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1649977179
transform -1 0 6164 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1649977179
transform 1 0 9016 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1649977179
transform -1 0 4784 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1649977179
transform 1 0 12880 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1649977179
transform 1 0 14444 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1649977179
transform -1 0 16468 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1649977179
transform 1 0 17480 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1649977179
transform 1 0 18032 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1649977179
transform -1 0 18308 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1649977179
transform -1 0 4692 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1649977179
transform 1 0 10672 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1649977179
transform -1 0 14076 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1649977179
transform -1 0 9660 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1649977179
transform -1 0 11408 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1649977179
transform 1 0 17388 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1649977179
transform 1 0 17020 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1649977179
transform -1 0 4600 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1649977179
transform -1 0 13156 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1649977179
transform -1 0 3496 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1649977179
transform -1 0 16560 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1649977179
transform -1 0 12420 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1649977179
transform -1 0 6716 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold32 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20976 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1649977179
transform -1 0 12144 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1649977179
transform -1 0 23184 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1649977179
transform -1 0 2484 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1649977179
transform -1 0 16928 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1649977179
transform 1 0 18584 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1649977179
transform -1 0 3680 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1649977179
transform -1 0 16376 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1649977179
transform -1 0 5428 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1649977179
transform 1 0 19044 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1649977179
transform -1 0 21436 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1649977179
transform 1 0 6348 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1649977179
transform 1 0 4968 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1649977179
transform -1 0 12144 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1649977179
transform -1 0 14812 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold49
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1649977179
transform -1 0 5520 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1649977179
transform -1 0 11408 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1649977179
transform 1 0 11684 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold53
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold54
timestamp 1649977179
transform -1 0 16008 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1649977179
transform -1 0 21436 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1649977179
transform 1 0 15824 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold57
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold58
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1649977179
transform 1 0 12052 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1649977179
transform 1 0 12880 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold61
timestamp 1649977179
transform -1 0 3680 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold62
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold63
timestamp 1649977179
transform -1 0 3956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold64
timestamp 1649977179
transform -1 0 15548 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold65
timestamp 1649977179
transform -1 0 7084 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold66
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold67
timestamp 1649977179
transform -1 0 3680 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold68
timestamp 1649977179
transform 1 0 4508 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold69
timestamp 1649977179
transform -1 0 8832 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold70
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold71
timestamp 1649977179
transform 1 0 2576 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold72
timestamp 1649977179
transform -1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold73
timestamp 1649977179
transform -1 0 20056 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold74
timestamp 1649977179
transform -1 0 10212 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold75
timestamp 1649977179
transform 1 0 15640 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold76
timestamp 1649977179
transform -1 0 8832 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold77
timestamp 1649977179
transform 1 0 15180 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold78
timestamp 1649977179
transform -1 0 14812 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold79
timestamp 1649977179
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold80
timestamp 1649977179
transform -1 0 2208 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold81
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold82
timestamp 1649977179
transform -1 0 4692 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold83
timestamp 1649977179
transform -1 0 8280 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold84
timestamp 1649977179
transform 1 0 17756 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold85
timestamp 1649977179
transform -1 0 3680 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold86
timestamp 1649977179
transform -1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold87
timestamp 1649977179
transform 1 0 13248 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold88
timestamp 1649977179
transform 1 0 1748 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold89
timestamp 1649977179
transform -1 0 4048 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold90
timestamp 1649977179
transform -1 0 10028 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold91
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold92
timestamp 1649977179
transform -1 0 2668 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold93
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold94
timestamp 1649977179
transform -1 0 7268 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold95
timestamp 1649977179
transform -1 0 7084 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold96
timestamp 1649977179
transform 1 0 20700 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold97
timestamp 1649977179
transform -1 0 3680 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold98
timestamp 1649977179
transform -1 0 15272 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold99
timestamp 1649977179
transform 1 0 15180 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold100
timestamp 1649977179
transform -1 0 12880 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold101
timestamp 1649977179
transform 1 0 12144 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold102
timestamp 1649977179
transform -1 0 17020 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold103
timestamp 1649977179
transform -1 0 20976 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold104
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold105
timestamp 1649977179
transform -1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold106
timestamp 1649977179
transform -1 0 21712 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold107
timestamp 1649977179
transform -1 0 19964 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold108
timestamp 1649977179
transform 1 0 4048 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold109
timestamp 1649977179
transform -1 0 16008 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold110
timestamp 1649977179
transform 1 0 6900 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold111
timestamp 1649977179
transform -1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold112
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold113
timestamp 1649977179
transform -1 0 7268 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold114
timestamp 1649977179
transform -1 0 4784 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold115
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold116
timestamp 1649977179
transform -1 0 6992 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold117
timestamp 1649977179
transform -1 0 10120 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold118
timestamp 1649977179
transform 1 0 3312 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold119
timestamp 1649977179
transform -1 0 6256 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold120
timestamp 1649977179
transform 1 0 18124 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold121
timestamp 1649977179
transform -1 0 4784 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold122
timestamp 1649977179
transform -1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold123
timestamp 1649977179
transform -1 0 6164 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold124
timestamp 1649977179
transform -1 0 22540 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold125
timestamp 1649977179
transform -1 0 13984 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold126
timestamp 1649977179
transform -1 0 9568 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold127
timestamp 1649977179
transform -1 0 18860 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold128
timestamp 1649977179
transform -1 0 9936 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold129
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold130
timestamp 1649977179
transform 1 0 10212 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold131
timestamp 1649977179
transform -1 0 3680 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold132
timestamp 1649977179
transform 1 0 18216 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold133
timestamp 1649977179
transform -1 0 4508 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold134
timestamp 1649977179
transform -1 0 7360 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold135
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold136
timestamp 1649977179
transform -1 0 4048 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold137
timestamp 1649977179
transform -1 0 2576 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold138
timestamp 1649977179
transform 1 0 15732 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold139
timestamp 1649977179
transform 1 0 3312 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold140
timestamp 1649977179
transform 1 0 11776 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold141
timestamp 1649977179
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold142
timestamp 1649977179
transform 1 0 1472 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold143
timestamp 1649977179
transform -1 0 15640 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold144
timestamp 1649977179
transform 1 0 17480 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold145
timestamp 1649977179
transform -1 0 2944 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold146
timestamp 1649977179
transform 1 0 7268 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold147
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold148
timestamp 1649977179
transform -1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold149
timestamp 1649977179
transform -1 0 3680 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold150
timestamp 1649977179
transform -1 0 2944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold151
timestamp 1649977179
transform -1 0 15548 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold152
timestamp 1649977179
transform 1 0 13892 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold153
timestamp 1649977179
transform -1 0 13248 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold154
timestamp 1649977179
transform -1 0 16560 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold155
timestamp 1649977179
transform -1 0 16744 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold156
timestamp 1649977179
transform -1 0 22540 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold157
timestamp 1649977179
transform -1 0 6348 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold158
timestamp 1649977179
transform -1 0 21712 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold159
timestamp 1649977179
transform -1 0 17664 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold160
timestamp 1649977179
transform -1 0 6256 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold161
timestamp 1649977179
transform 1 0 18952 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold162
timestamp 1649977179
transform -1 0 4232 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold163
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold164
timestamp 1649977179
transform -1 0 7084 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold165
timestamp 1649977179
transform 1 0 5888 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold166
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold167
timestamp 1649977179
transform -1 0 21712 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold168
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold169
timestamp 1649977179
transform 1 0 4232 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold170
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold171
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold172
timestamp 1649977179
transform -1 0 12236 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold173
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold174
timestamp 1649977179
transform -1 0 22724 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold175
timestamp 1649977179
transform -1 0 18952 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold176
timestamp 1649977179
transform 1 0 20884 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold177
timestamp 1649977179
transform -1 0 18492 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold178
timestamp 1649977179
transform 1 0 4048 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold179
timestamp 1649977179
transform -1 0 10396 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold180
timestamp 1649977179
transform -1 0 9660 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold181
timestamp 1649977179
transform -1 0 6256 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold182
timestamp 1649977179
transform 1 0 9108 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold183
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold184
timestamp 1649977179
transform -1 0 15640 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold185
timestamp 1649977179
transform -1 0 5428 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold186
timestamp 1649977179
transform -1 0 8740 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold187
timestamp 1649977179
transform -1 0 2668 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold188
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold189
timestamp 1649977179
transform -1 0 15640 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold190
timestamp 1649977179
transform -1 0 13984 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold191
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold192
timestamp 1649977179
transform 1 0 15456 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold193
timestamp 1649977179
transform -1 0 7360 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold194
timestamp 1649977179
transform -1 0 3680 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold195
timestamp 1649977179
transform -1 0 8004 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 8832 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23184 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 1656 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 11408 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 22908 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 22908 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform 1 0 22908 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform 1 0 22908 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform 1 0 22908 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform 1 0 22908 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 22908 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 23184 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 11408 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform -1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 21712 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform 1 0 5704 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform 1 0 11868 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 11868 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 12512 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform 1 0 20700 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform 1 0 21436 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 5520 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 1656 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform 1 0 22172 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform 1 0 10028 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform 1 0 9752 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 9108 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform 1 0 9108 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform 1 0 9384 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 9936 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9936 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform -1 0 8372 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4324 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3496 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4600 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 5336 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 6164 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 5152 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 3220 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4508 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3956 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3496 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4324 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 5428 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4416 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 4324 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 6164 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 3680 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 3772 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 3680 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform -1 0 4324 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 4324 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 5796 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 6624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5888 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3128 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2024 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 2208 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 4692 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 3956 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 4784 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform -1 0 6900 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 5520 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform -1 0 6256 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 4692 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform -1 0 6256 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform -1 0 3220 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 1748 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform -1 0 3220 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 2024 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 3312 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 2116 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4600 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__127
timestamp 1649977179
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2852 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4324 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4968 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7820 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7176 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9476 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5336 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__128
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6624 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__129
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 7176 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_0.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__130
timestamp 1649977179
transform 1 0 9476 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform -1 0 8648 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 7268 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform -1 0 3312 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform -1 0 3772 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 6072 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform -1 0 3772 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform -1 0 4600 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform -1 0 3312 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform -1 0 2208 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5796 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3220 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4784 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 4876 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4876 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 5152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 6992 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 1748 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 4048 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 3680 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 4876 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 6716 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 9476 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 2944 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform -1 0 5428 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 2852 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 1472 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 2852 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 3772 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 4600 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 4784 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 5060 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform -1 0 2944 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 2024 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform 1 0 3496 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 1656 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 1472 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform -1 0 3220 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform 1 0 2208 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 3404 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4324 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4784 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5980 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6808 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__131
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8280 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7268 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8832 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7268 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8648 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__132
timestamp 1649977179
transform -1 0 4048 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7268 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__133
timestamp 1649977179
transform 1 0 9660 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7820 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8188 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__134
timestamp 1649977179
transform -1 0 7268 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_1.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 10488 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9292 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9016 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform -1 0 7912 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 9752 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 10580 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 11592 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9292 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8740 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8740 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10120 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10212 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 10948 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10488 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 10488 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 11592 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 10212 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 8832 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 9200 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform -1 0 9384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 11316 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform 1 0 11960 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8464 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8188 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6716 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 8464 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform -1 0 8648 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 7360 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 7360 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 8280 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform 1 0 9108 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform 1 0 9844 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform -1 0 11408 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 9936 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform -1 0 11592 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform 1 0 10488 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13064 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11408 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10488 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__135
timestamp 1649977179
transform 1 0 11408 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10488 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11224 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11316 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11408 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11132 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10304 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__136
timestamp 1649977179
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11316 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10396 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__137
timestamp 1649977179
transform 1 0 11500 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9660 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_2.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__106
timestamp 1649977179
transform 1 0 10856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 17112 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13340 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13432 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform 1 0 14260 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 14444 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform -1 0 13800 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12972 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform -1 0 14996 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform -1 0 14076 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 14444 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 14996 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform -1 0 16560 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 17296 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 17664 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 17388 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 12880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 13984 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform 1 0 14904 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform -1 0 14076 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform 1 0 12512 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 16652 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform -1 0 17112 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11960 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13892 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 12236 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 14260 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 14812 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 15088 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform 1 0 15088 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform -1 0 17020 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform -1 0 15548 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform -1 0 13524 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 12144 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform 1 0 12512 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform -1 0 15548 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 14260 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15548 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17848 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18676 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__107
timestamp 1649977179
transform 1 0 21160 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18124 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21068 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19964 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 20240 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18216 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 19780 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19504 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__108
timestamp 1649977179
transform -1 0 19136 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 22632 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__109
timestamp 1649977179
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18216 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__110
timestamp 1649977179
transform 1 0 22908 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_3.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17296 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 19688 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17020 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform -1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 17020 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform -1 0 18676 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform -1 0 19688 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 20792 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform -1 0 17388 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform -1 0 20056 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform -1 0 21344 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18308 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform 1 0 19412 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 19412 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 20240 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 19136 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 17664 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 21712 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 23000 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 16560 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform 1 0 22632 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16008 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 17020 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 15088 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 16560 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 15088 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 15548 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform -1 0 16560 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform 1 0 16744 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform -1 0 21068 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 19320 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 20240 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform 1 0 20240 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 21712 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 21712 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17664 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18584 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 19136 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__111
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18216 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21344 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 21068 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18400 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19688 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 21344 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__112
timestamp 1649977179
transform -1 0 19688 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 22632 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 21896 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__113
timestamp 1649977179
transform 1 0 22908 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19688 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__114
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_4.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 19136 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 11408 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 12788 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8096 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform -1 0 7176 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform -1 0 6992 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform 1 0 6992 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 8004 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 9384 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8004 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform -1 0 7360 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7728 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10948 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 10304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 9568 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 8832 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 7360 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 7728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform -1 0 8096 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 10396 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 10764 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 10304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 10948 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform -1 0 12236 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 9384 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10396 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10396 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 6256 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 5428 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform -1 0 8372 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 4784 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 4784 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform 1 0 4784 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 5520 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 7084 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 7360 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform -1 0 10672 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 9568 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11040 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11408 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__115
timestamp 1649977179
transform -1 0 12052 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13064 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12236 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12512 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16284 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9936 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13892 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__116
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14536 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_2  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16560 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__117
timestamp 1649977179
transform -1 0 14996 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12052 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__118
timestamp 1649977179
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_5.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 17940 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12696 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13156 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform 1 0 15732 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform 1 0 14904 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform -1 0 14444 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform -1 0 13800 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform -1 0 14812 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13524 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform 1 0 13984 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform -1 0 14904 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform -1 0 14904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15732 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 15180 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform -1 0 16560 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 17848 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 17572 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 13708 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 14352 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform 1 0 15456 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform 1 0 15180 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 17388 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 15916 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform -1 0 16560 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10212 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13156 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 11960 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform -1 0 15548 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform 1 0 14352 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform -1 0 15824 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform -1 0 13432 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 12144 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform 1 0 12328 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform -1 0 13984 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform 1 0 12512 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform 1 0 13156 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform 1 0 14628 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 14720 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15640 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18584 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__119
timestamp 1649977179
transform 1 0 18584 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17572 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17112 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18584 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19320 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15824 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18768 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18768 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__120
timestamp 1649977179
transform -1 0 19504 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 20884 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 20700 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__121
timestamp 1649977179
transform -1 0 20148 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20792 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__122
timestamp 1649977179
transform -1 0 16560 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_6.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__sdfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_0.sky130_fd_sc_hd__sdfxtp_1_0_
timestamp 1649977179
transform 1 0 19964 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__sdfxtp_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_clb_fle_ff_1.sky130_fd_sc_hd__sdfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19688 0 1 11968
box -38 -48 2062 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_0_
timestamp 1649977179
transform -1 0 19136 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_1_
timestamp 1649977179
transform -1 0 19872 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_2_
timestamp 1649977179
transform -1 0 18952 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_3_
timestamp 1649977179
transform -1 0 18768 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_4_
timestamp 1649977179
transform -1 0 19688 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_5_
timestamp 1649977179
transform -1 0 19596 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_6_
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l1_in_7_
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_1_
timestamp 1649977179
transform -1 0 19228 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_2_
timestamp 1649977179
transform 1 0 19688 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l2_in_3_
timestamp 1649977179
transform 1 0 20792 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_0_
timestamp 1649977179
transform -1 0 20884 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l3_in_1_
timestamp 1649977179
transform -1 0 21160 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.mux_l4_in_0_
timestamp 1649977179
transform 1 0 20884 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform -1 0 21436 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform 1 0 20148 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform -1 0 21160 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform -1 0 20240 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_4_
timestamp 1649977179
transform -1 0 19136 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_5_
timestamp 1649977179
transform -1 0 19136 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.frac_lut4_mux_0_.sky130_fd_sc_hd__buf_2_6_
timestamp 1649977179
transform 1 0 20516 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_0_
timestamp 1649977179
transform 1 0 22908 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_1_
timestamp 1649977179
transform -1 0 23000 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_2_
timestamp 1649977179
transform 1 0 22632 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__buf_2_3_
timestamp 1649977179
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_0_.sky130_fd_sc_hd__or2_1_0_
timestamp 1649977179
transform 1 0 22540 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17480 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 18492 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 20700 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 18124 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_5_
timestamp 1649977179
transform 1 0 16100 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_6_
timestamp 1649977179
transform 1 0 16468 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_7_
timestamp 1649977179
transform -1 0 18400 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_8_
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_9_
timestamp 1649977179
transform -1 0 18860 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_10_
timestamp 1649977179
transform 1 0 17664 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_11_
timestamp 1649977179
transform -1 0 20700 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_12_
timestamp 1649977179
transform 1 0 19596 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_13_
timestamp 1649977179
transform -1 0 21988 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_14_
timestamp 1649977179
transform 1 0 21160 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_15_
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.ltile_frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_16_
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mem_frac_logic_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 21160 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 22632 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0__123
timestamp 1649977179
transform 1 0 22632 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.ltile_frac_logic_0.mux_frac_logic_out_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 22632 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 21252 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21712 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 21712 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_fabric_out_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 21068 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 20240 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mem_ff_0_D_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 21712 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0__124
timestamp 1649977179
transform 1 0 22632 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20424 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0__125
timestamp 1649977179
transform 1 0 22632 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_fabric_out_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20884 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 21896 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0__126
timestamp 1649977179
transform 1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  ltile_clb_mode__0.ltile_fle_7.ltile_phy_fabric_0.mux_ff_0_D_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  output38 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11316 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output39
timestamp 1649977179
transform 1 0 17664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output40
timestamp 1649977179
transform 1 0 22816 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output41
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1649977179
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output43
timestamp 1649977179
transform 1 0 22816 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output44
timestamp 1649977179
transform -1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output45
timestamp 1649977179
transform -1 0 12052 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output46
timestamp 1649977179
transform -1 0 15088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output47
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform -1 0 18860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform 1 0 22816 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform 1 0 22816 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform 1 0 18400 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform 1 0 15088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform 1 0 16376 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform 1 0 19504 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform 1 0 22540 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform 1 0 22540 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform -1 0 20240 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform -1 0 20700 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform 1 0 21344 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform 1 0 22816 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 1748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 21804 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 1748 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform 1 0 22632 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform 1 0 1748 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 21344 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform 1 0 2300 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 16744 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 12144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 19780 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform 1 0 4048 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 4416 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_E_FTB01 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22540 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01
timestamp 1649977179
transform -1 0 19780 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1649977179
transform 1 0 22632 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01
timestamp 1649977179
transform -1 0 2392 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  repeater80
timestamp 1649977179
transform -1 0 20148 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater81
timestamp 1649977179
transform -1 0 23000 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater82
timestamp 1649977179
transform -1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater83
timestamp 1649977179
transform -1 0 14536 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater84
timestamp 1649977179
transform 1 0 9476 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater85
timestamp 1649977179
transform -1 0 9476 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater86
timestamp 1649977179
transform -1 0 19044 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater87
timestamp 1649977179
transform -1 0 22908 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater88
timestamp 1649977179
transform 1 0 16008 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater89
timestamp 1649977179
transform -1 0 12144 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater90
timestamp 1649977179
transform -1 0 11316 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater91
timestamp 1649977179
transform -1 0 10488 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater92
timestamp 1649977179
transform -1 0 4140 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater93
timestamp 1649977179
transform -1 0 7176 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater94
timestamp 1649977179
transform -1 0 6716 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater95
timestamp 1649977179
transform -1 0 6624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater96
timestamp 1649977179
transform -1 0 9476 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater97 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17204 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater98
timestamp 1649977179
transform 1 0 18032 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater99
timestamp 1649977179
transform -1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater100
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater101
timestamp 1649977179
transform 1 0 5888 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater102
timestamp 1649977179
transform -1 0 8556 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater103
timestamp 1649977179
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater104
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 406 592
<< labels >>
rlabel metal2 s 17038 23800 17094 24600 6 SC_IN_TOP
port 0 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 SC_OUT_BOT
port 1 nsew signal tristate
rlabel metal2 s 17682 23800 17738 24600 6 SC_OUT_TOP
port 2 nsew signal tristate
rlabel metal3 s 23800 6808 24600 6928 6 Test_en_E_in
port 3 nsew signal input
rlabel metal3 s 23800 6264 24600 6384 6 Test_en_E_out
port 4 nsew signal tristate
rlabel metal3 s 0 21360 800 21480 6 Test_en_W_in
port 5 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 Test_en_W_out
port 6 nsew signal tristate
rlabel metal4 s 6542 2128 6862 22352 6 VGND
port 7 nsew ground input
rlabel metal4 s 12140 2128 12460 22352 6 VGND
port 7 nsew ground input
rlabel metal4 s 17738 2128 18058 22352 6 VGND
port 7 nsew ground input
rlabel metal4 s 3743 2128 4063 22352 6 VPWR
port 8 nsew power input
rlabel metal4 s 9341 2128 9661 22352 6 VPWR
port 8 nsew power input
rlabel metal4 s 14939 2128 15259 22352 6 VPWR
port 8 nsew power input
rlabel metal4 s 20537 2128 20857 22352 6 VPWR
port 8 nsew power input
rlabel metal2 s 2042 0 2098 800 6 bottom_width_0_height_0__pin_50_
port 9 nsew signal tristate
rlabel metal2 s 6090 0 6146 800 6 bottom_width_0_height_0__pin_51_
port 10 nsew signal tristate
rlabel metal3 s 0 9120 800 9240 6 ccff_head
port 11 nsew signal input
rlabel metal3 s 23800 5584 24600 5704 6 ccff_tail
port 12 nsew signal tristate
rlabel metal2 s 18326 23800 18382 24600 6 clk_0_N_in
port 13 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 clk_0_S_in
port 14 nsew signal input
rlabel metal3 s 23800 8168 24600 8288 6 prog_clk_0_E_out
port 15 nsew signal tristate
rlabel metal3 s 23800 7488 24600 7608 6 prog_clk_0_N_in
port 16 nsew signal input
rlabel metal2 s 18970 23800 19026 24600 6 prog_clk_0_N_out
port 17 nsew signal tristate
rlabel metal2 s 18418 0 18474 800 6 prog_clk_0_S_in
port 18 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 prog_clk_0_S_out
port 19 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 prog_clk_0_W_out
port 20 nsew signal tristate
rlabel metal3 s 23800 8848 24600 8968 6 right_width_0_height_0__pin_16_
port 21 nsew signal input
rlabel metal3 s 23800 9528 24600 9648 6 right_width_0_height_0__pin_17_
port 22 nsew signal input
rlabel metal3 s 23800 10208 24600 10328 6 right_width_0_height_0__pin_18_
port 23 nsew signal input
rlabel metal3 s 23800 10888 24600 11008 6 right_width_0_height_0__pin_19_
port 24 nsew signal input
rlabel metal3 s 23800 11568 24600 11688 6 right_width_0_height_0__pin_20_
port 25 nsew signal input
rlabel metal3 s 23800 12248 24600 12368 6 right_width_0_height_0__pin_21_
port 26 nsew signal input
rlabel metal3 s 23800 12792 24600 12912 6 right_width_0_height_0__pin_22_
port 27 nsew signal input
rlabel metal3 s 23800 13472 24600 13592 6 right_width_0_height_0__pin_23_
port 28 nsew signal input
rlabel metal3 s 23800 14152 24600 14272 6 right_width_0_height_0__pin_24_
port 29 nsew signal input
rlabel metal3 s 23800 14832 24600 14952 6 right_width_0_height_0__pin_25_
port 30 nsew signal input
rlabel metal3 s 23800 15512 24600 15632 6 right_width_0_height_0__pin_26_
port 31 nsew signal input
rlabel metal3 s 23800 16192 24600 16312 6 right_width_0_height_0__pin_27_
port 32 nsew signal input
rlabel metal3 s 23800 16872 24600 16992 6 right_width_0_height_0__pin_28_
port 33 nsew signal input
rlabel metal3 s 23800 17552 24600 17672 6 right_width_0_height_0__pin_29_
port 34 nsew signal input
rlabel metal3 s 23800 18232 24600 18352 6 right_width_0_height_0__pin_30_
port 35 nsew signal input
rlabel metal3 s 23800 18776 24600 18896 6 right_width_0_height_0__pin_31_
port 36 nsew signal input
rlabel metal3 s 23800 280 24600 400 6 right_width_0_height_0__pin_42_lower
port 37 nsew signal tristate
rlabel metal3 s 23800 19456 24600 19576 6 right_width_0_height_0__pin_42_upper
port 38 nsew signal tristate
rlabel metal3 s 23800 824 24600 944 6 right_width_0_height_0__pin_43_lower
port 39 nsew signal tristate
rlabel metal3 s 23800 20136 24600 20256 6 right_width_0_height_0__pin_43_upper
port 40 nsew signal tristate
rlabel metal3 s 23800 1504 24600 1624 6 right_width_0_height_0__pin_44_lower
port 41 nsew signal tristate
rlabel metal3 s 23800 20816 24600 20936 6 right_width_0_height_0__pin_44_upper
port 42 nsew signal tristate
rlabel metal3 s 23800 2184 24600 2304 6 right_width_0_height_0__pin_45_lower
port 43 nsew signal tristate
rlabel metal3 s 23800 21496 24600 21616 6 right_width_0_height_0__pin_45_upper
port 44 nsew signal tristate
rlabel metal3 s 23800 2864 24600 2984 6 right_width_0_height_0__pin_46_lower
port 45 nsew signal tristate
rlabel metal3 s 23800 22176 24600 22296 6 right_width_0_height_0__pin_46_upper
port 46 nsew signal tristate
rlabel metal3 s 23800 3544 24600 3664 6 right_width_0_height_0__pin_47_lower
port 47 nsew signal tristate
rlabel metal3 s 23800 22856 24600 22976 6 right_width_0_height_0__pin_47_upper
port 48 nsew signal tristate
rlabel metal3 s 23800 4224 24600 4344 6 right_width_0_height_0__pin_48_lower
port 49 nsew signal tristate
rlabel metal3 s 23800 23536 24600 23656 6 right_width_0_height_0__pin_48_upper
port 50 nsew signal tristate
rlabel metal3 s 23800 4904 24600 5024 6 right_width_0_height_0__pin_49_lower
port 51 nsew signal tristate
rlabel metal3 s 23800 24216 24600 24336 6 right_width_0_height_0__pin_49_upper
port 52 nsew signal tristate
rlabel metal2 s 5446 23800 5502 24600 6 top_width_0_height_0__pin_0_
port 53 nsew signal input
rlabel metal2 s 11886 23800 11942 24600 6 top_width_0_height_0__pin_10_
port 54 nsew signal input
rlabel metal2 s 12530 23800 12586 24600 6 top_width_0_height_0__pin_11_
port 55 nsew signal input
rlabel metal2 s 13174 23800 13230 24600 6 top_width_0_height_0__pin_12_
port 56 nsew signal input
rlabel metal2 s 13818 23800 13874 24600 6 top_width_0_height_0__pin_13_
port 57 nsew signal input
rlabel metal2 s 14462 23800 14518 24600 6 top_width_0_height_0__pin_14_
port 58 nsew signal input
rlabel metal2 s 15106 23800 15162 24600 6 top_width_0_height_0__pin_15_
port 59 nsew signal input
rlabel metal2 s 6090 23800 6146 24600 6 top_width_0_height_0__pin_1_
port 60 nsew signal input
rlabel metal2 s 6734 23800 6790 24600 6 top_width_0_height_0__pin_2_
port 61 nsew signal input
rlabel metal2 s 15750 23800 15806 24600 6 top_width_0_height_0__pin_32_
port 62 nsew signal input
rlabel metal2 s 16394 23800 16450 24600 6 top_width_0_height_0__pin_33_
port 63 nsew signal input
rlabel metal2 s 19614 23800 19670 24600 6 top_width_0_height_0__pin_34_lower
port 64 nsew signal tristate
rlabel metal2 s 294 23800 350 24600 6 top_width_0_height_0__pin_34_upper
port 65 nsew signal tristate
rlabel metal2 s 20258 23800 20314 24600 6 top_width_0_height_0__pin_35_lower
port 66 nsew signal tristate
rlabel metal2 s 938 23800 994 24600 6 top_width_0_height_0__pin_35_upper
port 67 nsew signal tristate
rlabel metal2 s 20902 23800 20958 24600 6 top_width_0_height_0__pin_36_lower
port 68 nsew signal tristate
rlabel metal2 s 1582 23800 1638 24600 6 top_width_0_height_0__pin_36_upper
port 69 nsew signal tristate
rlabel metal2 s 21546 23800 21602 24600 6 top_width_0_height_0__pin_37_lower
port 70 nsew signal tristate
rlabel metal2 s 2226 23800 2282 24600 6 top_width_0_height_0__pin_37_upper
port 71 nsew signal tristate
rlabel metal2 s 22190 23800 22246 24600 6 top_width_0_height_0__pin_38_lower
port 72 nsew signal tristate
rlabel metal2 s 2870 23800 2926 24600 6 top_width_0_height_0__pin_38_upper
port 73 nsew signal tristate
rlabel metal2 s 22834 23800 22890 24600 6 top_width_0_height_0__pin_39_lower
port 74 nsew signal tristate
rlabel metal2 s 3514 23800 3570 24600 6 top_width_0_height_0__pin_39_upper
port 75 nsew signal tristate
rlabel metal2 s 7378 23800 7434 24600 6 top_width_0_height_0__pin_3_
port 76 nsew signal input
rlabel metal2 s 23478 23800 23534 24600 6 top_width_0_height_0__pin_40_lower
port 77 nsew signal tristate
rlabel metal2 s 4158 23800 4214 24600 6 top_width_0_height_0__pin_40_upper
port 78 nsew signal tristate
rlabel metal2 s 24122 23800 24178 24600 6 top_width_0_height_0__pin_41_lower
port 79 nsew signal tristate
rlabel metal2 s 4802 23800 4858 24600 6 top_width_0_height_0__pin_41_upper
port 80 nsew signal tristate
rlabel metal2 s 8022 23800 8078 24600 6 top_width_0_height_0__pin_4_
port 81 nsew signal input
rlabel metal2 s 8666 23800 8722 24600 6 top_width_0_height_0__pin_5_
port 82 nsew signal input
rlabel metal2 s 9310 23800 9366 24600 6 top_width_0_height_0__pin_6_
port 83 nsew signal input
rlabel metal2 s 9954 23800 10010 24600 6 top_width_0_height_0__pin_7_
port 84 nsew signal input
rlabel metal2 s 10598 23800 10654 24600 6 top_width_0_height_0__pin_8_
port 85 nsew signal input
rlabel metal2 s 11242 23800 11298 24600 6 top_width_0_height_0__pin_9_
port 86 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 24600 24600
<< end >>
