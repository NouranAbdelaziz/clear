VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO cby_2__1_
  CLASS BLOCK ;
  FOREIGN cby_2__1_ ;
  ORIGIN 0.000 0.000 ;
  SIZE 86.000 BY 100.000 ;
  PIN IO_ISOL_N
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 96.000 1.290 100.000 ;
    END
  END IO_ISOL_N
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 23.460 10.640 25.060 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 42.200 10.640 43.800 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.940 10.640 62.540 87.280 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.090 10.640 15.690 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 32.830 10.640 34.430 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 51.570 10.640 53.170 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 70.310 10.640 71.910 87.280 ;
    END
  END VPWR
  PIN ccff_head
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END ccff_head
  PIN ccff_tail
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 82.000 9.560 86.000 10.160 ;
    END
  END ccff_tail
  PIN chany_bottom_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END chany_bottom_in[0]
  PIN chany_bottom_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END chany_bottom_in[10]
  PIN chany_bottom_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.870 0.000 66.150 4.000 ;
    END
  END chany_bottom_in[11]
  PIN chany_bottom_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END chany_bottom_in[12]
  PIN chany_bottom_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END chany_bottom_in[13]
  PIN chany_bottom_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 0.000 72.590 4.000 ;
    END
  END chany_bottom_in[14]
  PIN chany_bottom_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END chany_bottom_in[15]
  PIN chany_bottom_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END chany_bottom_in[16]
  PIN chany_bottom_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 4.000 ;
    END
  END chany_bottom_in[17]
  PIN chany_bottom_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END chany_bottom_in[18]
  PIN chany_bottom_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END chany_bottom_in[19]
  PIN chany_bottom_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END chany_bottom_in[1]
  PIN chany_bottom_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END chany_bottom_in[2]
  PIN chany_bottom_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END chany_bottom_in[3]
  PIN chany_bottom_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 4.000 ;
    END
  END chany_bottom_in[4]
  PIN chany_bottom_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END chany_bottom_in[5]
  PIN chany_bottom_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END chany_bottom_in[6]
  PIN chany_bottom_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END chany_bottom_in[7]
  PIN chany_bottom_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END chany_bottom_in[8]
  PIN chany_bottom_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 4.000 ;
    END
  END chany_bottom_in[9]
  PIN chany_bottom_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.010 0.000 1.290 4.000 ;
    END
  END chany_bottom_out[0]
  PIN chany_bottom_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.710 0.000 21.990 4.000 ;
    END
  END chany_bottom_out[10]
  PIN chany_bottom_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END chany_bottom_out[11]
  PIN chany_bottom_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END chany_bottom_out[12]
  PIN chany_bottom_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END chany_bottom_out[13]
  PIN chany_bottom_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END chany_bottom_out[14]
  PIN chany_bottom_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END chany_bottom_out[15]
  PIN chany_bottom_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END chany_bottom_out[16]
  PIN chany_bottom_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END chany_bottom_out[17]
  PIN chany_bottom_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END chany_bottom_out[18]
  PIN chany_bottom_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END chany_bottom_out[19]
  PIN chany_bottom_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END chany_bottom_out[1]
  PIN chany_bottom_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 0.000 5.430 4.000 ;
    END
  END chany_bottom_out[2]
  PIN chany_bottom_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END chany_bottom_out[3]
  PIN chany_bottom_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.290 0.000 9.570 4.000 ;
    END
  END chany_bottom_out[4]
  PIN chany_bottom_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END chany_bottom_out[5]
  PIN chany_bottom_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END chany_bottom_out[6]
  PIN chany_bottom_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 4.000 ;
    END
  END chany_bottom_out[7]
  PIN chany_bottom_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 0.000 17.850 4.000 ;
    END
  END chany_bottom_out[8]
  PIN chany_bottom_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END chany_bottom_out[9]
  PIN chany_top_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.790 96.000 44.070 100.000 ;
    END
  END chany_top_in[0]
  PIN chany_top_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 96.000 64.770 100.000 ;
    END
  END chany_top_in[10]
  PIN chany_top_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 96.000 66.610 100.000 ;
    END
  END chany_top_in[11]
  PIN chany_top_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 96.000 68.450 100.000 ;
    END
  END chany_top_in[12]
  PIN chany_top_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 96.000 70.750 100.000 ;
    END
  END chany_top_in[13]
  PIN chany_top_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.310 96.000 72.590 100.000 ;
    END
  END chany_top_in[14]
  PIN chany_top_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 96.000 74.890 100.000 ;
    END
  END chany_top_in[15]
  PIN chany_top_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 96.000 76.730 100.000 ;
    END
  END chany_top_in[16]
  PIN chany_top_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 96.000 79.030 100.000 ;
    END
  END chany_top_in[17]
  PIN chany_top_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 96.000 80.870 100.000 ;
    END
  END chany_top_in[18]
  PIN chany_top_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 96.000 83.170 100.000 ;
    END
  END chany_top_in[19]
  PIN chany_top_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 96.000 45.910 100.000 ;
    END
  END chany_top_in[1]
  PIN chany_top_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.930 96.000 48.210 100.000 ;
    END
  END chany_top_in[2]
  PIN chany_top_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.770 96.000 50.050 100.000 ;
    END
  END chany_top_in[3]
  PIN chany_top_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.070 96.000 52.350 100.000 ;
    END
  END chany_top_in[4]
  PIN chany_top_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.910 96.000 54.190 100.000 ;
    END
  END chany_top_in[5]
  PIN chany_top_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.210 96.000 56.490 100.000 ;
    END
  END chany_top_in[6]
  PIN chany_top_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 96.000 58.330 100.000 ;
    END
  END chany_top_in[7]
  PIN chany_top_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 96.000 60.630 100.000 ;
    END
  END chany_top_in[8]
  PIN chany_top_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 96.000 62.470 100.000 ;
    END
  END chany_top_in[9]
  PIN chany_top_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.850 96.000 3.130 100.000 ;
    END
  END chany_top_out[0]
  PIN chany_top_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 96.000 23.370 100.000 ;
    END
  END chany_top_out[10]
  PIN chany_top_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 96.000 25.670 100.000 ;
    END
  END chany_top_out[11]
  PIN chany_top_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 96.000 27.510 100.000 ;
    END
  END chany_top_out[12]
  PIN chany_top_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 96.000 29.810 100.000 ;
    END
  END chany_top_out[13]
  PIN chany_top_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 31.370 96.000 31.650 100.000 ;
    END
  END chany_top_out[14]
  PIN chany_top_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 96.000 33.950 100.000 ;
    END
  END chany_top_out[15]
  PIN chany_top_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 96.000 35.790 100.000 ;
    END
  END chany_top_out[16]
  PIN chany_top_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 96.000 38.090 100.000 ;
    END
  END chany_top_out[17]
  PIN chany_top_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 96.000 39.930 100.000 ;
    END
  END chany_top_out[18]
  PIN chany_top_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 96.000 42.230 100.000 ;
    END
  END chany_top_out[19]
  PIN chany_top_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 96.000 4.970 100.000 ;
    END
  END chany_top_out[1]
  PIN chany_top_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 96.000 7.270 100.000 ;
    END
  END chany_top_out[2]
  PIN chany_top_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 96.000 9.110 100.000 ;
    END
  END chany_top_out[3]
  PIN chany_top_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 96.000 11.410 100.000 ;
    END
  END chany_top_out[4]
  PIN chany_top_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 96.000 13.250 100.000 ;
    END
  END chany_top_out[5]
  PIN chany_top_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.270 96.000 15.550 100.000 ;
    END
  END chany_top_out[6]
  PIN chany_top_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 96.000 17.390 100.000 ;
    END
  END chany_top_out[7]
  PIN chany_top_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 96.000 19.690 100.000 ;
    END
  END chany_top_out[8]
  PIN chany_top_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 96.000 21.530 100.000 ;
    END
  END chany_top_out[9]
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 82.000 49.000 86.000 49.600 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 82.000 69.400 86.000 70.000 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_IN
  PIN gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 82.000 89.120 86.000 89.720 ;
    END
  END gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
  PIN left_grid_pin_16_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END left_grid_pin_16_
  PIN left_grid_pin_17_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END left_grid_pin_17_
  PIN left_grid_pin_18_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.880 4.000 26.480 ;
    END
  END left_grid_pin_18_
  PIN left_grid_pin_19_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END left_grid_pin_19_
  PIN left_grid_pin_20_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END left_grid_pin_20_
  PIN left_grid_pin_21_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END left_grid_pin_21_
  PIN left_grid_pin_22_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END left_grid_pin_22_
  PIN left_grid_pin_23_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.680 4.000 50.280 ;
    END
  END left_grid_pin_23_
  PIN left_grid_pin_24_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END left_grid_pin_24_
  PIN left_grid_pin_25_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.200 4.000 59.800 ;
    END
  END left_grid_pin_25_
  PIN left_grid_pin_26_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END left_grid_pin_26_
  PIN left_grid_pin_27_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END left_grid_pin_27_
  PIN left_grid_pin_28_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 73.480 4.000 74.080 ;
    END
  END left_grid_pin_28_
  PIN left_grid_pin_29_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END left_grid_pin_29_
  PIN left_grid_pin_30_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END left_grid_pin_30_
  PIN left_grid_pin_31_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END left_grid_pin_31_
  PIN left_width_0_height_0__pin_0_
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END left_width_0_height_0__pin_0_
  PIN left_width_0_height_0__pin_1_lower
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END left_width_0_height_0__pin_1_lower
  PIN left_width_0_height_0__pin_1_upper
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END left_width_0_height_0__pin_1_upper
  PIN prog_clk_0_N_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 96.000 85.010 100.000 ;
    END
  END prog_clk_0_N_out
  PIN prog_clk_0_S_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END prog_clk_0_S_out
  PIN prog_clk_0_W_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END prog_clk_0_W_in
  PIN right_grid_pin_0_
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 82.000 29.280 86.000 29.880 ;
    END
  END right_grid_pin_0_
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 80.040 87.125 ;
      LAYER met1 ;
        RECT 0.990 7.860 85.030 88.360 ;
      LAYER met2 ;
        RECT 1.570 95.720 2.570 96.290 ;
        RECT 3.410 95.720 4.410 96.290 ;
        RECT 5.250 95.720 6.710 96.290 ;
        RECT 7.550 95.720 8.550 96.290 ;
        RECT 9.390 95.720 10.850 96.290 ;
        RECT 11.690 95.720 12.690 96.290 ;
        RECT 13.530 95.720 14.990 96.290 ;
        RECT 15.830 95.720 16.830 96.290 ;
        RECT 17.670 95.720 19.130 96.290 ;
        RECT 19.970 95.720 20.970 96.290 ;
        RECT 21.810 95.720 22.810 96.290 ;
        RECT 23.650 95.720 25.110 96.290 ;
        RECT 25.950 95.720 26.950 96.290 ;
        RECT 27.790 95.720 29.250 96.290 ;
        RECT 30.090 95.720 31.090 96.290 ;
        RECT 31.930 95.720 33.390 96.290 ;
        RECT 34.230 95.720 35.230 96.290 ;
        RECT 36.070 95.720 37.530 96.290 ;
        RECT 38.370 95.720 39.370 96.290 ;
        RECT 40.210 95.720 41.670 96.290 ;
        RECT 42.510 95.720 43.510 96.290 ;
        RECT 44.350 95.720 45.350 96.290 ;
        RECT 46.190 95.720 47.650 96.290 ;
        RECT 48.490 95.720 49.490 96.290 ;
        RECT 50.330 95.720 51.790 96.290 ;
        RECT 52.630 95.720 53.630 96.290 ;
        RECT 54.470 95.720 55.930 96.290 ;
        RECT 56.770 95.720 57.770 96.290 ;
        RECT 58.610 95.720 60.070 96.290 ;
        RECT 60.910 95.720 61.910 96.290 ;
        RECT 62.750 95.720 64.210 96.290 ;
        RECT 65.050 95.720 66.050 96.290 ;
        RECT 66.890 95.720 67.890 96.290 ;
        RECT 68.730 95.720 70.190 96.290 ;
        RECT 71.030 95.720 72.030 96.290 ;
        RECT 72.870 95.720 74.330 96.290 ;
        RECT 75.170 95.720 76.170 96.290 ;
        RECT 77.010 95.720 78.470 96.290 ;
        RECT 79.310 95.720 80.310 96.290 ;
        RECT 81.150 95.720 82.610 96.290 ;
        RECT 83.450 95.720 84.450 96.290 ;
        RECT 1.020 4.280 85.000 95.720 ;
        RECT 1.570 2.195 2.570 4.280 ;
        RECT 3.410 2.195 4.870 4.280 ;
        RECT 5.710 2.195 6.710 4.280 ;
        RECT 7.550 2.195 9.010 4.280 ;
        RECT 9.850 2.195 10.850 4.280 ;
        RECT 11.690 2.195 13.150 4.280 ;
        RECT 13.990 2.195 14.990 4.280 ;
        RECT 15.830 2.195 17.290 4.280 ;
        RECT 18.130 2.195 19.590 4.280 ;
        RECT 20.430 2.195 21.430 4.280 ;
        RECT 22.270 2.195 23.730 4.280 ;
        RECT 24.570 2.195 25.570 4.280 ;
        RECT 26.410 2.195 27.870 4.280 ;
        RECT 28.710 2.195 29.710 4.280 ;
        RECT 30.550 2.195 32.010 4.280 ;
        RECT 32.850 2.195 33.850 4.280 ;
        RECT 34.690 2.195 36.150 4.280 ;
        RECT 36.990 2.195 38.450 4.280 ;
        RECT 39.290 2.195 40.290 4.280 ;
        RECT 41.130 2.195 42.590 4.280 ;
        RECT 43.430 2.195 44.430 4.280 ;
        RECT 45.270 2.195 46.730 4.280 ;
        RECT 47.570 2.195 48.570 4.280 ;
        RECT 49.410 2.195 50.870 4.280 ;
        RECT 51.710 2.195 53.170 4.280 ;
        RECT 54.010 2.195 55.010 4.280 ;
        RECT 55.850 2.195 57.310 4.280 ;
        RECT 58.150 2.195 59.150 4.280 ;
        RECT 59.990 2.195 61.450 4.280 ;
        RECT 62.290 2.195 63.290 4.280 ;
        RECT 64.130 2.195 65.590 4.280 ;
        RECT 66.430 2.195 67.430 4.280 ;
        RECT 68.270 2.195 69.730 4.280 ;
        RECT 70.570 2.195 72.030 4.280 ;
        RECT 72.870 2.195 73.870 4.280 ;
        RECT 74.710 2.195 76.170 4.280 ;
        RECT 77.010 2.195 78.010 4.280 ;
        RECT 78.850 2.195 80.310 4.280 ;
        RECT 81.150 2.195 82.150 4.280 ;
        RECT 82.990 2.195 84.450 4.280 ;
      LAYER met3 ;
        RECT 4.400 96.880 82.000 97.730 ;
        RECT 4.000 93.520 82.000 96.880 ;
        RECT 4.400 92.120 82.000 93.520 ;
        RECT 4.000 90.120 82.000 92.120 ;
        RECT 4.000 88.760 81.600 90.120 ;
        RECT 4.400 88.720 81.600 88.760 ;
        RECT 4.400 87.360 82.000 88.720 ;
        RECT 4.000 84.000 82.000 87.360 ;
        RECT 4.400 82.600 82.000 84.000 ;
        RECT 4.000 79.240 82.000 82.600 ;
        RECT 4.400 77.840 82.000 79.240 ;
        RECT 4.000 74.480 82.000 77.840 ;
        RECT 4.400 73.080 82.000 74.480 ;
        RECT 4.000 70.400 82.000 73.080 ;
        RECT 4.000 69.720 81.600 70.400 ;
        RECT 4.400 69.000 81.600 69.720 ;
        RECT 4.400 68.320 82.000 69.000 ;
        RECT 4.000 64.960 82.000 68.320 ;
        RECT 4.400 63.560 82.000 64.960 ;
        RECT 4.000 60.200 82.000 63.560 ;
        RECT 4.400 58.800 82.000 60.200 ;
        RECT 4.000 55.440 82.000 58.800 ;
        RECT 4.400 54.040 82.000 55.440 ;
        RECT 4.000 50.680 82.000 54.040 ;
        RECT 4.400 50.000 82.000 50.680 ;
        RECT 4.400 49.280 81.600 50.000 ;
        RECT 4.000 48.600 81.600 49.280 ;
        RECT 4.000 45.920 82.000 48.600 ;
        RECT 4.400 44.520 82.000 45.920 ;
        RECT 4.000 41.160 82.000 44.520 ;
        RECT 4.400 39.760 82.000 41.160 ;
        RECT 4.000 36.400 82.000 39.760 ;
        RECT 4.400 35.000 82.000 36.400 ;
        RECT 4.000 31.640 82.000 35.000 ;
        RECT 4.400 30.280 82.000 31.640 ;
        RECT 4.400 30.240 81.600 30.280 ;
        RECT 4.000 28.880 81.600 30.240 ;
        RECT 4.000 26.880 82.000 28.880 ;
        RECT 4.400 25.480 82.000 26.880 ;
        RECT 4.000 22.120 82.000 25.480 ;
        RECT 4.400 20.720 82.000 22.120 ;
        RECT 4.000 17.360 82.000 20.720 ;
        RECT 4.400 15.960 82.000 17.360 ;
        RECT 4.000 12.600 82.000 15.960 ;
        RECT 4.400 11.200 82.000 12.600 ;
        RECT 4.000 10.560 82.000 11.200 ;
        RECT 4.000 9.160 81.600 10.560 ;
        RECT 4.000 7.840 82.000 9.160 ;
        RECT 4.400 6.440 82.000 7.840 ;
        RECT 4.000 3.080 82.000 6.440 ;
        RECT 4.400 2.215 82.000 3.080 ;
      LAYER met4 ;
        RECT 7.655 11.735 13.690 86.185 ;
        RECT 16.090 11.735 23.060 86.185 ;
        RECT 25.460 11.735 32.430 86.185 ;
        RECT 34.830 11.735 41.800 86.185 ;
        RECT 44.200 11.735 51.170 86.185 ;
        RECT 53.570 11.735 60.540 86.185 ;
        RECT 62.940 11.735 69.910 86.185 ;
        RECT 72.310 11.735 75.145 86.185 ;
  END
END cby_2__1_
END LIBRARY

