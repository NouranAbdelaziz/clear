module sb_1__1_ (Test_en_N_out,
    Test_en_S_in,
    VGND,
    VPWR,
    bottom_left_grid_pin_42_,
    bottom_left_grid_pin_43_,
    bottom_left_grid_pin_44_,
    bottom_left_grid_pin_45_,
    bottom_left_grid_pin_46_,
    bottom_left_grid_pin_47_,
    bottom_left_grid_pin_48_,
    bottom_left_grid_pin_49_,
    ccff_head,
    ccff_tail,
    clk_1_E_out,
    clk_1_N_in,
    clk_1_W_out,
    clk_2_E_out,
    clk_2_N_in,
    clk_2_N_out,
    clk_2_S_out,
    clk_2_W_out,
    clk_3_E_out,
    clk_3_N_in,
    clk_3_N_out,
    clk_3_S_out,
    clk_3_W_out,
    left_bottom_grid_pin_34_,
    left_bottom_grid_pin_35_,
    left_bottom_grid_pin_36_,
    left_bottom_grid_pin_37_,
    left_bottom_grid_pin_38_,
    left_bottom_grid_pin_39_,
    left_bottom_grid_pin_40_,
    left_bottom_grid_pin_41_,
    prog_clk_0_N_in,
    prog_clk_1_E_out,
    prog_clk_1_N_in,
    prog_clk_1_W_out,
    prog_clk_2_E_out,
    prog_clk_2_N_in,
    prog_clk_2_N_out,
    prog_clk_2_S_out,
    prog_clk_2_W_out,
    prog_clk_3_E_out,
    prog_clk_3_N_in,
    prog_clk_3_N_out,
    prog_clk_3_S_out,
    prog_clk_3_W_out,
    right_bottom_grid_pin_34_,
    right_bottom_grid_pin_35_,
    right_bottom_grid_pin_36_,
    right_bottom_grid_pin_37_,
    right_bottom_grid_pin_38_,
    right_bottom_grid_pin_39_,
    right_bottom_grid_pin_40_,
    right_bottom_grid_pin_41_,
    top_left_grid_pin_42_,
    top_left_grid_pin_43_,
    top_left_grid_pin_44_,
    top_left_grid_pin_45_,
    top_left_grid_pin_46_,
    top_left_grid_pin_47_,
    top_left_grid_pin_48_,
    top_left_grid_pin_49_,
    chanx_left_in,
    chanx_left_out,
    chanx_right_in,
    chanx_right_out,
    chany_bottom_in,
    chany_bottom_out,
    chany_top_in,
    chany_top_out);
 output Test_en_N_out;
 inout Test_en_S_in;
 inout VGND;
 inout VPWR;
 inout bottom_left_grid_pin_42_;
 inout bottom_left_grid_pin_43_;
 inout bottom_left_grid_pin_44_;
 inout bottom_left_grid_pin_45_;
 inout bottom_left_grid_pin_46_;
 inout bottom_left_grid_pin_47_;
 inout bottom_left_grid_pin_48_;
 inout bottom_left_grid_pin_49_;
 inout ccff_head;
 output ccff_tail;
 output clk_1_E_out;
 inout clk_1_N_in;
 output clk_1_W_out;
 output clk_2_E_out;
 inout clk_2_N_in;
 output clk_2_N_out;
 output clk_2_S_out;
 output clk_2_W_out;
 output clk_3_E_out;
 inout clk_3_N_in;
 output clk_3_N_out;
 output clk_3_S_out;
 output clk_3_W_out;
 inout left_bottom_grid_pin_34_;
 inout left_bottom_grid_pin_35_;
 inout left_bottom_grid_pin_36_;
 inout left_bottom_grid_pin_37_;
 inout left_bottom_grid_pin_38_;
 inout left_bottom_grid_pin_39_;
 inout left_bottom_grid_pin_40_;
 inout left_bottom_grid_pin_41_;
 inout prog_clk_0_N_in;
 output prog_clk_1_E_out;
 inout prog_clk_1_N_in;
 output prog_clk_1_W_out;
 output prog_clk_2_E_out;
 inout prog_clk_2_N_in;
 output prog_clk_2_N_out;
 output prog_clk_2_S_out;
 output prog_clk_2_W_out;
 output prog_clk_3_E_out;
 inout prog_clk_3_N_in;
 output prog_clk_3_N_out;
 output prog_clk_3_S_out;
 output prog_clk_3_W_out;
 inout right_bottom_grid_pin_34_;
 inout right_bottom_grid_pin_35_;
 inout right_bottom_grid_pin_36_;
 inout right_bottom_grid_pin_37_;
 inout right_bottom_grid_pin_38_;
 inout right_bottom_grid_pin_39_;
 inout right_bottom_grid_pin_40_;
 inout right_bottom_grid_pin_41_;
 inout top_left_grid_pin_42_;
 inout top_left_grid_pin_43_;
 inout top_left_grid_pin_44_;
 inout top_left_grid_pin_45_;
 inout top_left_grid_pin_46_;
 inout top_left_grid_pin_47_;
 inout top_left_grid_pin_48_;
 inout top_left_grid_pin_49_;
 inout [19:0] chanx_left_in;
 output [19:0] chanx_left_out;
 inout [19:0] chanx_right_in;
 output [19:0] chanx_right_out;
 inout [19:0] chany_bottom_in;
 output [19:0] chany_bottom_out;
 inout [19:0] chany_top_in;
 output [19:0] chany_top_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire \clknet_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_1_0_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_1_1_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_2_0_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_2_1_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_2_2_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_2_3_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_0_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_1_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_2_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_3_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_4_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_5_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_6_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_7_0_mem_bottom_track_1.prog_clk ;
 wire \mem_bottom_track_1.ccff_head ;
 wire \mem_bottom_track_1.ccff_tail ;
 wire \mem_bottom_track_1.mem_out[0] ;
 wire \mem_bottom_track_1.mem_out[1] ;
 wire \mem_bottom_track_1.mem_out[2] ;
 wire \mem_bottom_track_1.prog_clk ;
 wire \mem_bottom_track_17.ccff_head ;
 wire \mem_bottom_track_17.ccff_tail ;
 wire \mem_bottom_track_17.mem_out[0] ;
 wire \mem_bottom_track_17.mem_out[1] ;
 wire \mem_bottom_track_17.mem_out[2] ;
 wire \mem_bottom_track_25.ccff_tail ;
 wire \mem_bottom_track_25.mem_out[0] ;
 wire \mem_bottom_track_25.mem_out[1] ;
 wire \mem_bottom_track_25.mem_out[2] ;
 wire \mem_bottom_track_3.ccff_tail ;
 wire \mem_bottom_track_3.mem_out[0] ;
 wire \mem_bottom_track_3.mem_out[1] ;
 wire \mem_bottom_track_3.mem_out[2] ;
 wire \mem_bottom_track_33.ccff_tail ;
 wire \mem_bottom_track_33.mem_out[0] ;
 wire \mem_bottom_track_33.mem_out[1] ;
 wire \mem_bottom_track_5.ccff_tail ;
 wire \mem_bottom_track_5.mem_out[0] ;
 wire \mem_bottom_track_5.mem_out[1] ;
 wire \mem_bottom_track_5.mem_out[2] ;
 wire \mem_bottom_track_5.mem_out[3] ;
 wire \mem_bottom_track_9.mem_out[0] ;
 wire \mem_bottom_track_9.mem_out[1] ;
 wire \mem_bottom_track_9.mem_out[2] ;
 wire \mem_left_track_1.ccff_tail ;
 wire \mem_left_track_1.mem_out[0] ;
 wire \mem_left_track_1.mem_out[1] ;
 wire \mem_left_track_1.mem_out[2] ;
 wire \mem_left_track_17.ccff_head ;
 wire \mem_left_track_17.ccff_tail ;
 wire \mem_left_track_17.mem_out[0] ;
 wire \mem_left_track_17.mem_out[1] ;
 wire \mem_left_track_17.mem_out[2] ;
 wire \mem_left_track_25.ccff_tail ;
 wire \mem_left_track_25.mem_out[0] ;
 wire \mem_left_track_25.mem_out[1] ;
 wire \mem_left_track_25.mem_out[2] ;
 wire \mem_left_track_3.ccff_tail ;
 wire \mem_left_track_3.mem_out[0] ;
 wire \mem_left_track_3.mem_out[1] ;
 wire \mem_left_track_3.mem_out[2] ;
 wire \mem_left_track_33.mem_out[0] ;
 wire \mem_left_track_33.mem_out[1] ;
 wire \mem_left_track_5.ccff_tail ;
 wire \mem_left_track_5.mem_out[0] ;
 wire \mem_left_track_5.mem_out[1] ;
 wire \mem_left_track_5.mem_out[2] ;
 wire \mem_left_track_5.mem_out[3] ;
 wire \mem_left_track_9.mem_out[0] ;
 wire \mem_left_track_9.mem_out[1] ;
 wire \mem_left_track_9.mem_out[2] ;
 wire \mem_right_track_0.ccff_head ;
 wire \mem_right_track_0.ccff_tail ;
 wire \mem_right_track_0.mem_out[0] ;
 wire \mem_right_track_0.mem_out[1] ;
 wire \mem_right_track_0.mem_out[2] ;
 wire \mem_right_track_16.ccff_head ;
 wire \mem_right_track_16.ccff_tail ;
 wire \mem_right_track_16.mem_out[0] ;
 wire \mem_right_track_16.mem_out[1] ;
 wire \mem_right_track_16.mem_out[2] ;
 wire \mem_right_track_2.ccff_tail ;
 wire \mem_right_track_2.mem_out[0] ;
 wire \mem_right_track_2.mem_out[1] ;
 wire \mem_right_track_2.mem_out[2] ;
 wire \mem_right_track_24.ccff_tail ;
 wire \mem_right_track_24.mem_out[0] ;
 wire \mem_right_track_24.mem_out[1] ;
 wire \mem_right_track_24.mem_out[2] ;
 wire \mem_right_track_32.mem_out[0] ;
 wire \mem_right_track_32.mem_out[1] ;
 wire \mem_right_track_4.ccff_tail ;
 wire \mem_right_track_4.mem_out[0] ;
 wire \mem_right_track_4.mem_out[1] ;
 wire \mem_right_track_4.mem_out[2] ;
 wire \mem_right_track_4.mem_out[3] ;
 wire \mem_right_track_8.mem_out[0] ;
 wire \mem_right_track_8.mem_out[1] ;
 wire \mem_right_track_8.mem_out[2] ;
 wire \mem_top_track_0.ccff_tail ;
 wire \mem_top_track_0.mem_out[0] ;
 wire \mem_top_track_0.mem_out[1] ;
 wire \mem_top_track_0.mem_out[2] ;
 wire \mem_top_track_16.ccff_head ;
 wire \mem_top_track_16.ccff_tail ;
 wire \mem_top_track_16.mem_out[0] ;
 wire \mem_top_track_16.mem_out[1] ;
 wire \mem_top_track_16.mem_out[2] ;
 wire \mem_top_track_2.ccff_tail ;
 wire \mem_top_track_2.mem_out[0] ;
 wire \mem_top_track_2.mem_out[1] ;
 wire \mem_top_track_2.mem_out[2] ;
 wire \mem_top_track_24.ccff_tail ;
 wire \mem_top_track_24.mem_out[0] ;
 wire \mem_top_track_24.mem_out[1] ;
 wire \mem_top_track_24.mem_out[2] ;
 wire \mem_top_track_32.mem_out[0] ;
 wire \mem_top_track_32.mem_out[1] ;
 wire \mem_top_track_4.ccff_tail ;
 wire \mem_top_track_4.mem_out[0] ;
 wire \mem_top_track_4.mem_out[1] ;
 wire \mem_top_track_4.mem_out[2] ;
 wire \mem_top_track_4.mem_out[3] ;
 wire \mem_top_track_8.mem_out[0] ;
 wire \mem_top_track_8.mem_out[1] ;
 wire \mem_top_track_8.mem_out[2] ;
 wire \mux_bottom_track_1.out ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_10_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_11_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_bottom_track_17.out ;
 wire \mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_bottom_track_25.out ;
 wire \mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_bottom_track_3.out ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_10_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_11_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_bottom_track_33.out ;
 wire \mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_bottom_track_5.out ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_10_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_11_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_12_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_13_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_14_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_15_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_bottom_track_9.out ;
 wire \mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_left_track_1.out ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_10_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_11_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_left_track_17.out ;
 wire \mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_17.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_left_track_17.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_left_track_17.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_left_track_17.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_left_track_17.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_left_track_17.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_left_track_17.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_left_track_17.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_left_track_25.out ;
 wire \mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_25.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_left_track_25.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_left_track_25.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_left_track_25.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_left_track_25.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_left_track_25.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_left_track_25.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_left_track_25.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_left_track_3.out ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_10_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_11_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_left_track_33.out ;
 wire \mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_33.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_left_track_33.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_left_track_33.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_left_track_33.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_left_track_33.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_left_track_5.out ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_10_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_11_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_12_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_13_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_14_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_15_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_left_track_9.out ;
 wire \mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_left_track_9.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_left_track_9.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_left_track_9.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_left_track_9.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_left_track_9.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_left_track_9.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_left_track_9.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_right_track_0.out ;
 wire \mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_right_track_0.sky130_fd_sc_hd__mux2_1_10_X ;
 wire \mux_right_track_0.sky130_fd_sc_hd__mux2_1_11_X ;
 wire \mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_right_track_0.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_right_track_0.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_right_track_0.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_right_track_0.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_right_track_16.out ;
 wire \mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_right_track_16.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_right_track_16.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_right_track_16.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_right_track_16.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_right_track_16.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_right_track_16.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_right_track_2.out ;
 wire \mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_right_track_2.sky130_fd_sc_hd__mux2_1_10_X ;
 wire \mux_right_track_2.sky130_fd_sc_hd__mux2_1_11_X ;
 wire \mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_right_track_2.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_right_track_2.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_right_track_2.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_right_track_2.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_right_track_24.out ;
 wire \mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_right_track_24.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_right_track_24.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_right_track_24.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_right_track_24.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_right_track_24.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_right_track_24.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_right_track_24.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_right_track_32.out ;
 wire \mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_right_track_32.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_right_track_32.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_right_track_32.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_right_track_32.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_right_track_4.out ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_10_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_11_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_12_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_13_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_14_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_15_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_right_track_4.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_right_track_8.out ;
 wire \mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_right_track_8.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_right_track_8.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_right_track_8.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_right_track_8.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_top_track_0.out ;
 wire \mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_top_track_0.sky130_fd_sc_hd__mux2_1_10_X ;
 wire \mux_top_track_0.sky130_fd_sc_hd__mux2_1_11_X ;
 wire \mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_top_track_0.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_top_track_0.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_top_track_0.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_top_track_16.out ;
 wire \mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_top_track_16.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_top_track_16.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_top_track_16.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_top_track_16.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_top_track_16.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_top_track_16.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_top_track_2.out ;
 wire \mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_top_track_2.sky130_fd_sc_hd__mux2_1_10_X ;
 wire \mux_top_track_2.sky130_fd_sc_hd__mux2_1_11_X ;
 wire \mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_top_track_2.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_top_track_2.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_top_track_2.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_top_track_2.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_top_track_24.out ;
 wire \mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_top_track_24.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_top_track_24.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_top_track_24.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_top_track_24.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_top_track_24.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_top_track_24.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_top_track_24.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_top_track_32.out ;
 wire \mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_top_track_32.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_top_track_32.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_top_track_32.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_top_track_32.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_top_track_32.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_top_track_4.out ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_10_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_11_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_12_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_13_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_14_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_15_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_top_track_4.sky130_fd_sc_hd__mux2_1_9_X ;
 wire \mux_top_track_8.out ;
 wire \mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_top_track_8.sky130_fd_sc_hd__mux2_1_6_X ;
 wire \mux_top_track_8.sky130_fd_sc_hd__mux2_1_7_X ;
 wire \mux_top_track_8.sky130_fd_sc_hd__mux2_1_8_X ;
 wire \mux_top_track_8.sky130_fd_sc_hd__mux2_1_9_X ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA__059__A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA__061__A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA__062__A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA__063__A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA__065__A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA__066__A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA__067__A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__069__A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__070__A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__071__A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__073__A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__074__A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__075__A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__079__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__081__A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__082__A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__083__A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__085__A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__086__A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__087__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__089__A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__090__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__091__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__093__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__094__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__095__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__099__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__101__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__102__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__103__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__105__A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__106__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__107__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__109__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__110__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__111__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__113__A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__114__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__115__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__119__A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA__121__A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__122__A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__123__A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__125__A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__126__A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__127__A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA__129__A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA__130__A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA__131__A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA__133__A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA__134__A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA__135__A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(left_bottom_grid_pin_40_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input101_A (.DIODE(left_bottom_grid_pin_41_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input102_A (.DIODE(prog_clk_0_N_in));
 sky130_fd_sc_hd__diode_2 ANTENNA_input103_A (.DIODE(prog_clk_1_N_in));
 sky130_fd_sc_hd__diode_2 ANTENNA_input104_A (.DIODE(prog_clk_3_N_in));
 sky130_fd_sc_hd__diode_2 ANTENNA_input105_A (.DIODE(right_bottom_grid_pin_34_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input106_A (.DIODE(right_bottom_grid_pin_35_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input107_A (.DIODE(right_bottom_grid_pin_36_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input108_A (.DIODE(right_bottom_grid_pin_37_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input109_A (.DIODE(right_bottom_grid_pin_38_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(ccff_head));
 sky130_fd_sc_hd__diode_2 ANTENNA_input110_A (.DIODE(right_bottom_grid_pin_39_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input111_A (.DIODE(right_bottom_grid_pin_40_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input112_A (.DIODE(right_bottom_grid_pin_41_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input113_A (.DIODE(top_left_grid_pin_42_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input114_A (.DIODE(top_left_grid_pin_43_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input115_A (.DIODE(top_left_grid_pin_44_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input116_A (.DIODE(top_left_grid_pin_45_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input117_A (.DIODE(top_left_grid_pin_46_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input118_A (.DIODE(top_left_grid_pin_47_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input119_A (.DIODE(top_left_grid_pin_48_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(chanx_left_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input120_A (.DIODE(top_left_grid_pin_49_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(chanx_left_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(chanx_left_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(chanx_left_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(chanx_left_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(chanx_left_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(chanx_left_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(chanx_left_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(chanx_left_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(Test_en_S_in));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(chanx_left_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(chanx_left_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(chanx_left_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(chanx_left_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(chanx_left_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(chanx_left_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(chanx_left_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(chanx_left_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(chanx_left_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(chanx_left_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(bottom_left_grid_pin_42_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(chanx_left_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(chanx_right_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(chanx_right_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(chanx_right_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(chanx_right_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(chanx_right_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(chanx_right_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(chanx_right_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(chanx_right_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(chanx_right_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(bottom_left_grid_pin_43_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(chanx_right_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(chanx_right_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(chanx_right_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(chanx_right_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(chanx_right_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(chanx_right_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(chanx_right_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(chanx_right_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(chanx_right_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(chanx_right_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(bottom_left_grid_pin_44_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(chanx_right_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(chany_bottom_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(chany_bottom_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(chany_bottom_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(chany_bottom_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(chany_bottom_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(chany_bottom_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(chany_bottom_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(chany_bottom_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(chany_bottom_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(bottom_left_grid_pin_45_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(chany_bottom_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(chany_bottom_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(chany_bottom_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(chany_bottom_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(chany_bottom_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(chany_bottom_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(chany_bottom_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(chany_bottom_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(chany_bottom_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(chany_bottom_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(bottom_left_grid_pin_46_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(chany_bottom_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(chany_top_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(chany_top_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(chany_top_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(chany_top_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(chany_top_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(chany_top_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(chany_top_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(chany_top_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(chany_top_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(bottom_left_grid_pin_47_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(chany_top_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(chany_top_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(chany_top_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(chany_top_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(chany_top_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(chany_top_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(chany_top_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(chany_top_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(chany_top_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(chany_top_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(bottom_left_grid_pin_48_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(chany_top_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(clk_1_N_in));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(clk_2_N_in));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(clk_3_N_in));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(left_bottom_grid_pin_34_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(left_bottom_grid_pin_35_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(left_bottom_grid_pin_36_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(left_bottom_grid_pin_37_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(left_bottom_grid_pin_38_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(left_bottom_grid_pin_39_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(bottom_left_grid_pin_49_));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0  (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1  (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1  (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1  (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1  (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_1.mux_l1_in_4__A0  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0  (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1  (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0  (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1  (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0  (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0  (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1  (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_17.mux_l2_in_2__A1  (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_17.mux_l2_in_3__A1  (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0  (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0  (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0  (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_25.mux_l2_in_2__A0  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_25.mux_l2_in_2__A1  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0  (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1  (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0  (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1  (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0  (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1  (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_3.mux_l1_in_4__A0  (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0  (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1  (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_33.mux_l1_in_3__A1  (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0  (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0  (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1  (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_5.mux_l2_in_6__A1  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_5.mux_l2_in_7__A1  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0  (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0  (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1  (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_1.mux_l1_in_0__A0  (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_1.mux_l1_in_0__A1  (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_1.mux_l1_in_1__A0  (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_1.mux_l1_in_1__A1  (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_1.mux_l1_in_2__A0  (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_1.mux_l1_in_2__A1  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_1.mux_l1_in_3__A1  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_17.mux_l1_in_0__A0  (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_17.mux_l1_in_0__A1  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_17.mux_l1_in_1__A0  (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_17.mux_l1_in_1__A1  (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_17.mux_l1_in_2__A1  (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_17.mux_l2_in_1__A0  (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_17.mux_l2_in_2__A1  (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_25.mux_l1_in_0__A0  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_25.mux_l1_in_0__A1  (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_25.mux_l1_in_1__A0  (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_25.mux_l1_in_1__A1  (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_25.mux_l1_in_2__A0  (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_25.mux_l1_in_2__A1  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_25.mux_l2_in_2__A1  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_3.mux_l1_in_0__A0  (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_3.mux_l1_in_0__A1  (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_3.mux_l1_in_1__A0  (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_3.mux_l1_in_1__A1  (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_3.mux_l1_in_2__A0  (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_3.mux_l1_in_2__A1  (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_3.mux_l1_in_3__A0  (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_3.mux_l1_in_3__A1  (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_33.mux_l1_in_0__A0  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_33.mux_l1_in_0__A1  (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_33.mux_l1_in_1__A0  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_33.mux_l1_in_1__A1  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_5.mux_l1_in_0__A0  (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_5.mux_l1_in_0__A1  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_5.mux_l2_in_0__A0  (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_5.mux_l2_in_1__A0  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_5.mux_l2_in_1__A1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_5.mux_l2_in_2__A0  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_5.mux_l2_in_2__A1  (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_5.mux_l2_in_3__A1  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_9.mux_l1_in_0__A1  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_9.mux_l1_in_1__A0  (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_9.mux_l1_in_1__A1  (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_9.mux_l1_in_2__A0  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_9.mux_l1_in_2__A1  (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_9.mux_l2_in_1__A0  (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_9.mux_l2_in_2__A1  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_0.mux_l1_in_0__A0  (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_0.mux_l1_in_0__A1  (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_0.mux_l1_in_1__A1  (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_0.mux_l1_in_3__A0  (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_0.mux_l1_in_4__A1  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_0.mux_l2_in_2__A0  (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_0.mux_l2_in_3__A1  (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_16.mux_l1_in_0__A0  (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_16.mux_l1_in_0__A1  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_16.mux_l1_in_1__A1  (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_16.mux_l1_in_2__A0  (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_16.mux_l2_in_1__A0  (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_16.mux_l2_in_2__A0  (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_16.mux_l2_in_2__A1  (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_16.mux_l2_in_3__A1  (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_2.mux_l1_in_0__A0  (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_2.mux_l1_in_0__A1  (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_2.mux_l1_in_1__A1  (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_2.mux_l1_in_3__A0  (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_2.mux_l1_in_4__A0  (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_2.mux_l2_in_2__A0  (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_2.mux_l2_in_3__A1  (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_24.mux_l1_in_0__A1  (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_24.mux_l1_in_1__A1  (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_24.mux_l1_in_2__A0  (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_24.mux_l2_in_1__A0  (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_24.mux_l2_in_2__A0  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_24.mux_l2_in_2__A1  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_24.mux_l2_in_3__A1  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_32.mux_l1_in_0__A0  (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_32.mux_l1_in_0__A1  (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_32.mux_l1_in_2__A1  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_32.mux_l1_in_3__A1  (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_4.mux_l1_in_0__A0  (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_4.mux_l1_in_0__A1  (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_4.mux_l2_in_0__A0  (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_4.mux_l2_in_5__A1  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_4.mux_l2_in_6__A0  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_4.mux_l2_in_6__A1  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_4.mux_l2_in_7__A1  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_8.mux_l1_in_0__A0  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_8.mux_l1_in_0__A1  (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_8.mux_l1_in_1__A1  (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_8.mux_l1_in_2__A0  (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_8.mux_l2_in_1__A0  (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_8.mux_l2_in_2__A0  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_8.mux_l2_in_2__A1  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_right_track_8.mux_l2_in_3__A1  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_0.mux_l1_in_2__A0  (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_0.mux_l1_in_2__A1  (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_0.mux_l1_in_3__A0  (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_0.mux_l1_in_3__A1  (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_0.mux_l1_in_4__A1  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_0.mux_l2_in_2__A0  (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_0.mux_l2_in_3__A1  (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_16.mux_l1_in_1__A0  (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_16.mux_l1_in_1__A1  (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_16.mux_l1_in_2__A0  (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_16.mux_l1_in_2__A1  (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_16.mux_l2_in_1__A0  (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_16.mux_l2_in_2__A0  (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_16.mux_l2_in_3__A1  (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_2.mux_l1_in_2__A0  (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_2.mux_l1_in_2__A1  (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_2.mux_l1_in_3__A0  (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_2.mux_l1_in_3__A1  (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_2.mux_l1_in_4__A0  (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_2.mux_l1_in_4__A1  (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_2.mux_l2_in_2__A0  (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_24.mux_l1_in_1__A0  (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_24.mux_l1_in_1__A1  (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_24.mux_l1_in_2__A0  (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_24.mux_l2_in_1__A0  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_24.mux_l2_in_2__A0  (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_24.mux_l2_in_2__A1  (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_24.mux_l2_in_3__A1  (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_32.mux_l1_in_1__A0  (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_32.mux_l1_in_2__A0  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_32.mux_l1_in_2__A1  (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_32.mux_l1_in_3__A1  (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_4.mux_l2_in_3__A0  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_4.mux_l2_in_4__A0  (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_4.mux_l2_in_4__A1  (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_4.mux_l2_in_5__A0  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_4.mux_l2_in_5__A1  (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_4.mux_l2_in_6__A0  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_4.mux_l2_in_6__A1  (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_8.mux_l1_in_1__A0  (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_8.mux_l1_in_1__A1  (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_8.mux_l1_in_2__A0  (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_8.mux_l1_in_2__A1  (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_8.mux_l2_in_1__A0  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_8.mux_l2_in_2__A1  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_top_track_8.mux_l2_in_3__A1  (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_prog_clk_2_E_FTB01_A (.DIODE(prog_clk_2_N_in));
 sky130_fd_sc_hd__diode_2 ANTENNA_prog_clk_2_N_FTB01_A (.DIODE(prog_clk_2_N_in));
 sky130_fd_sc_hd__diode_2 ANTENNA_prog_clk_2_S_FTB01_A (.DIODE(prog_clk_2_N_in));
 sky130_fd_sc_hd__diode_2 ANTENNA_prog_clk_2_W_FTB01_A (.DIODE(prog_clk_2_N_in));
 sky130_fd_sc_hd__fill_1 FILLER_0_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_142 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_172 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_160 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_172 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_171 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_183 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_143 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_127 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_142 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_149 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_7 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_99 ();
 sky130_fd_sc_hd__buf_1 Test_en_N_FTB01 (.A(net1),
    .X(net121));
 sky130_fd_sc_hd__conb_1 _028_ (.HI(_027_));
 sky130_fd_sc_hd__conb_1 _029_ (.HI(_000_));
 sky130_fd_sc_hd__conb_1 _030_ (.HI(_001_));
 sky130_fd_sc_hd__conb_1 _031_ (.HI(_002_));
 sky130_fd_sc_hd__conb_1 _032_ (.HI(_003_));
 sky130_fd_sc_hd__conb_1 _033_ (.HI(_004_));
 sky130_fd_sc_hd__conb_1 _034_ (.HI(_005_));
 sky130_fd_sc_hd__conb_1 _035_ (.HI(_006_));
 sky130_fd_sc_hd__conb_1 _036_ (.HI(_007_));
 sky130_fd_sc_hd__conb_1 _037_ (.HI(_008_));
 sky130_fd_sc_hd__conb_1 _038_ (.HI(_009_));
 sky130_fd_sc_hd__conb_1 _039_ (.HI(_010_));
 sky130_fd_sc_hd__conb_1 _040_ (.HI(_011_));
 sky130_fd_sc_hd__conb_1 _041_ (.HI(_012_));
 sky130_fd_sc_hd__conb_1 _042_ (.HI(_013_));
 sky130_fd_sc_hd__conb_1 _043_ (.HI(_014_));
 sky130_fd_sc_hd__conb_1 _044_ (.HI(_015_));
 sky130_fd_sc_hd__conb_1 _045_ (.HI(_016_));
 sky130_fd_sc_hd__conb_1 _046_ (.HI(_017_));
 sky130_fd_sc_hd__conb_1 _047_ (.HI(_018_));
 sky130_fd_sc_hd__conb_1 _048_ (.HI(_019_));
 sky130_fd_sc_hd__conb_1 _049_ (.HI(_020_));
 sky130_fd_sc_hd__conb_1 _050_ (.HI(_021_));
 sky130_fd_sc_hd__conb_1 _051_ (.HI(_022_));
 sky130_fd_sc_hd__conb_1 _052_ (.HI(_023_));
 sky130_fd_sc_hd__conb_1 _053_ (.HI(_024_));
 sky130_fd_sc_hd__conb_1 _054_ (.HI(_025_));
 sky130_fd_sc_hd__conb_1 _055_ (.HI(_026_));
 sky130_fd_sc_hd__clkbuf_1 _056_ (.A(\mux_left_track_1.out ),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 _057_ (.A(\mux_left_track_3.out ),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 _058_ (.A(\mux_left_track_5.out ),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 _059_ (.A(net43),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 _060_ (.A(\mux_left_track_9.out ),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 _061_ (.A(net45),
    .X(net138));
 sky130_fd_sc_hd__clkbuf_1 _062_ (.A(net46),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_1 _063_ (.A(net47),
    .X(net140));
 sky130_fd_sc_hd__clkbuf_1 _064_ (.A(\mux_left_track_17.out ),
    .X(net141));
 sky130_fd_sc_hd__clkbuf_1 _065_ (.A(net49),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 _066_ (.A(net50),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 _067_ (.A(net32),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_1 _068_ (.A(\mux_left_track_25.out ),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_1 _069_ (.A(net34),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 _070_ (.A(net35),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_1 _071_ (.A(net36),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_1 _072_ (.A(\mux_left_track_33.out ),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_1 _073_ (.A(net38),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_1 _074_ (.A(net39),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_1 _075_ (.A(net40),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_1 _076_ (.A(\mux_right_track_0.out ),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 _077_ (.A(\mux_right_track_2.out ),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_1 _078_ (.A(\mux_right_track_4.out ),
    .X(net155));
 sky130_fd_sc_hd__clkbuf_1 _079_ (.A(net23),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_1 _080_ (.A(\mux_right_track_8.out ),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_1 _081_ (.A(net25),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_1 _082_ (.A(net26),
    .X(net159));
 sky130_fd_sc_hd__clkbuf_1 _083_ (.A(net27),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_1 _084_ (.A(\mux_right_track_16.out ),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_1 _085_ (.A(net29),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_1 _086_ (.A(net30),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 _087_ (.A(net12),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 _088_ (.A(\mux_right_track_24.out ),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 _089_ (.A(net14),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 _090_ (.A(net15),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_1 _091_ (.A(net16),
    .X(net149));
 sky130_fd_sc_hd__clkbuf_1 _092_ (.A(\mux_right_track_32.out ),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 _093_ (.A(net18),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_1 _094_ (.A(net19),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_1 _095_ (.A(net20),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_1 _096_ (.A(\mux_bottom_track_1.out ),
    .X(net163));
 sky130_fd_sc_hd__clkbuf_1 _097_ (.A(\mux_bottom_track_3.out ),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 _098_ (.A(\mux_bottom_track_5.out ),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 _099_ (.A(net83),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 _100_ (.A(\mux_bottom_track_9.out ),
    .X(net177));
 sky130_fd_sc_hd__clkbuf_1 _101_ (.A(net85),
    .X(net178));
 sky130_fd_sc_hd__clkbuf_1 _102_ (.A(net86),
    .X(net179));
 sky130_fd_sc_hd__clkbuf_1 _103_ (.A(net87),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_1 _104_ (.A(\mux_bottom_track_17.out ),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_1 _105_ (.A(net89),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_1 _106_ (.A(net90),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_1 _107_ (.A(net72),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_1 _108_ (.A(\mux_bottom_track_25.out ),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 _109_ (.A(net74),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_1 _110_ (.A(net75),
    .X(net168));
 sky130_fd_sc_hd__clkbuf_1 _111_ (.A(net76),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_1 _112_ (.A(\mux_bottom_track_33.out ),
    .X(net170));
 sky130_fd_sc_hd__clkbuf_1 _113_ (.A(net78),
    .X(net171));
 sky130_fd_sc_hd__clkbuf_1 _114_ (.A(net79),
    .X(net172));
 sky130_fd_sc_hd__clkbuf_1 _115_ (.A(net80),
    .X(net173));
 sky130_fd_sc_hd__clkbuf_1 _116_ (.A(\mux_top_track_0.out ),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_1 _117_ (.A(\mux_top_track_2.out ),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_1 _118_ (.A(\mux_top_track_4.out ),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 _119_ (.A(net63),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 _120_ (.A(\mux_top_track_8.out ),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_1 _121_ (.A(net65),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_1 _122_ (.A(net66),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_1 _123_ (.A(net67),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_1 _124_ (.A(\mux_top_track_16.out ),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_1 _125_ (.A(net69),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_1 _126_ (.A(net70),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_1 _127_ (.A(net52),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_1 _128_ (.A(\mux_top_track_24.out ),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_1 _129_ (.A(net54),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_1 _130_ (.A(net55),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_1 _131_ (.A(net56),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_1 _132_ (.A(\mux_top_track_32.out ),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_1 _133_ (.A(net58),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_1 _134_ (.A(net59),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_1 _135_ (.A(net60),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 clk_1_E_FTB01 (.A(net91),
    .X(net203));
 sky130_fd_sc_hd__buf_1 clk_1_W_FTB01 (.A(net91),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_1 clk_2_E_FTB01 (.A(net92),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_1 clk_2_N_FTB01 (.A(net92),
    .X(net206));
 sky130_fd_sc_hd__buf_1 clk_2_S_FTB01 (.A(net92),
    .X(net207));
 sky130_fd_sc_hd__buf_1 clk_2_W_FTB01 (.A(net92),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_1 clk_3_E_FTB01 (.A(net93),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_1 clk_3_N_FTB01 (.A(net93),
    .X(net210));
 sky130_fd_sc_hd__buf_1 clk_3_S_FTB01 (.A(net93),
    .X(net211));
 sky130_fd_sc_hd__buf_1 clk_3_W_FTB01 (.A(net93),
    .X(net212));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_mem_bottom_track_1.prog_clk  (.A(\mem_bottom_track_1.prog_clk ),
    .X(\clknet_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_1_0_0_mem_bottom_track_1.prog_clk  (.A(\clknet_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_1_0_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_1_1_0_mem_bottom_track_1.prog_clk  (.A(\clknet_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_1_1_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_2_0_0_mem_bottom_track_1.prog_clk  (.A(\clknet_1_0_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_2_0_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_2_1_0_mem_bottom_track_1.prog_clk  (.A(\clknet_1_0_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_2_1_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_2_2_0_mem_bottom_track_1.prog_clk  (.A(\clknet_1_1_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_2_2_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_2_3_0_mem_bottom_track_1.prog_clk  (.A(\clknet_1_1_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_2_3_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_0_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_0_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_0_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_1_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_0_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_1_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_2_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_1_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_2_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_3_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_1_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_3_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_4_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_2_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_4_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_5_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_2_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_5_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_6_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_3_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_6_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_7_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_3_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_7_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__buf_1 input1 (.A(Test_en_S_in),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(ccff_head),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input100 (.A(left_bottom_grid_pin_40_),
    .X(net100));
 sky130_fd_sc_hd__buf_1 input101 (.A(left_bottom_grid_pin_41_),
    .X(net101));
 sky130_fd_sc_hd__buf_1 input102 (.A(prog_clk_0_N_in),
    .X(net102));
 sky130_fd_sc_hd__buf_1 input103 (.A(prog_clk_1_N_in),
    .X(net103));
 sky130_fd_sc_hd__buf_1 input104 (.A(prog_clk_3_N_in),
    .X(net104));
 sky130_fd_sc_hd__buf_1 input105 (.A(right_bottom_grid_pin_34_),
    .X(net105));
 sky130_fd_sc_hd__buf_1 input106 (.A(right_bottom_grid_pin_35_),
    .X(net106));
 sky130_fd_sc_hd__buf_1 input107 (.A(right_bottom_grid_pin_36_),
    .X(net107));
 sky130_fd_sc_hd__buf_1 input108 (.A(right_bottom_grid_pin_37_),
    .X(net108));
 sky130_fd_sc_hd__buf_1 input109 (.A(right_bottom_grid_pin_38_),
    .X(net109));
 sky130_fd_sc_hd__buf_1 input11 (.A(chanx_left_in[0]),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input110 (.A(right_bottom_grid_pin_39_),
    .X(net110));
 sky130_fd_sc_hd__buf_1 input111 (.A(right_bottom_grid_pin_40_),
    .X(net111));
 sky130_fd_sc_hd__buf_1 input112 (.A(right_bottom_grid_pin_41_),
    .X(net112));
 sky130_fd_sc_hd__buf_1 input113 (.A(top_left_grid_pin_42_),
    .X(net113));
 sky130_fd_sc_hd__buf_1 input114 (.A(top_left_grid_pin_43_),
    .X(net114));
 sky130_fd_sc_hd__buf_1 input115 (.A(top_left_grid_pin_44_),
    .X(net115));
 sky130_fd_sc_hd__buf_1 input116 (.A(top_left_grid_pin_45_),
    .X(net116));
 sky130_fd_sc_hd__buf_1 input117 (.A(top_left_grid_pin_46_),
    .X(net117));
 sky130_fd_sc_hd__buf_1 input118 (.A(top_left_grid_pin_47_),
    .X(net118));
 sky130_fd_sc_hd__buf_1 input119 (.A(top_left_grid_pin_48_),
    .X(net119));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(chanx_left_in[10]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input120 (.A(top_left_grid_pin_49_),
    .X(net120));
 sky130_fd_sc_hd__buf_1 input13 (.A(chanx_left_in[11]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(chanx_left_in[12]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 input15 (.A(chanx_left_in[13]),
    .X(net15));
 sky130_fd_sc_hd__buf_2 input16 (.A(chanx_left_in[14]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(chanx_left_in[15]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(chanx_left_in[16]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(chanx_left_in[17]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(bottom_left_grid_pin_42_),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(chanx_left_in[18]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(chanx_left_in[19]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(chanx_left_in[1]),
    .X(net22));
 sky130_fd_sc_hd__buf_2 input23 (.A(chanx_left_in[2]),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(chanx_left_in[3]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 input25 (.A(chanx_left_in[4]),
    .X(net25));
 sky130_fd_sc_hd__buf_2 input26 (.A(chanx_left_in[5]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(chanx_left_in[6]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(chanx_left_in[7]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 input29 (.A(chanx_left_in[8]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input3 (.A(bottom_left_grid_pin_43_),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input30 (.A(chanx_left_in[9]),
    .X(net30));
 sky130_fd_sc_hd__buf_1 input31 (.A(chanx_right_in[0]),
    .X(net31));
 sky130_fd_sc_hd__buf_2 input32 (.A(chanx_right_in[10]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(chanx_right_in[11]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(chanx_right_in[12]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input35 (.A(chanx_right_in[13]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(chanx_right_in[14]),
    .X(net36));
 sky130_fd_sc_hd__buf_1 input37 (.A(chanx_right_in[15]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(chanx_right_in[16]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_2 input39 (.A(chanx_right_in[17]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input4 (.A(bottom_left_grid_pin_44_),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input40 (.A(chanx_right_in[18]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(chanx_right_in[19]),
    .X(net41));
 sky130_fd_sc_hd__buf_1 input42 (.A(chanx_right_in[1]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(chanx_right_in[2]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(chanx_right_in[3]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 input45 (.A(chanx_right_in[4]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(chanx_right_in[5]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(chanx_right_in[6]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 input48 (.A(chanx_right_in[7]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(chanx_right_in[8]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input5 (.A(bottom_left_grid_pin_45_),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(chanx_right_in[9]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(chany_bottom_in[0]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(chany_bottom_in[10]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(chany_bottom_in[11]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(chany_bottom_in[12]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(chany_bottom_in[13]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 input56 (.A(chany_bottom_in[14]),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(chany_bottom_in[15]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(chany_bottom_in[16]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(chany_bottom_in[17]),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input6 (.A(bottom_left_grid_pin_46_),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(chany_bottom_in[18]),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input61 (.A(chany_bottom_in[19]),
    .X(net61));
 sky130_fd_sc_hd__buf_1 input62 (.A(chany_bottom_in[1]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_2 input63 (.A(chany_bottom_in[2]),
    .X(net63));
 sky130_fd_sc_hd__buf_1 input64 (.A(chany_bottom_in[3]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(chany_bottom_in[4]),
    .X(net65));
 sky130_fd_sc_hd__buf_2 input66 (.A(chany_bottom_in[5]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_2 input67 (.A(chany_bottom_in[6]),
    .X(net67));
 sky130_fd_sc_hd__buf_1 input68 (.A(chany_bottom_in[7]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_2 input69 (.A(chany_bottom_in[8]),
    .X(net69));
 sky130_fd_sc_hd__buf_1 input7 (.A(bottom_left_grid_pin_47_),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input70 (.A(chany_bottom_in[9]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_2 input71 (.A(chany_top_in[0]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 input72 (.A(chany_top_in[10]),
    .X(net72));
 sky130_fd_sc_hd__buf_1 input73 (.A(chany_top_in[11]),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_2 input74 (.A(chany_top_in[12]),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 input75 (.A(chany_top_in[13]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_2 input76 (.A(chany_top_in[14]),
    .X(net76));
 sky130_fd_sc_hd__buf_1 input77 (.A(chany_top_in[15]),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_2 input78 (.A(chany_top_in[16]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_2 input79 (.A(chany_top_in[17]),
    .X(net79));
 sky130_fd_sc_hd__buf_1 input8 (.A(bottom_left_grid_pin_48_),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input80 (.A(chany_top_in[18]),
    .X(net80));
 sky130_fd_sc_hd__buf_1 input81 (.A(chany_top_in[19]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_2 input82 (.A(chany_top_in[1]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_2 input83 (.A(chany_top_in[2]),
    .X(net83));
 sky130_fd_sc_hd__buf_1 input84 (.A(chany_top_in[3]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_2 input85 (.A(chany_top_in[4]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_2 input86 (.A(chany_top_in[5]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_2 input87 (.A(chany_top_in[6]),
    .X(net87));
 sky130_fd_sc_hd__buf_1 input88 (.A(chany_top_in[7]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_2 input89 (.A(chany_top_in[8]),
    .X(net89));
 sky130_fd_sc_hd__buf_1 input9 (.A(bottom_left_grid_pin_49_),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input90 (.A(chany_top_in[9]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 input91 (.A(clk_1_N_in),
    .X(net91));
 sky130_fd_sc_hd__buf_1 input92 (.A(clk_2_N_in),
    .X(net92));
 sky130_fd_sc_hd__buf_1 input93 (.A(clk_3_N_in),
    .X(net93));
 sky130_fd_sc_hd__buf_1 input94 (.A(left_bottom_grid_pin_34_),
    .X(net94));
 sky130_fd_sc_hd__buf_1 input95 (.A(left_bottom_grid_pin_35_),
    .X(net95));
 sky130_fd_sc_hd__buf_1 input96 (.A(left_bottom_grid_pin_36_),
    .X(net96));
 sky130_fd_sc_hd__buf_1 input97 (.A(left_bottom_grid_pin_37_),
    .X(net97));
 sky130_fd_sc_hd__buf_1 input98 (.A(left_bottom_grid_pin_38_),
    .X(net98));
 sky130_fd_sc_hd__buf_1 input99 (.A(left_bottom_grid_pin_39_),
    .X(net99));
 sky130_fd_sc_hd__dfxtp_2 \mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_1.ccff_head ),
    .Q(\mem_bottom_track_1.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_1.mem_out[0] ),
    .Q(\mem_bottom_track_1.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_1.mem_out[1] ),
    .Q(\mem_bottom_track_1.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_1.mem_out[2] ),
    .Q(\mem_bottom_track_1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_17.ccff_head ),
    .Q(\mem_bottom_track_17.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_17.mem_out[0] ),
    .Q(\mem_bottom_track_17.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_17.mem_out[1] ),
    .Q(\mem_bottom_track_17.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_17.mem_out[2] ),
    .Q(\mem_bottom_track_17.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_17.ccff_tail ),
    .Q(\mem_bottom_track_25.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_25.mem_out[0] ),
    .Q(\mem_bottom_track_25.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_25.mem_out[1] ),
    .Q(\mem_bottom_track_25.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_25.mem_out[2] ),
    .Q(\mem_bottom_track_25.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_2 \mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_1.ccff_tail ),
    .Q(\mem_bottom_track_3.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_3.mem_out[0] ),
    .Q(\mem_bottom_track_3.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_3.mem_out[1] ),
    .Q(\mem_bottom_track_3.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_3.mem_out[2] ),
    .Q(\mem_bottom_track_3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_25.ccff_tail ),
    .Q(\mem_bottom_track_33.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_33.mem_out[0] ),
    .Q(\mem_bottom_track_33.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_33.mem_out[1] ),
    .Q(\mem_bottom_track_33.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_3.ccff_tail ),
    .Q(\mem_bottom_track_5.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_2 \mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_5.mem_out[0] ),
    .Q(\mem_bottom_track_5.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_5.mem_out[1] ),
    .Q(\mem_bottom_track_5.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_5.mem_out[2] ),
    .Q(\mem_bottom_track_5.mem_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_5.mem_out[3] ),
    .Q(\mem_bottom_track_5.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_5.ccff_tail ),
    .Q(\mem_bottom_track_9.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_9.mem_out[0] ),
    .Q(\mem_bottom_track_9.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_9.mem_out[1] ),
    .Q(\mem_bottom_track_9.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_9.mem_out[2] ),
    .Q(\mem_bottom_track_17.ccff_head ));
 sky130_fd_sc_hd__dfxtp_2 \mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_33.ccff_tail ),
    .Q(\mem_left_track_1.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_1.mem_out[0] ),
    .Q(\mem_left_track_1.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_1.mem_out[1] ),
    .Q(\mem_left_track_1.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_1.mem_out[2] ),
    .Q(\mem_left_track_1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_17.ccff_head ),
    .Q(\mem_left_track_17.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_17.mem_out[0] ),
    .Q(\mem_left_track_17.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_17.mem_out[1] ),
    .Q(\mem_left_track_17.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_17.mem_out[2] ),
    .Q(\mem_left_track_17.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_17.ccff_tail ),
    .Q(\mem_left_track_25.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_25.mem_out[0] ),
    .Q(\mem_left_track_25.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_25.mem_out[1] ),
    .Q(\mem_left_track_25.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_25.mem_out[2] ),
    .Q(\mem_left_track_25.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_2 \mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_1.ccff_tail ),
    .Q(\mem_left_track_3.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_3.mem_out[0] ),
    .Q(\mem_left_track_3.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_3.mem_out[1] ),
    .Q(\mem_left_track_3.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_3.mem_out[2] ),
    .Q(\mem_left_track_3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_25.ccff_tail ),
    .Q(\mem_left_track_33.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_33.mem_out[0] ),
    .Q(\mem_left_track_33.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_33.mem_out[1] ),
    .Q(net122));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_3.ccff_tail ),
    .Q(\mem_left_track_5.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_2 \mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_5.mem_out[0] ),
    .Q(\mem_left_track_5.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_5.mem_out[1] ),
    .Q(\mem_left_track_5.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_5.mem_out[2] ),
    .Q(\mem_left_track_5.mem_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_5.mem_out[3] ),
    .Q(\mem_left_track_5.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_5.ccff_tail ),
    .Q(\mem_left_track_9.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_9.mem_out[0] ),
    .Q(\mem_left_track_9.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_9.mem_out[1] ),
    .Q(\mem_left_track_9.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_9.mem_out[2] ),
    .Q(\mem_left_track_17.ccff_head ));
 sky130_fd_sc_hd__dfxtp_2 \mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_0.ccff_head ),
    .Q(\mem_right_track_0.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_0.mem_out[0] ),
    .Q(\mem_right_track_0.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_0.mem_out[1] ),
    .Q(\mem_right_track_0.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_0.mem_out[2] ),
    .Q(\mem_right_track_0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_16.ccff_head ),
    .Q(\mem_right_track_16.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_16.mem_out[0] ),
    .Q(\mem_right_track_16.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_16.mem_out[1] ),
    .Q(\mem_right_track_16.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_16.mem_out[2] ),
    .Q(\mem_right_track_16.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_2 \mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_0.ccff_tail ),
    .Q(\mem_right_track_2.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_2.mem_out[0] ),
    .Q(\mem_right_track_2.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_2.mem_out[1] ),
    .Q(\mem_right_track_2.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_2.mem_out[2] ),
    .Q(\mem_right_track_2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_16.ccff_tail ),
    .Q(\mem_right_track_24.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_24.mem_out[0] ),
    .Q(\mem_right_track_24.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_24.mem_out[1] ),
    .Q(\mem_right_track_24.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_24.mem_out[2] ),
    .Q(\mem_right_track_24.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_24.ccff_tail ),
    .Q(\mem_right_track_32.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_32.mem_out[0] ),
    .Q(\mem_right_track_32.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_32.mem_out[1] ),
    .Q(\mem_bottom_track_1.ccff_head ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_2.ccff_tail ),
    .Q(\mem_right_track_4.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_2 \mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_4.mem_out[0] ),
    .Q(\mem_right_track_4.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_4.mem_out[1] ),
    .Q(\mem_right_track_4.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_4.mem_out[2] ),
    .Q(\mem_right_track_4.mem_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_4.mem_out[3] ),
    .Q(\mem_right_track_4.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_4.ccff_tail ),
    .Q(\mem_right_track_8.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_8.mem_out[0] ),
    .Q(\mem_right_track_8.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_8.mem_out[1] ),
    .Q(\mem_right_track_8.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_right_track_8.mem_out[2] ),
    .Q(\mem_right_track_16.ccff_head ));
 sky130_fd_sc_hd__dfxtp_2 \mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(net10),
    .Q(\mem_top_track_0.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_0.mem_out[0] ),
    .Q(\mem_top_track_0.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_0.mem_out[1] ),
    .Q(\mem_top_track_0.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_0.mem_out[2] ),
    .Q(\mem_top_track_0.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_16.ccff_head ),
    .Q(\mem_top_track_16.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_16.mem_out[0] ),
    .Q(\mem_top_track_16.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_16.mem_out[1] ),
    .Q(\mem_top_track_16.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_16.mem_out[2] ),
    .Q(\mem_top_track_16.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_2 \mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_0.ccff_tail ),
    .Q(\mem_top_track_2.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_2.mem_out[0] ),
    .Q(\mem_top_track_2.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_2.mem_out[1] ),
    .Q(\mem_top_track_2.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_2.mem_out[2] ),
    .Q(\mem_top_track_2.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_16.ccff_tail ),
    .Q(\mem_top_track_24.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_24.mem_out[0] ),
    .Q(\mem_top_track_24.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_24.mem_out[1] ),
    .Q(\mem_top_track_24.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_24.mem_out[2] ),
    .Q(\mem_top_track_24.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_24.ccff_tail ),
    .Q(\mem_top_track_32.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_32.mem_out[0] ),
    .Q(\mem_top_track_32.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_32.mem_out[1] ),
    .Q(\mem_right_track_0.ccff_head ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_2.ccff_tail ),
    .Q(\mem_top_track_4.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_2 \mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_4.mem_out[0] ),
    .Q(\mem_top_track_4.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_4.mem_out[1] ),
    .Q(\mem_top_track_4.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_4.mem_out[2] ),
    .Q(\mem_top_track_4.mem_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_4.mem_out[3] ),
    .Q(\mem_top_track_4.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_4.ccff_tail ),
    .Q(\mem_top_track_8.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_8.mem_out[0] ),
    .Q(\mem_top_track_8.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_8.mem_out[1] ),
    .Q(\mem_top_track_8.mem_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_top_track_8.mem_out[2] ),
    .Q(\mem_top_track_16.ccff_head ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l1_in_0_  (.A0(net74),
    .A1(net83),
    .S(\mem_bottom_track_1.mem_out[0] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l1_in_1_  (.A0(net34),
    .A1(net43),
    .S(\mem_bottom_track_1.mem_out[0] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l1_in_2_  (.A0(net2),
    .A1(net37),
    .S(\mem_bottom_track_1.mem_out[0] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l1_in_3_  (.A0(net6),
    .A1(net4),
    .S(\mem_bottom_track_1.mem_out[0] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l1_in_4_  (.A0(net22),
    .A1(net8),
    .S(\mem_bottom_track_1.mem_out[0] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l2_in_0_  (.A0(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_1.mem_out[1] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l2_in_1_  (.A0(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_bottom_track_1.mem_out[1] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l2_in_2_  (.A0(net23),
    .A1(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X ),
    .S(\mem_bottom_track_1.mem_out[1] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l2_in_3_  (.A0(_015_),
    .A1(net14),
    .S(\mem_bottom_track_1.mem_out[1] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l3_in_0_  (.A0(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_bottom_track_1.mem_out[2] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l3_in_1_  (.A0(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_bottom_track_1.mem_out[2] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_10_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l4_in_0_  (.A0(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_10_X ),
    .A1(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_9_X ),
    .S(\mem_bottom_track_1.ccff_tail ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_11_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_11_X ),
    .X(\mux_bottom_track_1.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_17.mux_l1_in_0_  (.A0(net79),
    .A1(net89),
    .S(\mem_bottom_track_17.mem_out[0] ),
    .X(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_17.mux_l1_in_1_  (.A0(net49),
    .A1(net42),
    .S(\mem_bottom_track_17.mem_out[0] ),
    .X(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_17.mux_l1_in_2_  (.A0(net3),
    .A1(net39),
    .S(\mem_bottom_track_17.mem_out[0] ),
    .X(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_17.mux_l2_in_0_  (.A0(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_17.mem_out[1] ),
    .X(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_17.mux_l2_in_1_  (.A0(net7),
    .A1(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_bottom_track_17.mem_out[1] ),
    .X(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_17.mux_l2_in_2_  (.A0(net17),
    .A1(net29),
    .S(\mem_bottom_track_17.mem_out[1] ),
    .X(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_17.mux_l2_in_3_  (.A0(_016_),
    .A1(net19),
    .S(\mem_bottom_track_17.mem_out[1] ),
    .X(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_17.mux_l3_in_0_  (.A0(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_bottom_track_17.mem_out[2] ),
    .X(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_17.mux_l3_in_1_  (.A0(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_bottom_track_17.mem_out[2] ),
    .X(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_17.mux_l4_in_0_  (.A0(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_bottom_track_17.ccff_tail ),
    .X(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_9_X ),
    .X(\mux_bottom_track_17.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_25.mux_l1_in_0_  (.A0(net80),
    .A1(net90),
    .S(\mem_bottom_track_25.mem_out[0] ),
    .X(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_25.mux_l1_in_1_  (.A0(net50),
    .A1(net31),
    .S(\mem_bottom_track_25.mem_out[0] ),
    .X(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_25.mux_l1_in_2_  (.A0(net4),
    .A1(net40),
    .S(\mem_bottom_track_25.mem_out[0] ),
    .X(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_25.mux_l2_in_0_  (.A0(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_25.mem_out[1] ),
    .X(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_25.mux_l2_in_1_  (.A0(net8),
    .A1(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_bottom_track_25.mem_out[1] ),
    .X(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_25.mux_l2_in_2_  (.A0(net20),
    .A1(net30),
    .S(\mem_bottom_track_25.mem_out[1] ),
    .X(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_25.mux_l2_in_3_  (.A0(_017_),
    .A1(net21),
    .S(\mem_bottom_track_25.mem_out[1] ),
    .X(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_25.mux_l3_in_0_  (.A0(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_bottom_track_25.mem_out[2] ),
    .X(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_25.mux_l3_in_1_  (.A0(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_bottom_track_25.mem_out[2] ),
    .X(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_25.mux_l4_in_0_  (.A0(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_bottom_track_25.ccff_tail ),
    .X(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_9_X ),
    .X(\mux_bottom_track_25.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l1_in_0_  (.A0(net75),
    .A1(net85),
    .S(\mem_bottom_track_3.mem_out[0] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l1_in_1_  (.A0(net33),
    .A1(net45),
    .S(\mem_bottom_track_3.mem_out[0] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l1_in_2_  (.A0(net3),
    .A1(net35),
    .S(\mem_bottom_track_3.mem_out[0] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l1_in_3_  (.A0(net7),
    .A1(net5),
    .S(\mem_bottom_track_3.mem_out[0] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l1_in_4_  (.A0(net24),
    .A1(net9),
    .S(\mem_bottom_track_3.mem_out[0] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l2_in_0_  (.A0(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_3.mem_out[1] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l2_in_1_  (.A0(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_bottom_track_3.mem_out[1] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l2_in_2_  (.A0(net25),
    .A1(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X ),
    .S(\mem_bottom_track_3.mem_out[1] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l2_in_3_  (.A0(_018_),
    .A1(net15),
    .S(\mem_bottom_track_3.mem_out[1] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l3_in_0_  (.A0(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_bottom_track_3.mem_out[2] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l3_in_1_  (.A0(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_bottom_track_3.mem_out[2] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_10_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l4_in_0_  (.A0(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_10_X ),
    .A1(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_9_X ),
    .S(\mem_bottom_track_3.ccff_tail ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_11_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_11_X ),
    .X(\mux_bottom_track_3.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_33.mux_l1_in_0_  (.A0(net32),
    .A1(net72),
    .S(\mem_bottom_track_33.mem_out[0] ),
    .X(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_33.mux_l1_in_1_  (.A0(net5),
    .A1(net41),
    .S(\mem_bottom_track_33.mem_out[0] ),
    .X(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_33.mux_l1_in_2_  (.A0(net11),
    .A1(net9),
    .S(\mem_bottom_track_33.mem_out[0] ),
    .X(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_33.mux_l1_in_3_  (.A0(_019_),
    .A1(net12),
    .S(\mem_bottom_track_33.mem_out[0] ),
    .X(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_33.mux_l2_in_0_  (.A0(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_33.mem_out[1] ),
    .X(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_33.mux_l2_in_1_  (.A0(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_bottom_track_33.mem_out[1] ),
    .X(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_33.mux_l3_in_0_  (.A0(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_5_X ),
    .A1(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_4_X ),
    .S(\mem_bottom_track_33.ccff_tail ),
    .X(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_33.sky130_fd_sc_hd__mux2_1_6_X ),
    .X(\mux_bottom_track_33.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l1_in_0_  (.A0(net76),
    .A1(net86),
    .S(\mem_bottom_track_5.mem_out[0] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l2_in_0_  (.A0(net46),
    .A1(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_5.mem_out[1] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l2_in_1_  (.A0(net36),
    .A1(net48),
    .S(\mem_bottom_track_5.mem_out[1] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l2_in_2_  (.A0(net3),
    .A1(net2),
    .S(\mem_bottom_track_5.mem_out[1] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l2_in_3_  (.A0(net5),
    .A1(net4),
    .S(\mem_bottom_track_5.mem_out[1] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l2_in_4_  (.A0(net7),
    .A1(net6),
    .S(\mem_bottom_track_5.mem_out[1] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l2_in_5_  (.A0(net9),
    .A1(net8),
    .S(\mem_bottom_track_5.mem_out[1] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l2_in_6_  (.A0(net28),
    .A1(net26),
    .S(\mem_bottom_track_5.mem_out[1] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l2_in_7_  (.A0(_020_),
    .A1(net16),
    .S(\mem_bottom_track_5.mem_out[1] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l3_in_0_  (.A0(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X ),
    .A1(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X ),
    .S(\mem_bottom_track_5.mem_out[2] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l3_in_1_  (.A0(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_bottom_track_5.mem_out[2] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_10_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l3_in_2_  (.A0(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_bottom_track_5.mem_out[2] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_11_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l3_in_3_  (.A0(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_bottom_track_5.mem_out[2] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_12_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l4_in_0_  (.A0(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_10_X ),
    .A1(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_9_X ),
    .S(\mem_bottom_track_5.mem_out[3] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_13_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l4_in_1_  (.A0(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_12_X ),
    .A1(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_11_X ),
    .S(\mem_bottom_track_5.mem_out[3] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_14_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l5_in_0_  (.A0(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_14_X ),
    .A1(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_13_X ),
    .S(\mem_bottom_track_5.ccff_tail ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_15_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_15_X ),
    .X(\mux_bottom_track_5.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_9.mux_l1_in_0_  (.A0(net78),
    .A1(net87),
    .S(\mem_bottom_track_9.mem_out[0] ),
    .X(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_9.mux_l1_in_1_  (.A0(net47),
    .A1(net44),
    .S(\mem_bottom_track_9.mem_out[0] ),
    .X(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_9.mux_l1_in_2_  (.A0(net2),
    .A1(net38),
    .S(\mem_bottom_track_9.mem_out[0] ),
    .X(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_9.mux_l2_in_0_  (.A0(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_9.mem_out[1] ),
    .X(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_9.mux_l2_in_1_  (.A0(net6),
    .A1(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_bottom_track_9.mem_out[1] ),
    .X(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_9.mux_l2_in_2_  (.A0(net13),
    .A1(net27),
    .S(\mem_bottom_track_9.mem_out[1] ),
    .X(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_9.mux_l2_in_3_  (.A0(_021_),
    .A1(net18),
    .S(\mem_bottom_track_9.mem_out[1] ),
    .X(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_9.mux_l3_in_0_  (.A0(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_bottom_track_9.mem_out[2] ),
    .X(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_9.mux_l3_in_1_  (.A0(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_bottom_track_9.mem_out[2] ),
    .X(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_9.mux_l4_in_0_  (.A0(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_bottom_track_17.ccff_head ),
    .X(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_9_X ),
    .X(\mux_bottom_track_9.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l1_in_0_  (.A0(net83),
    .A1(net71),
    .S(\mem_left_track_1.mem_out[0] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l1_in_1_  (.A0(net43),
    .A1(net74),
    .S(\mem_left_track_1.mem_out[0] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l1_in_2_  (.A0(net63),
    .A1(net34),
    .S(\mem_left_track_1.mem_out[0] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l1_in_3_  (.A0(net61),
    .A1(net54),
    .S(\mem_left_track_1.mem_out[0] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l1_in_4_  (.A0(net96),
    .A1(net94),
    .S(\mem_left_track_1.mem_out[0] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l2_in_0_  (.A0(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_1.mem_out[1] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l2_in_1_  (.A0(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_left_track_1.mem_out[1] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l2_in_2_  (.A0(net98),
    .A1(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X ),
    .S(\mem_left_track_1.mem_out[1] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l2_in_3_  (.A0(_022_),
    .A1(net100),
    .S(\mem_left_track_1.mem_out[1] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l3_in_0_  (.A0(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_left_track_1.mem_out[2] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l3_in_1_  (.A0(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_left_track_1.mem_out[2] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_10_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l4_in_0_  (.A0(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_10_X ),
    .A1(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_9_X ),
    .S(\mem_left_track_1.ccff_tail ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_11_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_1.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_11_X ),
    .X(\mux_left_track_1.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_17.mux_l1_in_0_  (.A0(net89),
    .A1(net88),
    .S(\mem_left_track_17.mem_out[0] ),
    .X(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_17.mux_l1_in_1_  (.A0(net49),
    .A1(net79),
    .S(\mem_left_track_17.mem_out[0] ),
    .X(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_17.mux_l1_in_2_  (.A0(net68),
    .A1(net39),
    .S(\mem_left_track_17.mem_out[0] ),
    .X(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_17.mux_l2_in_0_  (.A0(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_17.mem_out[1] ),
    .X(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_17.mux_l2_in_1_  (.A0(net69),
    .A1(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_left_track_17.mem_out[1] ),
    .X(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_17.mux_l2_in_2_  (.A0(net95),
    .A1(net59),
    .S(\mem_left_track_17.mem_out[1] ),
    .X(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_17.mux_l2_in_3_  (.A0(_023_),
    .A1(net99),
    .S(\mem_left_track_17.mem_out[1] ),
    .X(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_17.mux_l3_in_0_  (.A0(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_left_track_17.mem_out[2] ),
    .X(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_17.mux_l3_in_1_  (.A0(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_left_track_17.mem_out[2] ),
    .X(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_17.mux_l4_in_0_  (.A0(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_left_track_17.ccff_tail ),
    .X(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_17.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_9_X ),
    .X(\mux_left_track_17.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_25.mux_l1_in_0_  (.A0(net90),
    .A1(net84),
    .S(\mem_left_track_25.mem_out[0] ),
    .X(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_25.mux_l1_in_1_  (.A0(net50),
    .A1(net80),
    .S(\mem_left_track_25.mem_out[0] ),
    .X(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_25.mux_l1_in_2_  (.A0(net70),
    .A1(net40),
    .S(\mem_left_track_25.mem_out[0] ),
    .X(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_25.mux_l2_in_0_  (.A0(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_25.mem_out[1] ),
    .X(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_25.mux_l2_in_1_  (.A0(net53),
    .A1(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_left_track_25.mem_out[1] ),
    .X(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_25.mux_l2_in_2_  (.A0(net96),
    .A1(net60),
    .S(\mem_left_track_25.mem_out[1] ),
    .X(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_25.mux_l2_in_3_  (.A0(_024_),
    .A1(net100),
    .S(\mem_left_track_25.mem_out[1] ),
    .X(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_25.mux_l3_in_0_  (.A0(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_left_track_25.mem_out[2] ),
    .X(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_25.mux_l3_in_1_  (.A0(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_left_track_25.mem_out[2] ),
    .X(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_25.mux_l4_in_0_  (.A0(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_left_track_25.ccff_tail ),
    .X(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_25.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_9_X ),
    .X(\mux_left_track_25.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l1_in_0_  (.A0(net75),
    .A1(net85),
    .S(\mem_left_track_3.mem_out[0] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l1_in_1_  (.A0(net45),
    .A1(net81),
    .S(\mem_left_track_3.mem_out[0] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l1_in_2_  (.A0(net51),
    .A1(net35),
    .S(\mem_left_track_3.mem_out[0] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l1_in_3_  (.A0(net55),
    .A1(net65),
    .S(\mem_left_track_3.mem_out[0] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l1_in_4_  (.A0(net97),
    .A1(net95),
    .S(\mem_left_track_3.mem_out[0] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l2_in_0_  (.A0(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_3.mem_out[1] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l2_in_1_  (.A0(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_left_track_3.mem_out[1] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l2_in_2_  (.A0(net99),
    .A1(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X ),
    .S(\mem_left_track_3.mem_out[1] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l2_in_3_  (.A0(_025_),
    .A1(net101),
    .S(\mem_left_track_3.mem_out[1] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l3_in_0_  (.A0(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_left_track_3.mem_out[2] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l3_in_1_  (.A0(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_left_track_3.mem_out[2] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_10_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l4_in_0_  (.A0(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_10_X ),
    .A1(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_9_X ),
    .S(\mem_left_track_3.ccff_tail ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_11_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_3.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_11_X ),
    .X(\mux_left_track_3.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_33.mux_l1_in_0_  (.A0(net72),
    .A1(net82),
    .S(\mem_left_track_33.mem_out[0] ),
    .X(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_33.mux_l1_in_1_  (.A0(net52),
    .A1(net32),
    .S(\mem_left_track_33.mem_out[0] ),
    .X(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_33.mux_l1_in_2_  (.A0(net97),
    .A1(net57),
    .S(\mem_left_track_33.mem_out[0] ),
    .X(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_33.mux_l1_in_3_  (.A0(_026_),
    .A1(net101),
    .S(\mem_left_track_33.mem_out[0] ),
    .X(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_33.mux_l2_in_0_  (.A0(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_33.mem_out[1] ),
    .X(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_33.mux_l2_in_1_  (.A0(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_left_track_33.mem_out[1] ),
    .X(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_33.mux_l3_in_0_  (.A0(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_5_X ),
    .A1(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_4_X ),
    .S(net122),
    .X(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_33.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_6_X ),
    .X(\mux_left_track_33.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l1_in_0_  (.A0(net76),
    .A1(net86),
    .S(\mem_left_track_5.mem_out[0] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l2_in_0_  (.A0(net77),
    .A1(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_5.mem_out[1] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l2_in_1_  (.A0(net36),
    .A1(net46),
    .S(\mem_left_track_5.mem_out[1] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l2_in_2_  (.A0(net66),
    .A1(net62),
    .S(\mem_left_track_5.mem_out[1] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l2_in_3_  (.A0(net94),
    .A1(net56),
    .S(\mem_left_track_5.mem_out[1] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l2_in_4_  (.A0(net96),
    .A1(net95),
    .S(\mem_left_track_5.mem_out[1] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l2_in_5_  (.A0(net98),
    .A1(net97),
    .S(\mem_left_track_5.mem_out[1] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l2_in_6_  (.A0(net100),
    .A1(net99),
    .S(\mem_left_track_5.mem_out[1] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l2_in_7_  (.A0(_027_),
    .A1(net101),
    .S(\mem_left_track_5.mem_out[1] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l3_in_0_  (.A0(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X ),
    .A1(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X ),
    .S(\mem_left_track_5.mem_out[2] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l3_in_1_  (.A0(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_left_track_5.mem_out[2] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_10_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l3_in_2_  (.A0(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_left_track_5.mem_out[2] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_11_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l3_in_3_  (.A0(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_left_track_5.mem_out[2] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_12_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l4_in_0_  (.A0(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_10_X ),
    .A1(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_9_X ),
    .S(\mem_left_track_5.mem_out[3] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_13_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l4_in_1_  (.A0(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_12_X ),
    .A1(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_11_X ),
    .S(\mem_left_track_5.mem_out[3] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_14_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l5_in_0_  (.A0(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_14_X ),
    .A1(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_13_X ),
    .S(\mem_left_track_5.ccff_tail ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_15_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_5.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_15_X ),
    .X(\mux_left_track_5.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_9.mux_l1_in_0_  (.A0(net73),
    .A1(net87),
    .S(\mem_left_track_9.mem_out[0] ),
    .X(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_9.mux_l1_in_1_  (.A0(net47),
    .A1(net78),
    .S(\mem_left_track_9.mem_out[0] ),
    .X(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_9.mux_l1_in_2_  (.A0(net64),
    .A1(net38),
    .S(\mem_left_track_9.mem_out[0] ),
    .X(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_9.mux_l2_in_0_  (.A0(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_9.mem_out[1] ),
    .X(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_9.mux_l2_in_1_  (.A0(net67),
    .A1(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_left_track_9.mem_out[1] ),
    .X(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_9.mux_l2_in_2_  (.A0(net94),
    .A1(net58),
    .S(\mem_left_track_9.mem_out[1] ),
    .X(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_9.mux_l2_in_3_  (.A0(_000_),
    .A1(net98),
    .S(\mem_left_track_9.mem_out[1] ),
    .X(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_9.mux_l3_in_0_  (.A0(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_left_track_9.mem_out[2] ),
    .X(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_9.mux_l3_in_1_  (.A0(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_left_track_9.mem_out[2] ),
    .X(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_9.mux_l4_in_0_  (.A0(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_left_track_17.ccff_head ),
    .X(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_9.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_9_X ),
    .X(\mux_left_track_9.out ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_0.mux_l1_in_0_  (.A0(net74),
    .A1(net83),
    .S(\mem_right_track_0.mem_out[0] ),
    .X(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_0.mux_l1_in_1_  (.A0(net105),
    .A1(net81),
    .S(\mem_right_track_0.mem_out[0] ),
    .X(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_0.mux_l1_in_2_  (.A0(net109),
    .A1(net107),
    .S(\mem_right_track_0.mem_out[0] ),
    .X(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_0.mux_l1_in_3_  (.A0(net63),
    .A1(net111),
    .S(\mem_right_track_0.mem_out[0] ),
    .X(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_0.mux_l1_in_4_  (.A0(net57),
    .A1(net54),
    .S(\mem_right_track_0.mem_out[0] ),
    .X(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_0.mux_l2_in_0_  (.A0(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_right_track_0.mem_out[1] ),
    .X(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_0.mux_l2_in_1_  (.A0(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_right_track_0.mem_out[1] ),
    .X(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_0.mux_l2_in_2_  (.A0(net23),
    .A1(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_4_X ),
    .S(\mem_right_track_0.mem_out[1] ),
    .X(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_0.mux_l2_in_3_  (.A0(_001_),
    .A1(net14),
    .S(\mem_right_track_0.mem_out[1] ),
    .X(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_0.mux_l3_in_0_  (.A0(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_right_track_0.mem_out[2] ),
    .X(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_0.mux_l3_in_1_  (.A0(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_right_track_0.mem_out[2] ),
    .X(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_10_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_0.mux_l4_in_0_  (.A0(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_10_X ),
    .A1(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_9_X ),
    .S(\mem_right_track_0.ccff_tail ),
    .X(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_11_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_right_track_0.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_right_track_0.sky130_fd_sc_hd__mux2_1_11_X ),
    .X(\mux_right_track_0.out ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_16.mux_l1_in_0_  (.A0(net89),
    .A1(net88),
    .S(\mem_right_track_16.mem_out[0] ),
    .X(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_16.mux_l1_in_1_  (.A0(net106),
    .A1(net79),
    .S(\mem_right_track_16.mem_out[0] ),
    .X(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_16.mux_l1_in_2_  (.A0(net62),
    .A1(net110),
    .S(\mem_right_track_16.mem_out[0] ),
    .X(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_16.mux_l2_in_0_  (.A0(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_right_track_16.mem_out[1] ),
    .X(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_16.mux_l2_in_1_  (.A0(net69),
    .A1(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_right_track_16.mem_out[1] ),
    .X(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_16.mux_l2_in_2_  (.A0(net29),
    .A1(net59),
    .S(\mem_right_track_16.mem_out[1] ),
    .X(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_16.mux_l2_in_3_  (.A0(_002_),
    .A1(net19),
    .S(\mem_right_track_16.mem_out[1] ),
    .X(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_16.mux_l3_in_0_  (.A0(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_right_track_16.mem_out[2] ),
    .X(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_16.mux_l3_in_1_  (.A0(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_right_track_16.mem_out[2] ),
    .X(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_16.mux_l4_in_0_  (.A0(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_right_track_16.ccff_tail ),
    .X(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_right_track_16.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_right_track_16.sky130_fd_sc_hd__mux2_1_9_X ),
    .X(\mux_right_track_16.out ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_2.mux_l1_in_0_  (.A0(net85),
    .A1(net71),
    .S(\mem_right_track_2.mem_out[0] ),
    .X(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_2.mux_l1_in_1_  (.A0(net106),
    .A1(net75),
    .S(\mem_right_track_2.mem_out[0] ),
    .X(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_2.mux_l1_in_2_  (.A0(net110),
    .A1(net108),
    .S(\mem_right_track_2.mem_out[0] ),
    .X(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_2.mux_l1_in_3_  (.A0(net65),
    .A1(net112),
    .S(\mem_right_track_2.mem_out[0] ),
    .X(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_2.mux_l1_in_4_  (.A0(net55),
    .A1(net53),
    .S(\mem_right_track_2.mem_out[0] ),
    .X(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_2.mux_l2_in_0_  (.A0(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_right_track_2.mem_out[1] ),
    .X(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_2.mux_l2_in_1_  (.A0(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_right_track_2.mem_out[1] ),
    .X(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_2.mux_l2_in_2_  (.A0(net25),
    .A1(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_4_X ),
    .S(\mem_right_track_2.mem_out[1] ),
    .X(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_2.mux_l2_in_3_  (.A0(_003_),
    .A1(net15),
    .S(\mem_right_track_2.mem_out[1] ),
    .X(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_2.mux_l3_in_0_  (.A0(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_right_track_2.mem_out[2] ),
    .X(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_2.mux_l3_in_1_  (.A0(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_right_track_2.mem_out[2] ),
    .X(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_10_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_2.mux_l4_in_0_  (.A0(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_10_X ),
    .A1(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_9_X ),
    .S(\mem_right_track_2.ccff_tail ),
    .X(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_11_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_right_track_2.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_right_track_2.sky130_fd_sc_hd__mux2_1_11_X ),
    .X(\mux_right_track_2.out ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_24.mux_l1_in_0_  (.A0(net73),
    .A1(net90),
    .S(\mem_right_track_24.mem_out[0] ),
    .X(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_24.mux_l1_in_1_  (.A0(net107),
    .A1(net80),
    .S(\mem_right_track_24.mem_out[0] ),
    .X(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_24.mux_l1_in_2_  (.A0(net51),
    .A1(net111),
    .S(\mem_right_track_24.mem_out[0] ),
    .X(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_24.mux_l2_in_0_  (.A0(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_right_track_24.mem_out[1] ),
    .X(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_24.mux_l2_in_1_  (.A0(net70),
    .A1(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_right_track_24.mem_out[1] ),
    .X(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_24.mux_l2_in_2_  (.A0(net30),
    .A1(net60),
    .S(\mem_right_track_24.mem_out[1] ),
    .X(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_24.mux_l2_in_3_  (.A0(_004_),
    .A1(net20),
    .S(\mem_right_track_24.mem_out[1] ),
    .X(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_24.mux_l3_in_0_  (.A0(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_right_track_24.mem_out[2] ),
    .X(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_24.mux_l3_in_1_  (.A0(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_right_track_24.mem_out[2] ),
    .X(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_24.mux_l4_in_0_  (.A0(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_right_track_24.ccff_tail ),
    .X(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_right_track_24.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_right_track_24.sky130_fd_sc_hd__mux2_1_9_X ),
    .X(\mux_right_track_24.out ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_32.mux_l1_in_0_  (.A0(net77),
    .A1(net72),
    .S(\mem_right_track_32.mem_out[0] ),
    .X(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_32.mux_l1_in_1_  (.A0(net112),
    .A1(net108),
    .S(\mem_right_track_32.mem_out[0] ),
    .X(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_32.mux_l1_in_2_  (.A0(net61),
    .A1(net52),
    .S(\mem_right_track_32.mem_out[0] ),
    .X(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_32.mux_l1_in_3_  (.A0(_005_),
    .A1(net12),
    .S(\mem_right_track_32.mem_out[0] ),
    .X(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_32.mux_l2_in_0_  (.A0(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_right_track_32.mem_out[1] ),
    .X(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_32.mux_l2_in_1_  (.A0(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_right_track_32.mem_out[1] ),
    .X(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_32.mux_l3_in_0_  (.A0(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_5_X ),
    .A1(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_4_X ),
    .S(\mem_bottom_track_1.ccff_head ),
    .X(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_right_track_32.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_right_track_32.sky130_fd_sc_hd__mux2_1_6_X ),
    .X(\mux_right_track_32.out ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l1_in_0_  (.A0(net86),
    .A1(net82),
    .S(\mem_right_track_4.mem_out[0] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l2_in_0_  (.A0(net76),
    .A1(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_right_track_4.mem_out[1] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l2_in_1_  (.A0(net106),
    .A1(net105),
    .S(\mem_right_track_4.mem_out[1] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l2_in_2_  (.A0(net108),
    .A1(net107),
    .S(\mem_right_track_4.mem_out[1] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l2_in_3_  (.A0(net110),
    .A1(net109),
    .S(\mem_right_track_4.mem_out[1] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l2_in_4_  (.A0(net112),
    .A1(net111),
    .S(\mem_right_track_4.mem_out[1] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l2_in_5_  (.A0(net68),
    .A1(net66),
    .S(\mem_right_track_4.mem_out[1] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l2_in_6_  (.A0(net26),
    .A1(net56),
    .S(\mem_right_track_4.mem_out[1] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l2_in_7_  (.A0(_006_),
    .A1(net16),
    .S(\mem_right_track_4.mem_out[1] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l3_in_0_  (.A0(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_2_X ),
    .A1(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_1_X ),
    .S(\mem_right_track_4.mem_out[2] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l3_in_1_  (.A0(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_right_track_4.mem_out[2] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_10_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l3_in_2_  (.A0(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_right_track_4.mem_out[2] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_11_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l3_in_3_  (.A0(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_right_track_4.mem_out[2] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_12_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l4_in_0_  (.A0(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_10_X ),
    .A1(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_9_X ),
    .S(\mem_right_track_4.mem_out[3] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_13_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l4_in_1_  (.A0(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_12_X ),
    .A1(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_11_X ),
    .S(\mem_right_track_4.mem_out[3] ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_14_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_4.mux_l5_in_0_  (.A0(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_14_X ),
    .A1(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_13_X ),
    .S(\mem_right_track_4.ccff_tail ),
    .X(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_15_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_right_track_4.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_right_track_4.sky130_fd_sc_hd__mux2_1_15_X ),
    .X(\mux_right_track_4.out ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_8.mux_l1_in_0_  (.A0(net87),
    .A1(net84),
    .S(\mem_right_track_8.mem_out[0] ),
    .X(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_8.mux_l1_in_1_  (.A0(net105),
    .A1(net78),
    .S(\mem_right_track_8.mem_out[0] ),
    .X(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_8.mux_l1_in_2_  (.A0(net64),
    .A1(net109),
    .S(\mem_right_track_8.mem_out[0] ),
    .X(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_8.mux_l2_in_0_  (.A0(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_right_track_8.mem_out[1] ),
    .X(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_8.mux_l2_in_1_  (.A0(net67),
    .A1(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_right_track_8.mem_out[1] ),
    .X(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_8.mux_l2_in_2_  (.A0(net27),
    .A1(net58),
    .S(\mem_right_track_8.mem_out[1] ),
    .X(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_8.mux_l2_in_3_  (.A0(_007_),
    .A1(net18),
    .S(\mem_right_track_8.mem_out[1] ),
    .X(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_8.mux_l3_in_0_  (.A0(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_right_track_8.mem_out[2] ),
    .X(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_8.mux_l3_in_1_  (.A0(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_right_track_8.mem_out[2] ),
    .X(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_right_track_8.mux_l4_in_0_  (.A0(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_right_track_16.ccff_head ),
    .X(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_right_track_8.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_right_track_8.sky130_fd_sc_hd__mux2_1_9_X ),
    .X(\mux_right_track_8.out ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_0.mux_l1_in_0_  (.A0(net115),
    .A1(net113),
    .S(\mem_top_track_0.mem_out[0] ),
    .X(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_0.mux_l1_in_1_  (.A0(net119),
    .A1(net117),
    .S(\mem_top_track_0.mem_out[0] ),
    .X(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_0.mux_l1_in_2_  (.A0(net43),
    .A1(net42),
    .S(\mem_top_track_0.mem_out[0] ),
    .X(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_0.mux_l1_in_3_  (.A0(net63),
    .A1(net34),
    .S(\mem_top_track_0.mem_out[0] ),
    .X(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_0.mux_l1_in_4_  (.A0(net11),
    .A1(net54),
    .S(\mem_top_track_0.mem_out[0] ),
    .X(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_0.mux_l2_in_0_  (.A0(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_top_track_0.mem_out[1] ),
    .X(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_0.mux_l2_in_1_  (.A0(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_top_track_0.mem_out[1] ),
    .X(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_0.mux_l2_in_2_  (.A0(net23),
    .A1(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_4_X ),
    .S(\mem_top_track_0.mem_out[1] ),
    .X(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_0.mux_l2_in_3_  (.A0(_008_),
    .A1(net14),
    .S(\mem_top_track_0.mem_out[1] ),
    .X(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_0.mux_l3_in_0_  (.A0(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_top_track_0.mem_out[2] ),
    .X(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_0.mux_l3_in_1_  (.A0(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_top_track_0.mem_out[2] ),
    .X(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_10_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_0.mux_l4_in_0_  (.A0(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_10_X ),
    .A1(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_9_X ),
    .S(\mem_top_track_0.ccff_tail ),
    .X(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_11_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_top_track_0.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_top_track_0.sky130_fd_sc_hd__mux2_1_11_X ),
    .X(\mux_top_track_0.out ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_16.mux_l1_in_0_  (.A0(net118),
    .A1(net114),
    .S(\mem_top_track_16.mem_out[0] ),
    .X(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_16.mux_l1_in_1_  (.A0(net37),
    .A1(net49),
    .S(\mem_top_track_16.mem_out[0] ),
    .X(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_16.mux_l1_in_2_  (.A0(net69),
    .A1(net39),
    .S(\mem_top_track_16.mem_out[0] ),
    .X(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_16.mux_l2_in_0_  (.A0(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_top_track_16.mem_out[1] ),
    .X(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_16.mux_l2_in_1_  (.A0(net59),
    .A1(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_top_track_16.mem_out[1] ),
    .X(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_16.mux_l2_in_2_  (.A0(net29),
    .A1(net28),
    .S(\mem_top_track_16.mem_out[1] ),
    .X(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_16.mux_l2_in_3_  (.A0(_009_),
    .A1(net19),
    .S(\mem_top_track_16.mem_out[1] ),
    .X(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_16.mux_l3_in_0_  (.A0(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_top_track_16.mem_out[2] ),
    .X(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_16.mux_l3_in_1_  (.A0(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_top_track_16.mem_out[2] ),
    .X(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_16.mux_l4_in_0_  (.A0(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_top_track_16.ccff_tail ),
    .X(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_top_track_16.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_top_track_16.sky130_fd_sc_hd__mux2_1_9_X ),
    .X(\mux_top_track_16.out ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_2.mux_l1_in_0_  (.A0(net116),
    .A1(net114),
    .S(\mem_top_track_2.mem_out[0] ),
    .X(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_2.mux_l1_in_1_  (.A0(net120),
    .A1(net118),
    .S(\mem_top_track_2.mem_out[0] ),
    .X(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_2.mux_l1_in_2_  (.A0(net45),
    .A1(net44),
    .S(\mem_top_track_2.mem_out[0] ),
    .X(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_2.mux_l1_in_3_  (.A0(net65),
    .A1(net35),
    .S(\mem_top_track_2.mem_out[0] ),
    .X(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_2.mux_l1_in_4_  (.A0(net25),
    .A1(net55),
    .S(\mem_top_track_2.mem_out[0] ),
    .X(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_2.mux_l2_in_0_  (.A0(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_top_track_2.mem_out[1] ),
    .X(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_2.mux_l2_in_1_  (.A0(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_top_track_2.mem_out[1] ),
    .X(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_2.mux_l2_in_2_  (.A0(net15),
    .A1(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_4_X ),
    .S(\mem_top_track_2.mem_out[1] ),
    .X(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_2.mux_l2_in_3_  (.A0(_010_),
    .A1(net21),
    .S(\mem_top_track_2.mem_out[1] ),
    .X(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_2.mux_l3_in_0_  (.A0(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_top_track_2.mem_out[2] ),
    .X(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_2.mux_l3_in_1_  (.A0(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_top_track_2.mem_out[2] ),
    .X(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_10_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_2.mux_l4_in_0_  (.A0(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_10_X ),
    .A1(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_9_X ),
    .S(\mem_top_track_2.ccff_tail ),
    .X(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_11_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_top_track_2.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_top_track_2.sky130_fd_sc_hd__mux2_1_11_X ),
    .X(\mux_top_track_2.out ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_24.mux_l1_in_0_  (.A0(net119),
    .A1(net115),
    .S(\mem_top_track_24.mem_out[0] ),
    .X(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_24.mux_l1_in_1_  (.A0(net40),
    .A1(net50),
    .S(\mem_top_track_24.mem_out[0] ),
    .X(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_24.mux_l1_in_2_  (.A0(net70),
    .A1(net41),
    .S(\mem_top_track_24.mem_out[0] ),
    .X(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_24.mux_l2_in_0_  (.A0(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_top_track_24.mem_out[1] ),
    .X(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_24.mux_l2_in_1_  (.A0(net60),
    .A1(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_top_track_24.mem_out[1] ),
    .X(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_24.mux_l2_in_2_  (.A0(net30),
    .A1(net24),
    .S(\mem_top_track_24.mem_out[1] ),
    .X(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_24.mux_l2_in_3_  (.A0(_011_),
    .A1(net20),
    .S(\mem_top_track_24.mem_out[1] ),
    .X(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_24.mux_l3_in_0_  (.A0(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_top_track_24.mem_out[2] ),
    .X(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_24.mux_l3_in_1_  (.A0(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_top_track_24.mem_out[2] ),
    .X(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_24.mux_l4_in_0_  (.A0(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_top_track_24.ccff_tail ),
    .X(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_top_track_24.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_top_track_24.sky130_fd_sc_hd__mux2_1_9_X ),
    .X(\mux_top_track_24.out ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_32.mux_l1_in_0_  (.A0(net120),
    .A1(net116),
    .S(\mem_top_track_32.mem_out[0] ),
    .X(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_32.mux_l1_in_1_  (.A0(net32),
    .A1(net31),
    .S(\mem_top_track_32.mem_out[0] ),
    .X(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_32.mux_l1_in_2_  (.A0(net22),
    .A1(net52),
    .S(\mem_top_track_32.mem_out[0] ),
    .X(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_32.mux_l1_in_3_  (.A0(_012_),
    .A1(net12),
    .S(\mem_top_track_32.mem_out[0] ),
    .X(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_32.mux_l2_in_0_  (.A0(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_top_track_32.mem_out[1] ),
    .X(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_32.mux_l2_in_1_  (.A0(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_top_track_32.mem_out[1] ),
    .X(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_32.mux_l3_in_0_  (.A0(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_5_X ),
    .A1(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_4_X ),
    .S(\mem_right_track_0.ccff_head ),
    .X(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_top_track_32.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_top_track_32.sky130_fd_sc_hd__mux2_1_6_X ),
    .X(\mux_top_track_32.out ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l1_in_0_  (.A0(net114),
    .A1(net113),
    .S(\mem_top_track_4.mem_out[0] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l2_in_0_  (.A0(net115),
    .A1(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_top_track_4.mem_out[1] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l2_in_1_  (.A0(net117),
    .A1(net116),
    .S(\mem_top_track_4.mem_out[1] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l2_in_2_  (.A0(net119),
    .A1(net118),
    .S(\mem_top_track_4.mem_out[1] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l2_in_3_  (.A0(net46),
    .A1(net120),
    .S(\mem_top_track_4.mem_out[1] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l2_in_4_  (.A0(net36),
    .A1(net48),
    .S(\mem_top_track_4.mem_out[1] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l2_in_5_  (.A0(net56),
    .A1(net66),
    .S(\mem_top_track_4.mem_out[1] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l2_in_6_  (.A0(net16),
    .A1(net26),
    .S(\mem_top_track_4.mem_out[1] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l2_in_7_  (.A0(_013_),
    .A1(net17),
    .S(\mem_top_track_4.mem_out[1] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l3_in_0_  (.A0(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_2_X ),
    .A1(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_1_X ),
    .S(\mem_top_track_4.mem_out[2] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l3_in_1_  (.A0(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_top_track_4.mem_out[2] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_10_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l3_in_2_  (.A0(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_top_track_4.mem_out[2] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_11_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l3_in_3_  (.A0(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_top_track_4.mem_out[2] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_12_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l4_in_0_  (.A0(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_10_X ),
    .A1(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_9_X ),
    .S(\mem_top_track_4.mem_out[3] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_13_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l4_in_1_  (.A0(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_12_X ),
    .A1(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_11_X ),
    .S(\mem_top_track_4.mem_out[3] ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_14_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_4.mux_l5_in_0_  (.A0(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_14_X ),
    .A1(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_13_X ),
    .S(\mem_top_track_4.ccff_tail ),
    .X(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_15_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_top_track_4.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_top_track_4.sky130_fd_sc_hd__mux2_1_15_X ),
    .X(\mux_top_track_4.out ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_8.mux_l1_in_0_  (.A0(net117),
    .A1(net113),
    .S(\mem_top_track_8.mem_out[0] ),
    .X(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_8.mux_l1_in_1_  (.A0(net33),
    .A1(net47),
    .S(\mem_top_track_8.mem_out[0] ),
    .X(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_8.mux_l1_in_2_  (.A0(net67),
    .A1(net38),
    .S(\mem_top_track_8.mem_out[0] ),
    .X(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_8.mux_l2_in_0_  (.A0(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_top_track_8.mem_out[1] ),
    .X(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_8.mux_l2_in_1_  (.A0(net58),
    .A1(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_top_track_8.mem_out[1] ),
    .X(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_8.mux_l2_in_2_  (.A0(net13),
    .A1(net27),
    .S(\mem_top_track_8.mem_out[1] ),
    .X(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_8.mux_l2_in_3_  (.A0(_014_),
    .A1(net18),
    .S(\mem_top_track_8.mem_out[1] ),
    .X(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_6_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_8.mux_l3_in_0_  (.A0(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_top_track_8.mem_out[2] ),
    .X(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_7_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_8.mux_l3_in_1_  (.A0(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_6_X ),
    .A1(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_5_X ),
    .S(\mem_top_track_8.mem_out[2] ),
    .X(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_8_X ));
 sky130_fd_sc_hd__mux2_1 \mux_top_track_8.mux_l4_in_0_  (.A0(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_8_X ),
    .A1(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_7_X ),
    .S(\mem_top_track_16.ccff_head ),
    .X(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_9_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_top_track_8.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_top_track_8.sky130_fd_sc_hd__mux2_1_9_X ),
    .X(\mux_top_track_8.out ));
 sky130_fd_sc_hd__clkbuf_2 output121 (.A(net121),
    .X(Test_en_N_out));
 sky130_fd_sc_hd__clkbuf_2 output122 (.A(net122),
    .X(ccff_tail));
 sky130_fd_sc_hd__clkbuf_2 output123 (.A(net123),
    .X(chanx_left_out[0]));
 sky130_fd_sc_hd__clkbuf_2 output124 (.A(net124),
    .X(chanx_left_out[10]));
 sky130_fd_sc_hd__clkbuf_2 output125 (.A(net125),
    .X(chanx_left_out[11]));
 sky130_fd_sc_hd__clkbuf_2 output126 (.A(net126),
    .X(chanx_left_out[12]));
 sky130_fd_sc_hd__clkbuf_2 output127 (.A(net127),
    .X(chanx_left_out[13]));
 sky130_fd_sc_hd__clkbuf_2 output128 (.A(net128),
    .X(chanx_left_out[14]));
 sky130_fd_sc_hd__clkbuf_2 output129 (.A(net129),
    .X(chanx_left_out[15]));
 sky130_fd_sc_hd__clkbuf_2 output130 (.A(net130),
    .X(chanx_left_out[16]));
 sky130_fd_sc_hd__clkbuf_2 output131 (.A(net131),
    .X(chanx_left_out[17]));
 sky130_fd_sc_hd__clkbuf_2 output132 (.A(net132),
    .X(chanx_left_out[18]));
 sky130_fd_sc_hd__clkbuf_2 output133 (.A(net133),
    .X(chanx_left_out[19]));
 sky130_fd_sc_hd__clkbuf_2 output134 (.A(net134),
    .X(chanx_left_out[1]));
 sky130_fd_sc_hd__clkbuf_2 output135 (.A(net135),
    .X(chanx_left_out[2]));
 sky130_fd_sc_hd__clkbuf_2 output136 (.A(net136),
    .X(chanx_left_out[3]));
 sky130_fd_sc_hd__clkbuf_2 output137 (.A(net137),
    .X(chanx_left_out[4]));
 sky130_fd_sc_hd__clkbuf_2 output138 (.A(net138),
    .X(chanx_left_out[5]));
 sky130_fd_sc_hd__clkbuf_2 output139 (.A(net139),
    .X(chanx_left_out[6]));
 sky130_fd_sc_hd__clkbuf_2 output140 (.A(net140),
    .X(chanx_left_out[7]));
 sky130_fd_sc_hd__clkbuf_2 output141 (.A(net141),
    .X(chanx_left_out[8]));
 sky130_fd_sc_hd__clkbuf_2 output142 (.A(net142),
    .X(chanx_left_out[9]));
 sky130_fd_sc_hd__clkbuf_2 output143 (.A(net143),
    .X(chanx_right_out[0]));
 sky130_fd_sc_hd__clkbuf_2 output144 (.A(net144),
    .X(chanx_right_out[10]));
 sky130_fd_sc_hd__clkbuf_2 output145 (.A(net145),
    .X(chanx_right_out[11]));
 sky130_fd_sc_hd__clkbuf_2 output146 (.A(net146),
    .X(chanx_right_out[12]));
 sky130_fd_sc_hd__clkbuf_2 output147 (.A(net147),
    .X(chanx_right_out[13]));
 sky130_fd_sc_hd__clkbuf_2 output148 (.A(net148),
    .X(chanx_right_out[14]));
 sky130_fd_sc_hd__clkbuf_2 output149 (.A(net149),
    .X(chanx_right_out[15]));
 sky130_fd_sc_hd__clkbuf_2 output150 (.A(net150),
    .X(chanx_right_out[16]));
 sky130_fd_sc_hd__clkbuf_2 output151 (.A(net151),
    .X(chanx_right_out[17]));
 sky130_fd_sc_hd__clkbuf_2 output152 (.A(net152),
    .X(chanx_right_out[18]));
 sky130_fd_sc_hd__clkbuf_2 output153 (.A(net153),
    .X(chanx_right_out[19]));
 sky130_fd_sc_hd__clkbuf_2 output154 (.A(net154),
    .X(chanx_right_out[1]));
 sky130_fd_sc_hd__clkbuf_2 output155 (.A(net155),
    .X(chanx_right_out[2]));
 sky130_fd_sc_hd__clkbuf_2 output156 (.A(net156),
    .X(chanx_right_out[3]));
 sky130_fd_sc_hd__clkbuf_2 output157 (.A(net157),
    .X(chanx_right_out[4]));
 sky130_fd_sc_hd__clkbuf_2 output158 (.A(net158),
    .X(chanx_right_out[5]));
 sky130_fd_sc_hd__clkbuf_2 output159 (.A(net159),
    .X(chanx_right_out[6]));
 sky130_fd_sc_hd__clkbuf_2 output160 (.A(net160),
    .X(chanx_right_out[7]));
 sky130_fd_sc_hd__clkbuf_2 output161 (.A(net161),
    .X(chanx_right_out[8]));
 sky130_fd_sc_hd__clkbuf_2 output162 (.A(net162),
    .X(chanx_right_out[9]));
 sky130_fd_sc_hd__clkbuf_2 output163 (.A(net163),
    .X(chany_bottom_out[0]));
 sky130_fd_sc_hd__clkbuf_2 output164 (.A(net164),
    .X(chany_bottom_out[10]));
 sky130_fd_sc_hd__clkbuf_2 output165 (.A(net165),
    .X(chany_bottom_out[11]));
 sky130_fd_sc_hd__clkbuf_2 output166 (.A(net166),
    .X(chany_bottom_out[12]));
 sky130_fd_sc_hd__clkbuf_2 output167 (.A(net167),
    .X(chany_bottom_out[13]));
 sky130_fd_sc_hd__clkbuf_2 output168 (.A(net168),
    .X(chany_bottom_out[14]));
 sky130_fd_sc_hd__clkbuf_2 output169 (.A(net169),
    .X(chany_bottom_out[15]));
 sky130_fd_sc_hd__clkbuf_2 output170 (.A(net170),
    .X(chany_bottom_out[16]));
 sky130_fd_sc_hd__clkbuf_2 output171 (.A(net171),
    .X(chany_bottom_out[17]));
 sky130_fd_sc_hd__clkbuf_2 output172 (.A(net172),
    .X(chany_bottom_out[18]));
 sky130_fd_sc_hd__clkbuf_2 output173 (.A(net173),
    .X(chany_bottom_out[19]));
 sky130_fd_sc_hd__clkbuf_2 output174 (.A(net174),
    .X(chany_bottom_out[1]));
 sky130_fd_sc_hd__clkbuf_2 output175 (.A(net175),
    .X(chany_bottom_out[2]));
 sky130_fd_sc_hd__clkbuf_2 output176 (.A(net176),
    .X(chany_bottom_out[3]));
 sky130_fd_sc_hd__clkbuf_2 output177 (.A(net177),
    .X(chany_bottom_out[4]));
 sky130_fd_sc_hd__clkbuf_2 output178 (.A(net178),
    .X(chany_bottom_out[5]));
 sky130_fd_sc_hd__clkbuf_2 output179 (.A(net179),
    .X(chany_bottom_out[6]));
 sky130_fd_sc_hd__clkbuf_2 output180 (.A(net180),
    .X(chany_bottom_out[7]));
 sky130_fd_sc_hd__clkbuf_2 output181 (.A(net181),
    .X(chany_bottom_out[8]));
 sky130_fd_sc_hd__clkbuf_2 output182 (.A(net182),
    .X(chany_bottom_out[9]));
 sky130_fd_sc_hd__clkbuf_2 output183 (.A(net183),
    .X(chany_top_out[0]));
 sky130_fd_sc_hd__clkbuf_2 output184 (.A(net184),
    .X(chany_top_out[10]));
 sky130_fd_sc_hd__clkbuf_2 output185 (.A(net185),
    .X(chany_top_out[11]));
 sky130_fd_sc_hd__clkbuf_2 output186 (.A(net186),
    .X(chany_top_out[12]));
 sky130_fd_sc_hd__clkbuf_2 output187 (.A(net187),
    .X(chany_top_out[13]));
 sky130_fd_sc_hd__clkbuf_2 output188 (.A(net188),
    .X(chany_top_out[14]));
 sky130_fd_sc_hd__clkbuf_2 output189 (.A(net189),
    .X(chany_top_out[15]));
 sky130_fd_sc_hd__clkbuf_2 output190 (.A(net190),
    .X(chany_top_out[16]));
 sky130_fd_sc_hd__clkbuf_2 output191 (.A(net191),
    .X(chany_top_out[17]));
 sky130_fd_sc_hd__clkbuf_2 output192 (.A(net192),
    .X(chany_top_out[18]));
 sky130_fd_sc_hd__clkbuf_2 output193 (.A(net193),
    .X(chany_top_out[19]));
 sky130_fd_sc_hd__clkbuf_2 output194 (.A(net194),
    .X(chany_top_out[1]));
 sky130_fd_sc_hd__clkbuf_2 output195 (.A(net195),
    .X(chany_top_out[2]));
 sky130_fd_sc_hd__clkbuf_2 output196 (.A(net196),
    .X(chany_top_out[3]));
 sky130_fd_sc_hd__clkbuf_2 output197 (.A(net197),
    .X(chany_top_out[4]));
 sky130_fd_sc_hd__clkbuf_2 output198 (.A(net198),
    .X(chany_top_out[5]));
 sky130_fd_sc_hd__clkbuf_2 output199 (.A(net199),
    .X(chany_top_out[6]));
 sky130_fd_sc_hd__clkbuf_2 output200 (.A(net200),
    .X(chany_top_out[7]));
 sky130_fd_sc_hd__clkbuf_2 output201 (.A(net201),
    .X(chany_top_out[8]));
 sky130_fd_sc_hd__clkbuf_2 output202 (.A(net202),
    .X(chany_top_out[9]));
 sky130_fd_sc_hd__clkbuf_2 output203 (.A(net203),
    .X(clk_1_E_out));
 sky130_fd_sc_hd__clkbuf_2 output204 (.A(net204),
    .X(clk_1_W_out));
 sky130_fd_sc_hd__clkbuf_2 output205 (.A(net205),
    .X(clk_2_E_out));
 sky130_fd_sc_hd__clkbuf_2 output206 (.A(net206),
    .X(clk_2_N_out));
 sky130_fd_sc_hd__clkbuf_2 output207 (.A(net207),
    .X(clk_2_S_out));
 sky130_fd_sc_hd__clkbuf_2 output208 (.A(net208),
    .X(clk_2_W_out));
 sky130_fd_sc_hd__clkbuf_2 output209 (.A(net209),
    .X(clk_3_E_out));
 sky130_fd_sc_hd__clkbuf_2 output210 (.A(net210),
    .X(clk_3_N_out));
 sky130_fd_sc_hd__clkbuf_2 output211 (.A(net211),
    .X(clk_3_S_out));
 sky130_fd_sc_hd__clkbuf_2 output212 (.A(net212),
    .X(clk_3_W_out));
 sky130_fd_sc_hd__clkbuf_2 output213 (.A(net213),
    .X(prog_clk_1_E_out));
 sky130_fd_sc_hd__clkbuf_2 output214 (.A(net214),
    .X(prog_clk_1_W_out));
 sky130_fd_sc_hd__buf_1 output215 (.A(net215),
    .X(prog_clk_2_E_out));
 sky130_fd_sc_hd__buf_1 output216 (.A(net216),
    .X(prog_clk_2_N_out));
 sky130_fd_sc_hd__buf_1 output217 (.A(net217),
    .X(prog_clk_2_S_out));
 sky130_fd_sc_hd__buf_1 output218 (.A(net218),
    .X(prog_clk_2_W_out));
 sky130_fd_sc_hd__clkbuf_2 output219 (.A(net219),
    .X(prog_clk_3_E_out));
 sky130_fd_sc_hd__clkbuf_2 output220 (.A(net220),
    .X(prog_clk_3_N_out));
 sky130_fd_sc_hd__clkbuf_2 output221 (.A(net221),
    .X(prog_clk_3_S_out));
 sky130_fd_sc_hd__clkbuf_2 output222 (.A(net222),
    .X(prog_clk_3_W_out));
 sky130_fd_sc_hd__clkbuf_16 prog_clk_0_FTB00 (.A(net102),
    .X(\mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 prog_clk_1_E_FTB01 (.A(net103),
    .X(net213));
 sky130_fd_sc_hd__buf_1 prog_clk_1_W_FTB01 (.A(net103),
    .X(net214));
 sky130_fd_sc_hd__buf_4 prog_clk_2_E_FTB01 (.A(prog_clk_2_N_in),
    .X(net215));
 sky130_fd_sc_hd__buf_4 prog_clk_2_N_FTB01 (.A(prog_clk_2_N_in),
    .X(net216));
 sky130_fd_sc_hd__buf_4 prog_clk_2_S_FTB01 (.A(prog_clk_2_N_in),
    .X(net217));
 sky130_fd_sc_hd__buf_4 prog_clk_2_W_FTB01 (.A(prog_clk_2_N_in),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_1 prog_clk_3_E_FTB01 (.A(net104),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_1 prog_clk_3_N_FTB01 (.A(net104),
    .X(net220));
 sky130_fd_sc_hd__buf_1 prog_clk_3_S_FTB01 (.A(net104),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 prog_clk_3_W_FTB01 (.A(net104),
    .X(net222));
endmodule
