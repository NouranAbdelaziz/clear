magic
tech sky130A
magscale 1 2
timestamp 1650893984
<< viali >>
rect 10333 20553 10367 20587
rect 13277 20553 13311 20587
rect 13829 20553 13863 20587
rect 14289 20553 14323 20587
rect 14749 20553 14783 20587
rect 15209 20553 15243 20587
rect 15669 20553 15703 20587
rect 16129 20553 16163 20587
rect 16865 20553 16899 20587
rect 17601 20553 17635 20587
rect 17969 20553 18003 20587
rect 18429 20553 18463 20587
rect 18889 20553 18923 20587
rect 19441 20553 19475 20587
rect 19809 20553 19843 20587
rect 20269 20553 20303 20587
rect 20729 20553 20763 20587
rect 21189 20553 21223 20587
rect 3249 20485 3283 20519
rect 8033 20485 8067 20519
rect 11161 20485 11195 20519
rect 16405 20485 16439 20519
rect 2053 20417 2087 20451
rect 2973 20417 3007 20451
rect 3525 20417 3559 20451
rect 4353 20417 4387 20451
rect 4905 20417 4939 20451
rect 5457 20417 5491 20451
rect 6009 20417 6043 20451
rect 6377 20417 6411 20451
rect 7205 20417 7239 20451
rect 8769 20417 8803 20451
rect 10241 20417 10275 20451
rect 10885 20417 10919 20451
rect 11529 20417 11563 20451
rect 13093 20417 13127 20451
rect 13461 20417 13495 20451
rect 13645 20417 13679 20451
rect 14105 20417 14139 20451
rect 14565 20417 14599 20451
rect 15025 20417 15059 20451
rect 15485 20417 15519 20451
rect 15945 20417 15979 20451
rect 16681 20417 16715 20451
rect 17049 20417 17083 20451
rect 17417 20417 17451 20451
rect 17785 20417 17819 20451
rect 18245 20417 18279 20451
rect 18705 20417 18739 20451
rect 19257 20417 19291 20451
rect 19625 20417 19659 20451
rect 20085 20417 20119 20451
rect 20545 20417 20579 20451
rect 21005 20417 21039 20451
rect 21557 20417 21591 20451
rect 2697 20349 2731 20383
rect 4629 20349 4663 20383
rect 5549 20349 5583 20383
rect 5641 20349 5675 20383
rect 8953 20349 8987 20383
rect 9229 20349 9263 20383
rect 10425 20349 10459 20383
rect 10701 20349 10735 20383
rect 12817 20349 12851 20383
rect 1409 20281 1443 20315
rect 5089 20281 5123 20315
rect 7021 20281 7055 20315
rect 12173 20281 12207 20315
rect 17233 20281 17267 20315
rect 3433 20213 3467 20247
rect 4813 20213 4847 20247
rect 6101 20213 6135 20247
rect 7849 20213 7883 20247
rect 8125 20213 8159 20247
rect 9873 20213 9907 20247
rect 11253 20213 11287 20247
rect 21373 20213 21407 20247
rect 5641 20009 5675 20043
rect 10977 20009 11011 20043
rect 13553 20009 13587 20043
rect 14289 20009 14323 20043
rect 14841 20009 14875 20043
rect 15117 20009 15151 20043
rect 15393 20009 15427 20043
rect 16129 20009 16163 20043
rect 17693 20009 17727 20043
rect 17969 20009 18003 20043
rect 18245 20009 18279 20043
rect 18521 20009 18555 20043
rect 19441 20009 19475 20043
rect 19809 20009 19843 20043
rect 20821 20009 20855 20043
rect 21465 20009 21499 20043
rect 6469 19941 6503 19975
rect 10885 19941 10919 19975
rect 13829 19941 13863 19975
rect 14565 19941 14599 19975
rect 15853 19941 15887 19975
rect 21097 19941 21131 19975
rect 2237 19873 2271 19907
rect 2881 19873 2915 19907
rect 6193 19873 6227 19907
rect 7113 19873 7147 19907
rect 7941 19873 7975 19907
rect 12449 19873 12483 19907
rect 1961 19805 1995 19839
rect 3157 19805 3191 19839
rect 3525 19805 3559 19839
rect 3985 19805 4019 19839
rect 4077 19805 4111 19839
rect 6101 19805 6135 19839
rect 6837 19805 6871 19839
rect 8769 19805 8803 19839
rect 10066 19805 10100 19839
rect 10333 19805 10367 19839
rect 12357 19805 12391 19839
rect 12725 19805 12759 19839
rect 13369 19805 13403 19839
rect 13645 19805 13679 19839
rect 14105 19805 14139 19839
rect 14381 19805 14415 19839
rect 14657 19805 14691 19839
rect 14933 19805 14967 19839
rect 15209 19805 15243 19839
rect 15669 19805 15703 19839
rect 15945 19805 15979 19839
rect 17417 19805 17451 19839
rect 17509 19805 17543 19839
rect 17785 19805 17819 19839
rect 18061 19805 18095 19839
rect 18337 19805 18371 19839
rect 19257 19805 19291 19839
rect 19625 19805 19659 19839
rect 20913 19805 20947 19839
rect 21281 19805 21315 19839
rect 4322 19737 4356 19771
rect 7757 19737 7791 19771
rect 10609 19737 10643 19771
rect 12112 19737 12146 19771
rect 16221 19737 16255 19771
rect 16589 19737 16623 19771
rect 19901 19737 19935 19771
rect 3433 19669 3467 19703
rect 3801 19669 3835 19703
rect 5457 19669 5491 19703
rect 6009 19669 6043 19703
rect 6929 19669 6963 19703
rect 7297 19669 7331 19703
rect 7665 19669 7699 19703
rect 8125 19669 8159 19703
rect 8953 19669 8987 19703
rect 10517 19669 10551 19703
rect 15485 19669 15519 19703
rect 18613 19669 18647 19703
rect 2329 19465 2363 19499
rect 3157 19465 3191 19499
rect 4813 19465 4847 19499
rect 7113 19465 7147 19499
rect 8677 19465 8711 19499
rect 11069 19465 11103 19499
rect 11713 19465 11747 19499
rect 12725 19465 12759 19499
rect 12817 19465 12851 19499
rect 13277 19465 13311 19499
rect 13553 19465 13587 19499
rect 14381 19465 14415 19499
rect 14749 19465 14783 19499
rect 15209 19465 15243 19499
rect 16221 19465 16255 19499
rect 16865 19465 16899 19499
rect 17141 19465 17175 19499
rect 18889 19465 18923 19499
rect 2697 19397 2731 19431
rect 8226 19397 8260 19431
rect 9790 19397 9824 19431
rect 10241 19397 10275 19431
rect 10425 19397 10459 19431
rect 12173 19397 12207 19431
rect 4281 19329 4315 19363
rect 4537 19329 4571 19363
rect 5926 19329 5960 19363
rect 6186 19329 6220 19363
rect 6377 19329 6411 19363
rect 7021 19329 7055 19363
rect 10977 19329 11011 19363
rect 12081 19329 12115 19363
rect 12541 19329 12575 19363
rect 13001 19329 13035 19363
rect 13093 19329 13127 19363
rect 13369 19329 13403 19363
rect 14565 19329 14599 19363
rect 15025 19329 15059 19363
rect 16037 19329 16071 19363
rect 16681 19329 16715 19363
rect 16957 19329 16991 19363
rect 18705 19329 18739 19363
rect 2237 19261 2271 19295
rect 2789 19261 2823 19295
rect 2973 19261 3007 19295
rect 8493 19261 8527 19295
rect 10057 19261 10091 19295
rect 11253 19261 11287 19295
rect 12265 19261 12299 19295
rect 13829 19261 13863 19295
rect 17693 19261 17727 19295
rect 13645 19193 13679 19227
rect 14013 19193 14047 19227
rect 14841 19193 14875 19227
rect 15485 19193 15519 19227
rect 2007 19125 2041 19159
rect 4721 19125 4755 19159
rect 10609 19125 10643 19159
rect 11529 19125 11563 19159
rect 14289 19125 14323 19159
rect 15301 19125 15335 19159
rect 15669 19125 15703 19159
rect 15853 19125 15887 19159
rect 17233 19125 17267 19159
rect 17417 19125 17451 19159
rect 17785 19125 17819 19159
rect 18521 19125 18555 19159
rect 1501 18921 1535 18955
rect 2881 18921 2915 18955
rect 6653 18921 6687 18955
rect 12725 18921 12759 18955
rect 13001 18921 13035 18955
rect 13829 18921 13863 18955
rect 14657 18921 14691 18955
rect 1869 18853 1903 18887
rect 10517 18853 10551 18887
rect 11989 18853 12023 18887
rect 13093 18853 13127 18887
rect 13461 18853 13495 18887
rect 14289 18853 14323 18887
rect 3341 18785 3375 18819
rect 3525 18785 3559 18819
rect 4353 18785 4387 18819
rect 6561 18785 6595 18819
rect 9413 18785 9447 18819
rect 9505 18785 9539 18819
rect 9965 18785 9999 18819
rect 10609 18785 10643 18819
rect 14473 18785 14507 18819
rect 1685 18717 1719 18751
rect 2053 18717 2087 18751
rect 2789 18717 2823 18751
rect 4905 18717 4939 18751
rect 6305 18717 6339 18751
rect 6837 18717 6871 18751
rect 8309 18717 8343 18751
rect 8677 18717 8711 18751
rect 12081 18717 12115 18751
rect 12817 18717 12851 18751
rect 13369 18717 13403 18751
rect 4721 18649 4755 18683
rect 8042 18649 8076 18683
rect 10876 18649 10910 18683
rect 13645 18649 13679 18683
rect 14841 18649 14875 18683
rect 2145 18581 2179 18615
rect 3249 18581 3283 18615
rect 3801 18581 3835 18615
rect 4169 18581 4203 18615
rect 4261 18581 4295 18615
rect 5181 18581 5215 18615
rect 6929 18581 6963 18615
rect 8585 18581 8619 18615
rect 8953 18581 8987 18615
rect 9321 18581 9355 18615
rect 10057 18581 10091 18615
rect 10149 18581 10183 18615
rect 14105 18581 14139 18615
rect 1869 18377 1903 18411
rect 2237 18377 2271 18411
rect 2789 18377 2823 18411
rect 4445 18377 4479 18411
rect 4905 18377 4939 18411
rect 6377 18377 6411 18411
rect 7481 18377 7515 18411
rect 8401 18377 8435 18411
rect 8861 18377 8895 18411
rect 9505 18377 9539 18411
rect 10793 18377 10827 18411
rect 11161 18377 11195 18411
rect 11529 18377 11563 18411
rect 11805 18377 11839 18411
rect 13645 18377 13679 18411
rect 13921 18377 13955 18411
rect 3924 18309 3958 18343
rect 5273 18309 5307 18343
rect 14013 18309 14047 18343
rect 1685 18241 1719 18275
rect 2053 18241 2087 18275
rect 2421 18241 2455 18275
rect 2513 18241 2547 18275
rect 4169 18241 4203 18275
rect 4813 18241 4847 18275
rect 5917 18241 5951 18275
rect 6193 18241 6227 18275
rect 6561 18241 6595 18275
rect 7021 18241 7055 18275
rect 8125 18241 8159 18275
rect 8585 18241 8619 18275
rect 9137 18241 9171 18275
rect 9413 18241 9447 18275
rect 9781 18241 9815 18275
rect 10701 18241 10735 18275
rect 11713 18241 11747 18275
rect 12929 18241 12963 18275
rect 13185 18241 13219 18275
rect 13461 18241 13495 18275
rect 5089 18173 5123 18207
rect 6745 18173 6779 18207
rect 6929 18173 6963 18207
rect 6009 18105 6043 18139
rect 8309 18105 8343 18139
rect 8953 18105 8987 18139
rect 9229 18105 9263 18139
rect 1501 18037 1535 18071
rect 2697 18037 2731 18071
rect 4353 18037 4387 18071
rect 7389 18037 7423 18071
rect 10425 18037 10459 18071
rect 10517 18037 10551 18071
rect 13277 18037 13311 18071
rect 1869 17833 1903 17867
rect 2237 17833 2271 17867
rect 2605 17833 2639 17867
rect 3065 17833 3099 17867
rect 3433 17833 3467 17867
rect 10333 17833 10367 17867
rect 13277 17833 13311 17867
rect 13829 17833 13863 17867
rect 8769 17765 8803 17799
rect 7481 17697 7515 17731
rect 8401 17697 8435 17731
rect 9045 17697 9079 17731
rect 10977 17697 11011 17731
rect 1685 17629 1719 17663
rect 2053 17629 2087 17663
rect 2421 17629 2455 17663
rect 2789 17629 2823 17663
rect 2881 17629 2915 17663
rect 3249 17629 3283 17663
rect 3801 17629 3835 17663
rect 5273 17629 5307 17663
rect 6009 17629 6043 17663
rect 7205 17629 7239 17663
rect 7757 17629 7791 17663
rect 8309 17629 8343 17663
rect 10241 17629 10275 17663
rect 11161 17629 11195 17663
rect 12633 17629 12667 17663
rect 13645 17629 13679 17663
rect 21281 17629 21315 17663
rect 4046 17561 4080 17595
rect 7297 17561 7331 17595
rect 8217 17561 8251 17595
rect 9321 17561 9355 17595
rect 9781 17561 9815 17595
rect 10701 17561 10735 17595
rect 11428 17561 11462 17595
rect 1501 17493 1535 17527
rect 5181 17493 5215 17527
rect 5917 17493 5951 17527
rect 6653 17493 6687 17527
rect 6837 17493 6871 17527
rect 7849 17493 7883 17527
rect 9229 17493 9263 17527
rect 9689 17493 9723 17527
rect 10057 17493 10091 17527
rect 10793 17493 10827 17527
rect 12541 17493 12575 17527
rect 13369 17493 13403 17527
rect 21097 17493 21131 17527
rect 21465 17493 21499 17527
rect 3525 17289 3559 17323
rect 3893 17289 3927 17323
rect 6377 17289 6411 17323
rect 11621 17289 11655 17323
rect 12081 17289 12115 17323
rect 12633 17289 12667 17323
rect 13369 17289 13403 17323
rect 5856 17221 5890 17255
rect 1685 17153 1719 17187
rect 2053 17153 2087 17187
rect 2237 17153 2271 17187
rect 2513 17153 2547 17187
rect 3433 17153 3467 17187
rect 4261 17153 4295 17187
rect 6561 17153 6595 17187
rect 6837 17153 6871 17187
rect 7196 17153 7230 17187
rect 8401 17153 8435 17187
rect 8657 17153 8691 17187
rect 9873 17153 9907 17187
rect 10140 17153 10174 17187
rect 11989 17153 12023 17187
rect 13185 17153 13219 17187
rect 2973 17085 3007 17119
rect 3709 17085 3743 17119
rect 4353 17085 4387 17119
rect 4537 17085 4571 17119
rect 6101 17085 6135 17119
rect 6929 17085 6963 17119
rect 12173 17085 12207 17119
rect 12541 17085 12575 17119
rect 1869 17017 1903 17051
rect 2697 17017 2731 17051
rect 4721 17017 4755 17051
rect 9781 17017 9815 17051
rect 11253 17017 11287 17051
rect 1501 16949 1535 16983
rect 2421 16949 2455 16983
rect 3065 16949 3099 16983
rect 8309 16949 8343 16983
rect 1869 16745 1903 16779
rect 3249 16745 3283 16779
rect 3617 16745 3651 16779
rect 7849 16745 7883 16779
rect 8953 16745 8987 16779
rect 9229 16745 9263 16779
rect 11253 16745 11287 16779
rect 12265 16745 12299 16779
rect 13553 16745 13587 16779
rect 6377 16677 6411 16711
rect 9413 16677 9447 16711
rect 3801 16609 3835 16643
rect 4721 16609 4755 16643
rect 4997 16609 5031 16643
rect 8769 16609 8803 16643
rect 10149 16609 10183 16643
rect 10609 16609 10643 16643
rect 10701 16609 10735 16643
rect 11805 16609 11839 16643
rect 13001 16609 13035 16643
rect 1685 16541 1719 16575
rect 2053 16541 2087 16575
rect 2329 16541 2363 16575
rect 2421 16541 2455 16575
rect 2697 16541 2731 16575
rect 2973 16541 3007 16575
rect 3433 16541 3467 16575
rect 5264 16541 5298 16575
rect 6469 16541 6503 16575
rect 6736 16541 6770 16575
rect 7941 16541 7975 16575
rect 8585 16541 8619 16575
rect 10057 16541 10091 16575
rect 14105 16541 14139 16575
rect 4537 16473 4571 16507
rect 11621 16473 11655 16507
rect 1501 16405 1535 16439
rect 2145 16405 2179 16439
rect 2605 16405 2639 16439
rect 2881 16405 2915 16439
rect 3157 16405 3191 16439
rect 4077 16405 4111 16439
rect 4445 16405 4479 16439
rect 9597 16405 9631 16439
rect 9965 16405 9999 16439
rect 10793 16405 10827 16439
rect 11161 16405 11195 16439
rect 11713 16405 11747 16439
rect 12081 16405 12115 16439
rect 13093 16405 13127 16439
rect 13185 16405 13219 16439
rect 14749 16405 14783 16439
rect 1869 16201 1903 16235
rect 2421 16201 2455 16235
rect 2881 16201 2915 16235
rect 5273 16201 5307 16235
rect 6837 16201 6871 16235
rect 7389 16201 7423 16235
rect 8217 16201 8251 16235
rect 9505 16201 9539 16235
rect 9965 16201 9999 16235
rect 10149 16201 10183 16235
rect 11805 16201 11839 16235
rect 12265 16201 12299 16235
rect 13829 16201 13863 16235
rect 9413 16133 9447 16167
rect 1685 16065 1719 16099
rect 2053 16065 2087 16099
rect 2329 16065 2363 16099
rect 2605 16065 2639 16099
rect 2697 16065 2731 16099
rect 2973 16065 3007 16099
rect 3433 16065 3467 16099
rect 3893 16065 3927 16099
rect 4160 16065 4194 16099
rect 5457 16065 5491 16099
rect 6745 16065 6779 16099
rect 7205 16065 7239 16099
rect 7757 16065 7791 16099
rect 8585 16065 8619 16099
rect 11897 16065 11931 16099
rect 12705 16065 12739 16099
rect 3801 15997 3835 16031
rect 6929 15997 6963 16031
rect 7849 15997 7883 16031
rect 7941 15997 7975 16031
rect 8677 15997 8711 16031
rect 8769 15997 8803 16031
rect 9597 15997 9631 16031
rect 10977 15997 11011 16031
rect 11253 15997 11287 16031
rect 11713 15997 11747 16031
rect 12449 15997 12483 16031
rect 1501 15929 1535 15963
rect 2145 15929 2179 15963
rect 3249 15929 3283 15963
rect 6377 15929 6411 15963
rect 3157 15861 3191 15895
rect 6101 15861 6135 15895
rect 9045 15861 9079 15895
rect 10333 15861 10367 15895
rect 2145 15657 2179 15691
rect 2697 15657 2731 15691
rect 3433 15657 3467 15691
rect 3893 15657 3927 15691
rect 4721 15657 4755 15691
rect 5549 15657 5583 15691
rect 8493 15657 8527 15691
rect 13553 15657 13587 15691
rect 2421 15589 2455 15623
rect 2973 15589 3007 15623
rect 4905 15589 4939 15623
rect 9229 15589 9263 15623
rect 3525 15521 3559 15555
rect 4169 15521 4203 15555
rect 7113 15521 7147 15555
rect 9413 15521 9447 15555
rect 12173 15521 12207 15555
rect 13001 15521 13035 15555
rect 1685 15453 1719 15487
rect 2053 15453 2087 15487
rect 2329 15453 2363 15487
rect 2605 15453 2639 15487
rect 2881 15453 2915 15487
rect 3157 15453 3191 15487
rect 3249 15453 3283 15487
rect 4353 15453 4387 15487
rect 5089 15453 5123 15487
rect 8677 15453 8711 15487
rect 14105 15453 14139 15487
rect 14372 15453 14406 15487
rect 16221 15453 16255 15487
rect 7021 15385 7055 15419
rect 7358 15385 7392 15419
rect 10425 15385 10459 15419
rect 13093 15385 13127 15419
rect 1501 15317 1535 15351
rect 1869 15317 1903 15351
rect 4261 15317 4295 15351
rect 9137 15317 9171 15351
rect 13185 15317 13219 15351
rect 15485 15317 15519 15351
rect 15577 15317 15611 15351
rect 1869 15113 1903 15147
rect 2329 15113 2363 15147
rect 3157 15113 3191 15147
rect 3249 15113 3283 15147
rect 6377 15113 6411 15147
rect 8217 15113 8251 15147
rect 8585 15113 8619 15147
rect 9413 15113 9447 15147
rect 11253 15113 11287 15147
rect 12909 15113 12943 15147
rect 13001 15113 13035 15147
rect 13829 15113 13863 15147
rect 14289 15113 14323 15147
rect 14657 15113 14691 15147
rect 4322 15045 4356 15079
rect 1685 14977 1719 15011
rect 2053 14977 2087 15011
rect 2145 14977 2179 15011
rect 2605 14977 2639 15011
rect 2697 14977 2731 15011
rect 2973 14977 3007 15011
rect 3617 14977 3651 15011
rect 6193 14977 6227 15011
rect 7490 14977 7524 15011
rect 7757 14977 7791 15011
rect 8677 14977 8711 15011
rect 9321 14977 9355 15011
rect 9873 14977 9907 15011
rect 10140 14977 10174 15011
rect 11529 14977 11563 15011
rect 11796 14977 11830 15011
rect 13369 14977 13403 15011
rect 14197 14977 14231 15011
rect 15025 14977 15059 15011
rect 3709 14909 3743 14943
rect 3801 14909 3835 14943
rect 4077 14909 4111 14943
rect 7849 14909 7883 14943
rect 8769 14909 8803 14943
rect 9229 14909 9263 14943
rect 13461 14909 13495 14943
rect 13553 14909 13587 14943
rect 14381 14909 14415 14943
rect 15117 14909 15151 14943
rect 15209 14909 15243 14943
rect 2421 14841 2455 14875
rect 2881 14841 2915 14875
rect 5457 14841 5491 14875
rect 1501 14773 1535 14807
rect 5549 14773 5583 14807
rect 9781 14773 9815 14807
rect 15577 14773 15611 14807
rect 1961 14569 1995 14603
rect 4445 14569 4479 14603
rect 7665 14569 7699 14603
rect 9137 14569 9171 14603
rect 10241 14569 10275 14603
rect 11529 14569 11563 14603
rect 13737 14569 13771 14603
rect 6929 14501 6963 14535
rect 9229 14501 9263 14535
rect 3617 14433 3651 14467
rect 4997 14433 5031 14467
rect 8309 14433 8343 14467
rect 9689 14433 9723 14467
rect 11161 14433 11195 14467
rect 12081 14433 12115 14467
rect 12633 14433 12667 14467
rect 13093 14433 13127 14467
rect 16589 14433 16623 14467
rect 1685 14365 1719 14399
rect 2145 14365 2179 14399
rect 4261 14365 4295 14399
rect 5549 14365 5583 14399
rect 5816 14365 5850 14399
rect 7021 14365 7055 14399
rect 9781 14365 9815 14399
rect 15678 14365 15712 14399
rect 15945 14365 15979 14399
rect 1777 14297 1811 14331
rect 3350 14297 3384 14331
rect 4813 14297 4847 14331
rect 10425 14297 10459 14331
rect 11069 14297 11103 14331
rect 16497 14297 16531 14331
rect 1501 14229 1535 14263
rect 2237 14229 2271 14263
rect 3801 14229 3835 14263
rect 4077 14229 4111 14263
rect 4905 14229 4939 14263
rect 5273 14229 5307 14263
rect 7757 14229 7791 14263
rect 8125 14229 8159 14263
rect 8217 14229 8251 14263
rect 9873 14229 9907 14263
rect 10609 14229 10643 14263
rect 10977 14229 11011 14263
rect 11897 14229 11931 14263
rect 11989 14229 12023 14263
rect 12725 14229 12759 14263
rect 13277 14229 13311 14263
rect 13369 14229 13403 14263
rect 13829 14229 13863 14263
rect 14565 14229 14599 14263
rect 16037 14229 16071 14263
rect 16405 14229 16439 14263
rect 1869 14025 1903 14059
rect 2145 14025 2179 14059
rect 3157 14025 3191 14059
rect 3617 14025 3651 14059
rect 3985 14025 4019 14059
rect 4077 14025 4111 14059
rect 7573 14025 7607 14059
rect 9413 14025 9447 14059
rect 10701 14025 10735 14059
rect 11161 14025 11195 14059
rect 13185 14025 13219 14059
rect 13829 14025 13863 14059
rect 14933 14025 14967 14059
rect 15761 14025 15795 14059
rect 5212 13957 5246 13991
rect 6193 13957 6227 13991
rect 10793 13957 10827 13991
rect 13277 13957 13311 13991
rect 15025 13957 15059 13991
rect 1685 13889 1719 13923
rect 2053 13889 2087 13923
rect 2329 13889 2363 13923
rect 2513 13889 2547 13923
rect 5549 13889 5583 13923
rect 6377 13889 6411 13923
rect 7481 13889 7515 13923
rect 9065 13889 9099 13923
rect 9781 13889 9815 13923
rect 11529 13889 11563 13923
rect 13737 13889 13771 13923
rect 15853 13889 15887 13923
rect 3433 13821 3467 13855
rect 3525 13821 3559 13855
rect 5457 13821 5491 13855
rect 7665 13821 7699 13855
rect 9321 13821 9355 13855
rect 9873 13821 9907 13855
rect 10057 13821 10091 13855
rect 10609 13821 10643 13855
rect 11345 13821 11379 13855
rect 13461 13821 13495 13855
rect 14749 13821 14783 13855
rect 7021 13753 7055 13787
rect 12817 13753 12851 13787
rect 1501 13685 1535 13719
rect 7113 13685 7147 13719
rect 7941 13685 7975 13719
rect 12633 13685 12667 13719
rect 15393 13685 15427 13719
rect 1777 13481 1811 13515
rect 3157 13481 3191 13515
rect 3433 13481 3467 13515
rect 4077 13481 4111 13515
rect 5181 13481 5215 13515
rect 7941 13481 7975 13515
rect 9045 13481 9079 13515
rect 9321 13481 9355 13515
rect 16313 13481 16347 13515
rect 3801 13413 3835 13447
rect 8033 13413 8067 13447
rect 15761 13413 15795 13447
rect 2605 13345 2639 13379
rect 4629 13345 4663 13379
rect 7389 13345 7423 13379
rect 8677 13345 8711 13379
rect 9781 13345 9815 13379
rect 15117 13345 15151 13379
rect 1409 13277 1443 13311
rect 1961 13277 1995 13311
rect 2881 13277 2915 13311
rect 3341 13277 3375 13311
rect 4721 13277 4755 13311
rect 7021 13277 7055 13311
rect 10425 13277 10459 13311
rect 12357 13277 12391 13311
rect 14105 13277 14139 13311
rect 17693 13277 17727 13311
rect 4353 13209 4387 13243
rect 4813 13209 4847 13243
rect 7573 13209 7607 13243
rect 8493 13209 8527 13243
rect 12624 13209 12658 13243
rect 14749 13209 14783 13243
rect 15853 13209 15887 13243
rect 17448 13209 17482 13243
rect 1593 13141 1627 13175
rect 2053 13141 2087 13175
rect 2421 13141 2455 13175
rect 2513 13141 2547 13175
rect 3065 13141 3099 13175
rect 5733 13141 5767 13175
rect 7481 13141 7515 13175
rect 8401 13141 8435 13175
rect 9873 13141 9907 13175
rect 9965 13141 9999 13175
rect 10333 13141 10367 13175
rect 11713 13141 11747 13175
rect 13737 13141 13771 13175
rect 14933 13141 14967 13175
rect 15301 13141 15335 13175
rect 15393 13141 15427 13175
rect 1869 12937 1903 12971
rect 1961 12937 1995 12971
rect 2329 12937 2363 12971
rect 2421 12937 2455 12971
rect 2789 12937 2823 12971
rect 3249 12937 3283 12971
rect 3617 12937 3651 12971
rect 6377 12937 6411 12971
rect 6561 12937 6595 12971
rect 6929 12937 6963 12971
rect 12909 12937 12943 12971
rect 13369 12937 13403 12971
rect 13737 12937 13771 12971
rect 14289 12937 14323 12971
rect 14749 12937 14783 12971
rect 15117 12937 15151 12971
rect 15485 12937 15519 12971
rect 15577 12937 15611 12971
rect 4077 12869 4111 12903
rect 1409 12801 1443 12835
rect 1685 12801 1719 12835
rect 3157 12801 3191 12835
rect 3985 12801 4019 12835
rect 4813 12801 4847 12835
rect 5069 12801 5103 12835
rect 7645 12801 7679 12835
rect 9229 12801 9263 12835
rect 9496 12801 9530 12835
rect 11529 12801 11563 12835
rect 11796 12801 11830 12835
rect 14657 12801 14691 12835
rect 2605 12733 2639 12767
rect 3341 12733 3375 12767
rect 4169 12733 4203 12767
rect 7021 12733 7055 12767
rect 7205 12733 7239 12767
rect 7389 12733 7423 12767
rect 13185 12733 13219 12767
rect 13277 12733 13311 12767
rect 14841 12733 14875 12767
rect 15669 12733 15703 12767
rect 4537 12665 4571 12699
rect 6193 12665 6227 12699
rect 1593 12597 1627 12631
rect 4721 12597 4755 12631
rect 8769 12597 8803 12631
rect 10609 12597 10643 12631
rect 3433 12393 3467 12427
rect 5457 12393 5491 12427
rect 8585 12393 8619 12427
rect 9597 12393 9631 12427
rect 9689 12393 9723 12427
rect 10517 12393 10551 12427
rect 12725 12393 12759 12427
rect 5549 12257 5583 12291
rect 7941 12257 7975 12291
rect 10333 12257 10367 12291
rect 12173 12257 12207 12291
rect 13369 12257 13403 12291
rect 1409 12189 1443 12223
rect 1685 12189 1719 12223
rect 3341 12189 3375 12223
rect 4077 12189 4111 12223
rect 5917 12189 5951 12223
rect 8953 12189 8987 12223
rect 11897 12189 11931 12223
rect 14289 12189 14323 12223
rect 15761 12189 15795 12223
rect 3096 12121 3130 12155
rect 4322 12121 4356 12155
rect 6162 12121 6196 12155
rect 8033 12121 8067 12155
rect 10149 12121 10183 12155
rect 11630 12121 11664 12155
rect 13185 12121 13219 12155
rect 14556 12121 14590 12155
rect 1593 12053 1627 12087
rect 1869 12053 1903 12087
rect 1961 12053 1995 12087
rect 3801 12053 3835 12087
rect 7297 12053 7331 12087
rect 8125 12053 8159 12087
rect 8493 12053 8527 12087
rect 10057 12053 10091 12087
rect 12265 12053 12299 12087
rect 12357 12053 12391 12087
rect 12817 12053 12851 12087
rect 13277 12053 13311 12087
rect 15669 12053 15703 12087
rect 16405 12053 16439 12087
rect 1501 11849 1535 11883
rect 3709 11849 3743 11883
rect 4169 11849 4203 11883
rect 4813 11849 4847 11883
rect 5825 11849 5859 11883
rect 6837 11849 6871 11883
rect 7297 11849 7331 11883
rect 8217 11849 8251 11883
rect 8309 11849 8343 11883
rect 9045 11849 9079 11883
rect 9137 11849 9171 11883
rect 9505 11849 9539 11883
rect 10057 11849 10091 11883
rect 11897 11849 11931 11883
rect 13185 11849 13219 11883
rect 13553 11849 13587 11883
rect 14289 11849 14323 11883
rect 15761 11849 15795 11883
rect 2614 11781 2648 11815
rect 6929 11781 6963 11815
rect 11345 11781 11379 11815
rect 13737 11781 13771 11815
rect 2881 11713 2915 11747
rect 2973 11713 3007 11747
rect 4077 11713 4111 11747
rect 5457 11713 5491 11747
rect 12357 11713 12391 11747
rect 15413 11713 15447 11747
rect 15669 11713 15703 11747
rect 16129 11713 16163 11747
rect 4261 11645 4295 11679
rect 5181 11645 5215 11679
rect 5365 11645 5399 11679
rect 5917 11645 5951 11679
rect 6745 11645 6779 11679
rect 7389 11645 7423 11679
rect 8125 11645 8159 11679
rect 8861 11645 8895 11679
rect 12081 11645 12115 11679
rect 12265 11645 12299 11679
rect 12909 11645 12943 11679
rect 13093 11645 13127 11679
rect 16221 11645 16255 11679
rect 16313 11645 16347 11679
rect 3617 11509 3651 11543
rect 4629 11509 4663 11543
rect 4905 11509 4939 11543
rect 6377 11509 6411 11543
rect 8677 11509 8711 11543
rect 11529 11509 11563 11543
rect 12725 11509 12759 11543
rect 1409 11305 1443 11339
rect 2329 11305 2363 11339
rect 3893 11305 3927 11339
rect 5365 11305 5399 11339
rect 7021 11305 7055 11339
rect 8585 11305 8619 11339
rect 10517 11305 10551 11339
rect 14197 11305 14231 11339
rect 4445 11237 4479 11271
rect 6193 11237 6227 11271
rect 12081 11237 12115 11271
rect 13093 11237 13127 11271
rect 14749 11237 14783 11271
rect 1777 11169 1811 11203
rect 2881 11169 2915 11203
rect 3065 11169 3099 11203
rect 3617 11169 3651 11203
rect 4813 11169 4847 11203
rect 5641 11169 5675 11203
rect 6469 11169 6503 11203
rect 11069 11169 11103 11203
rect 11529 11169 11563 11203
rect 12817 11169 12851 11203
rect 13645 11169 13679 11203
rect 4997 11101 5031 11135
rect 6653 11101 6687 11135
rect 7205 11101 7239 11135
rect 8953 11101 8987 11135
rect 10977 11101 11011 11135
rect 11621 11101 11655 11135
rect 12633 11101 12667 11135
rect 13461 11101 13495 11135
rect 16129 11101 16163 11135
rect 1869 11033 1903 11067
rect 1961 11033 1995 11067
rect 3249 11033 3283 11067
rect 3985 11033 4019 11067
rect 4261 11033 4295 11067
rect 4905 11033 4939 11067
rect 5825 11033 5859 11067
rect 7472 11033 7506 11067
rect 9220 11033 9254 11067
rect 11713 11033 11747 11067
rect 12725 11033 12759 11067
rect 13553 11033 13587 11067
rect 15884 11033 15918 11067
rect 2421 10965 2455 10999
rect 2789 10965 2823 10999
rect 5733 10965 5767 10999
rect 6561 10965 6595 10999
rect 10333 10965 10367 10999
rect 10885 10965 10919 10999
rect 12265 10965 12299 10999
rect 14657 10965 14691 10999
rect 4077 10761 4111 10795
rect 4629 10761 4663 10795
rect 4997 10761 5031 10795
rect 7757 10761 7791 10795
rect 8493 10761 8527 10795
rect 8953 10761 8987 10795
rect 9781 10761 9815 10795
rect 10241 10761 10275 10795
rect 11253 10761 11287 10795
rect 12541 10761 12575 10795
rect 13001 10761 13035 10795
rect 14933 10761 14967 10795
rect 15301 10761 15335 10795
rect 3893 10693 3927 10727
rect 8861 10693 8895 10727
rect 14841 10693 14875 10727
rect 15393 10693 15427 10727
rect 1409 10625 1443 10659
rect 1685 10625 1719 10659
rect 1961 10625 1995 10659
rect 2677 10625 2711 10659
rect 5457 10625 5491 10659
rect 6377 10625 6411 10659
rect 6644 10625 6678 10659
rect 9689 10625 9723 10659
rect 10609 10625 10643 10659
rect 12633 10625 12667 10659
rect 14206 10625 14240 10659
rect 14473 10625 14507 10659
rect 2421 10557 2455 10591
rect 4445 10557 4479 10591
rect 4537 10557 4571 10591
rect 5549 10557 5583 10591
rect 5641 10557 5675 10591
rect 9045 10557 9079 10591
rect 9965 10557 9999 10591
rect 10701 10557 10735 10591
rect 10885 10557 10919 10591
rect 11805 10557 11839 10591
rect 12449 10557 12483 10591
rect 14749 10557 14783 10591
rect 1593 10489 1627 10523
rect 2145 10489 2179 10523
rect 3801 10489 3835 10523
rect 5089 10489 5123 10523
rect 13093 10489 13127 10523
rect 1869 10421 1903 10455
rect 2237 10421 2271 10455
rect 5917 10421 5951 10455
rect 6101 10421 6135 10455
rect 9321 10421 9355 10455
rect 11621 10421 11655 10455
rect 1501 10217 1535 10251
rect 1777 10217 1811 10251
rect 3801 10217 3835 10251
rect 6561 10217 6595 10251
rect 9597 10217 9631 10251
rect 13553 10217 13587 10251
rect 15025 10217 15059 10251
rect 7389 10149 7423 10183
rect 3433 10081 3467 10115
rect 5181 10081 5215 10115
rect 6009 10081 6043 10115
rect 7941 10081 7975 10115
rect 10333 10081 10367 10115
rect 14473 10081 14507 10115
rect 1593 10013 1627 10047
rect 3249 10013 3283 10047
rect 5273 10013 5307 10047
rect 6193 10013 6227 10047
rect 6653 10013 6687 10047
rect 8953 10013 8987 10047
rect 10701 10013 10735 10047
rect 12173 10013 12207 10047
rect 12440 10013 12474 10047
rect 14197 10013 14231 10047
rect 14565 10013 14599 10047
rect 2982 9945 3016 9979
rect 4936 9945 4970 9979
rect 7757 9945 7791 9979
rect 10968 9945 11002 9979
rect 1869 9877 1903 9911
rect 3617 9877 3651 9911
rect 5549 9877 5583 9911
rect 6101 9877 6135 9911
rect 7297 9877 7331 9911
rect 7849 9877 7883 9911
rect 10057 9877 10091 9911
rect 12081 9877 12115 9911
rect 14657 9877 14691 9911
rect 4629 9673 4663 9707
rect 6929 9673 6963 9707
rect 14197 9673 14231 9707
rect 4169 9605 4203 9639
rect 4537 9605 4571 9639
rect 9812 9605 9846 9639
rect 1501 9537 1535 9571
rect 2881 9537 2915 9571
rect 3157 9537 3191 9571
rect 3525 9537 3559 9571
rect 5733 9537 5767 9571
rect 5825 9537 5859 9571
rect 8042 9537 8076 9571
rect 8309 9537 8343 9571
rect 10057 9537 10091 9571
rect 10517 9537 10551 9571
rect 11897 9537 11931 9571
rect 13553 9537 13587 9571
rect 3249 9469 3283 9503
rect 4445 9469 4479 9503
rect 5917 9469 5951 9503
rect 6377 9469 6411 9503
rect 10609 9469 10643 9503
rect 10701 9469 10735 9503
rect 11713 9469 11747 9503
rect 11805 9469 11839 9503
rect 14473 9469 14507 9503
rect 2973 9401 3007 9435
rect 5365 9401 5399 9435
rect 12265 9401 12299 9435
rect 2145 9333 2179 9367
rect 2237 9333 2271 9367
rect 4997 9333 5031 9367
rect 5181 9333 5215 9367
rect 6653 9333 6687 9367
rect 8401 9333 8435 9367
rect 8677 9333 8711 9367
rect 10149 9333 10183 9367
rect 6009 9129 6043 9163
rect 7665 9129 7699 9163
rect 8677 9129 8711 9163
rect 12173 9129 12207 9163
rect 1961 8993 1995 9027
rect 3157 8993 3191 9027
rect 4353 8993 4387 9027
rect 6101 8993 6135 9027
rect 8217 8993 8251 9027
rect 9137 8993 9171 9027
rect 11529 8993 11563 9027
rect 13277 8993 13311 9027
rect 14197 8993 14231 9027
rect 15117 8993 15151 9027
rect 1409 8925 1443 8959
rect 2145 8925 2179 8959
rect 2973 8925 3007 8959
rect 4629 8925 4663 8959
rect 6368 8925 6402 8959
rect 8125 8925 8159 8959
rect 9229 8925 9263 8959
rect 10701 8925 10735 8959
rect 11805 8925 11839 8959
rect 13461 8925 13495 8959
rect 14473 8925 14507 8959
rect 15761 8925 15795 8959
rect 2053 8857 2087 8891
rect 3065 8857 3099 8891
rect 4896 8857 4930 8891
rect 9496 8857 9530 8891
rect 11345 8857 11379 8891
rect 13001 8857 13035 8891
rect 13369 8857 13403 8891
rect 15301 8857 15335 8891
rect 1593 8789 1627 8823
rect 2513 8789 2547 8823
rect 2605 8789 2639 8823
rect 3433 8789 3467 8823
rect 3801 8789 3835 8823
rect 4169 8789 4203 8823
rect 4261 8789 4295 8823
rect 7481 8789 7515 8823
rect 8033 8789 8067 8823
rect 8493 8789 8527 8823
rect 10609 8789 10643 8823
rect 11713 8789 11747 8823
rect 13829 8789 13863 8823
rect 14381 8789 14415 8823
rect 14841 8789 14875 8823
rect 15209 8789 15243 8823
rect 15669 8789 15703 8823
rect 16405 8789 16439 8823
rect 2145 8585 2179 8619
rect 4445 8585 4479 8619
rect 4721 8585 4755 8619
rect 6377 8585 6411 8619
rect 6745 8585 6779 8619
rect 7297 8585 7331 8619
rect 8125 8585 8159 8619
rect 8493 8585 8527 8619
rect 9045 8585 9079 8619
rect 9505 8585 9539 8619
rect 9873 8585 9907 8619
rect 9965 8585 9999 8619
rect 10977 8585 11011 8619
rect 11897 8585 11931 8619
rect 12265 8585 12299 8619
rect 15577 8585 15611 8619
rect 1409 8517 1443 8551
rect 3258 8517 3292 8551
rect 8217 8517 8251 8551
rect 2053 8449 2087 8483
rect 3525 8449 3559 8483
rect 4077 8449 4111 8483
rect 4537 8449 4571 8483
rect 4813 8449 4847 8483
rect 5069 8449 5103 8483
rect 6837 8449 6871 8483
rect 7481 8449 7515 8483
rect 9137 8449 9171 8483
rect 11069 8449 11103 8483
rect 12725 8449 12759 8483
rect 12992 8449 13026 8483
rect 14197 8449 14231 8483
rect 14453 8449 14487 8483
rect 3801 8381 3835 8415
rect 3985 8381 4019 8415
rect 6929 8381 6963 8415
rect 8861 8381 8895 8415
rect 9781 8381 9815 8415
rect 11161 8381 11195 8415
rect 11713 8381 11747 8415
rect 11805 8381 11839 8415
rect 6193 8313 6227 8347
rect 10333 8313 10367 8347
rect 14105 8313 14139 8347
rect 10609 8245 10643 8279
rect 1409 8041 1443 8075
rect 2881 8041 2915 8075
rect 3801 8041 3835 8075
rect 5181 8041 5215 8075
rect 5733 8041 5767 8075
rect 7113 8041 7147 8075
rect 9229 8041 9263 8075
rect 14841 8041 14875 8075
rect 15025 7973 15059 8007
rect 3433 7905 3467 7939
rect 4353 7905 4387 7939
rect 7665 7905 7699 7939
rect 9689 7905 9723 7939
rect 9873 7905 9907 7939
rect 14197 7905 14231 7939
rect 14381 7905 14415 7939
rect 15301 7905 15335 7939
rect 2522 7837 2556 7871
rect 2789 7837 2823 7871
rect 3249 7837 3283 7871
rect 3341 7837 3375 7871
rect 4169 7837 4203 7871
rect 4905 7837 4939 7871
rect 4997 7837 5031 7871
rect 7481 7837 7515 7871
rect 7941 7837 7975 7871
rect 10425 7837 10459 7871
rect 13378 7837 13412 7871
rect 13645 7837 13679 7871
rect 15568 7837 15602 7871
rect 7021 7769 7055 7803
rect 8677 7769 8711 7803
rect 12173 7769 12207 7803
rect 14473 7769 14507 7803
rect 4261 7701 4295 7735
rect 4721 7701 4755 7735
rect 7573 7701 7607 7735
rect 8585 7701 8619 7735
rect 9137 7701 9171 7735
rect 9597 7701 9631 7735
rect 10241 7701 10275 7735
rect 12265 7701 12299 7735
rect 16681 7701 16715 7735
rect 2329 7497 2363 7531
rect 2697 7497 2731 7531
rect 3157 7497 3191 7531
rect 3525 7497 3559 7531
rect 4353 7497 4387 7531
rect 4905 7497 4939 7531
rect 5457 7497 5491 7531
rect 5825 7497 5859 7531
rect 8677 7497 8711 7531
rect 9597 7497 9631 7531
rect 9965 7497 9999 7531
rect 10425 7497 10459 7531
rect 13277 7497 13311 7531
rect 13369 7497 13403 7531
rect 13829 7497 13863 7531
rect 14289 7497 14323 7531
rect 14841 7497 14875 7531
rect 15209 7497 15243 7531
rect 2237 7429 2271 7463
rect 7564 7429 7598 7463
rect 8953 7429 8987 7463
rect 11253 7429 11287 7463
rect 15301 7429 15335 7463
rect 1409 7361 1443 7395
rect 1685 7361 1719 7395
rect 3065 7361 3099 7395
rect 3985 7361 4019 7395
rect 4997 7361 5031 7395
rect 6745 7361 6779 7395
rect 10333 7361 10367 7395
rect 12642 7361 12676 7395
rect 12909 7361 12943 7395
rect 14381 7361 14415 7395
rect 2053 7293 2087 7327
rect 2973 7293 3007 7327
rect 3709 7293 3743 7327
rect 3893 7293 3927 7327
rect 4813 7293 4847 7327
rect 5917 7293 5951 7327
rect 6009 7293 6043 7327
rect 6561 7293 6595 7327
rect 6653 7293 6687 7327
rect 7297 7293 7331 7327
rect 9413 7293 9447 7327
rect 9505 7293 9539 7327
rect 10149 7293 10183 7327
rect 11069 7293 11103 7327
rect 13093 7293 13127 7327
rect 14105 7293 14139 7327
rect 15393 7293 15427 7327
rect 1593 7225 1627 7259
rect 5365 7225 5399 7259
rect 11529 7225 11563 7259
rect 13737 7225 13771 7259
rect 14749 7225 14783 7259
rect 1869 7157 1903 7191
rect 4445 7157 4479 7191
rect 7113 7157 7147 7191
rect 8861 7157 8895 7191
rect 10793 7157 10827 7191
rect 10885 7157 10919 7191
rect 2881 6953 2915 6987
rect 6101 6953 6135 6987
rect 7573 6953 7607 6987
rect 12725 6953 12759 6987
rect 2789 6885 2823 6919
rect 8953 6885 8987 6919
rect 10977 6885 11011 6919
rect 14105 6885 14139 6919
rect 2237 6817 2271 6851
rect 3433 6817 3467 6851
rect 4261 6817 4295 6851
rect 4445 6817 4479 6851
rect 4629 6817 4663 6851
rect 5457 6817 5491 6851
rect 8217 6817 8251 6851
rect 8677 6817 8711 6851
rect 9137 6817 9171 6851
rect 9505 6817 9539 6851
rect 10701 6817 10735 6851
rect 11529 6817 11563 6851
rect 12173 6817 12207 6851
rect 12817 6817 12851 6851
rect 15485 6817 15519 6851
rect 1409 6749 1443 6783
rect 1685 6749 1719 6783
rect 2329 6749 2363 6783
rect 5273 6749 5307 6783
rect 6193 6749 6227 6783
rect 9597 6749 9631 6783
rect 12265 6749 12299 6783
rect 12357 6749 12391 6783
rect 15577 6749 15611 6783
rect 6460 6681 6494 6715
rect 8033 6681 8067 6715
rect 8493 6681 8527 6715
rect 9689 6681 9723 6715
rect 10517 6681 10551 6715
rect 15240 6681 15274 6715
rect 16221 6681 16255 6715
rect 1593 6613 1627 6647
rect 1869 6613 1903 6647
rect 2421 6613 2455 6647
rect 3249 6613 3283 6647
rect 3341 6613 3375 6647
rect 3801 6613 3835 6647
rect 4169 6613 4203 6647
rect 5641 6613 5675 6647
rect 5733 6613 5767 6647
rect 7665 6613 7699 6647
rect 8125 6613 8159 6647
rect 10057 6613 10091 6647
rect 10149 6613 10183 6647
rect 10609 6613 10643 6647
rect 11345 6613 11379 6647
rect 11437 6613 11471 6647
rect 11805 6613 11839 6647
rect 13921 6613 13955 6647
rect 1777 6409 1811 6443
rect 3341 6409 3375 6443
rect 3801 6409 3835 6443
rect 6193 6409 6227 6443
rect 7113 6409 7147 6443
rect 7205 6409 7239 6443
rect 8309 6409 8343 6443
rect 9505 6409 9539 6443
rect 11253 6409 11287 6443
rect 12265 6409 12299 6443
rect 13001 6409 13035 6443
rect 16037 6409 16071 6443
rect 17141 6409 17175 6443
rect 21373 6409 21407 6443
rect 5080 6341 5114 6375
rect 11529 6341 11563 6375
rect 12081 6341 12115 6375
rect 12909 6341 12943 6375
rect 15209 6341 15243 6375
rect 16129 6341 16163 6375
rect 1409 6273 1443 6307
rect 1869 6273 1903 6307
rect 2125 6273 2159 6307
rect 3709 6273 3743 6307
rect 4169 6273 4203 6307
rect 4445 6273 4479 6307
rect 6377 6273 6411 6307
rect 7757 6273 7791 6307
rect 8401 6273 8435 6307
rect 8861 6273 8895 6307
rect 9597 6273 9631 6307
rect 9864 6273 9898 6307
rect 13369 6273 13403 6307
rect 13636 6273 13670 6307
rect 17049 6273 17083 6307
rect 17509 6273 17543 6307
rect 18061 6273 18095 6307
rect 21281 6273 21315 6307
rect 21557 6273 21591 6307
rect 3893 6205 3927 6239
rect 4813 6205 4847 6239
rect 7389 6205 7423 6239
rect 8585 6205 8619 6239
rect 12633 6205 12667 6239
rect 15301 6205 15335 6239
rect 15393 6205 15427 6239
rect 16221 6205 16255 6239
rect 17233 6205 17267 6239
rect 3249 6137 3283 6171
rect 1593 6069 1627 6103
rect 4629 6069 4663 6103
rect 6561 6069 6595 6103
rect 6745 6069 6779 6103
rect 7573 6069 7607 6103
rect 7941 6069 7975 6103
rect 10977 6069 11011 6103
rect 11161 6069 11195 6103
rect 11713 6069 11747 6103
rect 11897 6069 11931 6103
rect 12449 6069 12483 6103
rect 13185 6069 13219 6103
rect 14749 6069 14783 6103
rect 14841 6069 14875 6103
rect 15669 6069 15703 6103
rect 16681 6069 16715 6103
rect 18705 6069 18739 6103
rect 1869 5865 1903 5899
rect 3985 5865 4019 5899
rect 4445 5865 4479 5899
rect 7113 5865 7147 5899
rect 12265 5865 12299 5899
rect 1685 5797 1719 5831
rect 8585 5797 8619 5831
rect 15577 5797 15611 5831
rect 17049 5797 17083 5831
rect 3249 5729 3283 5763
rect 4905 5729 4939 5763
rect 4997 5729 5031 5763
rect 8493 5729 8527 5763
rect 12173 5729 12207 5763
rect 12541 5729 12575 5763
rect 14565 5729 14599 5763
rect 14749 5729 14783 5763
rect 2982 5661 3016 5695
rect 3341 5661 3375 5695
rect 3801 5661 3835 5695
rect 4077 5661 4111 5695
rect 5457 5661 5491 5695
rect 7021 5661 7055 5695
rect 8769 5661 8803 5695
rect 10333 5661 10367 5695
rect 12808 5661 12842 5695
rect 14473 5661 14507 5695
rect 15669 5661 15703 5695
rect 18521 5661 18555 5695
rect 19257 5661 19291 5695
rect 1501 5593 1535 5627
rect 8226 5593 8260 5627
rect 10088 5593 10122 5627
rect 10425 5593 10459 5627
rect 15936 5593 15970 5627
rect 18276 5593 18310 5627
rect 3525 5525 3559 5559
rect 4261 5525 4295 5559
rect 4813 5525 4847 5559
rect 8953 5525 8987 5559
rect 13921 5525 13955 5559
rect 14105 5525 14139 5559
rect 14933 5525 14967 5559
rect 17141 5525 17175 5559
rect 19441 5525 19475 5559
rect 1593 5321 1627 5355
rect 3985 5321 4019 5355
rect 4353 5321 4387 5355
rect 6193 5321 6227 5355
rect 7113 5321 7147 5355
rect 7573 5321 7607 5355
rect 8033 5321 8067 5355
rect 8585 5321 8619 5355
rect 10057 5321 10091 5355
rect 10425 5321 10459 5355
rect 11345 5321 11379 5355
rect 11805 5321 11839 5355
rect 12633 5321 12667 5355
rect 14105 5321 14139 5355
rect 15209 5321 15243 5355
rect 16037 5321 16071 5355
rect 18153 5321 18187 5355
rect 2206 5253 2240 5287
rect 9698 5253 9732 5287
rect 18521 5253 18555 5287
rect 1501 5185 1535 5219
rect 3433 5185 3467 5219
rect 3709 5185 3743 5219
rect 4445 5185 4479 5219
rect 4813 5185 4847 5219
rect 5080 5185 5114 5219
rect 6653 5185 6687 5219
rect 6745 5185 6779 5219
rect 7665 5185 7699 5219
rect 8125 5185 8159 5219
rect 9965 5185 9999 5219
rect 10241 5185 10275 5219
rect 10977 5185 11011 5219
rect 11897 5185 11931 5219
rect 12357 5185 12391 5219
rect 13277 5185 13311 5219
rect 16129 5185 16163 5219
rect 16681 5185 16715 5219
rect 16937 5185 16971 5219
rect 19993 5185 20027 5219
rect 1961 5117 1995 5151
rect 4629 5117 4663 5151
rect 6561 5117 6595 5151
rect 7389 5117 7423 5151
rect 8401 5117 8435 5151
rect 10701 5117 10735 5151
rect 10885 5117 10919 5151
rect 11621 5117 11655 5151
rect 13093 5117 13127 5151
rect 13185 5117 13219 5151
rect 13921 5117 13955 5151
rect 14013 5117 14047 5151
rect 14565 5117 14599 5151
rect 15945 5117 15979 5151
rect 18613 5117 18647 5151
rect 18705 5117 18739 5151
rect 3341 5049 3375 5083
rect 3617 5049 3651 5083
rect 3893 5049 3927 5083
rect 12541 5049 12575 5083
rect 13645 5049 13679 5083
rect 14933 5049 14967 5083
rect 1777 4981 1811 5015
rect 8309 4981 8343 5015
rect 12265 4981 12299 5015
rect 14473 4981 14507 5015
rect 14841 4981 14875 5015
rect 16497 4981 16531 5015
rect 18061 4981 18095 5015
rect 20177 4981 20211 5015
rect 1961 4777 1995 4811
rect 2789 4777 2823 4811
rect 3617 4777 3651 4811
rect 7389 4777 7423 4811
rect 7573 4777 7607 4811
rect 9597 4777 9631 4811
rect 11437 4777 11471 4811
rect 11529 4777 11563 4811
rect 13369 4777 13403 4811
rect 14105 4777 14139 4811
rect 1685 4709 1719 4743
rect 3801 4709 3835 4743
rect 13461 4709 13495 4743
rect 15485 4709 15519 4743
rect 17509 4709 17543 4743
rect 2237 4641 2271 4675
rect 2973 4641 3007 4675
rect 4445 4641 4479 4675
rect 6929 4641 6963 4675
rect 8217 4641 8251 4675
rect 9965 4641 9999 4675
rect 10885 4641 10919 4675
rect 10977 4641 11011 4675
rect 12081 4641 12115 4675
rect 12725 4641 12759 4675
rect 13829 4641 13863 4675
rect 14749 4641 14783 4675
rect 15669 4641 15703 4675
rect 16589 4641 16623 4675
rect 16773 4641 16807 4675
rect 17969 4641 18003 4675
rect 1501 4573 1535 4607
rect 1777 4573 1811 4607
rect 2421 4573 2455 4607
rect 6193 4573 6227 4607
rect 6653 4573 6687 4607
rect 7113 4573 7147 4607
rect 7941 4573 7975 4607
rect 8953 4573 8987 4607
rect 10241 4573 10275 4607
rect 11897 4573 11931 4607
rect 13645 4573 13679 4607
rect 16865 4573 16899 4607
rect 17325 4573 17359 4607
rect 2329 4505 2363 4539
rect 4169 4505 4203 4539
rect 4629 4505 4663 4539
rect 5926 4505 5960 4539
rect 8493 4505 8527 4539
rect 8677 4505 8711 4539
rect 11069 4505 11103 4539
rect 12909 4505 12943 4539
rect 13001 4505 13035 4539
rect 15117 4505 15151 4539
rect 17785 4505 17819 4539
rect 3157 4437 3191 4471
rect 3249 4437 3283 4471
rect 4261 4437 4295 4471
rect 4813 4437 4847 4471
rect 6285 4437 6319 4471
rect 6745 4437 6779 4471
rect 7297 4437 7331 4471
rect 8033 4437 8067 4471
rect 9689 4437 9723 4471
rect 10149 4437 10183 4471
rect 10609 4437 10643 4471
rect 11989 4437 12023 4471
rect 12449 4437 12483 4471
rect 14473 4437 14507 4471
rect 14565 4437 14599 4471
rect 14933 4437 14967 4471
rect 15393 4437 15427 4471
rect 15853 4437 15887 4471
rect 17233 4437 17267 4471
rect 2421 4233 2455 4267
rect 2513 4233 2547 4267
rect 2973 4233 3007 4267
rect 3801 4233 3835 4267
rect 7665 4233 7699 4267
rect 10885 4233 10919 4267
rect 12173 4233 12207 4267
rect 15393 4233 15427 4267
rect 3341 4165 3375 4199
rect 6193 4165 6227 4199
rect 6745 4165 6779 4199
rect 7573 4165 7607 4199
rect 10977 4165 11011 4199
rect 12081 4165 12115 4199
rect 2053 4097 2087 4131
rect 4169 4097 4203 4131
rect 5181 4097 5215 4131
rect 5733 4097 5767 4131
rect 8493 4097 8527 4131
rect 9321 4097 9355 4131
rect 10057 4097 10091 4131
rect 10149 4097 10183 4131
rect 12633 4097 12667 4131
rect 13553 4097 13587 4131
rect 14280 4097 14314 4131
rect 2329 4029 2363 4063
rect 3433 4029 3467 4063
rect 3525 4029 3559 4063
rect 4261 4029 4295 4063
rect 4353 4029 4387 4063
rect 5273 4029 5307 4063
rect 5457 4029 5491 4063
rect 6837 4029 6871 4063
rect 6929 4029 6963 4063
rect 7481 4029 7515 4063
rect 8585 4029 8619 4063
rect 8769 4029 8803 4063
rect 9045 4029 9079 4063
rect 9229 4029 9263 4063
rect 9873 4029 9907 4063
rect 10701 4029 10735 4063
rect 11529 4029 11563 4063
rect 11989 4029 12023 4063
rect 14013 4029 14047 4063
rect 15853 4029 15887 4063
rect 6377 3961 6411 3995
rect 9689 3961 9723 3995
rect 12541 3961 12575 3995
rect 15485 3961 15519 3995
rect 16405 3961 16439 3995
rect 1409 3893 1443 3927
rect 2881 3893 2915 3927
rect 4629 3893 4663 3927
rect 4813 3893 4847 3927
rect 5917 3893 5951 3927
rect 8033 3893 8067 3927
rect 8125 3893 8159 3927
rect 10517 3893 10551 3927
rect 11345 3893 11379 3927
rect 13277 3893 13311 3927
rect 13369 3893 13403 3927
rect 13645 3893 13679 3927
rect 13829 3893 13863 3927
rect 15669 3893 15703 3927
rect 16037 3893 16071 3927
rect 16313 3893 16347 3927
rect 16681 3893 16715 3927
rect 1409 3689 1443 3723
rect 1777 3689 1811 3723
rect 3341 3689 3375 3723
rect 3617 3689 3651 3723
rect 4629 3689 4663 3723
rect 6377 3689 6411 3723
rect 8953 3689 8987 3723
rect 10609 3689 10643 3723
rect 10793 3689 10827 3723
rect 13921 3689 13955 3723
rect 14289 3689 14323 3723
rect 15117 3689 15151 3723
rect 16221 3689 16255 3723
rect 17049 3689 17083 3723
rect 17417 3689 17451 3723
rect 21373 3689 21407 3723
rect 4721 3621 4755 3655
rect 12449 3621 12483 3655
rect 15853 3621 15887 3655
rect 16037 3621 16071 3655
rect 1961 3553 1995 3587
rect 4077 3553 4111 3587
rect 6745 3553 6779 3587
rect 14841 3553 14875 3587
rect 16589 3553 16623 3587
rect 17969 3553 18003 3587
rect 2228 3485 2262 3519
rect 3433 3485 3467 3519
rect 4261 3485 4295 3519
rect 6101 3485 6135 3519
rect 7389 3485 7423 3519
rect 7656 3485 7690 3519
rect 9137 3485 9171 3519
rect 9229 3485 9263 3519
rect 10883 3485 10917 3519
rect 11069 3485 11103 3519
rect 12541 3485 12575 3519
rect 15393 3485 15427 3519
rect 18153 3485 18187 3519
rect 21281 3485 21315 3519
rect 21557 3485 21591 3519
rect 1685 3417 1719 3451
rect 5834 3417 5868 3451
rect 6285 3417 6319 3451
rect 9496 3417 9530 3451
rect 11314 3417 11348 3451
rect 12808 3417 12842 3451
rect 14749 3417 14783 3451
rect 15669 3417 15703 3451
rect 4169 3349 4203 3383
rect 6837 3349 6871 3383
rect 6929 3349 6963 3383
rect 7297 3349 7331 3383
rect 8769 3349 8803 3383
rect 14197 3349 14231 3383
rect 14657 3349 14691 3383
rect 15577 3349 15611 3383
rect 16405 3349 16439 3383
rect 16865 3349 16899 3383
rect 18337 3349 18371 3383
rect 1685 3145 1719 3179
rect 4629 3145 4663 3179
rect 5365 3145 5399 3179
rect 5457 3145 5491 3179
rect 5917 3145 5951 3179
rect 6837 3145 6871 3179
rect 7389 3145 7423 3179
rect 8309 3145 8343 3179
rect 8677 3145 8711 3179
rect 9781 3145 9815 3179
rect 10149 3145 10183 3179
rect 10609 3145 10643 3179
rect 14565 3145 14599 3179
rect 14841 3145 14875 3179
rect 14933 3145 14967 3179
rect 17969 3145 18003 3179
rect 18337 3145 18371 3179
rect 18889 3145 18923 3179
rect 19257 3145 19291 3179
rect 20269 3145 20303 3179
rect 3494 3077 3528 3111
rect 6377 3077 6411 3111
rect 6929 3077 6963 3111
rect 7481 3077 7515 3111
rect 8217 3077 8251 3111
rect 8861 3077 8895 3111
rect 10241 3077 10275 3111
rect 11621 3077 11655 3111
rect 11805 3077 11839 3111
rect 1409 3009 1443 3043
rect 2809 3009 2843 3043
rect 3065 3009 3099 3043
rect 4721 3009 4755 3043
rect 5825 3009 5859 3043
rect 6561 3009 6595 3043
rect 9321 3009 9355 3043
rect 10977 3009 11011 3043
rect 11069 3009 11103 3043
rect 12449 3009 12483 3043
rect 12909 3009 12943 3043
rect 13185 3009 13219 3043
rect 13461 3009 13495 3043
rect 13921 3009 13955 3043
rect 14657 3009 14691 3043
rect 15117 3009 15151 3043
rect 15393 3009 15427 3043
rect 15485 3009 15519 3043
rect 15945 2993 15979 3027
rect 16037 3009 16071 3043
rect 16313 3009 16347 3043
rect 16865 3009 16899 3043
rect 16957 3009 16991 3043
rect 17233 3009 17267 3043
rect 17509 3009 17543 3043
rect 17785 3009 17819 3043
rect 18061 3009 18095 3043
rect 18613 3009 18647 3043
rect 19073 3009 19107 3043
rect 19349 3009 19383 3043
rect 19533 3009 19567 3043
rect 19809 3009 19843 3043
rect 20453 3009 20487 3043
rect 20913 3009 20947 3043
rect 21281 3009 21315 3043
rect 3249 2941 3283 2975
rect 6009 2941 6043 2975
rect 7297 2941 7331 2975
rect 8125 2941 8159 2975
rect 9045 2941 9079 2975
rect 9229 2941 9263 2975
rect 10425 2941 10459 2975
rect 11253 2941 11287 2975
rect 12265 2941 12299 2975
rect 12357 2941 12391 2975
rect 13737 2941 13771 2975
rect 9689 2873 9723 2907
rect 12817 2873 12851 2907
rect 13645 2873 13679 2907
rect 16497 2873 16531 2907
rect 17417 2873 17451 2907
rect 18797 2873 18831 2907
rect 19717 2873 19751 2907
rect 21097 2873 21131 2907
rect 1593 2805 1627 2839
rect 7849 2805 7883 2839
rect 11897 2805 11931 2839
rect 13093 2805 13127 2839
rect 13369 2805 13403 2839
rect 15209 2805 15243 2839
rect 15669 2805 15703 2839
rect 15761 2805 15795 2839
rect 16221 2805 16255 2839
rect 16681 2805 16715 2839
rect 17141 2805 17175 2839
rect 17693 2805 17727 2839
rect 18245 2805 18279 2839
rect 20637 2805 20671 2839
rect 21465 2805 21499 2839
rect 3525 2601 3559 2635
rect 4629 2601 4663 2635
rect 6469 2601 6503 2635
rect 6837 2601 6871 2635
rect 7849 2601 7883 2635
rect 9045 2601 9079 2635
rect 9413 2601 9447 2635
rect 10609 2601 10643 2635
rect 4905 2533 4939 2567
rect 14289 2533 14323 2567
rect 2237 2465 2271 2499
rect 2881 2465 2915 2499
rect 3985 2465 4019 2499
rect 4169 2465 4203 2499
rect 5549 2465 5583 2499
rect 7205 2465 7239 2499
rect 8493 2465 8527 2499
rect 10241 2465 10275 2499
rect 11069 2465 11103 2499
rect 11161 2465 11195 2499
rect 12081 2465 12115 2499
rect 1961 2397 1995 2431
rect 3157 2397 3191 2431
rect 4721 2397 4755 2431
rect 5825 2397 5859 2431
rect 7389 2397 7423 2431
rect 7481 2397 7515 2431
rect 8769 2397 8803 2431
rect 10517 2397 10551 2431
rect 10977 2397 11011 2431
rect 12311 2397 12345 2431
rect 13001 2397 13035 2431
rect 13277 2397 13311 2431
rect 13369 2397 13403 2431
rect 13737 2397 13771 2431
rect 14105 2397 14139 2431
rect 14473 2397 14507 2431
rect 15117 2397 15151 2431
rect 15577 2397 15611 2431
rect 15761 2397 15795 2431
rect 16221 2397 16255 2431
rect 16681 2397 16715 2431
rect 17141 2397 17175 2431
rect 17601 2397 17635 2431
rect 18061 2397 18095 2431
rect 18521 2397 18555 2431
rect 19257 2397 19291 2431
rect 19625 2397 19659 2431
rect 19993 2397 20027 2431
rect 20453 2397 20487 2431
rect 20913 2397 20947 2431
rect 21281 2397 21315 2431
rect 3433 2329 3467 2363
rect 4261 2329 4295 2363
rect 6101 2329 6135 2363
rect 6561 2329 6595 2363
rect 6929 2329 6963 2363
rect 9137 2329 9171 2363
rect 9505 2329 9539 2363
rect 6009 2261 6043 2295
rect 13553 2261 13587 2295
rect 13921 2261 13955 2295
rect 14657 2261 14691 2295
rect 14933 2261 14967 2295
rect 15393 2261 15427 2295
rect 15945 2261 15979 2295
rect 16405 2261 16439 2295
rect 16865 2261 16899 2295
rect 17325 2261 17359 2295
rect 17785 2261 17819 2295
rect 18245 2261 18279 2295
rect 18705 2261 18739 2295
rect 19441 2261 19475 2295
rect 19809 2261 19843 2295
rect 20177 2261 20211 2295
rect 20637 2261 20671 2295
rect 21097 2261 21131 2295
rect 21465 2261 21499 2295
<< metal1 >>
rect 10226 20748 10232 20800
rect 10284 20788 10290 20800
rect 11238 20788 11244 20800
rect 10284 20760 11244 20788
rect 10284 20748 10290 20760
rect 11238 20748 11244 20760
rect 11296 20748 11302 20800
rect 1104 20698 21896 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21896 20698
rect 1104 20624 21896 20646
rect 3050 20544 3056 20596
rect 3108 20584 3114 20596
rect 4614 20584 4620 20596
rect 3108 20556 4620 20584
rect 3108 20544 3114 20556
rect 4614 20544 4620 20556
rect 4672 20544 4678 20596
rect 4890 20544 4896 20596
rect 4948 20584 4954 20596
rect 6638 20584 6644 20596
rect 4948 20556 6644 20584
rect 4948 20544 4954 20556
rect 6638 20544 6644 20556
rect 6696 20544 6702 20596
rect 7558 20544 7564 20596
rect 7616 20584 7622 20596
rect 9306 20584 9312 20596
rect 7616 20556 9312 20584
rect 7616 20544 7622 20556
rect 9306 20544 9312 20556
rect 9364 20544 9370 20596
rect 10226 20584 10232 20596
rect 9508 20556 10232 20584
rect 3237 20519 3295 20525
rect 3237 20485 3249 20519
rect 3283 20516 3295 20519
rect 5166 20516 5172 20528
rect 3283 20488 5172 20516
rect 3283 20485 3295 20488
rect 3237 20479 3295 20485
rect 5166 20476 5172 20488
rect 5224 20476 5230 20528
rect 8021 20519 8079 20525
rect 8021 20485 8033 20519
rect 8067 20516 8079 20519
rect 9508 20516 9536 20556
rect 10226 20544 10232 20556
rect 10284 20544 10290 20596
rect 10321 20587 10379 20593
rect 10321 20553 10333 20587
rect 10367 20584 10379 20587
rect 12894 20584 12900 20596
rect 10367 20556 12900 20584
rect 10367 20553 10379 20556
rect 10321 20547 10379 20553
rect 12894 20544 12900 20556
rect 12952 20544 12958 20596
rect 13078 20544 13084 20596
rect 13136 20584 13142 20596
rect 13265 20587 13323 20593
rect 13265 20584 13277 20587
rect 13136 20556 13277 20584
rect 13136 20544 13142 20556
rect 13265 20553 13277 20556
rect 13311 20553 13323 20587
rect 13265 20547 13323 20553
rect 13538 20544 13544 20596
rect 13596 20584 13602 20596
rect 13817 20587 13875 20593
rect 13817 20584 13829 20587
rect 13596 20556 13829 20584
rect 13596 20544 13602 20556
rect 13817 20553 13829 20556
rect 13863 20553 13875 20587
rect 13817 20547 13875 20553
rect 13998 20544 14004 20596
rect 14056 20584 14062 20596
rect 14277 20587 14335 20593
rect 14277 20584 14289 20587
rect 14056 20556 14289 20584
rect 14056 20544 14062 20556
rect 14277 20553 14289 20556
rect 14323 20553 14335 20587
rect 14277 20547 14335 20553
rect 14458 20544 14464 20596
rect 14516 20584 14522 20596
rect 14737 20587 14795 20593
rect 14737 20584 14749 20587
rect 14516 20556 14749 20584
rect 14516 20544 14522 20556
rect 14737 20553 14749 20556
rect 14783 20553 14795 20587
rect 15194 20584 15200 20596
rect 15155 20556 15200 20584
rect 14737 20547 14795 20553
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 15378 20544 15384 20596
rect 15436 20584 15442 20596
rect 15657 20587 15715 20593
rect 15657 20584 15669 20587
rect 15436 20556 15669 20584
rect 15436 20544 15442 20556
rect 15657 20553 15669 20556
rect 15703 20553 15715 20587
rect 15657 20547 15715 20553
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 16117 20587 16175 20593
rect 16117 20584 16129 20587
rect 15896 20556 16129 20584
rect 15896 20544 15902 20556
rect 16117 20553 16129 20556
rect 16163 20553 16175 20587
rect 16117 20547 16175 20553
rect 16298 20544 16304 20596
rect 16356 20584 16362 20596
rect 16853 20587 16911 20593
rect 16853 20584 16865 20587
rect 16356 20556 16865 20584
rect 16356 20544 16362 20556
rect 16853 20553 16865 20556
rect 16899 20553 16911 20587
rect 16853 20547 16911 20553
rect 17218 20544 17224 20596
rect 17276 20584 17282 20596
rect 17589 20587 17647 20593
rect 17589 20584 17601 20587
rect 17276 20556 17601 20584
rect 17276 20544 17282 20556
rect 17589 20553 17601 20556
rect 17635 20553 17647 20587
rect 17954 20584 17960 20596
rect 17915 20556 17960 20584
rect 17589 20547 17647 20553
rect 17954 20544 17960 20556
rect 18012 20544 18018 20596
rect 18138 20544 18144 20596
rect 18196 20584 18202 20596
rect 18417 20587 18475 20593
rect 18417 20584 18429 20587
rect 18196 20556 18429 20584
rect 18196 20544 18202 20556
rect 18417 20553 18429 20556
rect 18463 20553 18475 20587
rect 18417 20547 18475 20553
rect 18598 20544 18604 20596
rect 18656 20584 18662 20596
rect 18877 20587 18935 20593
rect 18877 20584 18889 20587
rect 18656 20556 18889 20584
rect 18656 20544 18662 20556
rect 18877 20553 18889 20556
rect 18923 20553 18935 20587
rect 18877 20547 18935 20553
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 19429 20587 19487 20593
rect 19429 20584 19441 20587
rect 19392 20556 19441 20584
rect 19392 20544 19398 20556
rect 19429 20553 19441 20556
rect 19475 20553 19487 20587
rect 19429 20547 19487 20553
rect 19518 20544 19524 20596
rect 19576 20584 19582 20596
rect 19797 20587 19855 20593
rect 19797 20584 19809 20587
rect 19576 20556 19809 20584
rect 19576 20544 19582 20556
rect 19797 20553 19809 20556
rect 19843 20553 19855 20587
rect 19797 20547 19855 20553
rect 19978 20544 19984 20596
rect 20036 20584 20042 20596
rect 20257 20587 20315 20593
rect 20257 20584 20269 20587
rect 20036 20556 20269 20584
rect 20036 20544 20042 20556
rect 20257 20553 20269 20556
rect 20303 20553 20315 20587
rect 20257 20547 20315 20553
rect 20438 20544 20444 20596
rect 20496 20584 20502 20596
rect 20717 20587 20775 20593
rect 20717 20584 20729 20587
rect 20496 20556 20729 20584
rect 20496 20544 20502 20556
rect 20717 20553 20729 20556
rect 20763 20553 20775 20587
rect 20717 20547 20775 20553
rect 20898 20544 20904 20596
rect 20956 20584 20962 20596
rect 21177 20587 21235 20593
rect 21177 20584 21189 20587
rect 20956 20556 21189 20584
rect 20956 20544 20962 20556
rect 21177 20553 21189 20556
rect 21223 20553 21235 20587
rect 21177 20547 21235 20553
rect 8067 20488 9536 20516
rect 11149 20519 11207 20525
rect 8067 20485 8079 20488
rect 8021 20479 8079 20485
rect 11149 20485 11161 20519
rect 11195 20516 11207 20519
rect 11238 20516 11244 20528
rect 11195 20488 11244 20516
rect 11195 20485 11207 20488
rect 11149 20479 11207 20485
rect 11238 20476 11244 20488
rect 11296 20476 11302 20528
rect 16393 20519 16451 20525
rect 16393 20516 16405 20519
rect 11440 20488 16405 20516
rect 2038 20448 2044 20460
rect 1999 20420 2044 20448
rect 2038 20408 2044 20420
rect 2096 20408 2102 20460
rect 2130 20408 2136 20460
rect 2188 20448 2194 20460
rect 2961 20451 3019 20457
rect 2961 20448 2973 20451
rect 2188 20420 2973 20448
rect 2188 20408 2194 20420
rect 2961 20417 2973 20420
rect 3007 20417 3019 20451
rect 3510 20448 3516 20460
rect 3471 20420 3516 20448
rect 2961 20411 3019 20417
rect 3510 20408 3516 20420
rect 3568 20408 3574 20460
rect 4341 20451 4399 20457
rect 4341 20417 4353 20451
rect 4387 20448 4399 20451
rect 4387 20420 4844 20448
rect 4387 20417 4399 20420
rect 4341 20411 4399 20417
rect 2682 20380 2688 20392
rect 2643 20352 2688 20380
rect 2682 20340 2688 20352
rect 2740 20340 2746 20392
rect 4154 20380 4160 20392
rect 3252 20352 4160 20380
rect 1397 20315 1455 20321
rect 1397 20281 1409 20315
rect 1443 20312 1455 20315
rect 3252 20312 3280 20352
rect 4154 20340 4160 20352
rect 4212 20340 4218 20392
rect 4614 20380 4620 20392
rect 4575 20352 4620 20380
rect 4614 20340 4620 20352
rect 4672 20340 4678 20392
rect 4816 20380 4844 20420
rect 4890 20408 4896 20460
rect 4948 20448 4954 20460
rect 5442 20448 5448 20460
rect 4948 20420 4993 20448
rect 5403 20420 5448 20448
rect 4948 20408 4954 20420
rect 5442 20408 5448 20420
rect 5500 20408 5506 20460
rect 5997 20451 6055 20457
rect 5997 20417 6009 20451
rect 6043 20417 6055 20451
rect 6362 20448 6368 20460
rect 6323 20420 6368 20448
rect 5997 20411 6055 20417
rect 5166 20380 5172 20392
rect 4816 20352 5172 20380
rect 5166 20340 5172 20352
rect 5224 20340 5230 20392
rect 5534 20380 5540 20392
rect 5495 20352 5540 20380
rect 5534 20340 5540 20352
rect 5592 20340 5598 20392
rect 5626 20340 5632 20392
rect 5684 20380 5690 20392
rect 6012 20380 6040 20411
rect 6362 20408 6368 20420
rect 6420 20408 6426 20460
rect 7098 20408 7104 20460
rect 7156 20448 7162 20460
rect 7193 20451 7251 20457
rect 7193 20448 7205 20451
rect 7156 20420 7205 20448
rect 7156 20408 7162 20420
rect 7193 20417 7205 20420
rect 7239 20417 7251 20451
rect 7193 20411 7251 20417
rect 8757 20451 8815 20457
rect 8757 20417 8769 20451
rect 8803 20448 8815 20451
rect 9398 20448 9404 20460
rect 8803 20420 9404 20448
rect 8803 20417 8815 20420
rect 8757 20411 8815 20417
rect 9398 20408 9404 20420
rect 9456 20408 9462 20460
rect 10134 20408 10140 20460
rect 10192 20448 10198 20460
rect 10229 20451 10287 20457
rect 10229 20448 10241 20451
rect 10192 20420 10241 20448
rect 10192 20408 10198 20420
rect 10229 20417 10241 20420
rect 10275 20417 10287 20451
rect 10229 20411 10287 20417
rect 10873 20451 10931 20457
rect 10873 20417 10885 20451
rect 10919 20417 10931 20451
rect 11440 20448 11468 20488
rect 16393 20485 16405 20488
rect 16439 20485 16451 20519
rect 16393 20479 16451 20485
rect 10873 20411 10931 20417
rect 10980 20420 11468 20448
rect 11517 20451 11575 20457
rect 7558 20380 7564 20392
rect 5684 20352 5729 20380
rect 6012 20352 7564 20380
rect 5684 20340 5690 20352
rect 7558 20340 7564 20352
rect 7616 20340 7622 20392
rect 8294 20340 8300 20392
rect 8352 20380 8358 20392
rect 8941 20383 8999 20389
rect 8941 20380 8953 20383
rect 8352 20352 8953 20380
rect 8352 20340 8358 20352
rect 8941 20349 8953 20352
rect 8987 20349 8999 20383
rect 8941 20343 8999 20349
rect 9217 20383 9275 20389
rect 9217 20349 9229 20383
rect 9263 20349 9275 20383
rect 9217 20343 9275 20349
rect 5077 20315 5135 20321
rect 5077 20312 5089 20315
rect 1443 20284 3280 20312
rect 3344 20284 5089 20312
rect 1443 20281 1455 20284
rect 1397 20275 1455 20281
rect 1302 20204 1308 20256
rect 1360 20244 1366 20256
rect 3344 20244 3372 20284
rect 5077 20281 5089 20284
rect 5123 20281 5135 20315
rect 5077 20275 5135 20281
rect 5902 20272 5908 20324
rect 5960 20312 5966 20324
rect 7009 20315 7067 20321
rect 7009 20312 7021 20315
rect 5960 20284 7021 20312
rect 5960 20272 5966 20284
rect 7009 20281 7021 20284
rect 7055 20281 7067 20315
rect 7009 20275 7067 20281
rect 8662 20272 8668 20324
rect 8720 20312 8726 20324
rect 9232 20312 9260 20343
rect 9306 20340 9312 20392
rect 9364 20380 9370 20392
rect 10042 20380 10048 20392
rect 9364 20352 10048 20380
rect 9364 20340 9370 20352
rect 10042 20340 10048 20352
rect 10100 20340 10106 20392
rect 10410 20340 10416 20392
rect 10468 20380 10474 20392
rect 10468 20352 10513 20380
rect 10468 20340 10474 20352
rect 10594 20340 10600 20392
rect 10652 20380 10658 20392
rect 10689 20383 10747 20389
rect 10689 20380 10701 20383
rect 10652 20352 10701 20380
rect 10652 20340 10658 20352
rect 10689 20349 10701 20352
rect 10735 20349 10747 20383
rect 10689 20343 10747 20349
rect 10888 20324 10916 20411
rect 8720 20284 9260 20312
rect 8720 20272 8726 20284
rect 9674 20272 9680 20324
rect 9732 20312 9738 20324
rect 10870 20312 10876 20324
rect 9732 20284 10876 20312
rect 9732 20272 9738 20284
rect 10870 20272 10876 20284
rect 10928 20272 10934 20324
rect 1360 20216 3372 20244
rect 3421 20247 3479 20253
rect 1360 20204 1366 20216
rect 3421 20213 3433 20247
rect 3467 20244 3479 20247
rect 3970 20244 3976 20256
rect 3467 20216 3976 20244
rect 3467 20213 3479 20216
rect 3421 20207 3479 20213
rect 3970 20204 3976 20216
rect 4028 20204 4034 20256
rect 4798 20244 4804 20256
rect 4759 20216 4804 20244
rect 4798 20204 4804 20216
rect 4856 20204 4862 20256
rect 5810 20204 5816 20256
rect 5868 20244 5874 20256
rect 6089 20247 6147 20253
rect 6089 20244 6101 20247
rect 5868 20216 6101 20244
rect 5868 20204 5874 20216
rect 6089 20213 6101 20216
rect 6135 20213 6147 20247
rect 7834 20244 7840 20256
rect 7795 20216 7840 20244
rect 6089 20207 6147 20213
rect 7834 20204 7840 20216
rect 7892 20204 7898 20256
rect 8113 20247 8171 20253
rect 8113 20213 8125 20247
rect 8159 20244 8171 20247
rect 9306 20244 9312 20256
rect 8159 20216 9312 20244
rect 8159 20213 8171 20216
rect 8113 20207 8171 20213
rect 9306 20204 9312 20216
rect 9364 20204 9370 20256
rect 9398 20204 9404 20256
rect 9456 20244 9462 20256
rect 9861 20247 9919 20253
rect 9861 20244 9873 20247
rect 9456 20216 9873 20244
rect 9456 20204 9462 20216
rect 9861 20213 9873 20216
rect 9907 20213 9919 20247
rect 9861 20207 9919 20213
rect 10042 20204 10048 20256
rect 10100 20244 10106 20256
rect 10980 20244 11008 20420
rect 11517 20417 11529 20451
rect 11563 20417 11575 20451
rect 11517 20411 11575 20417
rect 11146 20340 11152 20392
rect 11204 20380 11210 20392
rect 11532 20380 11560 20411
rect 12434 20408 12440 20460
rect 12492 20448 12498 20460
rect 13081 20451 13139 20457
rect 13081 20448 13093 20451
rect 12492 20420 13093 20448
rect 12492 20408 12498 20420
rect 13081 20417 13093 20420
rect 13127 20448 13139 20451
rect 13262 20448 13268 20460
rect 13127 20420 13268 20448
rect 13127 20417 13139 20420
rect 13081 20411 13139 20417
rect 13262 20408 13268 20420
rect 13320 20408 13326 20460
rect 13449 20451 13507 20457
rect 13449 20417 13461 20451
rect 13495 20448 13507 20451
rect 13538 20448 13544 20460
rect 13495 20420 13544 20448
rect 13495 20417 13507 20420
rect 13449 20411 13507 20417
rect 13538 20408 13544 20420
rect 13596 20408 13602 20460
rect 13630 20408 13636 20460
rect 13688 20448 13694 20460
rect 13688 20420 13733 20448
rect 13688 20408 13694 20420
rect 13814 20408 13820 20460
rect 13872 20448 13878 20460
rect 14093 20451 14151 20457
rect 14093 20448 14105 20451
rect 13872 20420 14105 20448
rect 13872 20408 13878 20420
rect 14093 20417 14105 20420
rect 14139 20417 14151 20451
rect 14093 20411 14151 20417
rect 14274 20408 14280 20460
rect 14332 20448 14338 20460
rect 14553 20451 14611 20457
rect 14553 20448 14565 20451
rect 14332 20420 14565 20448
rect 14332 20408 14338 20420
rect 14553 20417 14565 20420
rect 14599 20417 14611 20451
rect 14553 20411 14611 20417
rect 14826 20408 14832 20460
rect 14884 20448 14890 20460
rect 15013 20451 15071 20457
rect 15013 20448 15025 20451
rect 14884 20420 15025 20448
rect 14884 20408 14890 20420
rect 15013 20417 15025 20420
rect 15059 20417 15071 20451
rect 15013 20411 15071 20417
rect 15102 20408 15108 20460
rect 15160 20448 15166 20460
rect 15473 20451 15531 20457
rect 15473 20448 15485 20451
rect 15160 20420 15485 20448
rect 15160 20408 15166 20420
rect 15473 20417 15485 20420
rect 15519 20417 15531 20451
rect 15930 20448 15936 20460
rect 15891 20420 15936 20448
rect 15473 20411 15531 20417
rect 15930 20408 15936 20420
rect 15988 20408 15994 20460
rect 16666 20448 16672 20460
rect 16627 20420 16672 20448
rect 16666 20408 16672 20420
rect 16724 20408 16730 20460
rect 17034 20448 17040 20460
rect 16995 20420 17040 20448
rect 17034 20408 17040 20420
rect 17092 20408 17098 20460
rect 17126 20408 17132 20460
rect 17184 20448 17190 20460
rect 17405 20451 17463 20457
rect 17405 20448 17417 20451
rect 17184 20420 17417 20448
rect 17184 20408 17190 20420
rect 17405 20417 17417 20420
rect 17451 20417 17463 20451
rect 17405 20411 17463 20417
rect 17678 20408 17684 20460
rect 17736 20448 17742 20460
rect 17773 20451 17831 20457
rect 17773 20448 17785 20451
rect 17736 20420 17785 20448
rect 17736 20408 17742 20420
rect 17773 20417 17785 20420
rect 17819 20417 17831 20451
rect 17773 20411 17831 20417
rect 17954 20408 17960 20460
rect 18012 20448 18018 20460
rect 18233 20451 18291 20457
rect 18233 20448 18245 20451
rect 18012 20420 18245 20448
rect 18012 20408 18018 20420
rect 18233 20417 18245 20420
rect 18279 20417 18291 20451
rect 18233 20411 18291 20417
rect 18322 20408 18328 20460
rect 18380 20448 18386 20460
rect 18693 20451 18751 20457
rect 18693 20448 18705 20451
rect 18380 20420 18705 20448
rect 18380 20408 18386 20420
rect 18693 20417 18705 20420
rect 18739 20417 18751 20451
rect 18693 20411 18751 20417
rect 18782 20408 18788 20460
rect 18840 20448 18846 20460
rect 19245 20451 19303 20457
rect 19245 20448 19257 20451
rect 18840 20420 19257 20448
rect 18840 20408 18846 20420
rect 19245 20417 19257 20420
rect 19291 20417 19303 20451
rect 19245 20411 19303 20417
rect 19613 20451 19671 20457
rect 19613 20417 19625 20451
rect 19659 20417 19671 20451
rect 19613 20411 19671 20417
rect 11204 20352 11560 20380
rect 12805 20383 12863 20389
rect 11204 20340 11210 20352
rect 12805 20349 12817 20383
rect 12851 20349 12863 20383
rect 19628 20380 19656 20411
rect 19702 20408 19708 20460
rect 19760 20448 19766 20460
rect 20073 20451 20131 20457
rect 20073 20448 20085 20451
rect 19760 20420 20085 20448
rect 19760 20408 19766 20420
rect 20073 20417 20085 20420
rect 20119 20417 20131 20451
rect 20530 20448 20536 20460
rect 20491 20420 20536 20448
rect 20073 20411 20131 20417
rect 20530 20408 20536 20420
rect 20588 20408 20594 20460
rect 20993 20451 21051 20457
rect 20993 20417 21005 20451
rect 21039 20417 21051 20451
rect 20993 20411 21051 20417
rect 12805 20343 12863 20349
rect 13464 20352 19656 20380
rect 11054 20272 11060 20324
rect 11112 20312 11118 20324
rect 12161 20315 12219 20321
rect 12161 20312 12173 20315
rect 11112 20284 12173 20312
rect 11112 20272 11118 20284
rect 12161 20281 12173 20284
rect 12207 20281 12219 20315
rect 12161 20275 12219 20281
rect 12434 20272 12440 20324
rect 12492 20312 12498 20324
rect 12820 20312 12848 20343
rect 13464 20324 13492 20352
rect 12492 20284 12848 20312
rect 12492 20272 12498 20284
rect 13446 20272 13452 20324
rect 13504 20272 13510 20324
rect 14366 20272 14372 20324
rect 14424 20312 14430 20324
rect 14424 20284 16574 20312
rect 14424 20272 14430 20284
rect 10100 20216 11008 20244
rect 11241 20247 11299 20253
rect 10100 20204 10106 20216
rect 11241 20213 11253 20247
rect 11287 20244 11299 20247
rect 11882 20244 11888 20256
rect 11287 20216 11888 20244
rect 11287 20213 11299 20216
rect 11241 20207 11299 20213
rect 11882 20204 11888 20216
rect 11940 20204 11946 20256
rect 16546 20244 16574 20284
rect 16942 20272 16948 20324
rect 17000 20312 17006 20324
rect 17221 20315 17279 20321
rect 17221 20312 17233 20315
rect 17000 20284 17233 20312
rect 17000 20272 17006 20284
rect 17221 20281 17233 20284
rect 17267 20281 17279 20315
rect 17221 20275 17279 20281
rect 18414 20272 18420 20324
rect 18472 20312 18478 20324
rect 21008 20312 21036 20411
rect 21174 20408 21180 20460
rect 21232 20448 21238 20460
rect 21545 20451 21603 20457
rect 21545 20448 21557 20451
rect 21232 20420 21557 20448
rect 21232 20408 21238 20420
rect 21545 20417 21557 20420
rect 21591 20448 21603 20451
rect 22738 20448 22744 20460
rect 21591 20420 22744 20448
rect 21591 20417 21603 20420
rect 21545 20411 21603 20417
rect 22738 20408 22744 20420
rect 22796 20408 22802 20460
rect 18472 20284 21036 20312
rect 18472 20272 18478 20284
rect 20898 20244 20904 20256
rect 16546 20216 20904 20244
rect 20898 20204 20904 20216
rect 20956 20204 20962 20256
rect 21358 20244 21364 20256
rect 21319 20216 21364 20244
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 3988 20012 5028 20040
rect 1118 19864 1124 19916
rect 1176 19904 1182 19916
rect 1762 19904 1768 19916
rect 1176 19876 1768 19904
rect 1176 19864 1182 19876
rect 1762 19864 1768 19876
rect 1820 19904 1826 19916
rect 2225 19907 2283 19913
rect 2225 19904 2237 19907
rect 1820 19876 2237 19904
rect 1820 19864 1826 19876
rect 2225 19873 2237 19876
rect 2271 19873 2283 19907
rect 2225 19867 2283 19873
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19873 2927 19907
rect 2869 19867 2927 19873
rect 1946 19836 1952 19848
rect 1907 19808 1952 19836
rect 1946 19796 1952 19808
rect 2004 19796 2010 19848
rect 2884 19768 2912 19867
rect 3145 19839 3203 19845
rect 3145 19805 3157 19839
rect 3191 19836 3203 19839
rect 3234 19836 3240 19848
rect 3191 19808 3240 19836
rect 3191 19805 3203 19808
rect 3145 19799 3203 19805
rect 3234 19796 3240 19808
rect 3292 19796 3298 19848
rect 3510 19836 3516 19848
rect 3471 19808 3516 19836
rect 3510 19796 3516 19808
rect 3568 19796 3574 19848
rect 3988 19845 4016 20012
rect 5000 19972 5028 20012
rect 5534 20000 5540 20052
rect 5592 20040 5598 20052
rect 5629 20043 5687 20049
rect 5629 20040 5641 20043
rect 5592 20012 5641 20040
rect 5592 20000 5598 20012
rect 5629 20009 5641 20012
rect 5675 20009 5687 20043
rect 5629 20003 5687 20009
rect 10134 20000 10140 20052
rect 10192 20040 10198 20052
rect 10686 20040 10692 20052
rect 10192 20012 10692 20040
rect 10192 20000 10198 20012
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 10965 20043 11023 20049
rect 10965 20040 10977 20043
rect 10796 20012 10977 20040
rect 6457 19975 6515 19981
rect 6457 19972 6469 19975
rect 5000 19944 6469 19972
rect 6457 19941 6469 19944
rect 6503 19941 6515 19975
rect 6457 19935 6515 19941
rect 10410 19932 10416 19984
rect 10468 19972 10474 19984
rect 10796 19972 10824 20012
rect 10965 20009 10977 20012
rect 11011 20040 11023 20043
rect 11146 20040 11152 20052
rect 11011 20012 11152 20040
rect 11011 20009 11023 20012
rect 10965 20003 11023 20009
rect 11146 20000 11152 20012
rect 11204 20000 11210 20052
rect 11698 20040 11704 20052
rect 11440 20012 11704 20040
rect 10468 19944 10824 19972
rect 10873 19975 10931 19981
rect 10468 19932 10474 19944
rect 10873 19941 10885 19975
rect 10919 19972 10931 19975
rect 11440 19972 11468 20012
rect 11698 20000 11704 20012
rect 11756 20040 11762 20052
rect 13538 20040 13544 20052
rect 11756 20012 12480 20040
rect 13499 20012 13544 20040
rect 11756 20000 11762 20012
rect 10919 19944 11468 19972
rect 10919 19941 10931 19944
rect 10873 19935 10931 19941
rect 6181 19907 6239 19913
rect 6181 19904 6193 19907
rect 5460 19876 6193 19904
rect 3973 19839 4031 19845
rect 3973 19805 3985 19839
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 4065 19839 4123 19845
rect 4065 19805 4077 19839
rect 4111 19836 4123 19839
rect 4111 19808 4568 19836
rect 4111 19805 4123 19808
rect 4065 19799 4123 19805
rect 4540 19780 4568 19808
rect 2884 19740 4108 19768
rect 3421 19703 3479 19709
rect 3421 19669 3433 19703
rect 3467 19700 3479 19703
rect 3694 19700 3700 19712
rect 3467 19672 3700 19700
rect 3467 19669 3479 19672
rect 3421 19663 3479 19669
rect 3694 19660 3700 19672
rect 3752 19660 3758 19712
rect 3789 19703 3847 19709
rect 3789 19669 3801 19703
rect 3835 19700 3847 19703
rect 3970 19700 3976 19712
rect 3835 19672 3976 19700
rect 3835 19669 3847 19672
rect 3789 19663 3847 19669
rect 3970 19660 3976 19672
rect 4028 19660 4034 19712
rect 4080 19700 4108 19740
rect 4154 19728 4160 19780
rect 4212 19768 4218 19780
rect 4310 19771 4368 19777
rect 4310 19768 4322 19771
rect 4212 19740 4322 19768
rect 4212 19728 4218 19740
rect 4310 19737 4322 19740
rect 4356 19737 4368 19771
rect 4310 19731 4368 19737
rect 4522 19728 4528 19780
rect 4580 19728 4586 19780
rect 5350 19700 5356 19712
rect 4080 19672 5356 19700
rect 5350 19660 5356 19672
rect 5408 19660 5414 19712
rect 5460 19709 5488 19876
rect 6181 19873 6193 19876
rect 6227 19904 6239 19907
rect 6362 19904 6368 19916
rect 6227 19876 6368 19904
rect 6227 19873 6239 19876
rect 6181 19867 6239 19873
rect 6362 19864 6368 19876
rect 6420 19864 6426 19916
rect 7098 19904 7104 19916
rect 7059 19876 7104 19904
rect 7098 19864 7104 19876
rect 7156 19864 7162 19916
rect 7929 19907 7987 19913
rect 7929 19873 7941 19907
rect 7975 19873 7987 19907
rect 11054 19904 11060 19916
rect 7929 19867 7987 19873
rect 10244 19876 11060 19904
rect 5994 19796 6000 19848
rect 6052 19836 6058 19848
rect 6089 19839 6147 19845
rect 6089 19836 6101 19839
rect 6052 19808 6101 19836
rect 6052 19796 6058 19808
rect 6089 19805 6101 19808
rect 6135 19805 6147 19839
rect 6822 19836 6828 19848
rect 6783 19808 6828 19836
rect 6089 19799 6147 19805
rect 6822 19796 6828 19808
rect 6880 19796 6886 19848
rect 7944 19836 7972 19867
rect 8662 19836 8668 19848
rect 7944 19808 8668 19836
rect 8662 19796 8668 19808
rect 8720 19836 8726 19848
rect 8757 19839 8815 19845
rect 8757 19836 8769 19839
rect 8720 19808 8769 19836
rect 8720 19796 8726 19808
rect 8757 19805 8769 19808
rect 8803 19805 8815 19839
rect 8757 19799 8815 19805
rect 10054 19839 10112 19845
rect 10054 19805 10066 19839
rect 10100 19836 10112 19839
rect 10244 19836 10272 19876
rect 11054 19864 11060 19876
rect 11112 19864 11118 19916
rect 12452 19913 12480 20012
rect 13538 20000 13544 20012
rect 13596 20000 13602 20052
rect 14274 20040 14280 20052
rect 14235 20012 14280 20040
rect 14274 20000 14280 20012
rect 14332 20000 14338 20052
rect 14826 20040 14832 20052
rect 14787 20012 14832 20040
rect 14826 20000 14832 20012
rect 14884 20000 14890 20052
rect 15102 20040 15108 20052
rect 15063 20012 15108 20040
rect 15102 20000 15108 20012
rect 15160 20000 15166 20052
rect 15381 20043 15439 20049
rect 15381 20009 15393 20043
rect 15427 20040 15439 20043
rect 15930 20040 15936 20052
rect 15427 20012 15936 20040
rect 15427 20009 15439 20012
rect 15381 20003 15439 20009
rect 15930 20000 15936 20012
rect 15988 20000 15994 20052
rect 16117 20043 16175 20049
rect 16117 20009 16129 20043
rect 16163 20040 16175 20043
rect 17034 20040 17040 20052
rect 16163 20012 17040 20040
rect 16163 20009 16175 20012
rect 16117 20003 16175 20009
rect 17034 20000 17040 20012
rect 17092 20000 17098 20052
rect 17678 20040 17684 20052
rect 17639 20012 17684 20040
rect 17678 20000 17684 20012
rect 17736 20000 17742 20052
rect 17954 20040 17960 20052
rect 17915 20012 17960 20040
rect 17954 20000 17960 20012
rect 18012 20000 18018 20052
rect 18233 20043 18291 20049
rect 18233 20009 18245 20043
rect 18279 20040 18291 20043
rect 18322 20040 18328 20052
rect 18279 20012 18328 20040
rect 18279 20009 18291 20012
rect 18233 20003 18291 20009
rect 18322 20000 18328 20012
rect 18380 20000 18386 20052
rect 18509 20043 18567 20049
rect 18509 20009 18521 20043
rect 18555 20040 18567 20043
rect 18782 20040 18788 20052
rect 18555 20012 18788 20040
rect 18555 20009 18567 20012
rect 18509 20003 18567 20009
rect 18782 20000 18788 20012
rect 18840 20000 18846 20052
rect 19429 20043 19487 20049
rect 19429 20009 19441 20043
rect 19475 20040 19487 20043
rect 19702 20040 19708 20052
rect 19475 20012 19708 20040
rect 19475 20009 19487 20012
rect 19429 20003 19487 20009
rect 19702 20000 19708 20012
rect 19760 20000 19766 20052
rect 19797 20043 19855 20049
rect 19797 20009 19809 20043
rect 19843 20040 19855 20043
rect 20530 20040 20536 20052
rect 19843 20012 20536 20040
rect 19843 20009 19855 20012
rect 19797 20003 19855 20009
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 20809 20043 20867 20049
rect 20809 20009 20821 20043
rect 20855 20040 20867 20043
rect 21174 20040 21180 20052
rect 20855 20012 21180 20040
rect 20855 20009 20867 20012
rect 20809 20003 20867 20009
rect 21174 20000 21180 20012
rect 21232 20000 21238 20052
rect 21450 20040 21456 20052
rect 21411 20012 21456 20040
rect 21450 20000 21456 20012
rect 21508 20000 21514 20052
rect 13817 19975 13875 19981
rect 13817 19941 13829 19975
rect 13863 19972 13875 19975
rect 14366 19972 14372 19984
rect 13863 19944 14372 19972
rect 13863 19941 13875 19944
rect 13817 19935 13875 19941
rect 14366 19932 14372 19944
rect 14424 19932 14430 19984
rect 14553 19975 14611 19981
rect 14553 19941 14565 19975
rect 14599 19941 14611 19975
rect 14553 19935 14611 19941
rect 15841 19975 15899 19981
rect 15841 19941 15853 19975
rect 15887 19972 15899 19975
rect 16666 19972 16672 19984
rect 15887 19944 16672 19972
rect 15887 19941 15899 19944
rect 15841 19935 15899 19941
rect 12437 19907 12495 19913
rect 12437 19873 12449 19907
rect 12483 19873 12495 19907
rect 14568 19904 14596 19935
rect 16666 19932 16672 19944
rect 16724 19932 16730 19984
rect 21085 19975 21143 19981
rect 21085 19941 21097 19975
rect 21131 19972 21143 19975
rect 21818 19972 21824 19984
rect 21131 19944 21824 19972
rect 21131 19941 21143 19944
rect 21085 19935 21143 19941
rect 21818 19932 21824 19944
rect 21876 19932 21882 19984
rect 14568 19876 21312 19904
rect 12437 19867 12495 19873
rect 10100 19808 10272 19836
rect 10321 19839 10379 19845
rect 10100 19805 10112 19808
rect 10054 19799 10112 19805
rect 10321 19805 10333 19839
rect 10367 19836 10379 19839
rect 12342 19836 12348 19848
rect 10367 19808 12348 19836
rect 10367 19805 10379 19808
rect 10321 19799 10379 19805
rect 12342 19796 12348 19808
rect 12400 19796 12406 19848
rect 12526 19796 12532 19848
rect 12584 19836 12590 19848
rect 12713 19839 12771 19845
rect 12713 19836 12725 19839
rect 12584 19808 12725 19836
rect 12584 19796 12590 19808
rect 12713 19805 12725 19808
rect 12759 19805 12771 19839
rect 13354 19836 13360 19848
rect 13315 19808 13360 19836
rect 12713 19799 12771 19805
rect 13354 19796 13360 19808
rect 13412 19796 13418 19848
rect 13633 19839 13691 19845
rect 13633 19805 13645 19839
rect 13679 19836 13691 19839
rect 13722 19836 13728 19848
rect 13679 19808 13728 19836
rect 13679 19805 13691 19808
rect 13633 19799 13691 19805
rect 13722 19796 13728 19808
rect 13780 19796 13786 19848
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19836 14151 19839
rect 14274 19836 14280 19848
rect 14139 19808 14280 19836
rect 14139 19805 14151 19808
rect 14093 19799 14151 19805
rect 14274 19796 14280 19808
rect 14332 19796 14338 19848
rect 14366 19796 14372 19848
rect 14424 19836 14430 19848
rect 14645 19839 14703 19845
rect 14424 19808 14469 19836
rect 14424 19796 14430 19808
rect 14645 19805 14657 19839
rect 14691 19836 14703 19839
rect 14734 19836 14740 19848
rect 14691 19808 14740 19836
rect 14691 19805 14703 19808
rect 14645 19799 14703 19805
rect 14734 19796 14740 19808
rect 14792 19796 14798 19848
rect 14921 19839 14979 19845
rect 14921 19805 14933 19839
rect 14967 19805 14979 19839
rect 14921 19799 14979 19805
rect 15197 19839 15255 19845
rect 15197 19805 15209 19839
rect 15243 19836 15255 19839
rect 15286 19836 15292 19848
rect 15243 19808 15292 19836
rect 15243 19805 15255 19808
rect 15197 19799 15255 19805
rect 5534 19728 5540 19780
rect 5592 19768 5598 19780
rect 7745 19771 7803 19777
rect 5592 19740 7420 19768
rect 5592 19728 5598 19740
rect 7392 19712 7420 19740
rect 7745 19737 7757 19771
rect 7791 19768 7803 19771
rect 9214 19768 9220 19780
rect 7791 19740 9220 19768
rect 7791 19737 7803 19740
rect 7745 19731 7803 19737
rect 9214 19728 9220 19740
rect 9272 19728 9278 19780
rect 9858 19728 9864 19780
rect 9916 19768 9922 19780
rect 10597 19771 10655 19777
rect 10597 19768 10609 19771
rect 9916 19740 10609 19768
rect 9916 19728 9922 19740
rect 10597 19737 10609 19740
rect 10643 19768 10655 19771
rect 10962 19768 10968 19780
rect 10643 19740 10968 19768
rect 10643 19737 10655 19740
rect 10597 19731 10655 19737
rect 10962 19728 10968 19740
rect 11020 19728 11026 19780
rect 12100 19771 12158 19777
rect 12100 19737 12112 19771
rect 12146 19768 12158 19771
rect 12618 19768 12624 19780
rect 12146 19740 12624 19768
rect 12146 19737 12158 19740
rect 12100 19731 12158 19737
rect 12618 19728 12624 19740
rect 12676 19728 12682 19780
rect 13538 19728 13544 19780
rect 13596 19768 13602 19780
rect 14936 19768 14964 19799
rect 15286 19796 15292 19808
rect 15344 19796 15350 19848
rect 15378 19796 15384 19848
rect 15436 19836 15442 19848
rect 15657 19839 15715 19845
rect 15657 19836 15669 19839
rect 15436 19808 15669 19836
rect 15436 19796 15442 19808
rect 15657 19805 15669 19808
rect 15703 19805 15715 19839
rect 15930 19836 15936 19848
rect 15891 19808 15936 19836
rect 15657 19799 15715 19805
rect 13596 19740 14964 19768
rect 15672 19768 15700 19799
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 17402 19836 17408 19848
rect 17363 19808 17408 19836
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 17494 19796 17500 19848
rect 17552 19836 17558 19848
rect 17770 19836 17776 19848
rect 17552 19808 17597 19836
rect 17731 19808 17776 19836
rect 17552 19796 17558 19808
rect 17770 19796 17776 19808
rect 17828 19796 17834 19848
rect 18049 19839 18107 19845
rect 18049 19805 18061 19839
rect 18095 19805 18107 19839
rect 18049 19799 18107 19805
rect 18325 19839 18383 19845
rect 18325 19805 18337 19839
rect 18371 19836 18383 19839
rect 18371 19808 18644 19836
rect 18371 19805 18383 19808
rect 18325 19799 18383 19805
rect 16209 19771 16267 19777
rect 16209 19768 16221 19771
rect 15672 19740 16221 19768
rect 13596 19728 13602 19740
rect 5445 19703 5503 19709
rect 5445 19669 5457 19703
rect 5491 19669 5503 19703
rect 5445 19663 5503 19669
rect 5997 19703 6055 19709
rect 5997 19669 6009 19703
rect 6043 19700 6055 19703
rect 6822 19700 6828 19712
rect 6043 19672 6828 19700
rect 6043 19669 6055 19672
rect 5997 19663 6055 19669
rect 6822 19660 6828 19672
rect 6880 19660 6886 19712
rect 6917 19703 6975 19709
rect 6917 19669 6929 19703
rect 6963 19700 6975 19703
rect 7285 19703 7343 19709
rect 7285 19700 7297 19703
rect 6963 19672 7297 19700
rect 6963 19669 6975 19672
rect 6917 19663 6975 19669
rect 7285 19669 7297 19672
rect 7331 19669 7343 19703
rect 7285 19663 7343 19669
rect 7374 19660 7380 19712
rect 7432 19700 7438 19712
rect 7653 19703 7711 19709
rect 7653 19700 7665 19703
rect 7432 19672 7665 19700
rect 7432 19660 7438 19672
rect 7653 19669 7665 19672
rect 7699 19669 7711 19703
rect 8110 19700 8116 19712
rect 8071 19672 8116 19700
rect 7653 19663 7711 19669
rect 8110 19660 8116 19672
rect 8168 19660 8174 19712
rect 8941 19703 8999 19709
rect 8941 19669 8953 19703
rect 8987 19700 8999 19703
rect 9490 19700 9496 19712
rect 8987 19672 9496 19700
rect 8987 19669 8999 19672
rect 8941 19663 8999 19669
rect 9490 19660 9496 19672
rect 9548 19660 9554 19712
rect 10134 19660 10140 19712
rect 10192 19700 10198 19712
rect 10505 19703 10563 19709
rect 10505 19700 10517 19703
rect 10192 19672 10517 19700
rect 10192 19660 10198 19672
rect 10505 19669 10517 19672
rect 10551 19669 10563 19703
rect 14936 19700 14964 19740
rect 16209 19737 16221 19740
rect 16255 19737 16267 19771
rect 16209 19731 16267 19737
rect 16574 19728 16580 19780
rect 16632 19768 16638 19780
rect 16632 19740 16677 19768
rect 16632 19728 16638 19740
rect 16942 19728 16948 19780
rect 17000 19768 17006 19780
rect 18064 19768 18092 19799
rect 17000 19740 18092 19768
rect 17000 19728 17006 19740
rect 18616 19712 18644 19808
rect 19058 19796 19064 19848
rect 19116 19836 19122 19848
rect 19245 19839 19303 19845
rect 19245 19836 19257 19839
rect 19116 19808 19257 19836
rect 19116 19796 19122 19808
rect 19245 19805 19257 19808
rect 19291 19805 19303 19839
rect 19610 19836 19616 19848
rect 19571 19808 19616 19836
rect 19245 19799 19303 19805
rect 19260 19768 19288 19799
rect 19610 19796 19616 19808
rect 19668 19796 19674 19848
rect 20898 19836 20904 19848
rect 20859 19808 20904 19836
rect 20898 19796 20904 19808
rect 20956 19796 20962 19848
rect 21284 19845 21312 19876
rect 21269 19839 21327 19845
rect 21269 19805 21281 19839
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 19889 19771 19947 19777
rect 19889 19768 19901 19771
rect 19260 19740 19901 19768
rect 19889 19737 19901 19740
rect 19935 19737 19947 19771
rect 19889 19731 19947 19737
rect 15473 19703 15531 19709
rect 15473 19700 15485 19703
rect 14936 19672 15485 19700
rect 10505 19663 10563 19669
rect 15473 19669 15485 19672
rect 15519 19669 15531 19703
rect 15473 19663 15531 19669
rect 16298 19660 16304 19712
rect 16356 19700 16362 19712
rect 18414 19700 18420 19712
rect 16356 19672 18420 19700
rect 16356 19660 16362 19672
rect 18414 19660 18420 19672
rect 18472 19660 18478 19712
rect 18598 19700 18604 19712
rect 18559 19672 18604 19700
rect 18598 19660 18604 19672
rect 18656 19660 18662 19712
rect 1104 19610 21896 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21896 19610
rect 1104 19536 21896 19558
rect 2317 19499 2375 19505
rect 2317 19465 2329 19499
rect 2363 19496 2375 19499
rect 2406 19496 2412 19508
rect 2363 19468 2412 19496
rect 2363 19465 2375 19468
rect 2317 19459 2375 19465
rect 2406 19456 2412 19468
rect 2464 19456 2470 19508
rect 3145 19499 3203 19505
rect 3145 19496 3157 19499
rect 2608 19468 3157 19496
rect 1394 19388 1400 19440
rect 1452 19428 1458 19440
rect 2498 19428 2504 19440
rect 1452 19400 2504 19428
rect 1452 19388 1458 19400
rect 2498 19388 2504 19400
rect 2556 19388 2562 19440
rect 2038 19320 2044 19372
rect 2096 19360 2102 19372
rect 2608 19360 2636 19468
rect 3145 19465 3157 19468
rect 3191 19465 3203 19499
rect 4430 19496 4436 19508
rect 3145 19459 3203 19465
rect 4284 19468 4436 19496
rect 2685 19431 2743 19437
rect 2685 19397 2697 19431
rect 2731 19428 2743 19431
rect 4154 19428 4160 19440
rect 2731 19400 4160 19428
rect 2731 19397 2743 19400
rect 2685 19391 2743 19397
rect 4154 19388 4160 19400
rect 4212 19388 4218 19440
rect 4284 19369 4312 19468
rect 4430 19456 4436 19468
rect 4488 19456 4494 19508
rect 4522 19456 4528 19508
rect 4580 19496 4586 19508
rect 4801 19499 4859 19505
rect 4580 19468 4660 19496
rect 4580 19456 4586 19468
rect 4632 19428 4660 19468
rect 4801 19465 4813 19499
rect 4847 19496 4859 19499
rect 5626 19496 5632 19508
rect 4847 19468 5632 19496
rect 4847 19465 4859 19468
rect 4801 19459 4859 19465
rect 5626 19456 5632 19468
rect 5684 19496 5690 19508
rect 7098 19496 7104 19508
rect 5684 19468 6408 19496
rect 7059 19468 7104 19496
rect 5684 19456 5690 19468
rect 4551 19400 6224 19428
rect 4269 19363 4327 19369
rect 2096 19332 3004 19360
rect 2096 19320 2102 19332
rect 198 19252 204 19304
rect 256 19292 262 19304
rect 2222 19292 2228 19304
rect 256 19264 2228 19292
rect 256 19252 262 19264
rect 2222 19252 2228 19264
rect 2280 19252 2286 19304
rect 2976 19301 3004 19332
rect 4269 19329 4281 19363
rect 4315 19329 4327 19363
rect 4269 19323 4327 19329
rect 4430 19320 4436 19372
rect 4488 19320 4494 19372
rect 4551 19369 4579 19400
rect 4525 19363 4583 19369
rect 4525 19329 4537 19363
rect 4571 19329 4583 19363
rect 5534 19360 5540 19372
rect 4724 19334 5540 19360
rect 4525 19323 4583 19329
rect 4632 19332 5540 19334
rect 2777 19295 2835 19301
rect 2777 19261 2789 19295
rect 2823 19261 2835 19295
rect 2777 19255 2835 19261
rect 2961 19295 3019 19301
rect 2961 19261 2973 19295
rect 3007 19261 3019 19295
rect 4448 19292 4476 19320
rect 4632 19306 4752 19332
rect 5534 19320 5540 19332
rect 5592 19320 5598 19372
rect 5902 19320 5908 19372
rect 5960 19369 5966 19372
rect 6196 19369 6224 19400
rect 6380 19369 6408 19468
rect 7098 19456 7104 19468
rect 7156 19456 7162 19508
rect 8662 19496 8668 19508
rect 8623 19468 8668 19496
rect 8662 19456 8668 19468
rect 8720 19456 8726 19508
rect 9858 19456 9864 19508
rect 9916 19496 9922 19508
rect 10502 19496 10508 19508
rect 9916 19468 10508 19496
rect 9916 19456 9922 19468
rect 10502 19456 10508 19468
rect 10560 19456 10566 19508
rect 11057 19499 11115 19505
rect 11057 19465 11069 19499
rect 11103 19496 11115 19499
rect 11701 19499 11759 19505
rect 11701 19496 11713 19499
rect 11103 19468 11713 19496
rect 11103 19465 11115 19468
rect 11057 19459 11115 19465
rect 11701 19465 11713 19468
rect 11747 19465 11759 19499
rect 11701 19459 11759 19465
rect 12713 19499 12771 19505
rect 12713 19465 12725 19499
rect 12759 19465 12771 19499
rect 12713 19459 12771 19465
rect 12805 19499 12863 19505
rect 12805 19465 12817 19499
rect 12851 19496 12863 19499
rect 12894 19496 12900 19508
rect 12851 19468 12900 19496
rect 12851 19465 12863 19468
rect 12805 19459 12863 19465
rect 8110 19388 8116 19440
rect 8168 19428 8174 19440
rect 8214 19431 8272 19437
rect 8214 19428 8226 19431
rect 8168 19400 8226 19428
rect 8168 19388 8174 19400
rect 8214 19397 8226 19400
rect 8260 19397 8272 19431
rect 8214 19391 8272 19397
rect 9306 19388 9312 19440
rect 9364 19428 9370 19440
rect 9778 19431 9836 19437
rect 9778 19428 9790 19431
rect 9364 19400 9790 19428
rect 9364 19388 9370 19400
rect 9778 19397 9790 19400
rect 9824 19397 9836 19431
rect 9778 19391 9836 19397
rect 10042 19388 10048 19440
rect 10100 19428 10106 19440
rect 10229 19431 10287 19437
rect 10229 19428 10241 19431
rect 10100 19400 10241 19428
rect 10100 19388 10106 19400
rect 10229 19397 10241 19400
rect 10275 19397 10287 19431
rect 10229 19391 10287 19397
rect 10318 19388 10324 19440
rect 10376 19428 10382 19440
rect 10413 19431 10471 19437
rect 10413 19428 10425 19431
rect 10376 19400 10425 19428
rect 10376 19388 10382 19400
rect 10413 19397 10425 19400
rect 10459 19397 10471 19431
rect 10413 19391 10471 19397
rect 12161 19431 12219 19437
rect 12161 19397 12173 19431
rect 12207 19428 12219 19431
rect 12434 19428 12440 19440
rect 12207 19400 12440 19428
rect 12207 19397 12219 19400
rect 12161 19391 12219 19397
rect 12434 19388 12440 19400
rect 12492 19388 12498 19440
rect 12728 19428 12756 19459
rect 12894 19456 12900 19468
rect 12952 19456 12958 19508
rect 13265 19499 13323 19505
rect 13265 19465 13277 19499
rect 13311 19496 13323 19499
rect 13446 19496 13452 19508
rect 13311 19468 13452 19496
rect 13311 19465 13323 19468
rect 13265 19459 13323 19465
rect 13446 19456 13452 19468
rect 13504 19456 13510 19508
rect 13541 19499 13599 19505
rect 13541 19465 13553 19499
rect 13587 19496 13599 19499
rect 13630 19496 13636 19508
rect 13587 19468 13636 19496
rect 13587 19465 13599 19468
rect 13541 19459 13599 19465
rect 13630 19456 13636 19468
rect 13688 19456 13694 19508
rect 14366 19496 14372 19508
rect 14327 19468 14372 19496
rect 14366 19456 14372 19468
rect 14424 19456 14430 19508
rect 14734 19496 14740 19508
rect 14695 19468 14740 19496
rect 14734 19456 14740 19468
rect 14792 19456 14798 19508
rect 15197 19499 15255 19505
rect 15197 19465 15209 19499
rect 15243 19496 15255 19499
rect 15930 19496 15936 19508
rect 15243 19468 15936 19496
rect 15243 19465 15255 19468
rect 15197 19459 15255 19465
rect 15930 19456 15936 19468
rect 15988 19456 15994 19508
rect 16209 19499 16267 19505
rect 16209 19465 16221 19499
rect 16255 19496 16267 19499
rect 16298 19496 16304 19508
rect 16255 19468 16304 19496
rect 16255 19465 16267 19468
rect 16209 19459 16267 19465
rect 16298 19456 16304 19468
rect 16356 19456 16362 19508
rect 16853 19499 16911 19505
rect 16853 19465 16865 19499
rect 16899 19496 16911 19499
rect 16942 19496 16948 19508
rect 16899 19468 16948 19496
rect 16899 19465 16911 19468
rect 16853 19459 16911 19465
rect 16942 19456 16948 19468
rect 17000 19456 17006 19508
rect 17126 19496 17132 19508
rect 17087 19468 17132 19496
rect 17126 19456 17132 19468
rect 17184 19456 17190 19508
rect 18877 19499 18935 19505
rect 18877 19465 18889 19499
rect 18923 19496 18935 19499
rect 19610 19496 19616 19508
rect 18923 19468 19616 19496
rect 18923 19465 18935 19468
rect 18877 19459 18935 19465
rect 19610 19456 19616 19468
rect 19668 19456 19674 19508
rect 17034 19428 17040 19440
rect 12728 19400 13400 19428
rect 5960 19360 5972 19369
rect 6174 19363 6232 19369
rect 5960 19332 6005 19360
rect 5960 19323 5972 19332
rect 6174 19329 6186 19363
rect 6220 19360 6232 19363
rect 6365 19363 6423 19369
rect 6220 19332 6322 19360
rect 6220 19329 6232 19332
rect 6174 19323 6232 19329
rect 6365 19329 6377 19363
rect 6411 19329 6423 19363
rect 6365 19323 6423 19329
rect 5960 19320 5966 19323
rect 4632 19292 4660 19306
rect 4448 19264 4660 19292
rect 6196 19292 6224 19323
rect 6454 19320 6460 19372
rect 6512 19360 6518 19372
rect 7009 19363 7067 19369
rect 7009 19360 7021 19363
rect 6512 19332 7021 19360
rect 6512 19320 6518 19332
rect 7009 19329 7021 19332
rect 7055 19329 7067 19363
rect 7009 19323 7067 19329
rect 10502 19320 10508 19372
rect 10560 19360 10566 19372
rect 10965 19363 11023 19369
rect 10965 19360 10977 19363
rect 10560 19332 10977 19360
rect 10560 19320 10566 19332
rect 10965 19329 10977 19332
rect 11011 19329 11023 19363
rect 12066 19360 12072 19372
rect 12027 19332 12072 19360
rect 10965 19323 11023 19329
rect 12066 19320 12072 19332
rect 12124 19360 12130 19372
rect 12529 19363 12587 19369
rect 12124 19332 12480 19360
rect 12124 19320 12130 19332
rect 6546 19292 6552 19304
rect 6196 19264 6552 19292
rect 2961 19255 3019 19261
rect 2792 19224 2820 19255
rect 6546 19252 6552 19264
rect 6604 19252 6610 19304
rect 8478 19292 8484 19304
rect 8439 19264 8484 19292
rect 8478 19252 8484 19264
rect 8536 19252 8542 19304
rect 10045 19295 10103 19301
rect 10045 19261 10057 19295
rect 10091 19292 10103 19295
rect 10318 19292 10324 19304
rect 10091 19264 10324 19292
rect 10091 19261 10103 19264
rect 10045 19255 10103 19261
rect 10318 19252 10324 19264
rect 10376 19252 10382 19304
rect 10410 19252 10416 19304
rect 10468 19292 10474 19304
rect 11054 19292 11060 19304
rect 10468 19264 11060 19292
rect 10468 19252 10474 19264
rect 11054 19252 11060 19264
rect 11112 19252 11118 19304
rect 11241 19295 11299 19301
rect 11241 19261 11253 19295
rect 11287 19292 11299 19295
rect 11974 19292 11980 19304
rect 11287 19264 11980 19292
rect 11287 19261 11299 19264
rect 11241 19255 11299 19261
rect 11974 19252 11980 19264
rect 12032 19252 12038 19304
rect 12250 19292 12256 19304
rect 12211 19264 12256 19292
rect 12250 19252 12256 19264
rect 12308 19252 12314 19304
rect 3142 19224 3148 19236
rect 2792 19196 3148 19224
rect 3142 19184 3148 19196
rect 3200 19184 3206 19236
rect 6178 19184 6184 19236
rect 6236 19224 6242 19236
rect 6236 19196 7604 19224
rect 6236 19184 6242 19196
rect 1995 19159 2053 19165
rect 1995 19125 2007 19159
rect 2041 19156 2053 19159
rect 2958 19156 2964 19168
rect 2041 19128 2964 19156
rect 2041 19125 2053 19128
rect 1995 19119 2053 19125
rect 2958 19116 2964 19128
rect 3016 19116 3022 19168
rect 4709 19159 4767 19165
rect 4709 19125 4721 19159
rect 4755 19156 4767 19159
rect 5442 19156 5448 19168
rect 4755 19128 5448 19156
rect 4755 19125 4767 19128
rect 4709 19119 4767 19125
rect 5442 19116 5448 19128
rect 5500 19116 5506 19168
rect 5534 19116 5540 19168
rect 5592 19156 5598 19168
rect 6822 19156 6828 19168
rect 5592 19128 6828 19156
rect 5592 19116 5598 19128
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 7576 19156 7604 19196
rect 10060 19196 10824 19224
rect 10060 19156 10088 19196
rect 7576 19128 10088 19156
rect 10597 19159 10655 19165
rect 10597 19125 10609 19159
rect 10643 19156 10655 19159
rect 10686 19156 10692 19168
rect 10643 19128 10692 19156
rect 10643 19125 10655 19128
rect 10597 19119 10655 19125
rect 10686 19116 10692 19128
rect 10744 19116 10750 19168
rect 10796 19156 10824 19196
rect 10870 19184 10876 19236
rect 10928 19224 10934 19236
rect 12158 19224 12164 19236
rect 10928 19196 12164 19224
rect 10928 19184 10934 19196
rect 12158 19184 12164 19196
rect 12216 19184 12222 19236
rect 12452 19224 12480 19332
rect 12529 19329 12541 19363
rect 12575 19360 12587 19363
rect 12710 19360 12716 19372
rect 12575 19332 12716 19360
rect 12575 19329 12587 19332
rect 12529 19323 12587 19329
rect 12710 19320 12716 19332
rect 12768 19320 12774 19372
rect 12802 19320 12808 19372
rect 12860 19360 12866 19372
rect 12989 19363 13047 19369
rect 12989 19360 13001 19363
rect 12860 19332 13001 19360
rect 12860 19320 12866 19332
rect 12989 19329 13001 19332
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 13078 19320 13084 19372
rect 13136 19360 13142 19372
rect 13372 19369 13400 19400
rect 16684 19400 17040 19428
rect 13357 19363 13415 19369
rect 13136 19332 13308 19360
rect 13136 19320 13142 19332
rect 13280 19292 13308 19332
rect 13357 19329 13369 19363
rect 13403 19329 13415 19363
rect 13357 19323 13415 19329
rect 14553 19363 14611 19369
rect 14553 19329 14565 19363
rect 14599 19360 14611 19363
rect 14734 19360 14740 19372
rect 14599 19332 14740 19360
rect 14599 19329 14611 19332
rect 14553 19323 14611 19329
rect 14734 19320 14740 19332
rect 14792 19320 14798 19372
rect 15010 19360 15016 19372
rect 14971 19332 15016 19360
rect 15010 19320 15016 19332
rect 15068 19320 15074 19372
rect 16684 19369 16712 19400
rect 17034 19388 17040 19400
rect 17092 19388 17098 19440
rect 16025 19363 16083 19369
rect 16025 19360 16037 19363
rect 15856 19332 16037 19360
rect 13817 19295 13875 19301
rect 13817 19292 13829 19295
rect 13280 19264 13829 19292
rect 13817 19261 13829 19264
rect 13863 19261 13875 19295
rect 13817 19255 13875 19261
rect 13633 19227 13691 19233
rect 13633 19224 13645 19227
rect 12452 19196 13645 19224
rect 13633 19193 13645 19196
rect 13679 19224 13691 19227
rect 13722 19224 13728 19236
rect 13679 19196 13728 19224
rect 13679 19193 13691 19196
rect 13633 19187 13691 19193
rect 13722 19184 13728 19196
rect 13780 19224 13786 19236
rect 14001 19227 14059 19233
rect 14001 19224 14013 19227
rect 13780 19196 14013 19224
rect 13780 19184 13786 19196
rect 14001 19193 14013 19196
rect 14047 19193 14059 19227
rect 14829 19227 14887 19233
rect 14829 19224 14841 19227
rect 14001 19187 14059 19193
rect 14108 19196 14841 19224
rect 11517 19159 11575 19165
rect 11517 19156 11529 19159
rect 10796 19128 11529 19156
rect 11517 19125 11529 19128
rect 11563 19156 11575 19159
rect 11698 19156 11704 19168
rect 11563 19128 11704 19156
rect 11563 19125 11575 19128
rect 11517 19119 11575 19125
rect 11698 19116 11704 19128
rect 11756 19116 11762 19168
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 12894 19156 12900 19168
rect 12492 19128 12900 19156
rect 12492 19116 12498 19128
rect 12894 19116 12900 19128
rect 12952 19116 12958 19168
rect 12986 19116 12992 19168
rect 13044 19156 13050 19168
rect 14108 19156 14136 19196
rect 14829 19193 14841 19196
rect 14875 19193 14887 19227
rect 15470 19224 15476 19236
rect 15431 19196 15476 19224
rect 14829 19187 14887 19193
rect 15470 19184 15476 19196
rect 15528 19184 15534 19236
rect 14274 19156 14280 19168
rect 13044 19128 14136 19156
rect 14235 19128 14280 19156
rect 13044 19116 13050 19128
rect 14274 19116 14280 19128
rect 14332 19116 14338 19168
rect 15286 19116 15292 19168
rect 15344 19156 15350 19168
rect 15654 19156 15660 19168
rect 15344 19128 15389 19156
rect 15615 19128 15660 19156
rect 15344 19116 15350 19128
rect 15654 19116 15660 19128
rect 15712 19116 15718 19168
rect 15746 19116 15752 19168
rect 15804 19156 15810 19168
rect 15856 19165 15884 19332
rect 16025 19329 16037 19332
rect 16071 19329 16083 19363
rect 16025 19323 16083 19329
rect 16669 19363 16727 19369
rect 16669 19329 16681 19363
rect 16715 19329 16727 19363
rect 16669 19323 16727 19329
rect 16945 19363 17003 19369
rect 16945 19329 16957 19363
rect 16991 19360 17003 19363
rect 17218 19360 17224 19372
rect 16991 19332 17224 19360
rect 16991 19329 17003 19332
rect 16945 19323 17003 19329
rect 17218 19320 17224 19332
rect 17276 19320 17282 19372
rect 18506 19320 18512 19372
rect 18564 19360 18570 19372
rect 18693 19363 18751 19369
rect 18693 19360 18705 19363
rect 18564 19332 18705 19360
rect 18564 19320 18570 19332
rect 18693 19329 18705 19332
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 17402 19252 17408 19304
rect 17460 19292 17466 19304
rect 17681 19295 17739 19301
rect 17681 19292 17693 19295
rect 17460 19264 17693 19292
rect 17460 19252 17466 19264
rect 17681 19261 17693 19264
rect 17727 19292 17739 19295
rect 22278 19292 22284 19304
rect 17727 19264 22284 19292
rect 17727 19261 17739 19264
rect 17681 19255 17739 19261
rect 22278 19252 22284 19264
rect 22336 19252 22342 19304
rect 15841 19159 15899 19165
rect 15841 19156 15853 19159
rect 15804 19128 15853 19156
rect 15804 19116 15810 19128
rect 15841 19125 15853 19128
rect 15887 19125 15899 19159
rect 15841 19119 15899 19125
rect 17218 19116 17224 19168
rect 17276 19156 17282 19168
rect 17402 19156 17408 19168
rect 17276 19128 17321 19156
rect 17363 19128 17408 19156
rect 17276 19116 17282 19128
rect 17402 19116 17408 19128
rect 17460 19116 17466 19168
rect 17770 19156 17776 19168
rect 17731 19128 17776 19156
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 18506 19156 18512 19168
rect 18467 19128 18512 19156
rect 18506 19116 18512 19128
rect 18564 19116 18570 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1486 18952 1492 18964
rect 1447 18924 1492 18952
rect 1486 18912 1492 18924
rect 1544 18912 1550 18964
rect 2869 18955 2927 18961
rect 2869 18921 2881 18955
rect 2915 18952 2927 18955
rect 3142 18952 3148 18964
rect 2915 18924 3148 18952
rect 2915 18921 2927 18924
rect 2869 18915 2927 18921
rect 3142 18912 3148 18924
rect 3200 18912 3206 18964
rect 6641 18955 6699 18961
rect 6641 18952 6653 18955
rect 3344 18924 6653 18952
rect 1857 18887 1915 18893
rect 1857 18853 1869 18887
rect 1903 18884 1915 18887
rect 2774 18884 2780 18896
rect 1903 18856 2780 18884
rect 1903 18853 1915 18856
rect 1857 18847 1915 18853
rect 2774 18844 2780 18856
rect 2832 18844 2838 18896
rect 3344 18884 3372 18924
rect 6641 18921 6653 18924
rect 6687 18921 6699 18955
rect 6641 18915 6699 18921
rect 6730 18912 6736 18964
rect 6788 18952 6794 18964
rect 10226 18952 10232 18964
rect 6788 18924 10232 18952
rect 6788 18912 6794 18924
rect 10226 18912 10232 18924
rect 10284 18912 10290 18964
rect 10318 18912 10324 18964
rect 10376 18952 10382 18964
rect 11238 18952 11244 18964
rect 10376 18924 11244 18952
rect 10376 18912 10382 18924
rect 10502 18884 10508 18896
rect 3160 18856 3372 18884
rect 3528 18856 5580 18884
rect 10463 18856 10508 18884
rect 3160 18816 3188 18856
rect 3326 18816 3332 18828
rect 2056 18788 3188 18816
rect 3287 18788 3332 18816
rect 1578 18708 1584 18760
rect 1636 18748 1642 18760
rect 2056 18757 2084 18788
rect 3326 18776 3332 18788
rect 3384 18776 3390 18828
rect 3528 18825 3556 18856
rect 3513 18819 3571 18825
rect 3513 18785 3525 18819
rect 3559 18785 3571 18819
rect 3513 18779 3571 18785
rect 4341 18819 4399 18825
rect 4341 18785 4353 18819
rect 4387 18785 4399 18819
rect 4341 18779 4399 18785
rect 1673 18751 1731 18757
rect 1673 18748 1685 18751
rect 1636 18720 1685 18748
rect 1636 18708 1642 18720
rect 1673 18717 1685 18720
rect 1719 18717 1731 18751
rect 1673 18711 1731 18717
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18717 2099 18751
rect 2041 18711 2099 18717
rect 2774 18708 2780 18760
rect 2832 18748 2838 18760
rect 4356 18748 4384 18779
rect 2832 18720 4384 18748
rect 4893 18751 4951 18757
rect 2832 18708 2838 18720
rect 4893 18717 4905 18751
rect 4939 18748 4951 18751
rect 4982 18748 4988 18760
rect 4939 18720 4988 18748
rect 4939 18717 4951 18720
rect 4893 18711 4951 18717
rect 4982 18708 4988 18720
rect 5040 18708 5046 18760
rect 2222 18640 2228 18692
rect 2280 18680 2286 18692
rect 4706 18680 4712 18692
rect 2280 18652 3832 18680
rect 4667 18652 4712 18680
rect 2280 18640 2286 18652
rect 2133 18615 2191 18621
rect 2133 18581 2145 18615
rect 2179 18612 2191 18615
rect 3142 18612 3148 18624
rect 2179 18584 3148 18612
rect 2179 18581 2191 18584
rect 2133 18575 2191 18581
rect 3142 18572 3148 18584
rect 3200 18572 3206 18624
rect 3237 18615 3295 18621
rect 3237 18581 3249 18615
rect 3283 18612 3295 18615
rect 3326 18612 3332 18624
rect 3283 18584 3332 18612
rect 3283 18581 3295 18584
rect 3237 18575 3295 18581
rect 3326 18572 3332 18584
rect 3384 18572 3390 18624
rect 3804 18621 3832 18652
rect 4706 18640 4712 18652
rect 4764 18640 4770 18692
rect 3789 18615 3847 18621
rect 3789 18581 3801 18615
rect 3835 18581 3847 18615
rect 4154 18612 4160 18624
rect 4115 18584 4160 18612
rect 3789 18575 3847 18581
rect 4154 18572 4160 18584
rect 4212 18572 4218 18624
rect 4249 18615 4307 18621
rect 4249 18581 4261 18615
rect 4295 18612 4307 18615
rect 4430 18612 4436 18624
rect 4295 18584 4436 18612
rect 4295 18581 4307 18584
rect 4249 18575 4307 18581
rect 4430 18572 4436 18584
rect 4488 18572 4494 18624
rect 5074 18572 5080 18624
rect 5132 18612 5138 18624
rect 5169 18615 5227 18621
rect 5169 18612 5181 18615
rect 5132 18584 5181 18612
rect 5132 18572 5138 18584
rect 5169 18581 5181 18584
rect 5215 18581 5227 18615
rect 5552 18612 5580 18856
rect 10502 18844 10508 18856
rect 10560 18844 10566 18896
rect 6546 18816 6552 18828
rect 6507 18788 6552 18816
rect 6546 18776 6552 18788
rect 6604 18816 6610 18828
rect 9398 18816 9404 18828
rect 6604 18788 7328 18816
rect 9359 18788 9404 18816
rect 6604 18776 6610 18788
rect 6293 18751 6351 18757
rect 6293 18717 6305 18751
rect 6339 18748 6351 18751
rect 6454 18748 6460 18760
rect 6339 18720 6460 18748
rect 6339 18717 6351 18720
rect 6293 18711 6351 18717
rect 6454 18708 6460 18720
rect 6512 18708 6518 18760
rect 6638 18708 6644 18760
rect 6696 18748 6702 18760
rect 6825 18751 6883 18757
rect 6825 18748 6837 18751
rect 6696 18720 6837 18748
rect 6696 18708 6702 18720
rect 6825 18717 6837 18720
rect 6871 18717 6883 18751
rect 7300 18748 7328 18788
rect 9398 18776 9404 18788
rect 9456 18776 9462 18828
rect 9490 18776 9496 18828
rect 9548 18816 9554 18828
rect 10612 18825 10640 18924
rect 11238 18912 11244 18924
rect 11296 18952 11302 18964
rect 12342 18952 12348 18964
rect 11296 18924 12348 18952
rect 11296 18912 11302 18924
rect 12342 18912 12348 18924
rect 12400 18912 12406 18964
rect 12618 18912 12624 18964
rect 12676 18952 12682 18964
rect 12713 18955 12771 18961
rect 12713 18952 12725 18955
rect 12676 18924 12725 18952
rect 12676 18912 12682 18924
rect 12713 18921 12725 18924
rect 12759 18921 12771 18955
rect 12713 18915 12771 18921
rect 12989 18955 13047 18961
rect 12989 18921 13001 18955
rect 13035 18952 13047 18955
rect 13354 18952 13360 18964
rect 13035 18924 13360 18952
rect 13035 18921 13047 18924
rect 12989 18915 13047 18921
rect 13354 18912 13360 18924
rect 13412 18912 13418 18964
rect 13630 18912 13636 18964
rect 13688 18952 13694 18964
rect 13817 18955 13875 18961
rect 13817 18952 13829 18955
rect 13688 18924 13829 18952
rect 13688 18912 13694 18924
rect 13817 18921 13829 18924
rect 13863 18921 13875 18955
rect 14642 18952 14648 18964
rect 14603 18924 14648 18952
rect 13817 18915 13875 18921
rect 14642 18912 14648 18924
rect 14700 18912 14706 18964
rect 11974 18884 11980 18896
rect 11935 18856 11980 18884
rect 11974 18844 11980 18856
rect 12032 18844 12038 18896
rect 12802 18844 12808 18896
rect 12860 18884 12866 18896
rect 13081 18887 13139 18893
rect 13081 18884 13093 18887
rect 12860 18856 13093 18884
rect 12860 18844 12866 18856
rect 13081 18853 13093 18856
rect 13127 18853 13139 18887
rect 13081 18847 13139 18853
rect 13262 18844 13268 18896
rect 13320 18884 13326 18896
rect 13449 18887 13507 18893
rect 13449 18884 13461 18887
rect 13320 18856 13461 18884
rect 13320 18844 13326 18856
rect 13449 18853 13461 18856
rect 13495 18853 13507 18887
rect 13449 18847 13507 18853
rect 13906 18844 13912 18896
rect 13964 18884 13970 18896
rect 14277 18887 14335 18893
rect 14277 18884 14289 18887
rect 13964 18856 14289 18884
rect 13964 18844 13970 18856
rect 14277 18853 14289 18856
rect 14323 18853 14335 18887
rect 14277 18847 14335 18853
rect 9953 18819 10011 18825
rect 9548 18788 9593 18816
rect 9548 18776 9554 18788
rect 9953 18785 9965 18819
rect 9999 18785 10011 18819
rect 9953 18779 10011 18785
rect 10597 18819 10655 18825
rect 10597 18785 10609 18819
rect 10643 18785 10655 18819
rect 10597 18779 10655 18785
rect 8297 18751 8355 18757
rect 8297 18748 8309 18751
rect 7300 18720 8309 18748
rect 6825 18711 6883 18717
rect 8297 18717 8309 18720
rect 8343 18748 8355 18751
rect 8478 18748 8484 18760
rect 8343 18720 8484 18748
rect 8343 18717 8355 18720
rect 8297 18711 8355 18717
rect 8478 18708 8484 18720
rect 8536 18708 8542 18760
rect 8570 18708 8576 18760
rect 8628 18748 8634 18760
rect 8665 18751 8723 18757
rect 8665 18748 8677 18751
rect 8628 18720 8677 18748
rect 8628 18708 8634 18720
rect 8665 18717 8677 18720
rect 8711 18717 8723 18751
rect 8665 18711 8723 18717
rect 6546 18640 6552 18692
rect 6604 18680 6610 18692
rect 7006 18680 7012 18692
rect 6604 18652 7012 18680
rect 6604 18640 6610 18652
rect 7006 18640 7012 18652
rect 7064 18640 7070 18692
rect 7834 18640 7840 18692
rect 7892 18680 7898 18692
rect 8030 18683 8088 18689
rect 8030 18680 8042 18683
rect 7892 18652 8042 18680
rect 7892 18640 7898 18652
rect 8030 18649 8042 18652
rect 8076 18649 8088 18683
rect 9398 18680 9404 18692
rect 8030 18643 8088 18649
rect 8588 18652 9404 18680
rect 6917 18615 6975 18621
rect 6917 18612 6929 18615
rect 5552 18584 6929 18612
rect 5169 18575 5227 18581
rect 6917 18581 6929 18584
rect 6963 18612 6975 18615
rect 8110 18612 8116 18624
rect 6963 18584 8116 18612
rect 6963 18581 6975 18584
rect 6917 18575 6975 18581
rect 8110 18572 8116 18584
rect 8168 18572 8174 18624
rect 8588 18621 8616 18652
rect 9398 18640 9404 18652
rect 9456 18640 9462 18692
rect 9968 18680 9996 18779
rect 11606 18776 11612 18828
rect 11664 18816 11670 18828
rect 14461 18819 14519 18825
rect 14461 18816 14473 18819
rect 11664 18788 14473 18816
rect 11664 18776 11670 18788
rect 14461 18785 14473 18788
rect 14507 18785 14519 18819
rect 14461 18779 14519 18785
rect 11974 18708 11980 18760
rect 12032 18748 12038 18760
rect 12069 18751 12127 18757
rect 12069 18748 12081 18751
rect 12032 18720 12081 18748
rect 12032 18708 12038 18720
rect 12069 18717 12081 18720
rect 12115 18717 12127 18751
rect 12069 18711 12127 18717
rect 12158 18708 12164 18760
rect 12216 18748 12222 18760
rect 12802 18748 12808 18760
rect 12216 18720 12388 18748
rect 12763 18720 12808 18748
rect 12216 18708 12222 18720
rect 10864 18683 10922 18689
rect 10864 18680 10876 18683
rect 9968 18652 10876 18680
rect 10864 18649 10876 18652
rect 10910 18680 10922 18683
rect 10910 18652 11284 18680
rect 10910 18649 10922 18652
rect 10864 18643 10922 18649
rect 8573 18615 8631 18621
rect 8573 18581 8585 18615
rect 8619 18581 8631 18615
rect 8938 18612 8944 18624
rect 8899 18584 8944 18612
rect 8573 18575 8631 18581
rect 8938 18572 8944 18584
rect 8996 18572 9002 18624
rect 9306 18612 9312 18624
rect 9267 18584 9312 18612
rect 9306 18572 9312 18584
rect 9364 18572 9370 18624
rect 9950 18572 9956 18624
rect 10008 18612 10014 18624
rect 10045 18615 10103 18621
rect 10045 18612 10057 18615
rect 10008 18584 10057 18612
rect 10008 18572 10014 18584
rect 10045 18581 10057 18584
rect 10091 18581 10103 18615
rect 10045 18575 10103 18581
rect 10137 18615 10195 18621
rect 10137 18581 10149 18615
rect 10183 18612 10195 18615
rect 11146 18612 11152 18624
rect 10183 18584 11152 18612
rect 10183 18581 10195 18584
rect 10137 18575 10195 18581
rect 11146 18572 11152 18584
rect 11204 18572 11210 18624
rect 11256 18612 11284 18652
rect 12250 18612 12256 18624
rect 11256 18584 12256 18612
rect 12250 18572 12256 18584
rect 12308 18572 12314 18624
rect 12360 18612 12388 18720
rect 12802 18708 12808 18720
rect 12860 18708 12866 18760
rect 12894 18708 12900 18760
rect 12952 18748 12958 18760
rect 13357 18751 13415 18757
rect 13357 18748 13369 18751
rect 12952 18720 13369 18748
rect 12952 18708 12958 18720
rect 13357 18717 13369 18720
rect 13403 18748 13415 18751
rect 13403 18720 16574 18748
rect 13403 18717 13415 18720
rect 13357 18711 13415 18717
rect 12618 18640 12624 18692
rect 12676 18680 12682 18692
rect 13633 18683 13691 18689
rect 13633 18680 13645 18683
rect 12676 18652 13645 18680
rect 12676 18640 12682 18652
rect 13633 18649 13645 18652
rect 13679 18649 13691 18683
rect 14826 18680 14832 18692
rect 14787 18652 14832 18680
rect 13633 18643 13691 18649
rect 14826 18640 14832 18652
rect 14884 18640 14890 18692
rect 16546 18680 16574 18720
rect 17954 18680 17960 18692
rect 16546 18652 17960 18680
rect 17954 18640 17960 18652
rect 18012 18640 18018 18692
rect 14093 18615 14151 18621
rect 14093 18612 14105 18615
rect 12360 18584 14105 18612
rect 14093 18581 14105 18584
rect 14139 18581 14151 18615
rect 14093 18575 14151 18581
rect 1104 18522 21896 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21896 18522
rect 1104 18448 21896 18470
rect 1857 18411 1915 18417
rect 1857 18377 1869 18411
rect 1903 18377 1915 18411
rect 1857 18371 1915 18377
rect 2225 18411 2283 18417
rect 2225 18377 2237 18411
rect 2271 18408 2283 18411
rect 2314 18408 2320 18420
rect 2271 18380 2320 18408
rect 2271 18377 2283 18380
rect 2225 18371 2283 18377
rect 1872 18340 1900 18371
rect 2314 18368 2320 18380
rect 2372 18368 2378 18420
rect 2774 18368 2780 18420
rect 2832 18408 2838 18420
rect 3786 18408 3792 18420
rect 2832 18380 2877 18408
rect 2976 18380 3792 18408
rect 2832 18368 2838 18380
rect 2866 18340 2872 18352
rect 1872 18312 2872 18340
rect 2866 18300 2872 18312
rect 2924 18300 2930 18352
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 1946 18272 1952 18284
rect 1719 18244 1952 18272
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 2041 18275 2099 18281
rect 2041 18241 2053 18275
rect 2087 18241 2099 18275
rect 2041 18235 2099 18241
rect 2056 18204 2084 18235
rect 2314 18232 2320 18284
rect 2372 18272 2378 18284
rect 2409 18275 2467 18281
rect 2409 18272 2421 18275
rect 2372 18244 2421 18272
rect 2372 18232 2378 18244
rect 2409 18241 2421 18244
rect 2455 18241 2467 18275
rect 2409 18235 2467 18241
rect 2501 18275 2559 18281
rect 2682 18276 2688 18284
rect 2501 18241 2513 18275
rect 2547 18272 2559 18275
rect 2608 18272 2688 18276
rect 2547 18248 2688 18272
rect 2547 18244 2636 18248
rect 2547 18241 2559 18244
rect 2501 18235 2559 18241
rect 2682 18232 2688 18248
rect 2740 18232 2746 18284
rect 2774 18232 2780 18284
rect 2832 18272 2838 18284
rect 2976 18272 3004 18380
rect 3786 18368 3792 18380
rect 3844 18408 3850 18420
rect 4246 18408 4252 18420
rect 3844 18380 4252 18408
rect 3844 18368 3850 18380
rect 4246 18368 4252 18380
rect 4304 18368 4310 18420
rect 4430 18408 4436 18420
rect 4391 18380 4436 18408
rect 4430 18368 4436 18380
rect 4488 18368 4494 18420
rect 4893 18411 4951 18417
rect 4893 18377 4905 18411
rect 4939 18408 4951 18411
rect 4939 18380 5948 18408
rect 4939 18377 4951 18380
rect 4893 18371 4951 18377
rect 3912 18343 3970 18349
rect 3912 18309 3924 18343
rect 3958 18340 3970 18343
rect 5261 18343 5319 18349
rect 5261 18340 5273 18343
rect 3958 18312 5273 18340
rect 3958 18309 3970 18312
rect 3912 18303 3970 18309
rect 5261 18309 5273 18312
rect 5307 18309 5319 18343
rect 5920 18340 5948 18380
rect 5994 18368 6000 18420
rect 6052 18408 6058 18420
rect 6365 18411 6423 18417
rect 6365 18408 6377 18411
rect 6052 18380 6377 18408
rect 6052 18368 6058 18380
rect 6365 18377 6377 18380
rect 6411 18377 6423 18411
rect 6365 18371 6423 18377
rect 6822 18368 6828 18420
rect 6880 18408 6886 18420
rect 7469 18411 7527 18417
rect 7469 18408 7481 18411
rect 6880 18380 7481 18408
rect 6880 18368 6886 18380
rect 7469 18377 7481 18380
rect 7515 18377 7527 18411
rect 7469 18371 7527 18377
rect 8294 18368 8300 18420
rect 8352 18408 8358 18420
rect 8389 18411 8447 18417
rect 8389 18408 8401 18411
rect 8352 18380 8401 18408
rect 8352 18368 8358 18380
rect 8389 18377 8401 18380
rect 8435 18377 8447 18411
rect 8389 18371 8447 18377
rect 8849 18411 8907 18417
rect 8849 18377 8861 18411
rect 8895 18408 8907 18411
rect 9306 18408 9312 18420
rect 8895 18380 9312 18408
rect 8895 18377 8907 18380
rect 8849 18371 8907 18377
rect 9306 18368 9312 18380
rect 9364 18368 9370 18420
rect 9493 18411 9551 18417
rect 9493 18377 9505 18411
rect 9539 18408 9551 18411
rect 9582 18408 9588 18420
rect 9539 18380 9588 18408
rect 9539 18377 9551 18380
rect 9493 18371 9551 18377
rect 9582 18368 9588 18380
rect 9640 18368 9646 18420
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 10781 18411 10839 18417
rect 10781 18408 10793 18411
rect 9732 18380 10793 18408
rect 9732 18368 9738 18380
rect 10781 18377 10793 18380
rect 10827 18377 10839 18411
rect 11146 18408 11152 18420
rect 11107 18380 11152 18408
rect 10781 18371 10839 18377
rect 11146 18368 11152 18380
rect 11204 18368 11210 18420
rect 11517 18411 11575 18417
rect 11517 18377 11529 18411
rect 11563 18377 11575 18411
rect 11517 18371 11575 18377
rect 11793 18411 11851 18417
rect 11793 18377 11805 18411
rect 11839 18408 11851 18411
rect 12158 18408 12164 18420
rect 11839 18380 12164 18408
rect 11839 18377 11851 18380
rect 11793 18371 11851 18377
rect 11532 18340 11560 18371
rect 12158 18368 12164 18380
rect 12216 18368 12222 18420
rect 13633 18411 13691 18417
rect 13633 18408 13645 18411
rect 12268 18380 13645 18408
rect 5920 18312 11560 18340
rect 5261 18303 5319 18309
rect 11606 18300 11612 18352
rect 11664 18340 11670 18352
rect 12268 18340 12296 18380
rect 13633 18377 13645 18380
rect 13679 18377 13691 18411
rect 13633 18371 13691 18377
rect 13909 18411 13967 18417
rect 13909 18377 13921 18411
rect 13955 18408 13967 18411
rect 14458 18408 14464 18420
rect 13955 18380 14464 18408
rect 13955 18377 13967 18380
rect 13909 18371 13967 18377
rect 14458 18368 14464 18380
rect 14516 18368 14522 18420
rect 11664 18312 12296 18340
rect 11664 18300 11670 18312
rect 12342 18300 12348 18352
rect 12400 18340 12406 18352
rect 12400 18312 13216 18340
rect 12400 18300 12406 18312
rect 2832 18244 3004 18272
rect 2832 18232 2838 18244
rect 3418 18232 3424 18284
rect 3476 18272 3482 18284
rect 4157 18275 4215 18281
rect 3476 18244 4108 18272
rect 3476 18232 3482 18244
rect 4080 18204 4108 18244
rect 4157 18241 4169 18275
rect 4203 18272 4215 18275
rect 4522 18272 4528 18284
rect 4203 18244 4528 18272
rect 4203 18241 4215 18244
rect 4157 18235 4215 18241
rect 4522 18232 4528 18244
rect 4580 18232 4586 18284
rect 4798 18272 4804 18284
rect 4759 18244 4804 18272
rect 4798 18232 4804 18244
rect 4856 18232 4862 18284
rect 5905 18275 5963 18281
rect 5905 18272 5917 18275
rect 5092 18244 5917 18272
rect 5092 18216 5120 18244
rect 5905 18241 5917 18244
rect 5951 18241 5963 18275
rect 5905 18235 5963 18241
rect 6181 18275 6239 18281
rect 6181 18241 6193 18275
rect 6227 18241 6239 18275
rect 6546 18272 6552 18284
rect 6507 18244 6552 18272
rect 6181 18235 6239 18241
rect 4890 18204 4896 18216
rect 2056 18176 2820 18204
rect 4080 18176 4896 18204
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 2314 18028 2320 18080
rect 2372 18068 2378 18080
rect 2498 18068 2504 18080
rect 2372 18040 2504 18068
rect 2372 18028 2378 18040
rect 2498 18028 2504 18040
rect 2556 18028 2562 18080
rect 2682 18068 2688 18080
rect 2643 18040 2688 18068
rect 2682 18028 2688 18040
rect 2740 18028 2746 18080
rect 2792 18068 2820 18176
rect 4890 18164 4896 18176
rect 4948 18164 4954 18216
rect 5074 18204 5080 18216
rect 5035 18176 5080 18204
rect 5074 18164 5080 18176
rect 5132 18164 5138 18216
rect 5626 18164 5632 18216
rect 5684 18204 5690 18216
rect 6196 18204 6224 18235
rect 6546 18232 6552 18244
rect 6604 18232 6610 18284
rect 6822 18232 6828 18284
rect 6880 18272 6886 18284
rect 7009 18275 7067 18281
rect 7009 18272 7021 18275
rect 6880 18244 7021 18272
rect 6880 18232 6886 18244
rect 7009 18241 7021 18244
rect 7055 18241 7067 18275
rect 8110 18272 8116 18284
rect 8071 18244 8116 18272
rect 7009 18235 7067 18241
rect 8110 18232 8116 18244
rect 8168 18232 8174 18284
rect 8573 18275 8631 18281
rect 8573 18241 8585 18275
rect 8619 18272 8631 18275
rect 8938 18272 8944 18284
rect 8619 18244 8944 18272
rect 8619 18241 8631 18244
rect 8573 18235 8631 18241
rect 8938 18232 8944 18244
rect 8996 18232 9002 18284
rect 9122 18272 9128 18284
rect 9083 18244 9128 18272
rect 9122 18232 9128 18244
rect 9180 18232 9186 18284
rect 9401 18275 9459 18281
rect 9401 18241 9413 18275
rect 9447 18241 9459 18275
rect 9766 18272 9772 18284
rect 9727 18244 9772 18272
rect 9401 18235 9459 18241
rect 5684 18176 6224 18204
rect 6733 18207 6791 18213
rect 5684 18164 5690 18176
rect 6733 18173 6745 18207
rect 6779 18173 6791 18207
rect 6914 18204 6920 18216
rect 6875 18176 6920 18204
rect 6733 18167 6791 18173
rect 5997 18139 6055 18145
rect 5997 18136 6009 18139
rect 4163 18108 6009 18136
rect 4163 18068 4191 18108
rect 5997 18105 6009 18108
rect 6043 18105 6055 18139
rect 6748 18136 6776 18167
rect 6914 18164 6920 18176
rect 6972 18164 6978 18216
rect 9416 18204 9444 18235
rect 9766 18232 9772 18244
rect 9824 18232 9830 18284
rect 10686 18272 10692 18284
rect 10647 18244 10692 18272
rect 10686 18232 10692 18244
rect 10744 18232 10750 18284
rect 11698 18272 11704 18284
rect 11659 18244 11704 18272
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 12618 18272 12624 18284
rect 11799 18244 12624 18272
rect 10594 18204 10600 18216
rect 7116 18176 8984 18204
rect 7006 18136 7012 18148
rect 6748 18108 7012 18136
rect 5997 18099 6055 18105
rect 7006 18096 7012 18108
rect 7064 18096 7070 18148
rect 2792 18040 4191 18068
rect 4341 18071 4399 18077
rect 4341 18037 4353 18071
rect 4387 18068 4399 18071
rect 4614 18068 4620 18080
rect 4387 18040 4620 18068
rect 4387 18037 4399 18040
rect 4341 18031 4399 18037
rect 4614 18028 4620 18040
rect 4672 18028 4678 18080
rect 4890 18028 4896 18080
rect 4948 18068 4954 18080
rect 7116 18068 7144 18176
rect 8956 18145 8984 18176
rect 9416 18176 10600 18204
rect 8297 18139 8355 18145
rect 8297 18105 8309 18139
rect 8343 18105 8355 18139
rect 8297 18099 8355 18105
rect 8941 18139 8999 18145
rect 8941 18105 8953 18139
rect 8987 18105 8999 18139
rect 9214 18136 9220 18148
rect 9175 18108 9220 18136
rect 8941 18099 8999 18105
rect 4948 18040 7144 18068
rect 4948 18028 4954 18040
rect 7190 18028 7196 18080
rect 7248 18068 7254 18080
rect 7377 18071 7435 18077
rect 7377 18068 7389 18071
rect 7248 18040 7389 18068
rect 7248 18028 7254 18040
rect 7377 18037 7389 18040
rect 7423 18037 7435 18071
rect 8312 18068 8340 18099
rect 9214 18096 9220 18108
rect 9272 18096 9278 18148
rect 9416 18068 9444 18176
rect 10594 18164 10600 18176
rect 10652 18164 10658 18216
rect 11054 18164 11060 18216
rect 11112 18204 11118 18216
rect 11799 18204 11827 18244
rect 12618 18232 12624 18244
rect 12676 18232 12682 18284
rect 12917 18275 12975 18281
rect 12917 18241 12929 18275
rect 12963 18272 12975 18275
rect 13078 18272 13084 18284
rect 12963 18244 13084 18272
rect 12963 18241 12975 18244
rect 12917 18235 12975 18241
rect 13078 18232 13084 18244
rect 13136 18232 13142 18284
rect 13188 18281 13216 18312
rect 13262 18300 13268 18352
rect 13320 18340 13326 18352
rect 14001 18343 14059 18349
rect 14001 18340 14013 18343
rect 13320 18312 14013 18340
rect 13320 18300 13326 18312
rect 14001 18309 14013 18312
rect 14047 18309 14059 18343
rect 14001 18303 14059 18309
rect 13173 18275 13231 18281
rect 13173 18241 13185 18275
rect 13219 18241 13231 18275
rect 13446 18272 13452 18284
rect 13407 18244 13452 18272
rect 13173 18235 13231 18241
rect 13446 18232 13452 18244
rect 13504 18232 13510 18284
rect 11112 18176 11827 18204
rect 11112 18164 11118 18176
rect 10410 18068 10416 18080
rect 8312 18040 9444 18068
rect 10371 18040 10416 18068
rect 7377 18031 7435 18037
rect 10410 18028 10416 18040
rect 10468 18028 10474 18080
rect 10502 18028 10508 18080
rect 10560 18068 10566 18080
rect 10560 18040 10605 18068
rect 10560 18028 10566 18040
rect 10962 18028 10968 18080
rect 11020 18068 11026 18080
rect 13265 18071 13323 18077
rect 13265 18068 13277 18071
rect 11020 18040 13277 18068
rect 11020 18028 11026 18040
rect 13265 18037 13277 18040
rect 13311 18037 13323 18071
rect 13265 18031 13323 18037
rect 14826 18028 14832 18080
rect 14884 18068 14890 18080
rect 17770 18068 17776 18080
rect 14884 18040 17776 18068
rect 14884 18028 14890 18040
rect 17770 18028 17776 18040
rect 17828 18028 17834 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 1854 17864 1860 17876
rect 1815 17836 1860 17864
rect 1854 17824 1860 17836
rect 1912 17824 1918 17876
rect 2222 17864 2228 17876
rect 2183 17836 2228 17864
rect 2222 17824 2228 17836
rect 2280 17824 2286 17876
rect 2590 17864 2596 17876
rect 2551 17836 2596 17864
rect 2590 17824 2596 17836
rect 2648 17824 2654 17876
rect 3050 17864 3056 17876
rect 3011 17836 3056 17864
rect 3050 17824 3056 17836
rect 3108 17824 3114 17876
rect 3418 17864 3424 17876
rect 3379 17836 3424 17864
rect 3418 17824 3424 17836
rect 3476 17824 3482 17876
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 10321 17867 10379 17873
rect 10321 17864 10333 17867
rect 4120 17836 10333 17864
rect 4120 17824 4126 17836
rect 10321 17833 10333 17836
rect 10367 17833 10379 17867
rect 10321 17827 10379 17833
rect 10778 17824 10784 17876
rect 10836 17864 10842 17876
rect 12986 17864 12992 17876
rect 10836 17836 12992 17864
rect 10836 17824 10842 17836
rect 12986 17824 12992 17836
rect 13044 17824 13050 17876
rect 13078 17824 13084 17876
rect 13136 17864 13142 17876
rect 13265 17867 13323 17873
rect 13265 17864 13277 17867
rect 13136 17836 13277 17864
rect 13136 17824 13142 17836
rect 13265 17833 13277 17836
rect 13311 17833 13323 17867
rect 13814 17864 13820 17876
rect 13775 17836 13820 17864
rect 13265 17827 13323 17833
rect 13814 17824 13820 17836
rect 13872 17824 13878 17876
rect 4798 17756 4804 17808
rect 4856 17796 4862 17808
rect 8757 17799 8815 17805
rect 4856 17768 7328 17796
rect 4856 17756 4862 17768
rect 5534 17688 5540 17740
rect 5592 17728 5598 17740
rect 6638 17728 6644 17740
rect 5592 17700 6644 17728
rect 5592 17688 5598 17700
rect 6638 17688 6644 17700
rect 6696 17688 6702 17740
rect 1670 17660 1676 17672
rect 1631 17632 1676 17660
rect 1670 17620 1676 17632
rect 1728 17620 1734 17672
rect 2041 17663 2099 17669
rect 2041 17629 2053 17663
rect 2087 17660 2099 17663
rect 2222 17660 2228 17672
rect 2087 17632 2228 17660
rect 2087 17629 2099 17632
rect 2041 17623 2099 17629
rect 2222 17620 2228 17632
rect 2280 17620 2286 17672
rect 2409 17663 2467 17669
rect 2409 17629 2421 17663
rect 2455 17660 2467 17663
rect 2590 17660 2596 17672
rect 2455 17632 2596 17660
rect 2455 17629 2467 17632
rect 2409 17623 2467 17629
rect 2590 17620 2596 17632
rect 2648 17620 2654 17672
rect 2777 17663 2835 17669
rect 2777 17629 2789 17663
rect 2823 17629 2835 17663
rect 2777 17623 2835 17629
rect 2792 17592 2820 17623
rect 2866 17620 2872 17672
rect 2924 17660 2930 17672
rect 3234 17660 3240 17672
rect 2924 17632 2969 17660
rect 3195 17632 3240 17660
rect 2924 17620 2930 17632
rect 3234 17620 3240 17632
rect 3292 17620 3298 17672
rect 3789 17663 3847 17669
rect 3789 17629 3801 17663
rect 3835 17660 3847 17663
rect 4522 17660 4528 17672
rect 3835 17632 4528 17660
rect 3835 17629 3847 17632
rect 3789 17623 3847 17629
rect 4522 17620 4528 17632
rect 4580 17620 4586 17672
rect 5258 17660 5264 17672
rect 5219 17632 5264 17660
rect 5258 17620 5264 17632
rect 5316 17620 5322 17672
rect 5997 17663 6055 17669
rect 5997 17629 6009 17663
rect 6043 17629 6055 17663
rect 7190 17660 7196 17672
rect 7151 17632 7196 17660
rect 5997 17623 6055 17629
rect 3050 17592 3056 17604
rect 2792 17564 3056 17592
rect 3050 17552 3056 17564
rect 3108 17552 3114 17604
rect 3142 17552 3148 17604
rect 3200 17592 3206 17604
rect 4034 17595 4092 17601
rect 4034 17592 4046 17595
rect 3200 17564 4046 17592
rect 3200 17552 3206 17564
rect 4034 17561 4046 17564
rect 4080 17561 4092 17595
rect 6012 17592 6040 17623
rect 7190 17620 7196 17632
rect 7248 17620 7254 17672
rect 7300 17660 7328 17768
rect 8757 17765 8769 17799
rect 8803 17796 8815 17799
rect 10042 17796 10048 17808
rect 8803 17768 10048 17796
rect 8803 17765 8815 17768
rect 8757 17759 8815 17765
rect 7466 17728 7472 17740
rect 7427 17700 7472 17728
rect 7466 17688 7472 17700
rect 7524 17688 7530 17740
rect 7558 17688 7564 17740
rect 7616 17728 7622 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 7616 17700 8401 17728
rect 7616 17688 7622 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 7745 17663 7803 17669
rect 7745 17660 7757 17663
rect 7300 17632 7757 17660
rect 7745 17629 7757 17632
rect 7791 17660 7803 17663
rect 8297 17663 8355 17669
rect 7791 17632 7972 17660
rect 7791 17629 7803 17632
rect 7745 17623 7803 17629
rect 4034 17555 4092 17561
rect 5184 17564 6040 17592
rect 7285 17595 7343 17601
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 5074 17484 5080 17536
rect 5132 17524 5138 17536
rect 5184 17533 5212 17564
rect 7285 17561 7297 17595
rect 7331 17592 7343 17595
rect 7331 17564 7880 17592
rect 7331 17561 7343 17564
rect 7285 17555 7343 17561
rect 5169 17527 5227 17533
rect 5169 17524 5181 17527
rect 5132 17496 5181 17524
rect 5132 17484 5138 17496
rect 5169 17493 5181 17496
rect 5215 17493 5227 17527
rect 5169 17487 5227 17493
rect 5534 17484 5540 17536
rect 5592 17524 5598 17536
rect 5905 17527 5963 17533
rect 5905 17524 5917 17527
rect 5592 17496 5917 17524
rect 5592 17484 5598 17496
rect 5905 17493 5917 17496
rect 5951 17493 5963 17527
rect 6638 17524 6644 17536
rect 6599 17496 6644 17524
rect 5905 17487 5963 17493
rect 6638 17484 6644 17496
rect 6696 17484 6702 17536
rect 6730 17484 6736 17536
rect 6788 17524 6794 17536
rect 6825 17527 6883 17533
rect 6825 17524 6837 17527
rect 6788 17496 6837 17524
rect 6788 17484 6794 17496
rect 6825 17493 6837 17496
rect 6871 17493 6883 17527
rect 6825 17487 6883 17493
rect 7006 17484 7012 17536
rect 7064 17524 7070 17536
rect 7558 17524 7564 17536
rect 7064 17496 7564 17524
rect 7064 17484 7070 17496
rect 7558 17484 7564 17496
rect 7616 17484 7622 17536
rect 7852 17533 7880 17564
rect 7837 17527 7895 17533
rect 7837 17493 7849 17527
rect 7883 17493 7895 17527
rect 7944 17524 7972 17632
rect 8297 17629 8309 17663
rect 8343 17660 8355 17663
rect 8772 17660 8800 17759
rect 10042 17756 10048 17768
rect 10100 17796 10106 17808
rect 10870 17796 10876 17808
rect 10100 17768 10876 17796
rect 10100 17756 10106 17768
rect 10870 17756 10876 17768
rect 10928 17756 10934 17808
rect 9030 17728 9036 17740
rect 8991 17700 9036 17728
rect 9030 17688 9036 17700
rect 9088 17688 9094 17740
rect 9674 17688 9680 17740
rect 9732 17728 9738 17740
rect 10778 17728 10784 17740
rect 9732 17700 10784 17728
rect 9732 17688 9738 17700
rect 10778 17688 10784 17700
rect 10836 17688 10842 17740
rect 10965 17731 11023 17737
rect 10965 17697 10977 17731
rect 11011 17728 11023 17731
rect 11011 17700 11100 17728
rect 11011 17697 11023 17700
rect 10965 17691 11023 17697
rect 10226 17660 10232 17672
rect 8343 17632 8800 17660
rect 10187 17632 10232 17660
rect 8343 17629 8355 17632
rect 8297 17623 8355 17629
rect 10226 17620 10232 17632
rect 10284 17620 10290 17672
rect 8205 17595 8263 17601
rect 8205 17561 8217 17595
rect 8251 17592 8263 17595
rect 8478 17592 8484 17604
rect 8251 17564 8484 17592
rect 8251 17561 8263 17564
rect 8205 17555 8263 17561
rect 8478 17552 8484 17564
rect 8536 17552 8542 17604
rect 9309 17595 9367 17601
rect 9309 17561 9321 17595
rect 9355 17592 9367 17595
rect 9769 17595 9827 17601
rect 9769 17592 9781 17595
rect 9355 17564 9781 17592
rect 9355 17561 9367 17564
rect 9309 17555 9367 17561
rect 9769 17561 9781 17564
rect 9815 17561 9827 17595
rect 9769 17555 9827 17561
rect 10689 17595 10747 17601
rect 10689 17561 10701 17595
rect 10735 17592 10747 17595
rect 11072 17592 11100 17700
rect 11149 17663 11207 17669
rect 11149 17629 11161 17663
rect 11195 17660 11207 17663
rect 11238 17660 11244 17672
rect 11195 17632 11244 17660
rect 11195 17629 11207 17632
rect 11149 17623 11207 17629
rect 11238 17620 11244 17632
rect 11296 17620 11302 17672
rect 12621 17663 12679 17669
rect 12621 17660 12633 17663
rect 11348 17632 12633 17660
rect 11348 17592 11376 17632
rect 10735 17564 11008 17592
rect 11072 17564 11376 17592
rect 11416 17595 11474 17601
rect 10735 17561 10747 17564
rect 10689 17555 10747 17561
rect 9217 17527 9275 17533
rect 9217 17524 9229 17527
rect 7944 17496 9229 17524
rect 7837 17487 7895 17493
rect 9217 17493 9229 17496
rect 9263 17493 9275 17527
rect 9217 17487 9275 17493
rect 9398 17484 9404 17536
rect 9456 17524 9462 17536
rect 9677 17527 9735 17533
rect 9677 17524 9689 17527
rect 9456 17496 9689 17524
rect 9456 17484 9462 17496
rect 9677 17493 9689 17496
rect 9723 17493 9735 17527
rect 10042 17524 10048 17536
rect 10003 17496 10048 17524
rect 9677 17487 9735 17493
rect 10042 17484 10048 17496
rect 10100 17484 10106 17536
rect 10778 17484 10784 17536
rect 10836 17524 10842 17536
rect 10980 17524 11008 17564
rect 11416 17561 11428 17595
rect 11462 17592 11474 17595
rect 11698 17592 11704 17604
rect 11462 17564 11704 17592
rect 11462 17561 11474 17564
rect 11416 17555 11474 17561
rect 11698 17552 11704 17564
rect 11756 17552 11762 17604
rect 11146 17524 11152 17536
rect 10836 17496 10881 17524
rect 10980 17496 11152 17524
rect 10836 17484 10842 17496
rect 11146 17484 11152 17496
rect 11204 17484 11210 17536
rect 12544 17533 12572 17632
rect 12621 17629 12633 17632
rect 12667 17629 12679 17663
rect 12621 17623 12679 17629
rect 13354 17620 13360 17672
rect 13412 17660 13418 17672
rect 13633 17663 13691 17669
rect 13633 17660 13645 17663
rect 13412 17632 13645 17660
rect 13412 17620 13418 17632
rect 13633 17629 13645 17632
rect 13679 17629 13691 17663
rect 21269 17663 21327 17669
rect 21269 17660 21281 17663
rect 13633 17623 13691 17629
rect 21100 17632 21281 17660
rect 21100 17536 21128 17632
rect 21269 17629 21281 17632
rect 21315 17629 21327 17663
rect 21269 17623 21327 17629
rect 12529 17527 12587 17533
rect 12529 17493 12541 17527
rect 12575 17493 12587 17527
rect 12529 17487 12587 17493
rect 12618 17484 12624 17536
rect 12676 17524 12682 17536
rect 13357 17527 13415 17533
rect 13357 17524 13369 17527
rect 12676 17496 13369 17524
rect 12676 17484 12682 17496
rect 13357 17493 13369 17496
rect 13403 17493 13415 17527
rect 21082 17524 21088 17536
rect 21043 17496 21088 17524
rect 13357 17487 13415 17493
rect 21082 17484 21088 17496
rect 21140 17484 21146 17536
rect 21450 17524 21456 17536
rect 21411 17496 21456 17524
rect 21450 17484 21456 17496
rect 21508 17484 21514 17536
rect 1104 17434 21896 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21896 17434
rect 1104 17360 21896 17382
rect 1762 17280 1768 17332
rect 1820 17320 1826 17332
rect 3326 17320 3332 17332
rect 1820 17292 3332 17320
rect 1820 17280 1826 17292
rect 3326 17280 3332 17292
rect 3384 17280 3390 17332
rect 3513 17323 3571 17329
rect 3513 17289 3525 17323
rect 3559 17320 3571 17323
rect 3881 17323 3939 17329
rect 3881 17320 3893 17323
rect 3559 17292 3893 17320
rect 3559 17289 3571 17292
rect 3513 17283 3571 17289
rect 3881 17289 3893 17292
rect 3927 17289 3939 17323
rect 6365 17323 6423 17329
rect 6365 17320 6377 17323
rect 3881 17283 3939 17289
rect 3988 17292 6377 17320
rect 3988 17252 4016 17292
rect 6365 17289 6377 17292
rect 6411 17289 6423 17323
rect 6365 17283 6423 17289
rect 7098 17280 7104 17332
rect 7156 17320 7162 17332
rect 7156 17292 10456 17320
rect 7156 17280 7162 17292
rect 2884 17224 4016 17252
rect 5844 17255 5902 17261
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17184 1731 17187
rect 1762 17184 1768 17196
rect 1719 17156 1768 17184
rect 1719 17153 1731 17156
rect 1673 17147 1731 17153
rect 1762 17144 1768 17156
rect 1820 17144 1826 17196
rect 2038 17184 2044 17196
rect 1999 17156 2044 17184
rect 2038 17144 2044 17156
rect 2096 17144 2102 17196
rect 2130 17144 2136 17196
rect 2188 17184 2194 17196
rect 2225 17187 2283 17193
rect 2225 17184 2237 17187
rect 2188 17156 2237 17184
rect 2188 17144 2194 17156
rect 2225 17153 2237 17156
rect 2271 17153 2283 17187
rect 2225 17147 2283 17153
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17184 2559 17187
rect 2774 17184 2780 17196
rect 2547 17156 2780 17184
rect 2547 17153 2559 17156
rect 2501 17147 2559 17153
rect 2774 17144 2780 17156
rect 2832 17144 2838 17196
rect 1578 17076 1584 17128
rect 1636 17116 1642 17128
rect 2884 17116 2912 17224
rect 5844 17221 5856 17255
rect 5890 17252 5902 17255
rect 6638 17252 6644 17264
rect 5890 17224 6644 17252
rect 5890 17221 5902 17224
rect 5844 17215 5902 17221
rect 6638 17212 6644 17224
rect 6696 17212 6702 17264
rect 10318 17252 10324 17264
rect 7024 17224 8432 17252
rect 3418 17184 3424 17196
rect 3379 17156 3424 17184
rect 3418 17144 3424 17156
rect 3476 17144 3482 17196
rect 4154 17184 4160 17196
rect 3528 17156 4160 17184
rect 1636 17088 2912 17116
rect 2961 17119 3019 17125
rect 1636 17076 1642 17088
rect 2961 17085 2973 17119
rect 3007 17116 3019 17119
rect 3528 17116 3556 17156
rect 4154 17144 4160 17156
rect 4212 17144 4218 17196
rect 4249 17187 4307 17193
rect 4249 17153 4261 17187
rect 4295 17184 4307 17187
rect 4614 17184 4620 17196
rect 4295 17156 4620 17184
rect 4295 17153 4307 17156
rect 4249 17147 4307 17153
rect 4614 17144 4620 17156
rect 4672 17184 4678 17196
rect 6178 17184 6184 17196
rect 4672 17156 6184 17184
rect 4672 17144 4678 17156
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 6270 17144 6276 17196
rect 6328 17184 6334 17196
rect 6549 17187 6607 17193
rect 6549 17184 6561 17187
rect 6328 17156 6561 17184
rect 6328 17144 6334 17156
rect 6549 17153 6561 17156
rect 6595 17153 6607 17187
rect 6549 17147 6607 17153
rect 6822 17144 6828 17196
rect 6880 17184 6886 17196
rect 6880 17156 6925 17184
rect 6880 17144 6886 17156
rect 3007 17088 3556 17116
rect 3697 17119 3755 17125
rect 3007 17085 3019 17088
rect 2961 17079 3019 17085
rect 3697 17085 3709 17119
rect 3743 17085 3755 17119
rect 4338 17116 4344 17128
rect 4299 17088 4344 17116
rect 3697 17079 3755 17085
rect 1210 17008 1216 17060
rect 1268 17048 1274 17060
rect 1857 17051 1915 17057
rect 1857 17048 1869 17051
rect 1268 17020 1869 17048
rect 1268 17008 1274 17020
rect 1857 17017 1869 17020
rect 1903 17017 1915 17051
rect 1857 17011 1915 17017
rect 2314 17008 2320 17060
rect 2372 17048 2378 17060
rect 2685 17051 2743 17057
rect 2685 17048 2697 17051
rect 2372 17020 2697 17048
rect 2372 17008 2378 17020
rect 2685 17017 2697 17020
rect 2731 17017 2743 17051
rect 3712 17048 3740 17079
rect 4338 17076 4344 17088
rect 4396 17076 4402 17128
rect 4525 17119 4583 17125
rect 4525 17085 4537 17119
rect 4571 17116 4583 17119
rect 5074 17116 5080 17128
rect 4571 17088 5080 17116
rect 4571 17085 4583 17088
rect 4525 17079 4583 17085
rect 5074 17076 5080 17088
rect 5132 17076 5138 17128
rect 6086 17116 6092 17128
rect 6047 17088 6092 17116
rect 6086 17076 6092 17088
rect 6144 17116 6150 17128
rect 6917 17119 6975 17125
rect 6917 17116 6929 17119
rect 6144 17088 6929 17116
rect 6144 17076 6150 17088
rect 6917 17085 6929 17088
rect 6963 17116 6975 17119
rect 7024 17116 7052 17224
rect 7184 17187 7242 17193
rect 7184 17153 7196 17187
rect 7230 17184 7242 17187
rect 8294 17184 8300 17196
rect 7230 17156 8300 17184
rect 7230 17153 7242 17156
rect 7184 17147 7242 17153
rect 8294 17144 8300 17156
rect 8352 17144 8358 17196
rect 8404 17193 8432 17224
rect 9876 17224 10324 17252
rect 8389 17187 8447 17193
rect 8389 17153 8401 17187
rect 8435 17153 8447 17187
rect 8645 17187 8703 17193
rect 8645 17184 8657 17187
rect 8389 17147 8447 17153
rect 8496 17156 8657 17184
rect 8496 17116 8524 17156
rect 8645 17153 8657 17156
rect 8691 17184 8703 17187
rect 9030 17184 9036 17196
rect 8691 17156 9036 17184
rect 8691 17153 8703 17156
rect 8645 17147 8703 17153
rect 9030 17144 9036 17156
rect 9088 17144 9094 17196
rect 9876 17193 9904 17224
rect 10318 17212 10324 17224
rect 10376 17212 10382 17264
rect 10428 17252 10456 17292
rect 10778 17280 10784 17332
rect 10836 17320 10842 17332
rect 11609 17323 11667 17329
rect 11609 17320 11621 17323
rect 10836 17292 11621 17320
rect 10836 17280 10842 17292
rect 11609 17289 11621 17292
rect 11655 17289 11667 17323
rect 11609 17283 11667 17289
rect 12069 17323 12127 17329
rect 12069 17289 12081 17323
rect 12115 17320 12127 17323
rect 12526 17320 12532 17332
rect 12115 17292 12532 17320
rect 12115 17289 12127 17292
rect 12069 17283 12127 17289
rect 12526 17280 12532 17292
rect 12584 17320 12590 17332
rect 12621 17323 12679 17329
rect 12621 17320 12633 17323
rect 12584 17292 12633 17320
rect 12584 17280 12590 17292
rect 12621 17289 12633 17292
rect 12667 17289 12679 17323
rect 13354 17320 13360 17332
rect 13315 17292 13360 17320
rect 12621 17283 12679 17289
rect 13354 17280 13360 17292
rect 13412 17280 13418 17332
rect 11790 17252 11796 17264
rect 10428 17224 11796 17252
rect 11790 17212 11796 17224
rect 11848 17212 11854 17264
rect 9861 17187 9919 17193
rect 9861 17153 9873 17187
rect 9907 17153 9919 17187
rect 9861 17147 9919 17153
rect 10128 17187 10186 17193
rect 10128 17153 10140 17187
rect 10174 17184 10186 17187
rect 10410 17184 10416 17196
rect 10174 17156 10416 17184
rect 10174 17153 10186 17156
rect 10128 17147 10186 17153
rect 10410 17144 10416 17156
rect 10468 17144 10474 17196
rect 11977 17187 12035 17193
rect 11977 17153 11989 17187
rect 12023 17184 12035 17187
rect 13170 17184 13176 17196
rect 12023 17156 12572 17184
rect 13131 17156 13176 17184
rect 12023 17153 12035 17156
rect 11977 17147 12035 17153
rect 12544 17125 12572 17156
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 6963 17088 7052 17116
rect 8404 17088 8524 17116
rect 12161 17119 12219 17125
rect 6963 17085 6975 17088
rect 6917 17079 6975 17085
rect 4154 17048 4160 17060
rect 2685 17011 2743 17017
rect 2884 17020 3188 17048
rect 3712 17020 4160 17048
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 2409 16983 2467 16989
rect 2409 16949 2421 16983
rect 2455 16980 2467 16983
rect 2884 16980 2912 17020
rect 2455 16952 2912 16980
rect 2455 16949 2467 16952
rect 2409 16943 2467 16949
rect 2958 16940 2964 16992
rect 3016 16980 3022 16992
rect 3053 16983 3111 16989
rect 3053 16980 3065 16983
rect 3016 16952 3065 16980
rect 3016 16940 3022 16952
rect 3053 16949 3065 16952
rect 3099 16949 3111 16983
rect 3160 16980 3188 17020
rect 4154 17008 4160 17020
rect 4212 17048 4218 17060
rect 4709 17051 4767 17057
rect 4709 17048 4721 17051
rect 4212 17020 4721 17048
rect 4212 17008 4218 17020
rect 4709 17017 4721 17020
rect 4755 17048 4767 17051
rect 4798 17048 4804 17060
rect 4755 17020 4804 17048
rect 4755 17017 4767 17020
rect 4709 17011 4767 17017
rect 4798 17008 4804 17020
rect 4856 17008 4862 17060
rect 5442 16980 5448 16992
rect 3160 16952 5448 16980
rect 3053 16943 3111 16949
rect 5442 16940 5448 16952
rect 5500 16940 5506 16992
rect 6178 16940 6184 16992
rect 6236 16980 6242 16992
rect 7098 16980 7104 16992
rect 6236 16952 7104 16980
rect 6236 16940 6242 16952
rect 7098 16940 7104 16952
rect 7156 16940 7162 16992
rect 8297 16983 8355 16989
rect 8297 16949 8309 16983
rect 8343 16980 8355 16983
rect 8404 16980 8432 17088
rect 12161 17085 12173 17119
rect 12207 17085 12219 17119
rect 12161 17079 12219 17085
rect 12529 17119 12587 17125
rect 12529 17085 12541 17119
rect 12575 17116 12587 17119
rect 14366 17116 14372 17128
rect 12575 17088 14372 17116
rect 12575 17085 12587 17088
rect 12529 17079 12587 17085
rect 9766 17048 9772 17060
rect 9727 17020 9772 17048
rect 9766 17008 9772 17020
rect 9824 17008 9830 17060
rect 11241 17051 11299 17057
rect 11241 17017 11253 17051
rect 11287 17048 11299 17051
rect 11698 17048 11704 17060
rect 11287 17020 11704 17048
rect 11287 17017 11299 17020
rect 11241 17011 11299 17017
rect 11698 17008 11704 17020
rect 11756 17048 11762 17060
rect 12176 17048 12204 17079
rect 14366 17076 14372 17088
rect 14424 17076 14430 17128
rect 11756 17020 12204 17048
rect 11756 17008 11762 17020
rect 10134 16980 10140 16992
rect 8343 16952 10140 16980
rect 8343 16949 8355 16952
rect 8297 16943 8355 16949
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 1857 16779 1915 16785
rect 1857 16776 1869 16779
rect 1728 16748 1869 16776
rect 1728 16736 1734 16748
rect 1857 16745 1869 16748
rect 1903 16745 1915 16779
rect 3234 16776 3240 16788
rect 3195 16748 3240 16776
rect 1857 16739 1915 16745
rect 3234 16736 3240 16748
rect 3292 16736 3298 16788
rect 3605 16779 3663 16785
rect 3605 16745 3617 16779
rect 3651 16776 3663 16779
rect 4154 16776 4160 16788
rect 3651 16748 4160 16776
rect 3651 16745 3663 16748
rect 3605 16739 3663 16745
rect 4154 16736 4160 16748
rect 4212 16736 4218 16788
rect 6086 16776 6092 16788
rect 5000 16748 6092 16776
rect 3418 16668 3424 16720
rect 3476 16708 3482 16720
rect 3476 16680 3832 16708
rect 3476 16668 3482 16680
rect 3804 16649 3832 16680
rect 3878 16668 3884 16720
rect 3936 16708 3942 16720
rect 4522 16708 4528 16720
rect 3936 16680 4528 16708
rect 3936 16668 3942 16680
rect 4522 16668 4528 16680
rect 4580 16708 4586 16720
rect 5000 16708 5028 16748
rect 6086 16736 6092 16748
rect 6144 16736 6150 16788
rect 7466 16736 7472 16788
rect 7524 16776 7530 16788
rect 7837 16779 7895 16785
rect 7837 16776 7849 16779
rect 7524 16748 7849 16776
rect 7524 16736 7530 16748
rect 7837 16745 7849 16748
rect 7883 16745 7895 16779
rect 7837 16739 7895 16745
rect 4580 16680 5028 16708
rect 4580 16668 4586 16680
rect 3789 16643 3847 16649
rect 1964 16612 2636 16640
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 1854 16572 1860 16584
rect 1719 16544 1860 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 1854 16532 1860 16544
rect 1912 16532 1918 16584
rect 1302 16464 1308 16516
rect 1360 16504 1366 16516
rect 1964 16504 1992 16612
rect 2041 16575 2099 16581
rect 2041 16541 2053 16575
rect 2087 16541 2099 16575
rect 2041 16535 2099 16541
rect 2317 16575 2375 16581
rect 2317 16541 2329 16575
rect 2363 16541 2375 16575
rect 2317 16535 2375 16541
rect 1360 16476 1992 16504
rect 1360 16464 1366 16476
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 2056 16436 2084 16535
rect 2332 16504 2360 16535
rect 2406 16532 2412 16584
rect 2464 16572 2470 16584
rect 2608 16572 2636 16612
rect 3789 16609 3801 16643
rect 3835 16609 3847 16643
rect 3789 16603 3847 16609
rect 4709 16643 4767 16649
rect 4709 16609 4721 16643
rect 4755 16640 4767 16643
rect 4798 16640 4804 16652
rect 4755 16612 4804 16640
rect 4755 16609 4767 16612
rect 4709 16603 4767 16609
rect 4798 16600 4804 16612
rect 4856 16600 4862 16652
rect 5000 16649 5028 16680
rect 6365 16711 6423 16717
rect 6365 16677 6377 16711
rect 6411 16677 6423 16711
rect 6365 16671 6423 16677
rect 4985 16643 5043 16649
rect 4985 16609 4997 16643
rect 5031 16609 5043 16643
rect 6380 16640 6408 16671
rect 6380 16612 6592 16640
rect 4985 16603 5043 16609
rect 2685 16575 2743 16581
rect 2685 16572 2697 16575
rect 2464 16544 2509 16572
rect 2608 16544 2697 16572
rect 2464 16532 2470 16544
rect 2685 16541 2697 16544
rect 2731 16541 2743 16575
rect 2685 16535 2743 16541
rect 2961 16575 3019 16581
rect 2961 16541 2973 16575
rect 3007 16572 3019 16575
rect 3050 16572 3056 16584
rect 3007 16544 3056 16572
rect 3007 16541 3019 16544
rect 2961 16535 3019 16541
rect 3050 16532 3056 16544
rect 3108 16532 3114 16584
rect 3421 16575 3479 16581
rect 3421 16541 3433 16575
rect 3467 16572 3479 16575
rect 3970 16572 3976 16584
rect 3467 16544 3976 16572
rect 3467 16541 3479 16544
rect 3421 16535 3479 16541
rect 3970 16532 3976 16544
rect 4028 16532 4034 16584
rect 5000 16572 5028 16603
rect 5074 16572 5080 16584
rect 5000 16544 5080 16572
rect 5074 16532 5080 16544
rect 5132 16532 5138 16584
rect 5252 16575 5310 16581
rect 5252 16541 5264 16575
rect 5298 16572 5310 16575
rect 5534 16572 5540 16584
rect 5298 16544 5540 16572
rect 5298 16541 5310 16544
rect 5252 16535 5310 16541
rect 5534 16532 5540 16544
rect 5592 16532 5598 16584
rect 6086 16532 6092 16584
rect 6144 16572 6150 16584
rect 6457 16575 6515 16581
rect 6457 16572 6469 16575
rect 6144 16544 6469 16572
rect 6144 16532 6150 16544
rect 6457 16541 6469 16544
rect 6503 16541 6515 16575
rect 6564 16572 6592 16612
rect 6724 16575 6782 16581
rect 6724 16572 6736 16575
rect 6564 16544 6736 16572
rect 6457 16535 6515 16541
rect 6724 16541 6736 16544
rect 6770 16572 6782 16575
rect 7006 16572 7012 16584
rect 6770 16544 7012 16572
rect 6770 16541 6782 16544
rect 6724 16535 6782 16541
rect 7006 16532 7012 16544
rect 7064 16532 7070 16584
rect 7852 16572 7880 16739
rect 8570 16736 8576 16788
rect 8628 16776 8634 16788
rect 8941 16779 8999 16785
rect 8941 16776 8953 16779
rect 8628 16748 8953 16776
rect 8628 16736 8634 16748
rect 8941 16745 8953 16748
rect 8987 16745 8999 16779
rect 8941 16739 8999 16745
rect 9122 16736 9128 16788
rect 9180 16776 9186 16788
rect 9217 16779 9275 16785
rect 9217 16776 9229 16779
rect 9180 16748 9229 16776
rect 9180 16736 9186 16748
rect 9217 16745 9229 16748
rect 9263 16745 9275 16779
rect 9217 16739 9275 16745
rect 10520 16748 11100 16776
rect 8386 16668 8392 16720
rect 8444 16708 8450 16720
rect 9401 16711 9459 16717
rect 9401 16708 9413 16711
rect 8444 16680 9413 16708
rect 8444 16668 8450 16680
rect 9401 16677 9413 16680
rect 9447 16677 9459 16711
rect 9401 16671 9459 16677
rect 8478 16600 8484 16652
rect 8536 16640 8542 16652
rect 8754 16640 8760 16652
rect 8536 16612 8760 16640
rect 8536 16600 8542 16612
rect 8754 16600 8760 16612
rect 8812 16600 8818 16652
rect 10134 16640 10140 16652
rect 10095 16612 10140 16640
rect 10134 16600 10140 16612
rect 10192 16600 10198 16652
rect 10520 16640 10548 16748
rect 11072 16708 11100 16748
rect 11146 16736 11152 16788
rect 11204 16776 11210 16788
rect 11241 16779 11299 16785
rect 11241 16776 11253 16779
rect 11204 16748 11253 16776
rect 11204 16736 11210 16748
rect 11241 16745 11253 16748
rect 11287 16745 11299 16779
rect 11241 16739 11299 16745
rect 11882 16736 11888 16788
rect 11940 16776 11946 16788
rect 12253 16779 12311 16785
rect 12253 16776 12265 16779
rect 11940 16748 12265 16776
rect 11940 16736 11946 16748
rect 12253 16745 12265 16748
rect 12299 16776 12311 16779
rect 12299 16748 12434 16776
rect 12299 16745 12311 16748
rect 12253 16739 12311 16745
rect 11900 16708 11928 16736
rect 11072 16680 11928 16708
rect 12406 16708 12434 16748
rect 13170 16736 13176 16788
rect 13228 16776 13234 16788
rect 13541 16779 13599 16785
rect 13541 16776 13553 16779
rect 13228 16748 13553 16776
rect 13228 16736 13234 16748
rect 13541 16745 13553 16748
rect 13587 16745 13599 16779
rect 13541 16739 13599 16745
rect 14458 16708 14464 16720
rect 12406 16680 14464 16708
rect 14458 16668 14464 16680
rect 14516 16668 14522 16720
rect 10244 16612 10548 16640
rect 10597 16643 10655 16649
rect 7929 16575 7987 16581
rect 7929 16572 7941 16575
rect 7852 16544 7941 16572
rect 7929 16541 7941 16544
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 8294 16532 8300 16584
rect 8352 16572 8358 16584
rect 8573 16575 8631 16581
rect 8573 16572 8585 16575
rect 8352 16544 8585 16572
rect 8352 16532 8358 16544
rect 8573 16541 8585 16544
rect 8619 16541 8631 16575
rect 8573 16535 8631 16541
rect 10045 16575 10103 16581
rect 10045 16541 10057 16575
rect 10091 16572 10103 16575
rect 10244 16572 10272 16612
rect 10597 16609 10609 16643
rect 10643 16609 10655 16643
rect 10597 16603 10655 16609
rect 10689 16643 10747 16649
rect 10689 16609 10701 16643
rect 10735 16640 10747 16643
rect 11238 16640 11244 16652
rect 10735 16612 11244 16640
rect 10735 16609 10747 16612
rect 10689 16603 10747 16609
rect 10091 16544 10272 16572
rect 10612 16572 10640 16603
rect 11238 16600 11244 16612
rect 11296 16600 11302 16652
rect 11698 16600 11704 16652
rect 11756 16640 11762 16652
rect 11793 16643 11851 16649
rect 11793 16640 11805 16643
rect 11756 16612 11805 16640
rect 11756 16600 11762 16612
rect 11793 16609 11805 16612
rect 11839 16609 11851 16643
rect 11793 16603 11851 16609
rect 12989 16643 13047 16649
rect 12989 16609 13001 16643
rect 13035 16640 13047 16643
rect 13814 16640 13820 16652
rect 13035 16612 13820 16640
rect 13035 16609 13047 16612
rect 12989 16603 13047 16609
rect 13814 16600 13820 16612
rect 13872 16640 13878 16652
rect 13872 16612 14136 16640
rect 13872 16600 13878 16612
rect 11054 16572 11060 16584
rect 10612 16544 11060 16572
rect 10091 16541 10103 16544
rect 10045 16535 10103 16541
rect 11054 16532 11060 16544
rect 11112 16532 11118 16584
rect 14108 16581 14136 16612
rect 14093 16575 14151 16581
rect 14093 16541 14105 16575
rect 14139 16574 14151 16575
rect 14139 16546 14173 16574
rect 14139 16541 14151 16546
rect 14093 16535 14151 16541
rect 4525 16507 4583 16513
rect 2332 16476 4108 16504
rect 2133 16439 2191 16445
rect 2133 16436 2145 16439
rect 2056 16408 2145 16436
rect 2133 16405 2145 16408
rect 2179 16405 2191 16439
rect 2133 16399 2191 16405
rect 2593 16439 2651 16445
rect 2593 16405 2605 16439
rect 2639 16436 2651 16439
rect 2682 16436 2688 16448
rect 2639 16408 2688 16436
rect 2639 16405 2651 16408
rect 2593 16399 2651 16405
rect 2682 16396 2688 16408
rect 2740 16396 2746 16448
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 2869 16439 2927 16445
rect 2869 16436 2881 16439
rect 2832 16408 2881 16436
rect 2832 16396 2838 16408
rect 2869 16405 2881 16408
rect 2915 16405 2927 16439
rect 2869 16399 2927 16405
rect 3145 16439 3203 16445
rect 3145 16405 3157 16439
rect 3191 16436 3203 16439
rect 3970 16436 3976 16448
rect 3191 16408 3976 16436
rect 3191 16405 3203 16408
rect 3145 16399 3203 16405
rect 3970 16396 3976 16408
rect 4028 16396 4034 16448
rect 4080 16445 4108 16476
rect 4525 16473 4537 16507
rect 4571 16473 4583 16507
rect 4525 16467 4583 16473
rect 4065 16439 4123 16445
rect 4065 16405 4077 16439
rect 4111 16405 4123 16439
rect 4430 16436 4436 16448
rect 4391 16408 4436 16436
rect 4065 16399 4123 16405
rect 4430 16396 4436 16408
rect 4488 16396 4494 16448
rect 4540 16436 4568 16467
rect 6822 16464 6828 16516
rect 6880 16504 6886 16516
rect 10134 16504 10140 16516
rect 6880 16476 10140 16504
rect 6880 16464 6886 16476
rect 10134 16464 10140 16476
rect 10192 16464 10198 16516
rect 11609 16507 11667 16513
rect 11609 16473 11621 16507
rect 11655 16504 11667 16507
rect 12618 16504 12624 16516
rect 11655 16476 12624 16504
rect 11655 16473 11667 16476
rect 11609 16467 11667 16473
rect 12618 16464 12624 16476
rect 12676 16464 12682 16516
rect 8202 16436 8208 16448
rect 4540 16408 8208 16436
rect 8202 16396 8208 16408
rect 8260 16396 8266 16448
rect 9490 16396 9496 16448
rect 9548 16436 9554 16448
rect 9585 16439 9643 16445
rect 9585 16436 9597 16439
rect 9548 16408 9597 16436
rect 9548 16396 9554 16408
rect 9585 16405 9597 16408
rect 9631 16405 9643 16439
rect 9950 16436 9956 16448
rect 9911 16408 9956 16436
rect 9585 16399 9643 16405
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 10778 16396 10784 16448
rect 10836 16436 10842 16448
rect 11146 16436 11152 16448
rect 10836 16408 10881 16436
rect 11107 16408 11152 16436
rect 10836 16396 10842 16408
rect 11146 16396 11152 16408
rect 11204 16396 11210 16448
rect 11701 16439 11759 16445
rect 11701 16405 11713 16439
rect 11747 16436 11759 16439
rect 11790 16436 11796 16448
rect 11747 16408 11796 16436
rect 11747 16405 11759 16408
rect 11701 16399 11759 16405
rect 11790 16396 11796 16408
rect 11848 16436 11854 16448
rect 12069 16439 12127 16445
rect 12069 16436 12081 16439
rect 11848 16408 12081 16436
rect 11848 16396 11854 16408
rect 12069 16405 12081 16408
rect 12115 16405 12127 16439
rect 13078 16436 13084 16448
rect 13039 16408 13084 16436
rect 12069 16399 12127 16405
rect 13078 16396 13084 16408
rect 13136 16396 13142 16448
rect 13173 16439 13231 16445
rect 13173 16405 13185 16439
rect 13219 16436 13231 16439
rect 13538 16436 13544 16448
rect 13219 16408 13544 16436
rect 13219 16405 13231 16408
rect 13173 16399 13231 16405
rect 13538 16396 13544 16408
rect 13596 16396 13602 16448
rect 14734 16436 14740 16448
rect 14695 16408 14740 16436
rect 14734 16396 14740 16408
rect 14792 16396 14798 16448
rect 1104 16346 21896 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21896 16346
rect 1104 16272 21896 16294
rect 1854 16232 1860 16244
rect 1815 16204 1860 16232
rect 1854 16192 1860 16204
rect 1912 16192 1918 16244
rect 2038 16192 2044 16244
rect 2096 16232 2102 16244
rect 2409 16235 2467 16241
rect 2409 16232 2421 16235
rect 2096 16204 2421 16232
rect 2096 16192 2102 16204
rect 2409 16201 2421 16204
rect 2455 16201 2467 16235
rect 2866 16232 2872 16244
rect 2827 16204 2872 16232
rect 2409 16195 2467 16201
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 4798 16192 4804 16244
rect 4856 16232 4862 16244
rect 5258 16232 5264 16244
rect 4856 16204 5264 16232
rect 4856 16192 4862 16204
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 6825 16235 6883 16241
rect 6825 16201 6837 16235
rect 6871 16232 6883 16235
rect 7377 16235 7435 16241
rect 7377 16232 7389 16235
rect 6871 16204 7389 16232
rect 6871 16201 6883 16204
rect 6825 16195 6883 16201
rect 7377 16201 7389 16204
rect 7423 16201 7435 16235
rect 8202 16232 8208 16244
rect 8163 16204 8208 16232
rect 7377 16195 7435 16201
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 9490 16232 9496 16244
rect 9451 16204 9496 16232
rect 9490 16192 9496 16204
rect 9548 16192 9554 16244
rect 9953 16235 10011 16241
rect 9953 16201 9965 16235
rect 9999 16232 10011 16235
rect 10042 16232 10048 16244
rect 9999 16204 10048 16232
rect 9999 16201 10011 16204
rect 9953 16195 10011 16201
rect 1946 16124 1952 16176
rect 2004 16164 2010 16176
rect 2004 16136 2636 16164
rect 2004 16124 2010 16136
rect 1670 16096 1676 16108
rect 1631 16068 1676 16096
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 2041 16099 2099 16105
rect 2041 16065 2053 16099
rect 2087 16096 2099 16099
rect 2130 16096 2136 16108
rect 2087 16068 2136 16096
rect 2087 16065 2099 16068
rect 2041 16059 2099 16065
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 2314 16096 2320 16108
rect 2275 16068 2320 16096
rect 2314 16056 2320 16068
rect 2372 16056 2378 16108
rect 2608 16105 2636 16136
rect 2774 16124 2780 16176
rect 2832 16164 2838 16176
rect 5626 16164 5632 16176
rect 2832 16136 5632 16164
rect 2832 16124 2838 16136
rect 5626 16124 5632 16136
rect 5684 16124 5690 16176
rect 6546 16124 6552 16176
rect 6604 16164 6610 16176
rect 8294 16164 8300 16176
rect 6604 16136 8300 16164
rect 6604 16124 6610 16136
rect 8294 16124 8300 16136
rect 8352 16124 8358 16176
rect 9398 16164 9404 16176
rect 9359 16136 9404 16164
rect 9398 16124 9404 16136
rect 9456 16124 9462 16176
rect 2593 16099 2651 16105
rect 2593 16065 2605 16099
rect 2639 16065 2651 16099
rect 2593 16059 2651 16065
rect 2682 16056 2688 16108
rect 2740 16096 2746 16108
rect 2740 16068 2785 16096
rect 2740 16056 2746 16068
rect 2866 16056 2872 16108
rect 2924 16096 2930 16108
rect 2961 16099 3019 16105
rect 2961 16096 2973 16099
rect 2924 16068 2973 16096
rect 2924 16056 2930 16068
rect 2961 16065 2973 16068
rect 3007 16065 3019 16099
rect 3418 16096 3424 16108
rect 3379 16068 3424 16096
rect 2961 16059 3019 16065
rect 2976 16028 3004 16059
rect 3418 16056 3424 16068
rect 3476 16056 3482 16108
rect 3878 16096 3884 16108
rect 3839 16068 3884 16096
rect 3878 16056 3884 16068
rect 3936 16056 3942 16108
rect 4154 16105 4160 16108
rect 4148 16096 4160 16105
rect 4067 16068 4160 16096
rect 4148 16059 4160 16068
rect 4212 16096 4218 16108
rect 4212 16068 5396 16096
rect 4154 16056 4160 16059
rect 4212 16056 4218 16068
rect 3326 16028 3332 16040
rect 2976 16000 3332 16028
rect 3326 15988 3332 16000
rect 3384 15988 3390 16040
rect 3789 16031 3847 16037
rect 3789 15997 3801 16031
rect 3835 15997 3847 16031
rect 5368 16028 5396 16068
rect 5442 16056 5448 16108
rect 5500 16096 5506 16108
rect 6730 16096 6736 16108
rect 5500 16068 5545 16096
rect 6691 16068 6736 16096
rect 5500 16056 5506 16068
rect 6730 16056 6736 16068
rect 6788 16056 6794 16108
rect 7006 16056 7012 16108
rect 7064 16096 7070 16108
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 7064 16068 7205 16096
rect 7064 16056 7070 16068
rect 7193 16065 7205 16068
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 7745 16099 7803 16105
rect 7745 16065 7757 16099
rect 7791 16096 7803 16099
rect 8202 16096 8208 16108
rect 7791 16068 8208 16096
rect 7791 16065 7803 16068
rect 7745 16059 7803 16065
rect 8202 16056 8208 16068
rect 8260 16056 8266 16108
rect 8570 16096 8576 16108
rect 8531 16068 8576 16096
rect 8570 16056 8576 16068
rect 8628 16056 8634 16108
rect 9968 16096 9996 16195
rect 10042 16192 10048 16204
rect 10100 16192 10106 16244
rect 10134 16192 10140 16244
rect 10192 16232 10198 16244
rect 10192 16204 10237 16232
rect 10192 16192 10198 16204
rect 11146 16192 11152 16244
rect 11204 16232 11210 16244
rect 11793 16235 11851 16241
rect 11793 16232 11805 16235
rect 11204 16204 11805 16232
rect 11204 16192 11210 16204
rect 11793 16201 11805 16204
rect 11839 16201 11851 16235
rect 11793 16195 11851 16201
rect 12253 16235 12311 16241
rect 12253 16201 12265 16235
rect 12299 16232 12311 16235
rect 13078 16232 13084 16244
rect 12299 16204 13084 16232
rect 12299 16201 12311 16204
rect 12253 16195 12311 16201
rect 13078 16192 13084 16204
rect 13136 16192 13142 16244
rect 13814 16232 13820 16244
rect 13775 16204 13820 16232
rect 13814 16192 13820 16204
rect 13872 16192 13878 16244
rect 10318 16124 10324 16176
rect 10376 16164 10382 16176
rect 17402 16164 17408 16176
rect 10376 16136 17408 16164
rect 10376 16124 10382 16136
rect 17402 16124 17408 16136
rect 17460 16124 17466 16176
rect 11882 16096 11888 16108
rect 8680 16068 9996 16096
rect 11843 16068 11888 16096
rect 5368 16000 6500 16028
rect 3789 15991 3847 15997
rect 1486 15960 1492 15972
rect 1447 15932 1492 15960
rect 1486 15920 1492 15932
rect 1544 15920 1550 15972
rect 1762 15920 1768 15972
rect 1820 15960 1826 15972
rect 2133 15963 2191 15969
rect 2133 15960 2145 15963
rect 1820 15932 2145 15960
rect 1820 15920 1826 15932
rect 2133 15929 2145 15932
rect 2179 15929 2191 15963
rect 2133 15923 2191 15929
rect 2222 15920 2228 15972
rect 2280 15960 2286 15972
rect 3237 15963 3295 15969
rect 3237 15960 3249 15963
rect 2280 15932 3249 15960
rect 2280 15920 2286 15932
rect 3237 15929 3249 15932
rect 3283 15929 3295 15963
rect 3804 15960 3832 15991
rect 3878 15960 3884 15972
rect 3804 15932 3884 15960
rect 3237 15923 3295 15929
rect 3878 15920 3884 15932
rect 3936 15920 3942 15972
rect 6365 15963 6423 15969
rect 6365 15960 6377 15963
rect 4816 15932 6377 15960
rect 3142 15892 3148 15904
rect 3103 15864 3148 15892
rect 3142 15852 3148 15864
rect 3200 15852 3206 15904
rect 3326 15852 3332 15904
rect 3384 15892 3390 15904
rect 4816 15892 4844 15932
rect 6365 15929 6377 15932
rect 6411 15929 6423 15963
rect 6472 15960 6500 16000
rect 6546 15988 6552 16040
rect 6604 16028 6610 16040
rect 6917 16031 6975 16037
rect 6917 16028 6929 16031
rect 6604 16000 6929 16028
rect 6604 15988 6610 16000
rect 6917 15997 6929 16000
rect 6963 15997 6975 16031
rect 7834 16028 7840 16040
rect 7795 16000 7840 16028
rect 6917 15991 6975 15997
rect 7834 15988 7840 16000
rect 7892 15988 7898 16040
rect 7926 15988 7932 16040
rect 7984 16028 7990 16040
rect 7984 16000 8029 16028
rect 7984 15988 7990 16000
rect 8386 15988 8392 16040
rect 8444 16028 8450 16040
rect 8680 16037 8708 16068
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 12693 16099 12751 16105
rect 12693 16096 12705 16099
rect 11992 16068 12705 16096
rect 8665 16031 8723 16037
rect 8665 16028 8677 16031
rect 8444 16000 8677 16028
rect 8444 15988 8450 16000
rect 8665 15997 8677 16000
rect 8711 15997 8723 16031
rect 8665 15991 8723 15997
rect 8757 16031 8815 16037
rect 8757 15997 8769 16031
rect 8803 15997 8815 16031
rect 8757 15991 8815 15997
rect 9585 16031 9643 16037
rect 9585 15997 9597 16031
rect 9631 16028 9643 16031
rect 9766 16028 9772 16040
rect 9631 16000 9772 16028
rect 9631 15997 9643 16000
rect 9585 15991 9643 15997
rect 8478 15960 8484 15972
rect 6472 15932 8484 15960
rect 6365 15923 6423 15929
rect 8478 15920 8484 15932
rect 8536 15960 8542 15972
rect 8772 15960 8800 15991
rect 9766 15988 9772 16000
rect 9824 15988 9830 16040
rect 10134 15988 10140 16040
rect 10192 16028 10198 16040
rect 10965 16031 11023 16037
rect 10965 16028 10977 16031
rect 10192 16000 10977 16028
rect 10192 15988 10198 16000
rect 10965 15997 10977 16000
rect 11011 15997 11023 16031
rect 10965 15991 11023 15997
rect 11146 15988 11152 16040
rect 11204 16028 11210 16040
rect 11241 16031 11299 16037
rect 11241 16028 11253 16031
rect 11204 16000 11253 16028
rect 11204 15988 11210 16000
rect 11241 15997 11253 16000
rect 11287 15997 11299 16031
rect 11241 15991 11299 15997
rect 11701 16031 11759 16037
rect 11701 15997 11713 16031
rect 11747 15997 11759 16031
rect 11701 15991 11759 15997
rect 8536 15932 8800 15960
rect 8536 15920 8542 15932
rect 9950 15920 9956 15972
rect 10008 15960 10014 15972
rect 11716 15960 11744 15991
rect 11992 15960 12020 16068
rect 12693 16065 12705 16068
rect 12739 16096 12751 16099
rect 12986 16096 12992 16108
rect 12739 16068 12992 16096
rect 12739 16065 12751 16068
rect 12693 16059 12751 16065
rect 12986 16056 12992 16068
rect 13044 16056 13050 16108
rect 12437 16031 12495 16037
rect 12437 15997 12449 16031
rect 12483 15997 12495 16031
rect 12437 15991 12495 15997
rect 10008 15932 10364 15960
rect 11716 15932 12020 15960
rect 10008 15920 10014 15932
rect 3384 15864 4844 15892
rect 3384 15852 3390 15864
rect 5810 15852 5816 15904
rect 5868 15892 5874 15904
rect 6089 15895 6147 15901
rect 6089 15892 6101 15895
rect 5868 15864 6101 15892
rect 5868 15852 5874 15864
rect 6089 15861 6101 15864
rect 6135 15861 6147 15895
rect 6089 15855 6147 15861
rect 7466 15852 7472 15904
rect 7524 15892 7530 15904
rect 10336 15901 10364 15932
rect 12342 15920 12348 15972
rect 12400 15960 12406 15972
rect 12452 15960 12480 15991
rect 12400 15932 12480 15960
rect 12400 15920 12406 15932
rect 9033 15895 9091 15901
rect 9033 15892 9045 15895
rect 7524 15864 9045 15892
rect 7524 15852 7530 15864
rect 9033 15861 9045 15864
rect 9079 15861 9091 15895
rect 9033 15855 9091 15861
rect 10321 15895 10379 15901
rect 10321 15861 10333 15895
rect 10367 15892 10379 15895
rect 15746 15892 15752 15904
rect 10367 15864 15752 15892
rect 10367 15861 10379 15864
rect 10321 15855 10379 15861
rect 15746 15852 15752 15864
rect 15804 15852 15810 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 2130 15688 2136 15700
rect 2091 15660 2136 15688
rect 2130 15648 2136 15660
rect 2188 15648 2194 15700
rect 2314 15648 2320 15700
rect 2372 15688 2378 15700
rect 2685 15691 2743 15697
rect 2685 15688 2697 15691
rect 2372 15660 2697 15688
rect 2372 15648 2378 15660
rect 2685 15657 2697 15660
rect 2731 15657 2743 15691
rect 3418 15688 3424 15700
rect 3379 15660 3424 15688
rect 2685 15651 2743 15657
rect 3418 15648 3424 15660
rect 3476 15648 3482 15700
rect 3881 15691 3939 15697
rect 3881 15657 3893 15691
rect 3927 15688 3939 15691
rect 4246 15688 4252 15700
rect 3927 15660 4252 15688
rect 3927 15657 3939 15660
rect 3881 15651 3939 15657
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 4430 15648 4436 15700
rect 4488 15688 4494 15700
rect 4709 15691 4767 15697
rect 4709 15688 4721 15691
rect 4488 15660 4721 15688
rect 4488 15648 4494 15660
rect 4709 15657 4721 15660
rect 4755 15657 4767 15691
rect 4709 15651 4767 15657
rect 5074 15648 5080 15700
rect 5132 15688 5138 15700
rect 5534 15688 5540 15700
rect 5132 15660 5540 15688
rect 5132 15648 5138 15660
rect 5534 15648 5540 15660
rect 5592 15648 5598 15700
rect 8478 15688 8484 15700
rect 5828 15660 8064 15688
rect 8439 15660 8484 15688
rect 1670 15580 1676 15632
rect 1728 15620 1734 15632
rect 2409 15623 2467 15629
rect 2409 15620 2421 15623
rect 1728 15592 2421 15620
rect 1728 15580 1734 15592
rect 2409 15589 2421 15592
rect 2455 15589 2467 15623
rect 2409 15583 2467 15589
rect 2590 15580 2596 15632
rect 2648 15620 2654 15632
rect 2961 15623 3019 15629
rect 2961 15620 2973 15623
rect 2648 15592 2973 15620
rect 2648 15580 2654 15592
rect 2961 15589 2973 15592
rect 3007 15589 3019 15623
rect 2961 15583 3019 15589
rect 3326 15552 3332 15564
rect 2884 15524 3332 15552
rect 1670 15484 1676 15496
rect 1631 15456 1676 15484
rect 1670 15444 1676 15456
rect 1728 15444 1734 15496
rect 2038 15484 2044 15496
rect 1999 15456 2044 15484
rect 2038 15444 2044 15456
rect 2096 15444 2102 15496
rect 2317 15487 2375 15493
rect 2317 15453 2329 15487
rect 2363 15484 2375 15487
rect 2406 15484 2412 15496
rect 2363 15456 2412 15484
rect 2363 15453 2375 15456
rect 2317 15447 2375 15453
rect 2406 15444 2412 15456
rect 2464 15444 2470 15496
rect 2590 15484 2596 15496
rect 2551 15456 2596 15484
rect 2590 15444 2596 15456
rect 2648 15444 2654 15496
rect 2884 15493 2912 15524
rect 3326 15512 3332 15524
rect 3384 15512 3390 15564
rect 3510 15552 3516 15564
rect 3471 15524 3516 15552
rect 3510 15512 3516 15524
rect 3568 15512 3574 15564
rect 4154 15552 4160 15564
rect 4115 15524 4160 15552
rect 4154 15512 4160 15524
rect 4212 15512 4218 15564
rect 4264 15552 4292 15648
rect 4338 15580 4344 15632
rect 4396 15620 4402 15632
rect 4893 15623 4951 15629
rect 4893 15620 4905 15623
rect 4396 15592 4905 15620
rect 4396 15580 4402 15592
rect 4893 15589 4905 15592
rect 4939 15589 4951 15623
rect 4893 15583 4951 15589
rect 4982 15580 4988 15632
rect 5040 15620 5046 15632
rect 5828 15620 5856 15660
rect 5040 15592 5856 15620
rect 8036 15620 8064 15660
rect 8478 15648 8484 15660
rect 8536 15648 8542 15700
rect 13538 15688 13544 15700
rect 13499 15660 13544 15688
rect 13538 15648 13544 15660
rect 13596 15648 13602 15700
rect 9217 15623 9275 15629
rect 9217 15620 9229 15623
rect 8036 15592 9229 15620
rect 5040 15580 5046 15592
rect 9217 15589 9229 15592
rect 9263 15589 9275 15623
rect 9217 15583 9275 15589
rect 4264 15524 5120 15552
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15453 2927 15487
rect 3142 15484 3148 15496
rect 3103 15456 3148 15484
rect 2869 15447 2927 15453
rect 3142 15444 3148 15456
rect 3200 15444 3206 15496
rect 3237 15487 3295 15493
rect 3237 15453 3249 15487
rect 3283 15453 3295 15487
rect 3237 15447 3295 15453
rect 1394 15376 1400 15428
rect 1452 15416 1458 15428
rect 3050 15416 3056 15428
rect 1452 15388 3056 15416
rect 1452 15376 1458 15388
rect 3050 15376 3056 15388
rect 3108 15376 3114 15428
rect 3252 15416 3280 15447
rect 3878 15444 3884 15496
rect 3936 15484 3942 15496
rect 5092 15493 5120 15524
rect 5534 15512 5540 15564
rect 5592 15552 5598 15564
rect 7101 15555 7159 15561
rect 7101 15552 7113 15555
rect 5592 15524 7113 15552
rect 5592 15512 5598 15524
rect 7101 15521 7113 15524
rect 7147 15521 7159 15555
rect 7101 15515 7159 15521
rect 4341 15487 4399 15493
rect 4341 15484 4353 15487
rect 3936 15456 4353 15484
rect 3936 15444 3942 15456
rect 4341 15453 4353 15456
rect 4387 15453 4399 15487
rect 4341 15447 4399 15453
rect 5077 15487 5135 15493
rect 5077 15453 5089 15487
rect 5123 15453 5135 15487
rect 7116 15484 7144 15515
rect 8294 15512 8300 15564
rect 8352 15552 8358 15564
rect 9401 15555 9459 15561
rect 9401 15552 9413 15555
rect 8352 15524 9413 15552
rect 8352 15512 8358 15524
rect 9401 15521 9413 15524
rect 9447 15521 9459 15555
rect 9401 15515 9459 15521
rect 12161 15555 12219 15561
rect 12161 15521 12173 15555
rect 12207 15552 12219 15555
rect 12342 15552 12348 15564
rect 12207 15524 12348 15552
rect 12207 15521 12219 15524
rect 12161 15515 12219 15521
rect 12342 15512 12348 15524
rect 12400 15552 12406 15564
rect 12986 15552 12992 15564
rect 12400 15512 12434 15552
rect 12947 15524 12992 15552
rect 12986 15512 12992 15524
rect 13044 15512 13050 15564
rect 7742 15484 7748 15496
rect 7116 15456 7748 15484
rect 5077 15447 5135 15453
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 8202 15444 8208 15496
rect 8260 15484 8266 15496
rect 8665 15487 8723 15493
rect 8665 15484 8677 15487
rect 8260 15456 8677 15484
rect 8260 15444 8266 15456
rect 8665 15453 8677 15456
rect 8711 15484 8723 15487
rect 11698 15484 11704 15496
rect 8711 15456 11704 15484
rect 8711 15453 8723 15456
rect 8665 15447 8723 15453
rect 11698 15444 11704 15456
rect 11756 15444 11762 15496
rect 12406 15484 12434 15512
rect 14093 15487 14151 15493
rect 14093 15484 14105 15487
rect 12406 15456 14105 15484
rect 14093 15453 14105 15456
rect 14139 15453 14151 15487
rect 14093 15447 14151 15453
rect 14360 15487 14418 15493
rect 14360 15453 14372 15487
rect 14406 15484 14418 15487
rect 14734 15484 14740 15496
rect 14406 15456 14740 15484
rect 14406 15453 14418 15456
rect 14360 15447 14418 15453
rect 14734 15444 14740 15456
rect 14792 15444 14798 15496
rect 16206 15484 16212 15496
rect 15488 15456 16212 15484
rect 4062 15416 4068 15428
rect 3252 15388 4068 15416
rect 4062 15376 4068 15388
rect 4120 15376 4126 15428
rect 6822 15416 6828 15428
rect 4172 15388 6828 15416
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 1854 15348 1860 15360
rect 1815 15320 1860 15348
rect 1854 15308 1860 15320
rect 1912 15308 1918 15360
rect 3970 15308 3976 15360
rect 4028 15348 4034 15360
rect 4172 15348 4200 15388
rect 6822 15376 6828 15388
rect 6880 15376 6886 15428
rect 7006 15416 7012 15428
rect 6967 15388 7012 15416
rect 7006 15376 7012 15388
rect 7064 15376 7070 15428
rect 7098 15376 7104 15428
rect 7156 15416 7162 15428
rect 7346 15419 7404 15425
rect 7346 15416 7358 15419
rect 7156 15388 7358 15416
rect 7156 15376 7162 15388
rect 7346 15385 7358 15388
rect 7392 15385 7404 15419
rect 10410 15416 10416 15428
rect 10371 15388 10416 15416
rect 7346 15379 7404 15385
rect 10410 15376 10416 15388
rect 10468 15376 10474 15428
rect 13081 15419 13139 15425
rect 13081 15385 13093 15419
rect 13127 15416 13139 15419
rect 13814 15416 13820 15428
rect 13127 15388 13820 15416
rect 13127 15385 13139 15388
rect 13081 15379 13139 15385
rect 13814 15376 13820 15388
rect 13872 15376 13878 15428
rect 4028 15320 4200 15348
rect 4028 15308 4034 15320
rect 4246 15308 4252 15360
rect 4304 15348 4310 15360
rect 4304 15320 4349 15348
rect 4304 15308 4310 15320
rect 5994 15308 6000 15360
rect 6052 15348 6058 15360
rect 7466 15348 7472 15360
rect 6052 15320 7472 15348
rect 6052 15308 6058 15320
rect 7466 15308 7472 15320
rect 7524 15308 7530 15360
rect 8570 15308 8576 15360
rect 8628 15348 8634 15360
rect 9125 15351 9183 15357
rect 9125 15348 9137 15351
rect 8628 15320 9137 15348
rect 8628 15308 8634 15320
rect 9125 15317 9137 15320
rect 9171 15348 9183 15351
rect 12250 15348 12256 15360
rect 9171 15320 12256 15348
rect 9171 15317 9183 15320
rect 9125 15311 9183 15317
rect 12250 15308 12256 15320
rect 12308 15308 12314 15360
rect 13170 15308 13176 15360
rect 13228 15348 13234 15360
rect 15488 15357 15516 15456
rect 16206 15444 16212 15456
rect 16264 15444 16270 15496
rect 15473 15351 15531 15357
rect 13228 15320 13273 15348
rect 13228 15308 13234 15320
rect 15473 15317 15485 15351
rect 15519 15317 15531 15351
rect 15473 15311 15531 15317
rect 15565 15351 15623 15357
rect 15565 15317 15577 15351
rect 15611 15348 15623 15351
rect 15654 15348 15660 15360
rect 15611 15320 15660 15348
rect 15611 15317 15623 15320
rect 15565 15311 15623 15317
rect 15654 15308 15660 15320
rect 15712 15308 15718 15360
rect 1104 15258 21896 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21896 15258
rect 1104 15184 21896 15206
rect 1670 15104 1676 15156
rect 1728 15144 1734 15156
rect 1857 15147 1915 15153
rect 1857 15144 1869 15147
rect 1728 15116 1869 15144
rect 1728 15104 1734 15116
rect 1857 15113 1869 15116
rect 1903 15113 1915 15147
rect 1857 15107 1915 15113
rect 2317 15147 2375 15153
rect 2317 15113 2329 15147
rect 2363 15144 2375 15147
rect 2590 15144 2596 15156
rect 2363 15116 2596 15144
rect 2363 15113 2375 15116
rect 2317 15107 2375 15113
rect 2590 15104 2596 15116
rect 2648 15104 2654 15156
rect 3142 15144 3148 15156
rect 3103 15116 3148 15144
rect 3142 15104 3148 15116
rect 3200 15104 3206 15156
rect 3237 15147 3295 15153
rect 3237 15113 3249 15147
rect 3283 15113 3295 15147
rect 5994 15144 6000 15156
rect 3237 15107 3295 15113
rect 3344 15116 6000 15144
rect 2406 15036 2412 15088
rect 2464 15076 2470 15088
rect 3252 15076 3280 15107
rect 2464 15048 3280 15076
rect 2464 15036 2470 15048
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 1854 15008 1860 15020
rect 1719 14980 1860 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 1854 14968 1860 14980
rect 1912 14968 1918 15020
rect 1946 14968 1952 15020
rect 2004 15008 2010 15020
rect 2041 15011 2099 15017
rect 2041 15008 2053 15011
rect 2004 14980 2053 15008
rect 2004 14968 2010 14980
rect 2041 14977 2053 14980
rect 2087 14977 2099 15011
rect 2041 14971 2099 14977
rect 2133 15011 2191 15017
rect 2133 14977 2145 15011
rect 2179 15008 2191 15011
rect 2222 15008 2228 15020
rect 2179 14980 2228 15008
rect 2179 14977 2191 14980
rect 2133 14971 2191 14977
rect 2222 14968 2228 14980
rect 2280 14968 2286 15020
rect 2593 15011 2651 15017
rect 2593 14977 2605 15011
rect 2639 14977 2651 15011
rect 2593 14971 2651 14977
rect 2685 15011 2743 15017
rect 2685 14977 2697 15011
rect 2731 14977 2743 15011
rect 2685 14971 2743 14977
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 15008 3019 15011
rect 3344 15008 3372 15116
rect 5994 15104 6000 15116
rect 6052 15104 6058 15156
rect 6365 15147 6423 15153
rect 6365 15113 6377 15147
rect 6411 15144 6423 15147
rect 6546 15144 6552 15156
rect 6411 15116 6552 15144
rect 6411 15113 6423 15116
rect 6365 15107 6423 15113
rect 3418 15036 3424 15088
rect 3476 15076 3482 15088
rect 4310 15079 4368 15085
rect 4310 15076 4322 15079
rect 3476 15048 4322 15076
rect 3476 15036 3482 15048
rect 4310 15045 4322 15048
rect 4356 15045 4368 15079
rect 4310 15039 4368 15045
rect 3007 14980 3372 15008
rect 3605 15011 3663 15017
rect 3007 14977 3019 14980
rect 2961 14971 3019 14977
rect 3605 14977 3617 15011
rect 3651 15008 3663 15011
rect 3970 15008 3976 15020
rect 3651 14980 3976 15008
rect 3651 14977 3663 14980
rect 3605 14971 3663 14977
rect 1762 14900 1768 14952
rect 1820 14940 1826 14952
rect 2608 14940 2636 14971
rect 1820 14912 2636 14940
rect 2700 14940 2728 14971
rect 3970 14968 3976 14980
rect 4028 14968 4034 15020
rect 6181 15011 6239 15017
rect 6181 14977 6193 15011
rect 6227 15008 6239 15011
rect 6380 15008 6408 15107
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 7834 15104 7840 15156
rect 7892 15144 7898 15156
rect 8205 15147 8263 15153
rect 8205 15144 8217 15147
rect 7892 15116 8217 15144
rect 7892 15104 7898 15116
rect 8205 15113 8217 15116
rect 8251 15113 8263 15147
rect 8205 15107 8263 15113
rect 8573 15147 8631 15153
rect 8573 15113 8585 15147
rect 8619 15144 8631 15147
rect 9122 15144 9128 15156
rect 8619 15116 9128 15144
rect 8619 15113 8631 15116
rect 8573 15107 8631 15113
rect 9122 15104 9128 15116
rect 9180 15104 9186 15156
rect 9306 15104 9312 15156
rect 9364 15144 9370 15156
rect 9401 15147 9459 15153
rect 9401 15144 9413 15147
rect 9364 15116 9413 15144
rect 9364 15104 9370 15116
rect 9401 15113 9413 15116
rect 9447 15144 9459 15147
rect 9582 15144 9588 15156
rect 9447 15116 9588 15144
rect 9447 15113 9459 15116
rect 9401 15107 9459 15113
rect 9582 15104 9588 15116
rect 9640 15104 9646 15156
rect 11054 15104 11060 15156
rect 11112 15144 11118 15156
rect 11241 15147 11299 15153
rect 11241 15144 11253 15147
rect 11112 15116 11253 15144
rect 11112 15104 11118 15116
rect 11241 15113 11253 15116
rect 11287 15144 11299 15147
rect 11790 15144 11796 15156
rect 11287 15116 11796 15144
rect 11287 15113 11299 15116
rect 11241 15107 11299 15113
rect 11790 15104 11796 15116
rect 11848 15104 11854 15156
rect 12894 15144 12900 15156
rect 12855 15116 12900 15144
rect 12894 15104 12900 15116
rect 12952 15104 12958 15156
rect 12989 15147 13047 15153
rect 12989 15113 13001 15147
rect 13035 15144 13047 15147
rect 13170 15144 13176 15156
rect 13035 15116 13176 15144
rect 13035 15113 13047 15116
rect 12989 15107 13047 15113
rect 13170 15104 13176 15116
rect 13228 15104 13234 15156
rect 13814 15144 13820 15156
rect 13775 15116 13820 15144
rect 13814 15104 13820 15116
rect 13872 15104 13878 15156
rect 14277 15147 14335 15153
rect 14277 15113 14289 15147
rect 14323 15144 14335 15147
rect 14645 15147 14703 15153
rect 14645 15144 14657 15147
rect 14323 15116 14657 15144
rect 14323 15113 14335 15116
rect 14277 15107 14335 15113
rect 14645 15113 14657 15116
rect 14691 15113 14703 15147
rect 14645 15107 14703 15113
rect 12342 15076 12348 15088
rect 9876 15048 12348 15076
rect 7466 15008 7472 15020
rect 7524 15017 7530 15020
rect 6227 14980 6408 15008
rect 7436 14980 7472 15008
rect 6227 14977 6239 14980
rect 6181 14971 6239 14977
rect 7466 14968 7472 14980
rect 7524 14971 7536 15017
rect 7742 15008 7748 15020
rect 7703 14980 7748 15008
rect 7524 14968 7530 14971
rect 7742 14968 7748 14980
rect 7800 14968 7806 15020
rect 8570 14968 8576 15020
rect 8628 15008 8634 15020
rect 8665 15011 8723 15017
rect 8665 15008 8677 15011
rect 8628 14980 8677 15008
rect 8628 14968 8634 14980
rect 8665 14977 8677 14980
rect 8711 14977 8723 15011
rect 8665 14971 8723 14977
rect 9030 14968 9036 15020
rect 9088 15008 9094 15020
rect 9309 15011 9367 15017
rect 9309 15008 9321 15011
rect 9088 14980 9321 15008
rect 9088 14968 9094 14980
rect 9309 14977 9321 14980
rect 9355 15008 9367 15011
rect 9490 15008 9496 15020
rect 9355 14980 9496 15008
rect 9355 14977 9367 14980
rect 9309 14971 9367 14977
rect 9490 14968 9496 14980
rect 9548 14968 9554 15020
rect 9876 15017 9904 15048
rect 10134 15017 10140 15020
rect 9861 15011 9919 15017
rect 9861 14977 9873 15011
rect 9907 14977 9919 15011
rect 10128 15008 10140 15017
rect 9861 14971 9919 14977
rect 9968 14980 10140 15008
rect 3326 14940 3332 14952
rect 2700 14912 3332 14940
rect 1820 14900 1826 14912
rect 3326 14900 3332 14912
rect 3384 14900 3390 14952
rect 3694 14940 3700 14952
rect 3655 14912 3700 14940
rect 3694 14900 3700 14912
rect 3752 14900 3758 14952
rect 3789 14943 3847 14949
rect 3789 14909 3801 14943
rect 3835 14909 3847 14943
rect 4062 14940 4068 14952
rect 4023 14912 4068 14940
rect 3789 14903 3847 14909
rect 2038 14832 2044 14884
rect 2096 14872 2102 14884
rect 2409 14875 2467 14881
rect 2409 14872 2421 14875
rect 2096 14844 2421 14872
rect 2096 14832 2102 14844
rect 2409 14841 2421 14844
rect 2455 14841 2467 14875
rect 2409 14835 2467 14841
rect 2869 14875 2927 14881
rect 2869 14841 2881 14875
rect 2915 14872 2927 14875
rect 3510 14872 3516 14884
rect 2915 14844 3516 14872
rect 2915 14841 2927 14844
rect 2869 14835 2927 14841
rect 3510 14832 3516 14844
rect 3568 14832 3574 14884
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 3234 14764 3240 14816
rect 3292 14804 3298 14816
rect 3804 14804 3832 14903
rect 4062 14900 4068 14912
rect 4120 14900 4126 14952
rect 7837 14943 7895 14949
rect 7837 14909 7849 14943
rect 7883 14940 7895 14943
rect 8018 14940 8024 14952
rect 7883 14912 8024 14940
rect 7883 14909 7895 14912
rect 7837 14903 7895 14909
rect 8018 14900 8024 14912
rect 8076 14900 8082 14952
rect 8754 14940 8760 14952
rect 8715 14912 8760 14940
rect 8754 14900 8760 14912
rect 8812 14900 8818 14952
rect 9217 14943 9275 14949
rect 9217 14909 9229 14943
rect 9263 14940 9275 14943
rect 9968 14940 9996 14980
rect 10128 14971 10140 14980
rect 10134 14968 10140 14971
rect 10192 14968 10198 15020
rect 11532 15017 11560 15048
rect 12342 15036 12348 15048
rect 12400 15036 12406 15088
rect 11790 15017 11796 15020
rect 11517 15011 11575 15017
rect 11517 14977 11529 15011
rect 11563 14977 11575 15011
rect 11784 15008 11796 15017
rect 11751 14980 11796 15008
rect 11517 14971 11575 14977
rect 11784 14971 11796 14980
rect 11848 15008 11854 15020
rect 11848 14980 12572 15008
rect 11790 14968 11796 14971
rect 11848 14968 11854 14980
rect 9263 14912 9996 14940
rect 9263 14909 9275 14912
rect 9217 14903 9275 14909
rect 5442 14872 5448 14884
rect 5403 14844 5448 14872
rect 5442 14832 5448 14844
rect 5500 14832 5506 14884
rect 12544 14872 12572 14980
rect 12618 14968 12624 15020
rect 12676 15008 12682 15020
rect 13357 15011 13415 15017
rect 13357 15008 13369 15011
rect 12676 14980 13369 15008
rect 12676 14968 12682 14980
rect 13357 14977 13369 14980
rect 13403 14977 13415 15011
rect 13357 14971 13415 14977
rect 13722 14968 13728 15020
rect 13780 15008 13786 15020
rect 14185 15011 14243 15017
rect 14185 15008 14197 15011
rect 13780 14980 14197 15008
rect 13780 14968 13786 14980
rect 14185 14977 14197 14980
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 15013 15011 15071 15017
rect 15013 14977 15025 15011
rect 15059 15008 15071 15011
rect 15286 15008 15292 15020
rect 15059 14980 15292 15008
rect 15059 14977 15071 14980
rect 15013 14971 15071 14977
rect 15286 14968 15292 14980
rect 15344 15008 15350 15020
rect 15562 15008 15568 15020
rect 15344 14980 15568 15008
rect 15344 14968 15350 14980
rect 15562 14968 15568 14980
rect 15620 14968 15626 15020
rect 13446 14940 13452 14952
rect 13407 14912 13452 14940
rect 13446 14900 13452 14912
rect 13504 14900 13510 14952
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14940 13599 14943
rect 14369 14943 14427 14949
rect 14369 14940 14381 14943
rect 13587 14912 14381 14940
rect 13587 14909 13599 14912
rect 13541 14903 13599 14909
rect 14369 14909 14381 14912
rect 14415 14909 14427 14943
rect 15102 14940 15108 14952
rect 15063 14912 15108 14940
rect 14369 14903 14427 14909
rect 13556 14872 13584 14903
rect 15102 14900 15108 14912
rect 15160 14900 15166 14952
rect 15197 14943 15255 14949
rect 15197 14909 15209 14943
rect 15243 14909 15255 14943
rect 15197 14903 15255 14909
rect 12544 14844 13584 14872
rect 13814 14832 13820 14884
rect 13872 14872 13878 14884
rect 15212 14872 15240 14903
rect 13872 14844 15240 14872
rect 13872 14832 13878 14844
rect 3292 14776 3832 14804
rect 5537 14807 5595 14813
rect 3292 14764 3298 14776
rect 5537 14773 5549 14807
rect 5583 14804 5595 14807
rect 7098 14804 7104 14816
rect 5583 14776 7104 14804
rect 5583 14773 5595 14776
rect 5537 14767 5595 14773
rect 7098 14764 7104 14776
rect 7156 14764 7162 14816
rect 7466 14764 7472 14816
rect 7524 14804 7530 14816
rect 9674 14804 9680 14816
rect 7524 14776 9680 14804
rect 7524 14764 7530 14776
rect 9674 14764 9680 14776
rect 9732 14764 9738 14816
rect 9769 14807 9827 14813
rect 9769 14773 9781 14807
rect 9815 14804 9827 14807
rect 10594 14804 10600 14816
rect 9815 14776 10600 14804
rect 9815 14773 9827 14776
rect 9769 14767 9827 14773
rect 10594 14764 10600 14776
rect 10652 14764 10658 14816
rect 15562 14804 15568 14816
rect 15523 14776 15568 14804
rect 15562 14764 15568 14776
rect 15620 14764 15626 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 1946 14600 1952 14612
rect 1907 14572 1952 14600
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 3326 14560 3332 14612
rect 3384 14600 3390 14612
rect 3384 14572 3648 14600
rect 3384 14560 3390 14572
rect 3620 14532 3648 14572
rect 3878 14560 3884 14612
rect 3936 14600 3942 14612
rect 4433 14603 4491 14609
rect 4433 14600 4445 14603
rect 3936 14572 4445 14600
rect 3936 14560 3942 14572
rect 4433 14569 4445 14572
rect 4479 14569 4491 14603
rect 6638 14600 6644 14612
rect 4433 14563 4491 14569
rect 4540 14572 6644 14600
rect 4540 14532 4568 14572
rect 6638 14560 6644 14572
rect 6696 14560 6702 14612
rect 7466 14600 7472 14612
rect 6748 14572 7472 14600
rect 3620 14504 4568 14532
rect 1302 14424 1308 14476
rect 1360 14464 1366 14476
rect 3605 14467 3663 14473
rect 1360 14436 2176 14464
rect 1360 14424 1366 14436
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 2038 14396 2044 14408
rect 1719 14368 2044 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 2038 14356 2044 14368
rect 2096 14356 2102 14408
rect 2148 14405 2176 14436
rect 3605 14433 3617 14467
rect 3651 14464 3663 14467
rect 4062 14464 4068 14476
rect 3651 14436 4068 14464
rect 3651 14433 3663 14436
rect 3605 14427 3663 14433
rect 4062 14424 4068 14436
rect 4120 14464 4126 14476
rect 4120 14436 4936 14464
rect 4120 14424 4126 14436
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14365 2191 14399
rect 2133 14359 2191 14365
rect 2222 14356 2228 14408
rect 2280 14396 2286 14408
rect 4249 14399 4307 14405
rect 2280 14368 4200 14396
rect 2280 14356 2286 14368
rect 1394 14288 1400 14340
rect 1452 14328 1458 14340
rect 1765 14331 1823 14337
rect 1765 14328 1777 14331
rect 1452 14300 1777 14328
rect 1452 14288 1458 14300
rect 1765 14297 1777 14300
rect 1811 14297 1823 14331
rect 1765 14291 1823 14297
rect 3326 14288 3332 14340
rect 3384 14337 3390 14340
rect 3384 14328 3396 14337
rect 4172 14328 4200 14368
rect 4249 14365 4261 14399
rect 4295 14396 4307 14399
rect 4522 14396 4528 14408
rect 4295 14368 4528 14396
rect 4295 14365 4307 14368
rect 4249 14359 4307 14365
rect 4522 14356 4528 14368
rect 4580 14356 4586 14408
rect 4908 14396 4936 14436
rect 4982 14424 4988 14476
rect 5040 14464 5046 14476
rect 5040 14436 5085 14464
rect 5040 14424 5046 14436
rect 5537 14399 5595 14405
rect 5537 14396 5549 14399
rect 4908 14368 5549 14396
rect 5537 14365 5549 14368
rect 5583 14396 5595 14399
rect 5626 14396 5632 14408
rect 5583 14368 5632 14396
rect 5583 14365 5595 14368
rect 5537 14359 5595 14365
rect 5626 14356 5632 14368
rect 5684 14356 5690 14408
rect 5810 14405 5816 14408
rect 5804 14396 5816 14405
rect 5771 14368 5816 14396
rect 5804 14359 5816 14368
rect 5810 14356 5816 14359
rect 5868 14356 5874 14408
rect 4614 14328 4620 14340
rect 3384 14300 3429 14328
rect 4172 14300 4620 14328
rect 3384 14291 3396 14300
rect 3384 14288 3390 14291
rect 4614 14288 4620 14300
rect 4672 14288 4678 14340
rect 4801 14331 4859 14337
rect 4801 14297 4813 14331
rect 4847 14328 4859 14331
rect 4847 14300 5304 14328
rect 4847 14297 4859 14300
rect 4801 14291 4859 14297
rect 5276 14272 5304 14300
rect 5442 14288 5448 14340
rect 5500 14328 5506 14340
rect 6748 14328 6776 14572
rect 7466 14560 7472 14572
rect 7524 14560 7530 14612
rect 7558 14560 7564 14612
rect 7616 14600 7622 14612
rect 7653 14603 7711 14609
rect 7653 14600 7665 14603
rect 7616 14572 7665 14600
rect 7616 14560 7622 14572
rect 7653 14569 7665 14572
rect 7699 14569 7711 14603
rect 7653 14563 7711 14569
rect 7742 14560 7748 14612
rect 7800 14600 7806 14612
rect 8018 14600 8024 14612
rect 7800 14572 8024 14600
rect 7800 14560 7806 14572
rect 8018 14560 8024 14572
rect 8076 14560 8082 14612
rect 9122 14600 9128 14612
rect 9083 14572 9128 14600
rect 9122 14560 9128 14572
rect 9180 14560 9186 14612
rect 9858 14600 9864 14612
rect 9232 14572 9864 14600
rect 6917 14535 6975 14541
rect 6917 14501 6929 14535
rect 6963 14532 6975 14535
rect 7190 14532 7196 14544
rect 6963 14504 7196 14532
rect 6963 14501 6975 14504
rect 6917 14495 6975 14501
rect 6932 14396 6960 14495
rect 7190 14492 7196 14504
rect 7248 14532 7254 14544
rect 7926 14532 7932 14544
rect 7248 14504 7932 14532
rect 7248 14492 7254 14504
rect 7926 14492 7932 14504
rect 7984 14492 7990 14544
rect 8570 14492 8576 14544
rect 8628 14532 8634 14544
rect 9232 14541 9260 14572
rect 9858 14560 9864 14572
rect 9916 14560 9922 14612
rect 10229 14603 10287 14609
rect 10229 14569 10241 14603
rect 10275 14600 10287 14603
rect 10778 14600 10784 14612
rect 10275 14572 10784 14600
rect 10275 14569 10287 14572
rect 10229 14563 10287 14569
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 11238 14560 11244 14612
rect 11296 14600 11302 14612
rect 11517 14603 11575 14609
rect 11517 14600 11529 14603
rect 11296 14572 11529 14600
rect 11296 14560 11302 14572
rect 11517 14569 11529 14572
rect 11563 14569 11575 14603
rect 13722 14600 13728 14612
rect 13683 14572 13728 14600
rect 11517 14563 11575 14569
rect 13722 14560 13728 14572
rect 13780 14560 13786 14612
rect 19058 14600 19064 14612
rect 13832 14572 19064 14600
rect 9217 14535 9275 14541
rect 9217 14532 9229 14535
rect 8628 14504 9229 14532
rect 8628 14492 8634 14504
rect 9217 14501 9229 14504
rect 9263 14501 9275 14535
rect 10042 14532 10048 14544
rect 9217 14495 9275 14501
rect 9600 14504 10048 14532
rect 8018 14424 8024 14476
rect 8076 14464 8082 14476
rect 8297 14467 8355 14473
rect 8297 14464 8309 14467
rect 8076 14436 8309 14464
rect 8076 14424 8082 14436
rect 8297 14433 8309 14436
rect 8343 14433 8355 14467
rect 8297 14427 8355 14433
rect 7009 14399 7067 14405
rect 7009 14396 7021 14399
rect 6932 14368 7021 14396
rect 7009 14365 7021 14368
rect 7055 14365 7067 14399
rect 7009 14359 7067 14365
rect 5500 14300 6776 14328
rect 5500 14288 5506 14300
rect 6822 14288 6828 14340
rect 6880 14328 6886 14340
rect 9600 14328 9628 14504
rect 10042 14492 10048 14504
rect 10100 14532 10106 14544
rect 10962 14532 10968 14544
rect 10100 14504 10968 14532
rect 10100 14492 10106 14504
rect 10962 14492 10968 14504
rect 11020 14492 11026 14544
rect 11164 14504 13124 14532
rect 11164 14476 11192 14504
rect 9677 14467 9735 14473
rect 9677 14433 9689 14467
rect 9723 14464 9735 14467
rect 10134 14464 10140 14476
rect 9723 14436 10140 14464
rect 9723 14433 9735 14436
rect 9677 14427 9735 14433
rect 10134 14424 10140 14436
rect 10192 14464 10198 14476
rect 11146 14464 11152 14476
rect 10192 14436 10456 14464
rect 11107 14436 11152 14464
rect 10192 14424 10198 14436
rect 9766 14356 9772 14408
rect 9824 14396 9830 14408
rect 10428 14396 10456 14436
rect 11146 14424 11152 14436
rect 11204 14424 11210 14476
rect 12069 14467 12127 14473
rect 12069 14433 12081 14467
rect 12115 14433 12127 14467
rect 12618 14464 12624 14476
rect 12579 14436 12624 14464
rect 12069 14427 12127 14433
rect 12084 14396 12112 14427
rect 12618 14424 12624 14436
rect 12676 14424 12682 14476
rect 13096 14473 13124 14504
rect 13262 14492 13268 14544
rect 13320 14532 13326 14544
rect 13832 14532 13860 14572
rect 19058 14560 19064 14572
rect 19116 14560 19122 14612
rect 13320 14504 13860 14532
rect 13320 14492 13326 14504
rect 13081 14467 13139 14473
rect 13081 14433 13093 14467
rect 13127 14464 13139 14467
rect 13814 14464 13820 14476
rect 13127 14436 13820 14464
rect 13127 14433 13139 14436
rect 13081 14427 13139 14433
rect 13814 14424 13820 14436
rect 13872 14424 13878 14476
rect 16206 14424 16212 14476
rect 16264 14464 16270 14476
rect 16577 14467 16635 14473
rect 16577 14464 16589 14467
rect 16264 14436 16589 14464
rect 16264 14424 16270 14436
rect 16577 14433 16589 14436
rect 16623 14433 16635 14467
rect 16577 14427 16635 14433
rect 9824 14368 9869 14396
rect 10428 14368 12112 14396
rect 9824 14356 9830 14368
rect 12342 14356 12348 14408
rect 12400 14396 12406 14408
rect 14274 14396 14280 14408
rect 12400 14368 14280 14396
rect 12400 14356 12406 14368
rect 14274 14356 14280 14368
rect 14332 14356 14338 14408
rect 15654 14356 15660 14408
rect 15712 14405 15718 14408
rect 15712 14396 15724 14405
rect 15933 14399 15991 14405
rect 15712 14368 15757 14396
rect 15712 14359 15724 14368
rect 15933 14365 15945 14399
rect 15979 14396 15991 14399
rect 16942 14396 16948 14408
rect 15979 14368 16948 14396
rect 15979 14365 15991 14368
rect 15933 14359 15991 14365
rect 15712 14356 15718 14359
rect 16942 14356 16948 14368
rect 17000 14356 17006 14408
rect 6880 14300 9628 14328
rect 6880 14288 6886 14300
rect 9674 14288 9680 14340
rect 9732 14328 9738 14340
rect 10413 14331 10471 14337
rect 10413 14328 10425 14331
rect 9732 14300 10425 14328
rect 9732 14288 9738 14300
rect 10413 14297 10425 14300
rect 10459 14328 10471 14331
rect 11057 14331 11115 14337
rect 11057 14328 11069 14331
rect 10459 14300 11069 14328
rect 10459 14297 10471 14300
rect 10413 14291 10471 14297
rect 11057 14297 11069 14300
rect 11103 14328 11115 14331
rect 16482 14328 16488 14340
rect 11103 14300 16160 14328
rect 16443 14300 16488 14328
rect 11103 14297 11115 14300
rect 11057 14291 11115 14297
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 2225 14263 2283 14269
rect 2225 14229 2237 14263
rect 2271 14260 2283 14263
rect 2498 14260 2504 14272
rect 2271 14232 2504 14260
rect 2271 14229 2283 14232
rect 2225 14223 2283 14229
rect 2498 14220 2504 14232
rect 2556 14260 2562 14272
rect 3234 14260 3240 14272
rect 2556 14232 3240 14260
rect 2556 14220 2562 14232
rect 3234 14220 3240 14232
rect 3292 14220 3298 14272
rect 3602 14220 3608 14272
rect 3660 14260 3666 14272
rect 3789 14263 3847 14269
rect 3789 14260 3801 14263
rect 3660 14232 3801 14260
rect 3660 14220 3666 14232
rect 3789 14229 3801 14232
rect 3835 14229 3847 14263
rect 3789 14223 3847 14229
rect 3878 14220 3884 14272
rect 3936 14260 3942 14272
rect 4065 14263 4123 14269
rect 4065 14260 4077 14263
rect 3936 14232 4077 14260
rect 3936 14220 3942 14232
rect 4065 14229 4077 14232
rect 4111 14229 4123 14263
rect 4065 14223 4123 14229
rect 4890 14220 4896 14272
rect 4948 14260 4954 14272
rect 5258 14260 5264 14272
rect 4948 14232 4993 14260
rect 5219 14232 5264 14260
rect 4948 14220 4954 14232
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 5350 14220 5356 14272
rect 5408 14260 5414 14272
rect 7466 14260 7472 14272
rect 5408 14232 7472 14260
rect 5408 14220 5414 14232
rect 7466 14220 7472 14232
rect 7524 14220 7530 14272
rect 7558 14220 7564 14272
rect 7616 14260 7622 14272
rect 7745 14263 7803 14269
rect 7745 14260 7757 14263
rect 7616 14232 7757 14260
rect 7616 14220 7622 14232
rect 7745 14229 7757 14232
rect 7791 14229 7803 14263
rect 8110 14260 8116 14272
rect 8071 14232 8116 14260
rect 7745 14223 7803 14229
rect 8110 14220 8116 14232
rect 8168 14220 8174 14272
rect 8202 14220 8208 14272
rect 8260 14260 8266 14272
rect 8260 14232 8305 14260
rect 8260 14220 8266 14232
rect 8386 14220 8392 14272
rect 8444 14260 8450 14272
rect 8662 14260 8668 14272
rect 8444 14232 8668 14260
rect 8444 14220 8450 14232
rect 8662 14220 8668 14232
rect 8720 14220 8726 14272
rect 9858 14220 9864 14272
rect 9916 14260 9922 14272
rect 10597 14263 10655 14269
rect 9916 14232 9961 14260
rect 9916 14220 9922 14232
rect 10597 14229 10609 14263
rect 10643 14260 10655 14263
rect 10686 14260 10692 14272
rect 10643 14232 10692 14260
rect 10643 14229 10655 14232
rect 10597 14223 10655 14229
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 10962 14260 10968 14272
rect 10923 14232 10968 14260
rect 10962 14220 10968 14232
rect 11020 14220 11026 14272
rect 11790 14220 11796 14272
rect 11848 14260 11854 14272
rect 11885 14263 11943 14269
rect 11885 14260 11897 14263
rect 11848 14232 11897 14260
rect 11848 14220 11854 14232
rect 11885 14229 11897 14232
rect 11931 14229 11943 14263
rect 11885 14223 11943 14229
rect 11977 14263 12035 14269
rect 11977 14229 11989 14263
rect 12023 14260 12035 14263
rect 12066 14260 12072 14272
rect 12023 14232 12072 14260
rect 12023 14229 12035 14232
rect 11977 14223 12035 14229
rect 12066 14220 12072 14232
rect 12124 14220 12130 14272
rect 12618 14220 12624 14272
rect 12676 14260 12682 14272
rect 12713 14263 12771 14269
rect 12713 14260 12725 14263
rect 12676 14232 12725 14260
rect 12676 14220 12682 14232
rect 12713 14229 12725 14232
rect 12759 14260 12771 14263
rect 13262 14260 13268 14272
rect 12759 14232 13268 14260
rect 12759 14229 12771 14232
rect 12713 14223 12771 14229
rect 13262 14220 13268 14232
rect 13320 14220 13326 14272
rect 13357 14263 13415 14269
rect 13357 14229 13369 14263
rect 13403 14260 13415 14263
rect 13630 14260 13636 14272
rect 13403 14232 13636 14260
rect 13403 14229 13415 14232
rect 13357 14223 13415 14229
rect 13630 14220 13636 14232
rect 13688 14260 13694 14272
rect 13817 14263 13875 14269
rect 13817 14260 13829 14263
rect 13688 14232 13829 14260
rect 13688 14220 13694 14232
rect 13817 14229 13829 14232
rect 13863 14229 13875 14263
rect 13817 14223 13875 14229
rect 14553 14263 14611 14269
rect 14553 14229 14565 14263
rect 14599 14260 14611 14263
rect 14734 14260 14740 14272
rect 14599 14232 14740 14260
rect 14599 14229 14611 14232
rect 14553 14223 14611 14229
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 14918 14220 14924 14272
rect 14976 14260 14982 14272
rect 16025 14263 16083 14269
rect 16025 14260 16037 14263
rect 14976 14232 16037 14260
rect 14976 14220 14982 14232
rect 16025 14229 16037 14232
rect 16071 14229 16083 14263
rect 16132 14260 16160 14300
rect 16482 14288 16488 14300
rect 16540 14288 16546 14340
rect 16390 14260 16396 14272
rect 16132 14232 16396 14260
rect 16025 14223 16083 14229
rect 16390 14220 16396 14232
rect 16448 14220 16454 14272
rect 1104 14170 21896 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21896 14170
rect 1104 14096 21896 14118
rect 1854 14056 1860 14068
rect 1815 14028 1860 14056
rect 1854 14016 1860 14028
rect 1912 14016 1918 14068
rect 2038 14016 2044 14068
rect 2096 14056 2102 14068
rect 2133 14059 2191 14065
rect 2133 14056 2145 14059
rect 2096 14028 2145 14056
rect 2096 14016 2102 14028
rect 2133 14025 2145 14028
rect 2179 14025 2191 14059
rect 2133 14019 2191 14025
rect 3145 14059 3203 14065
rect 3145 14025 3157 14059
rect 3191 14056 3203 14059
rect 3418 14056 3424 14068
rect 3191 14028 3424 14056
rect 3191 14025 3203 14028
rect 3145 14019 3203 14025
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 3602 14056 3608 14068
rect 3563 14028 3608 14056
rect 3602 14016 3608 14028
rect 3660 14016 3666 14068
rect 3970 14056 3976 14068
rect 3931 14028 3976 14056
rect 3970 14016 3976 14028
rect 4028 14016 4034 14068
rect 4065 14059 4123 14065
rect 4065 14025 4077 14059
rect 4111 14056 4123 14059
rect 4154 14056 4160 14068
rect 4111 14028 4160 14056
rect 4111 14025 4123 14028
rect 4065 14019 4123 14025
rect 4154 14016 4160 14028
rect 4212 14056 4218 14068
rect 4982 14056 4988 14068
rect 4212 14028 4988 14056
rect 4212 14016 4218 14028
rect 4982 14016 4988 14028
rect 5040 14016 5046 14068
rect 7558 14056 7564 14068
rect 7519 14028 7564 14056
rect 7558 14016 7564 14028
rect 7616 14016 7622 14068
rect 7650 14016 7656 14068
rect 7708 14016 7714 14068
rect 8110 14016 8116 14068
rect 8168 14056 8174 14068
rect 9401 14059 9459 14065
rect 9401 14056 9413 14059
rect 8168 14028 9413 14056
rect 8168 14016 8174 14028
rect 9401 14025 9413 14028
rect 9447 14025 9459 14059
rect 10686 14056 10692 14068
rect 10647 14028 10692 14056
rect 9401 14019 9459 14025
rect 10686 14016 10692 14028
rect 10744 14016 10750 14068
rect 11149 14059 11207 14065
rect 11149 14025 11161 14059
rect 11195 14056 11207 14059
rect 11882 14056 11888 14068
rect 11195 14028 11888 14056
rect 11195 14025 11207 14028
rect 11149 14019 11207 14025
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 12342 14016 12348 14068
rect 12400 14056 12406 14068
rect 13173 14059 13231 14065
rect 13173 14056 13185 14059
rect 12400 14028 13185 14056
rect 12400 14016 12406 14028
rect 13173 14025 13185 14028
rect 13219 14025 13231 14059
rect 13814 14056 13820 14068
rect 13775 14028 13820 14056
rect 13173 14019 13231 14025
rect 13814 14016 13820 14028
rect 13872 14016 13878 14068
rect 14918 14056 14924 14068
rect 14879 14028 14924 14056
rect 14918 14016 14924 14028
rect 14976 14016 14982 14068
rect 15749 14059 15807 14065
rect 15749 14025 15761 14059
rect 15795 14056 15807 14059
rect 16390 14056 16396 14068
rect 15795 14028 16396 14056
rect 15795 14025 15807 14028
rect 15749 14019 15807 14025
rect 16390 14016 16396 14028
rect 16448 14016 16454 14068
rect 5200 13991 5258 13997
rect 5200 13957 5212 13991
rect 5246 13988 5258 13991
rect 6181 13991 6239 13997
rect 6181 13988 6193 13991
rect 5246 13960 6193 13988
rect 5246 13957 5258 13960
rect 5200 13951 5258 13957
rect 6181 13957 6193 13960
rect 6227 13957 6239 13991
rect 7668 13988 7696 14016
rect 9306 13988 9312 14000
rect 7668 13960 9312 13988
rect 6181 13951 6239 13957
rect 9306 13948 9312 13960
rect 9364 13988 9370 14000
rect 9858 13988 9864 14000
rect 9364 13960 9864 13988
rect 9364 13948 9370 13960
rect 9858 13948 9864 13960
rect 9916 13948 9922 14000
rect 10594 13948 10600 14000
rect 10652 13988 10658 14000
rect 10781 13991 10839 13997
rect 10781 13988 10793 13991
rect 10652 13960 10793 13988
rect 10652 13948 10658 13960
rect 10781 13957 10793 13960
rect 10827 13957 10839 13991
rect 12802 13988 12808 14000
rect 10781 13951 10839 13957
rect 10888 13960 12808 13988
rect 1670 13920 1676 13932
rect 1631 13892 1676 13920
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 2038 13920 2044 13932
rect 1999 13892 2044 13920
rect 2038 13880 2044 13892
rect 2096 13880 2102 13932
rect 2317 13923 2375 13929
rect 2317 13889 2329 13923
rect 2363 13889 2375 13923
rect 2498 13920 2504 13932
rect 2459 13892 2504 13920
rect 2317 13883 2375 13889
rect 2332 13852 2360 13883
rect 2498 13880 2504 13892
rect 2556 13880 2562 13932
rect 3326 13880 3332 13932
rect 3384 13920 3390 13932
rect 4154 13920 4160 13932
rect 3384 13892 4160 13920
rect 3384 13880 3390 13892
rect 2682 13852 2688 13864
rect 2332 13824 2688 13852
rect 2682 13812 2688 13824
rect 2740 13812 2746 13864
rect 3436 13861 3464 13892
rect 4154 13880 4160 13892
rect 4212 13880 4218 13932
rect 5350 13920 5356 13932
rect 4448 13892 5356 13920
rect 3421 13855 3479 13861
rect 3421 13821 3433 13855
rect 3467 13821 3479 13855
rect 3421 13815 3479 13821
rect 3510 13812 3516 13864
rect 3568 13852 3574 13864
rect 4448 13852 4476 13892
rect 5350 13880 5356 13892
rect 5408 13880 5414 13932
rect 5534 13920 5540 13932
rect 5495 13892 5540 13920
rect 5534 13880 5540 13892
rect 5592 13880 5598 13932
rect 6365 13923 6423 13929
rect 6365 13889 6377 13923
rect 6411 13920 6423 13923
rect 7282 13920 7288 13932
rect 6411 13892 7288 13920
rect 6411 13889 6423 13892
rect 6365 13883 6423 13889
rect 7282 13880 7288 13892
rect 7340 13880 7346 13932
rect 7469 13923 7527 13929
rect 7469 13889 7481 13923
rect 7515 13920 7527 13923
rect 8018 13920 8024 13932
rect 7515 13892 8024 13920
rect 7515 13889 7527 13892
rect 7469 13883 7527 13889
rect 8018 13880 8024 13892
rect 8076 13880 8082 13932
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 9053 13923 9111 13929
rect 9053 13920 9065 13923
rect 8352 13892 9065 13920
rect 8352 13880 8358 13892
rect 9053 13889 9065 13892
rect 9099 13920 9111 13923
rect 9099 13892 9444 13920
rect 9099 13889 9111 13892
rect 9053 13883 9111 13889
rect 3568 13824 4476 13852
rect 5445 13855 5503 13861
rect 3568 13812 3574 13824
rect 5445 13821 5457 13855
rect 5491 13852 5503 13855
rect 5718 13852 5724 13864
rect 5491 13824 5724 13852
rect 5491 13821 5503 13824
rect 5445 13815 5503 13821
rect 5718 13812 5724 13824
rect 5776 13812 5782 13864
rect 7653 13855 7711 13861
rect 7653 13852 7665 13855
rect 6932 13824 7665 13852
rect 6546 13744 6552 13796
rect 6604 13784 6610 13796
rect 6932 13784 6960 13824
rect 7653 13821 7665 13824
rect 7699 13821 7711 13855
rect 9306 13852 9312 13864
rect 9267 13824 9312 13852
rect 7653 13815 7711 13821
rect 9306 13812 9312 13824
rect 9364 13812 9370 13864
rect 6604 13756 6960 13784
rect 7009 13787 7067 13793
rect 6604 13744 6610 13756
rect 7009 13753 7021 13787
rect 7055 13784 7067 13787
rect 7466 13784 7472 13796
rect 7055 13756 7472 13784
rect 7055 13753 7067 13756
rect 7009 13747 7067 13753
rect 7466 13744 7472 13756
rect 7524 13744 7530 13796
rect 7558 13744 7564 13796
rect 7616 13784 7622 13796
rect 9416 13784 9444 13892
rect 9490 13880 9496 13932
rect 9548 13920 9554 13932
rect 9769 13923 9827 13929
rect 9769 13920 9781 13923
rect 9548 13892 9781 13920
rect 9548 13880 9554 13892
rect 9769 13889 9781 13892
rect 9815 13889 9827 13923
rect 9769 13883 9827 13889
rect 10226 13880 10232 13932
rect 10284 13920 10290 13932
rect 10888 13920 10916 13960
rect 12802 13948 12808 13960
rect 12860 13948 12866 14000
rect 13265 13991 13323 13997
rect 13265 13957 13277 13991
rect 13311 13988 13323 13991
rect 15013 13991 15071 13997
rect 15013 13988 15025 13991
rect 13311 13960 15025 13988
rect 13311 13957 13323 13960
rect 13265 13951 13323 13957
rect 15013 13957 15025 13960
rect 15059 13988 15071 13991
rect 15102 13988 15108 14000
rect 15059 13960 15108 13988
rect 15059 13957 15071 13960
rect 15013 13951 15071 13957
rect 15102 13948 15108 13960
rect 15160 13988 15166 14000
rect 15160 13960 16574 13988
rect 15160 13948 15166 13960
rect 10284 13892 10916 13920
rect 10284 13880 10290 13892
rect 11146 13880 11152 13932
rect 11204 13920 11210 13932
rect 11517 13923 11575 13929
rect 11517 13920 11529 13923
rect 11204 13892 11529 13920
rect 11204 13880 11210 13892
rect 11517 13889 11529 13892
rect 11563 13920 11575 13923
rect 12066 13920 12072 13932
rect 11563 13892 12072 13920
rect 11563 13889 11575 13892
rect 11517 13883 11575 13889
rect 12066 13880 12072 13892
rect 12124 13920 12130 13932
rect 13722 13920 13728 13932
rect 12124 13892 13032 13920
rect 12124 13880 12130 13892
rect 9858 13852 9864 13864
rect 9819 13824 9864 13852
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 10045 13855 10103 13861
rect 10045 13821 10057 13855
rect 10091 13821 10103 13855
rect 10045 13815 10103 13821
rect 10597 13855 10655 13861
rect 10597 13821 10609 13855
rect 10643 13852 10655 13855
rect 11054 13852 11060 13864
rect 10643 13824 11060 13852
rect 10643 13821 10655 13824
rect 10597 13815 10655 13821
rect 10060 13784 10088 13815
rect 11054 13812 11060 13824
rect 11112 13812 11118 13864
rect 11333 13855 11391 13861
rect 11333 13821 11345 13855
rect 11379 13852 11391 13855
rect 11790 13852 11796 13864
rect 11379 13824 11796 13852
rect 11379 13821 11391 13824
rect 11333 13815 11391 13821
rect 11790 13812 11796 13824
rect 11848 13812 11854 13864
rect 13004 13852 13032 13892
rect 13280 13892 13584 13920
rect 13683 13892 13728 13920
rect 13280 13852 13308 13892
rect 12452 13824 12940 13852
rect 13004 13824 13308 13852
rect 13449 13855 13507 13861
rect 12452 13784 12480 13824
rect 12802 13784 12808 13796
rect 7616 13756 8064 13784
rect 9416 13756 12480 13784
rect 12763 13756 12808 13784
rect 7616 13744 7622 13756
rect 1486 13716 1492 13728
rect 1447 13688 1492 13716
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 7098 13676 7104 13728
rect 7156 13716 7162 13728
rect 7926 13716 7932 13728
rect 7156 13688 7201 13716
rect 7887 13688 7932 13716
rect 7156 13676 7162 13688
rect 7926 13676 7932 13688
rect 7984 13676 7990 13728
rect 8036 13716 8064 13756
rect 12802 13744 12808 13756
rect 12860 13744 12866 13796
rect 12912 13784 12940 13824
rect 13449 13821 13461 13855
rect 13495 13821 13507 13855
rect 13556 13852 13584 13892
rect 13722 13880 13728 13892
rect 13780 13880 13786 13932
rect 15841 13923 15899 13929
rect 15841 13920 15853 13923
rect 13832 13892 15853 13920
rect 13832 13852 13860 13892
rect 15841 13889 15853 13892
rect 15887 13920 15899 13923
rect 16298 13920 16304 13932
rect 15887 13892 16304 13920
rect 15887 13889 15899 13892
rect 15841 13883 15899 13889
rect 16298 13880 16304 13892
rect 16356 13880 16362 13932
rect 16546 13920 16574 13960
rect 21358 13920 21364 13932
rect 16546 13892 21364 13920
rect 21358 13880 21364 13892
rect 21416 13880 21422 13932
rect 14734 13852 14740 13864
rect 13556 13824 13860 13852
rect 14695 13824 14740 13852
rect 13449 13815 13507 13821
rect 13464 13784 13492 13815
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 16298 13784 16304 13796
rect 12912 13756 16304 13784
rect 16298 13744 16304 13756
rect 16356 13744 16362 13796
rect 9766 13716 9772 13728
rect 8036 13688 9772 13716
rect 9766 13676 9772 13688
rect 9824 13676 9830 13728
rect 11882 13676 11888 13728
rect 11940 13716 11946 13728
rect 12342 13716 12348 13728
rect 11940 13688 12348 13716
rect 11940 13676 11946 13688
rect 12342 13676 12348 13688
rect 12400 13716 12406 13728
rect 12621 13719 12679 13725
rect 12621 13716 12633 13719
rect 12400 13688 12633 13716
rect 12400 13676 12406 13688
rect 12621 13685 12633 13688
rect 12667 13685 12679 13719
rect 12621 13679 12679 13685
rect 15381 13719 15439 13725
rect 15381 13685 15393 13719
rect 15427 13716 15439 13719
rect 15562 13716 15568 13728
rect 15427 13688 15568 13716
rect 15427 13685 15439 13688
rect 15381 13679 15439 13685
rect 15562 13676 15568 13688
rect 15620 13676 15626 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 1670 13472 1676 13524
rect 1728 13512 1734 13524
rect 1765 13515 1823 13521
rect 1765 13512 1777 13515
rect 1728 13484 1777 13512
rect 1728 13472 1734 13484
rect 1765 13481 1777 13484
rect 1811 13481 1823 13515
rect 1765 13475 1823 13481
rect 2590 13472 2596 13524
rect 2648 13512 2654 13524
rect 3145 13515 3203 13521
rect 3145 13512 3157 13515
rect 2648 13484 3157 13512
rect 2648 13472 2654 13484
rect 3145 13481 3157 13484
rect 3191 13481 3203 13515
rect 3418 13512 3424 13524
rect 3379 13484 3424 13512
rect 3145 13475 3203 13481
rect 3418 13472 3424 13484
rect 3476 13472 3482 13524
rect 4065 13515 4123 13521
rect 4065 13481 4077 13515
rect 4111 13512 4123 13515
rect 4430 13512 4436 13524
rect 4111 13484 4436 13512
rect 4111 13481 4123 13484
rect 4065 13475 4123 13481
rect 4430 13472 4436 13484
rect 4488 13472 4494 13524
rect 4890 13472 4896 13524
rect 4948 13512 4954 13524
rect 5169 13515 5227 13521
rect 5169 13512 5181 13515
rect 4948 13484 5181 13512
rect 4948 13472 4954 13484
rect 5169 13481 5181 13484
rect 5215 13481 5227 13515
rect 5169 13475 5227 13481
rect 7929 13515 7987 13521
rect 7929 13481 7941 13515
rect 7975 13512 7987 13515
rect 8202 13512 8208 13524
rect 7975 13484 8208 13512
rect 7975 13481 7987 13484
rect 7929 13475 7987 13481
rect 8202 13472 8208 13484
rect 8260 13472 8266 13524
rect 9033 13515 9091 13521
rect 9033 13481 9045 13515
rect 9079 13512 9091 13515
rect 9122 13512 9128 13524
rect 9079 13484 9128 13512
rect 9079 13481 9091 13484
rect 9033 13475 9091 13481
rect 9122 13472 9128 13484
rect 9180 13472 9186 13524
rect 9309 13515 9367 13521
rect 9309 13481 9321 13515
rect 9355 13512 9367 13515
rect 9674 13512 9680 13524
rect 9355 13484 9680 13512
rect 9355 13481 9367 13484
rect 9309 13475 9367 13481
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 11698 13472 11704 13524
rect 11756 13512 11762 13524
rect 15102 13512 15108 13524
rect 11756 13484 15108 13512
rect 11756 13472 11762 13484
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 16298 13512 16304 13524
rect 16259 13484 16304 13512
rect 16298 13472 16304 13484
rect 16356 13472 16362 13524
rect 16390 13472 16396 13524
rect 16448 13512 16454 13524
rect 17034 13512 17040 13524
rect 16448 13484 17040 13512
rect 16448 13472 16454 13484
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 2866 13404 2872 13456
rect 2924 13444 2930 13456
rect 3789 13447 3847 13453
rect 3789 13444 3801 13447
rect 2924 13416 3801 13444
rect 2924 13404 2930 13416
rect 3789 13413 3801 13416
rect 3835 13413 3847 13447
rect 8018 13444 8024 13456
rect 7979 13416 8024 13444
rect 3789 13407 3847 13413
rect 8018 13404 8024 13416
rect 8076 13404 8082 13456
rect 8570 13404 8576 13456
rect 8628 13444 8634 13456
rect 9490 13444 9496 13456
rect 8628 13416 9496 13444
rect 8628 13404 8634 13416
rect 9490 13404 9496 13416
rect 9548 13404 9554 13456
rect 15470 13404 15476 13456
rect 15528 13444 15534 13456
rect 15749 13447 15807 13453
rect 15749 13444 15761 13447
rect 15528 13416 15761 13444
rect 15528 13404 15534 13416
rect 15749 13413 15761 13416
rect 15795 13413 15807 13447
rect 15749 13407 15807 13413
rect 2222 13336 2228 13388
rect 2280 13376 2286 13388
rect 2593 13379 2651 13385
rect 2593 13376 2605 13379
rect 2280 13348 2605 13376
rect 2280 13336 2286 13348
rect 2593 13345 2605 13348
rect 2639 13345 2651 13379
rect 2593 13339 2651 13345
rect 2774 13336 2780 13388
rect 2832 13376 2838 13388
rect 3418 13376 3424 13388
rect 2832 13348 3424 13376
rect 2832 13336 2838 13348
rect 3418 13336 3424 13348
rect 3476 13336 3482 13388
rect 4617 13379 4675 13385
rect 4617 13345 4629 13379
rect 4663 13376 4675 13379
rect 5534 13376 5540 13388
rect 4663 13348 5540 13376
rect 4663 13345 4675 13348
rect 4617 13339 4675 13345
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 7377 13379 7435 13385
rect 7377 13345 7389 13379
rect 7423 13376 7435 13379
rect 8202 13376 8208 13388
rect 7423 13348 8208 13376
rect 7423 13345 7435 13348
rect 7377 13339 7435 13345
rect 8202 13336 8208 13348
rect 8260 13336 8266 13388
rect 8662 13376 8668 13388
rect 8623 13348 8668 13376
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 9030 13336 9036 13388
rect 9088 13376 9094 13388
rect 9398 13376 9404 13388
rect 9088 13348 9404 13376
rect 9088 13336 9094 13348
rect 9398 13336 9404 13348
rect 9456 13336 9462 13388
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13376 9827 13379
rect 10502 13376 10508 13388
rect 9815 13348 10508 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 10502 13336 10508 13348
rect 10560 13336 10566 13388
rect 10612 13348 12480 13376
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13268 1458 13320
rect 1854 13268 1860 13320
rect 1912 13308 1918 13320
rect 1949 13311 2007 13317
rect 1949 13308 1961 13311
rect 1912 13280 1961 13308
rect 1912 13268 1918 13280
rect 1949 13277 1961 13280
rect 1995 13277 2007 13311
rect 1949 13271 2007 13277
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13308 2927 13311
rect 2958 13308 2964 13320
rect 2915 13280 2964 13308
rect 2915 13277 2927 13280
rect 2869 13271 2927 13277
rect 2958 13268 2964 13280
rect 3016 13268 3022 13320
rect 3329 13311 3387 13317
rect 3329 13308 3341 13311
rect 3068 13280 3341 13308
rect 1578 13172 1584 13184
rect 1539 13144 1584 13172
rect 1578 13132 1584 13144
rect 1636 13132 1642 13184
rect 2041 13175 2099 13181
rect 2041 13141 2053 13175
rect 2087 13172 2099 13175
rect 2130 13172 2136 13184
rect 2087 13144 2136 13172
rect 2087 13141 2099 13144
rect 2041 13135 2099 13141
rect 2130 13132 2136 13144
rect 2188 13132 2194 13184
rect 2406 13172 2412 13184
rect 2367 13144 2412 13172
rect 2406 13132 2412 13144
rect 2464 13132 2470 13184
rect 2498 13132 2504 13184
rect 2556 13172 2562 13184
rect 3068 13181 3096 13280
rect 3329 13277 3341 13280
rect 3375 13277 3387 13311
rect 3329 13271 3387 13277
rect 4709 13311 4767 13317
rect 4709 13277 4721 13311
rect 4755 13308 4767 13311
rect 5442 13308 5448 13320
rect 4755 13280 5448 13308
rect 4755 13277 4767 13280
rect 4709 13271 4767 13277
rect 5442 13268 5448 13280
rect 5500 13308 5506 13320
rect 6638 13308 6644 13320
rect 5500 13280 6644 13308
rect 5500 13268 5506 13280
rect 6638 13268 6644 13280
rect 6696 13268 6702 13320
rect 7006 13308 7012 13320
rect 6967 13280 7012 13308
rect 7006 13268 7012 13280
rect 7064 13308 7070 13320
rect 10410 13308 10416 13320
rect 7064 13280 10416 13308
rect 7064 13268 7070 13280
rect 10410 13268 10416 13280
rect 10468 13268 10474 13320
rect 4341 13243 4399 13249
rect 4341 13209 4353 13243
rect 4387 13240 4399 13243
rect 4801 13243 4859 13249
rect 4801 13240 4813 13243
rect 4387 13212 4813 13240
rect 4387 13209 4399 13212
rect 4341 13203 4399 13209
rect 4801 13209 4813 13212
rect 4847 13240 4859 13243
rect 5626 13240 5632 13252
rect 4847 13212 5632 13240
rect 4847 13209 4859 13212
rect 4801 13203 4859 13209
rect 5626 13200 5632 13212
rect 5684 13200 5690 13252
rect 7558 13240 7564 13252
rect 7519 13212 7564 13240
rect 7558 13200 7564 13212
rect 7616 13200 7622 13252
rect 8481 13243 8539 13249
rect 8481 13209 8493 13243
rect 8527 13240 8539 13243
rect 10612 13240 10640 13348
rect 12345 13311 12403 13317
rect 12345 13308 12357 13311
rect 8527 13212 10640 13240
rect 11716 13280 12357 13308
rect 8527 13209 8539 13212
rect 8481 13203 8539 13209
rect 11716 13184 11744 13280
rect 12345 13277 12357 13280
rect 12391 13277 12403 13311
rect 12345 13271 12403 13277
rect 3053 13175 3111 13181
rect 2556 13144 2601 13172
rect 2556 13132 2562 13144
rect 3053 13141 3065 13175
rect 3099 13141 3111 13175
rect 5718 13172 5724 13184
rect 5679 13144 5724 13172
rect 3053 13135 3111 13141
rect 5718 13132 5724 13144
rect 5776 13132 5782 13184
rect 5810 13132 5816 13184
rect 5868 13172 5874 13184
rect 7469 13175 7527 13181
rect 7469 13172 7481 13175
rect 5868 13144 7481 13172
rect 5868 13132 5874 13144
rect 7469 13141 7481 13144
rect 7515 13172 7527 13175
rect 7834 13172 7840 13184
rect 7515 13144 7840 13172
rect 7515 13141 7527 13144
rect 7469 13135 7527 13141
rect 7834 13132 7840 13144
rect 7892 13132 7898 13184
rect 8389 13175 8447 13181
rect 8389 13141 8401 13175
rect 8435 13172 8447 13175
rect 9122 13172 9128 13184
rect 8435 13144 9128 13172
rect 8435 13141 8447 13144
rect 8389 13135 8447 13141
rect 9122 13132 9128 13144
rect 9180 13172 9186 13184
rect 9398 13172 9404 13184
rect 9180 13144 9404 13172
rect 9180 13132 9186 13144
rect 9398 13132 9404 13144
rect 9456 13132 9462 13184
rect 9858 13172 9864 13184
rect 9819 13144 9864 13172
rect 9858 13132 9864 13144
rect 9916 13132 9922 13184
rect 9950 13132 9956 13184
rect 10008 13172 10014 13184
rect 10321 13175 10379 13181
rect 10008 13144 10053 13172
rect 10008 13132 10014 13144
rect 10321 13141 10333 13175
rect 10367 13172 10379 13175
rect 11238 13172 11244 13184
rect 10367 13144 11244 13172
rect 10367 13141 10379 13144
rect 10321 13135 10379 13141
rect 11238 13132 11244 13144
rect 11296 13132 11302 13184
rect 11698 13172 11704 13184
rect 11659 13144 11704 13172
rect 11698 13132 11704 13144
rect 11756 13132 11762 13184
rect 12452 13172 12480 13348
rect 14734 13336 14740 13388
rect 14792 13376 14798 13388
rect 15105 13379 15163 13385
rect 15105 13376 15117 13379
rect 14792 13348 15117 13376
rect 14792 13336 14798 13348
rect 15105 13345 15117 13348
rect 15151 13345 15163 13379
rect 15105 13339 15163 13345
rect 12894 13268 12900 13320
rect 12952 13308 12958 13320
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 12952 13280 14105 13308
rect 12952 13268 12958 13280
rect 14093 13277 14105 13280
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 15746 13268 15752 13320
rect 15804 13268 15810 13320
rect 16942 13268 16948 13320
rect 17000 13308 17006 13320
rect 17681 13311 17739 13317
rect 17681 13308 17693 13311
rect 17000 13280 17693 13308
rect 17000 13268 17006 13280
rect 17681 13277 17693 13280
rect 17727 13277 17739 13311
rect 17681 13271 17739 13277
rect 12612 13243 12670 13249
rect 12612 13209 12624 13243
rect 12658 13240 12670 13243
rect 14737 13243 14795 13249
rect 14737 13240 14749 13243
rect 12658 13212 14749 13240
rect 12658 13209 12670 13212
rect 12612 13203 12670 13209
rect 14737 13209 14749 13212
rect 14783 13209 14795 13243
rect 15764 13240 15792 13268
rect 15841 13243 15899 13249
rect 15841 13240 15853 13243
rect 14737 13203 14795 13209
rect 15396 13212 15853 13240
rect 15396 13184 15424 13212
rect 15841 13209 15853 13212
rect 15887 13209 15899 13243
rect 15841 13203 15899 13209
rect 17436 13243 17494 13249
rect 17436 13209 17448 13243
rect 17482 13240 17494 13243
rect 21358 13240 21364 13252
rect 17482 13212 21364 13240
rect 17482 13209 17494 13212
rect 17436 13203 17494 13209
rect 21358 13200 21364 13212
rect 21416 13200 21422 13252
rect 12802 13172 12808 13184
rect 12452 13144 12808 13172
rect 12802 13132 12808 13144
rect 12860 13132 12866 13184
rect 13170 13132 13176 13184
rect 13228 13172 13234 13184
rect 13722 13172 13728 13184
rect 13228 13144 13728 13172
rect 13228 13132 13234 13144
rect 13722 13132 13728 13144
rect 13780 13132 13786 13184
rect 14921 13175 14979 13181
rect 14921 13141 14933 13175
rect 14967 13172 14979 13175
rect 15194 13172 15200 13184
rect 14967 13144 15200 13172
rect 14967 13141 14979 13144
rect 14921 13135 14979 13141
rect 15194 13132 15200 13144
rect 15252 13172 15258 13184
rect 15289 13175 15347 13181
rect 15289 13172 15301 13175
rect 15252 13144 15301 13172
rect 15252 13132 15258 13144
rect 15289 13141 15301 13144
rect 15335 13141 15347 13175
rect 15289 13135 15347 13141
rect 15378 13132 15384 13184
rect 15436 13172 15442 13184
rect 15436 13144 15481 13172
rect 15436 13132 15442 13144
rect 1104 13082 21896 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21896 13082
rect 1104 13008 21896 13030
rect 1854 12968 1860 12980
rect 1815 12940 1860 12968
rect 1854 12928 1860 12940
rect 1912 12928 1918 12980
rect 1949 12971 2007 12977
rect 1949 12937 1961 12971
rect 1995 12937 2007 12971
rect 1949 12931 2007 12937
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 1964 12832 1992 12931
rect 2130 12928 2136 12980
rect 2188 12968 2194 12980
rect 2317 12971 2375 12977
rect 2317 12968 2329 12971
rect 2188 12940 2329 12968
rect 2188 12928 2194 12940
rect 2317 12937 2329 12940
rect 2363 12937 2375 12971
rect 2317 12931 2375 12937
rect 2409 12971 2467 12977
rect 2409 12937 2421 12971
rect 2455 12968 2467 12971
rect 2777 12971 2835 12977
rect 2777 12968 2789 12971
rect 2455 12940 2789 12968
rect 2455 12937 2467 12940
rect 2409 12931 2467 12937
rect 2777 12937 2789 12940
rect 2823 12937 2835 12971
rect 2777 12931 2835 12937
rect 3237 12971 3295 12977
rect 3237 12937 3249 12971
rect 3283 12968 3295 12971
rect 3605 12971 3663 12977
rect 3605 12968 3617 12971
rect 3283 12940 3617 12968
rect 3283 12937 3295 12940
rect 3237 12931 3295 12937
rect 3605 12937 3617 12940
rect 3651 12937 3663 12971
rect 3605 12931 3663 12937
rect 5810 12928 5816 12980
rect 5868 12968 5874 12980
rect 6365 12971 6423 12977
rect 6365 12968 6377 12971
rect 5868 12940 6377 12968
rect 5868 12928 5874 12940
rect 6365 12937 6377 12940
rect 6411 12937 6423 12971
rect 6365 12931 6423 12937
rect 6549 12971 6607 12977
rect 6549 12937 6561 12971
rect 6595 12968 6607 12971
rect 6730 12968 6736 12980
rect 6595 12940 6736 12968
rect 6595 12937 6607 12940
rect 6549 12931 6607 12937
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 6917 12971 6975 12977
rect 6917 12937 6929 12971
rect 6963 12968 6975 12971
rect 7742 12968 7748 12980
rect 6963 12940 7748 12968
rect 6963 12937 6975 12940
rect 6917 12931 6975 12937
rect 7742 12928 7748 12940
rect 7800 12928 7806 12980
rect 7834 12928 7840 12980
rect 7892 12968 7898 12980
rect 11146 12968 11152 12980
rect 7892 12940 11152 12968
rect 7892 12928 7898 12940
rect 11146 12928 11152 12940
rect 11204 12928 11210 12980
rect 11698 12968 11704 12980
rect 11532 12940 11704 12968
rect 2590 12860 2596 12912
rect 2648 12900 2654 12912
rect 4065 12903 4123 12909
rect 4065 12900 4077 12903
rect 2648 12872 4077 12900
rect 2648 12860 2654 12872
rect 4065 12869 4077 12872
rect 4111 12869 4123 12903
rect 5718 12900 5724 12912
rect 4065 12863 4123 12869
rect 4816 12872 5724 12900
rect 3142 12832 3148 12844
rect 1719 12804 1992 12832
rect 3103 12804 3148 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 3142 12792 3148 12804
rect 3200 12792 3206 12844
rect 4816 12841 4844 12872
rect 5718 12860 5724 12872
rect 5776 12860 5782 12912
rect 7926 12900 7932 12912
rect 7392 12872 7932 12900
rect 3973 12835 4031 12841
rect 3973 12801 3985 12835
rect 4019 12832 4031 12835
rect 4801 12835 4859 12841
rect 4019 12804 4568 12832
rect 4019 12801 4031 12804
rect 3973 12795 4031 12801
rect 2590 12764 2596 12776
rect 2551 12736 2596 12764
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 3329 12767 3387 12773
rect 3329 12733 3341 12767
rect 3375 12733 3387 12767
rect 3329 12727 3387 12733
rect 4157 12767 4215 12773
rect 4157 12733 4169 12767
rect 4203 12733 4215 12767
rect 4157 12727 4215 12733
rect 2222 12656 2228 12708
rect 2280 12696 2286 12708
rect 3344 12696 3372 12727
rect 4172 12696 4200 12727
rect 4540 12705 4568 12804
rect 4801 12801 4813 12835
rect 4847 12801 4859 12835
rect 4801 12795 4859 12801
rect 4890 12792 4896 12844
rect 4948 12832 4954 12844
rect 5057 12835 5115 12841
rect 5057 12832 5069 12835
rect 4948 12804 5069 12832
rect 4948 12792 4954 12804
rect 5057 12801 5069 12804
rect 5103 12832 5115 12835
rect 7392 12832 7420 12872
rect 7926 12860 7932 12872
rect 7984 12900 7990 12912
rect 8662 12900 8668 12912
rect 7984 12872 8668 12900
rect 7984 12860 7990 12872
rect 8662 12860 8668 12872
rect 8720 12860 8726 12912
rect 11330 12900 11336 12912
rect 9324 12872 11336 12900
rect 9324 12844 9352 12872
rect 11330 12860 11336 12872
rect 11388 12900 11394 12912
rect 11532 12900 11560 12940
rect 11698 12928 11704 12940
rect 11756 12928 11762 12980
rect 12894 12968 12900 12980
rect 12855 12940 12900 12968
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 13354 12968 13360 12980
rect 13315 12940 13360 12968
rect 13354 12928 13360 12940
rect 13412 12928 13418 12980
rect 13446 12928 13452 12980
rect 13504 12968 13510 12980
rect 13725 12971 13783 12977
rect 13725 12968 13737 12971
rect 13504 12940 13737 12968
rect 13504 12928 13510 12940
rect 13725 12937 13737 12940
rect 13771 12937 13783 12971
rect 13725 12931 13783 12937
rect 14277 12971 14335 12977
rect 14277 12937 14289 12971
rect 14323 12968 14335 12971
rect 14642 12968 14648 12980
rect 14323 12940 14648 12968
rect 14323 12937 14335 12940
rect 14277 12931 14335 12937
rect 14642 12928 14648 12940
rect 14700 12928 14706 12980
rect 14737 12971 14795 12977
rect 14737 12937 14749 12971
rect 14783 12968 14795 12971
rect 15105 12971 15163 12977
rect 15105 12968 15117 12971
rect 14783 12940 15117 12968
rect 14783 12937 14795 12940
rect 14737 12931 14795 12937
rect 15105 12937 15117 12940
rect 15151 12937 15163 12971
rect 15470 12968 15476 12980
rect 15431 12940 15476 12968
rect 15105 12931 15163 12937
rect 15470 12928 15476 12940
rect 15528 12928 15534 12980
rect 15562 12928 15568 12980
rect 15620 12968 15626 12980
rect 15620 12940 15665 12968
rect 15620 12928 15626 12940
rect 16390 12900 16396 12912
rect 11388 12872 11560 12900
rect 11388 12860 11394 12872
rect 5103 12804 7420 12832
rect 5103 12801 5115 12804
rect 5057 12795 5115 12801
rect 7466 12792 7472 12844
rect 7524 12832 7530 12844
rect 7633 12835 7691 12841
rect 7633 12832 7645 12835
rect 7524 12804 7645 12832
rect 7524 12792 7530 12804
rect 7633 12801 7645 12804
rect 7679 12801 7691 12835
rect 7633 12795 7691 12801
rect 8202 12792 8208 12844
rect 8260 12832 8266 12844
rect 8478 12832 8484 12844
rect 8260 12804 8484 12832
rect 8260 12792 8266 12804
rect 8478 12792 8484 12804
rect 8536 12792 8542 12844
rect 9217 12835 9275 12841
rect 9217 12801 9229 12835
rect 9263 12832 9275 12835
rect 9306 12832 9312 12844
rect 9263 12804 9312 12832
rect 9263 12801 9275 12804
rect 9217 12795 9275 12801
rect 9306 12792 9312 12804
rect 9364 12792 9370 12844
rect 9490 12841 9496 12844
rect 9484 12795 9496 12841
rect 9548 12832 9554 12844
rect 11532 12841 11560 12872
rect 11624 12872 16396 12900
rect 11517 12835 11575 12841
rect 9548 12804 9584 12832
rect 9490 12792 9496 12795
rect 9548 12792 9554 12804
rect 11517 12801 11529 12835
rect 11563 12801 11575 12835
rect 11517 12795 11575 12801
rect 7006 12764 7012 12776
rect 6967 12736 7012 12764
rect 7006 12724 7012 12736
rect 7064 12724 7070 12776
rect 7190 12764 7196 12776
rect 7151 12736 7196 12764
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 7377 12767 7435 12773
rect 7377 12733 7389 12767
rect 7423 12733 7435 12767
rect 7377 12727 7435 12733
rect 2280 12668 3372 12696
rect 4080 12668 4200 12696
rect 4525 12699 4583 12705
rect 2280 12656 2286 12668
rect 4080 12640 4108 12668
rect 4525 12665 4537 12699
rect 4571 12696 4583 12699
rect 4798 12696 4804 12708
rect 4571 12668 4804 12696
rect 4571 12665 4583 12668
rect 4525 12659 4583 12665
rect 4798 12656 4804 12668
rect 4856 12656 4862 12708
rect 6181 12699 6239 12705
rect 6181 12665 6193 12699
rect 6227 12696 6239 12699
rect 6546 12696 6552 12708
rect 6227 12668 6552 12696
rect 6227 12665 6239 12668
rect 6181 12659 6239 12665
rect 6546 12656 6552 12668
rect 6604 12656 6610 12708
rect 6822 12656 6828 12708
rect 6880 12696 6886 12708
rect 7392 12696 7420 12727
rect 11054 12724 11060 12776
rect 11112 12764 11118 12776
rect 11624 12764 11652 12872
rect 16390 12860 16396 12872
rect 16448 12860 16454 12912
rect 11784 12835 11842 12841
rect 11784 12801 11796 12835
rect 11830 12832 11842 12835
rect 12066 12832 12072 12844
rect 11830 12804 12072 12832
rect 11830 12801 11842 12804
rect 11784 12795 11842 12801
rect 12066 12792 12072 12804
rect 12124 12792 12130 12844
rect 14645 12835 14703 12841
rect 14645 12801 14657 12835
rect 14691 12832 14703 12835
rect 15746 12832 15752 12844
rect 14691 12804 15752 12832
rect 14691 12801 14703 12804
rect 14645 12795 14703 12801
rect 15746 12792 15752 12804
rect 15804 12792 15810 12844
rect 13170 12764 13176 12776
rect 11112 12736 11652 12764
rect 13131 12736 13176 12764
rect 11112 12724 11118 12736
rect 13170 12724 13176 12736
rect 13228 12724 13234 12776
rect 13265 12767 13323 12773
rect 13265 12733 13277 12767
rect 13311 12764 13323 12767
rect 13446 12764 13452 12776
rect 13311 12736 13452 12764
rect 13311 12733 13323 12736
rect 13265 12727 13323 12733
rect 13446 12724 13452 12736
rect 13504 12724 13510 12776
rect 14458 12724 14464 12776
rect 14516 12764 14522 12776
rect 14829 12767 14887 12773
rect 14829 12764 14841 12767
rect 14516 12736 14841 12764
rect 14516 12724 14522 12736
rect 14829 12733 14841 12736
rect 14875 12733 14887 12767
rect 14829 12727 14887 12733
rect 15562 12724 15568 12776
rect 15620 12764 15626 12776
rect 15657 12767 15715 12773
rect 15657 12764 15669 12767
rect 15620 12736 15669 12764
rect 15620 12724 15626 12736
rect 15657 12733 15669 12736
rect 15703 12733 15715 12767
rect 15657 12727 15715 12733
rect 9214 12696 9220 12708
rect 6880 12668 7420 12696
rect 8312 12668 9220 12696
rect 6880 12656 6886 12668
rect 1578 12628 1584 12640
rect 1539 12600 1584 12628
rect 1578 12588 1584 12600
rect 1636 12588 1642 12640
rect 4062 12588 4068 12640
rect 4120 12588 4126 12640
rect 4709 12631 4767 12637
rect 4709 12597 4721 12631
rect 4755 12628 4767 12631
rect 5074 12628 5080 12640
rect 4755 12600 5080 12628
rect 4755 12597 4767 12600
rect 4709 12591 4767 12597
rect 5074 12588 5080 12600
rect 5132 12588 5138 12640
rect 6638 12588 6644 12640
rect 6696 12628 6702 12640
rect 8312 12628 8340 12668
rect 9214 12656 9220 12668
rect 9272 12656 9278 12708
rect 15194 12696 15200 12708
rect 13280 12668 15200 12696
rect 6696 12600 8340 12628
rect 6696 12588 6702 12600
rect 8662 12588 8668 12640
rect 8720 12628 8726 12640
rect 8757 12631 8815 12637
rect 8757 12628 8769 12631
rect 8720 12600 8769 12628
rect 8720 12588 8726 12600
rect 8757 12597 8769 12600
rect 8803 12597 8815 12631
rect 10594 12628 10600 12640
rect 10555 12600 10600 12628
rect 8757 12591 8815 12597
rect 10594 12588 10600 12600
rect 10652 12588 10658 12640
rect 11698 12588 11704 12640
rect 11756 12628 11762 12640
rect 13280 12628 13308 12668
rect 15194 12656 15200 12668
rect 15252 12656 15258 12708
rect 11756 12600 13308 12628
rect 11756 12588 11762 12600
rect 13354 12588 13360 12640
rect 13412 12628 13418 12640
rect 14826 12628 14832 12640
rect 13412 12600 14832 12628
rect 13412 12588 13418 12600
rect 14826 12588 14832 12600
rect 14884 12588 14890 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 2958 12424 2964 12436
rect 1688 12396 2964 12424
rect 1688 12232 1716 12396
rect 2958 12384 2964 12396
rect 3016 12384 3022 12436
rect 3326 12384 3332 12436
rect 3384 12424 3390 12436
rect 3421 12427 3479 12433
rect 3421 12424 3433 12427
rect 3384 12396 3433 12424
rect 3384 12384 3390 12396
rect 3421 12393 3433 12396
rect 3467 12393 3479 12427
rect 5445 12427 5503 12433
rect 3421 12387 3479 12393
rect 4080 12396 5396 12424
rect 4080 12288 4108 12396
rect 5368 12356 5396 12396
rect 5445 12393 5457 12427
rect 5491 12424 5503 12427
rect 5534 12424 5540 12436
rect 5491 12396 5540 12424
rect 5491 12393 5503 12396
rect 5445 12387 5503 12393
rect 5534 12384 5540 12396
rect 5592 12384 5598 12436
rect 6638 12424 6644 12436
rect 5920 12396 6644 12424
rect 5920 12356 5948 12396
rect 6638 12384 6644 12396
rect 6696 12384 6702 12436
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 7374 12424 7380 12436
rect 7064 12396 7380 12424
rect 7064 12384 7070 12396
rect 7374 12384 7380 12396
rect 7432 12384 7438 12436
rect 7650 12384 7656 12436
rect 7708 12424 7714 12436
rect 8573 12427 8631 12433
rect 8573 12424 8585 12427
rect 7708 12396 8585 12424
rect 7708 12384 7714 12396
rect 8573 12393 8585 12396
rect 8619 12424 8631 12427
rect 8619 12396 9076 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 9048 12368 9076 12396
rect 9490 12384 9496 12436
rect 9548 12424 9554 12436
rect 9585 12427 9643 12433
rect 9585 12424 9597 12427
rect 9548 12396 9597 12424
rect 9548 12384 9554 12396
rect 9585 12393 9597 12396
rect 9631 12393 9643 12427
rect 9585 12387 9643 12393
rect 9677 12427 9735 12433
rect 9677 12393 9689 12427
rect 9723 12424 9735 12427
rect 9858 12424 9864 12436
rect 9723 12396 9864 12424
rect 9723 12393 9735 12396
rect 9677 12387 9735 12393
rect 9858 12384 9864 12396
rect 9916 12384 9922 12436
rect 10502 12424 10508 12436
rect 10463 12396 10508 12424
rect 10502 12384 10508 12396
rect 10560 12424 10566 12436
rect 12066 12424 12072 12436
rect 10560 12396 12072 12424
rect 10560 12384 10566 12396
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 12710 12424 12716 12436
rect 12671 12396 12716 12424
rect 12710 12384 12716 12396
rect 12768 12384 12774 12436
rect 14642 12384 14648 12436
rect 14700 12424 14706 12436
rect 15010 12424 15016 12436
rect 14700 12396 15016 12424
rect 14700 12384 14706 12396
rect 15010 12384 15016 12396
rect 15068 12384 15074 12436
rect 5368 12328 5948 12356
rect 8386 12316 8392 12368
rect 8444 12356 8450 12368
rect 8754 12356 8760 12368
rect 8444 12328 8760 12356
rect 8444 12316 8450 12328
rect 8754 12316 8760 12328
rect 8812 12316 8818 12368
rect 9030 12316 9036 12368
rect 9088 12316 9094 12368
rect 10778 12356 10784 12368
rect 10244 12328 10784 12356
rect 5534 12288 5540 12300
rect 3252 12260 4108 12288
rect 5495 12260 5540 12288
rect 1397 12223 1455 12229
rect 1397 12189 1409 12223
rect 1443 12220 1455 12223
rect 1486 12220 1492 12232
rect 1443 12192 1492 12220
rect 1443 12189 1455 12192
rect 1397 12183 1455 12189
rect 1486 12180 1492 12192
rect 1544 12180 1550 12232
rect 1670 12220 1676 12232
rect 1631 12192 1676 12220
rect 1670 12180 1676 12192
rect 1728 12180 1734 12232
rect 3252 12220 3280 12260
rect 5534 12248 5540 12260
rect 5592 12248 5598 12300
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12288 7987 12291
rect 8478 12288 8484 12300
rect 7975 12260 8484 12288
rect 7975 12257 7987 12260
rect 7929 12251 7987 12257
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 10244 12288 10272 12328
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 12084 12356 12112 12384
rect 12084 12328 13400 12356
rect 8588 12260 10272 12288
rect 10321 12291 10379 12297
rect 2746 12192 3280 12220
rect 2746 12152 2774 12192
rect 3326 12180 3332 12232
rect 3384 12220 3390 12232
rect 4065 12223 4123 12229
rect 4065 12220 4077 12223
rect 3384 12192 4077 12220
rect 3384 12180 3390 12192
rect 4065 12189 4077 12192
rect 4111 12220 4123 12223
rect 5718 12220 5724 12232
rect 4111 12192 5724 12220
rect 4111 12189 4123 12192
rect 4065 12183 4123 12189
rect 5718 12180 5724 12192
rect 5776 12220 5782 12232
rect 5905 12223 5963 12229
rect 5905 12220 5917 12223
rect 5776 12192 5917 12220
rect 5776 12180 5782 12192
rect 5905 12189 5917 12192
rect 5951 12220 5963 12223
rect 8588 12220 8616 12260
rect 10321 12257 10333 12291
rect 10367 12288 10379 12291
rect 10594 12288 10600 12300
rect 10367 12260 10600 12288
rect 10367 12257 10379 12260
rect 10321 12251 10379 12257
rect 10594 12248 10600 12260
rect 10652 12248 10658 12300
rect 12161 12291 12219 12297
rect 12161 12257 12173 12291
rect 12207 12288 12219 12291
rect 12894 12288 12900 12300
rect 12207 12260 12900 12288
rect 12207 12257 12219 12260
rect 12161 12251 12219 12257
rect 12894 12248 12900 12260
rect 12952 12248 12958 12300
rect 13372 12297 13400 12328
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12257 13415 12291
rect 13357 12251 13415 12257
rect 5951 12192 6868 12220
rect 5951 12189 5963 12192
rect 5905 12183 5963 12189
rect 6840 12164 6868 12192
rect 7116 12192 8616 12220
rect 1596 12124 2774 12152
rect 3084 12155 3142 12161
rect 1596 12093 1624 12124
rect 3084 12121 3096 12155
rect 3130 12152 3142 12155
rect 3130 12124 4108 12152
rect 3130 12121 3142 12124
rect 3084 12115 3142 12121
rect 4080 12096 4108 12124
rect 4154 12112 4160 12164
rect 4212 12152 4218 12164
rect 4310 12155 4368 12161
rect 4310 12152 4322 12155
rect 4212 12124 4322 12152
rect 4212 12112 4218 12124
rect 4310 12121 4322 12124
rect 4356 12121 4368 12155
rect 4310 12115 4368 12121
rect 5626 12112 5632 12164
rect 5684 12152 5690 12164
rect 6150 12155 6208 12161
rect 6150 12152 6162 12155
rect 5684 12124 6162 12152
rect 5684 12112 5690 12124
rect 6150 12121 6162 12124
rect 6196 12152 6208 12155
rect 6546 12152 6552 12164
rect 6196 12124 6552 12152
rect 6196 12121 6208 12124
rect 6150 12115 6208 12121
rect 6546 12112 6552 12124
rect 6604 12112 6610 12164
rect 6822 12112 6828 12164
rect 6880 12112 6886 12164
rect 1581 12087 1639 12093
rect 1581 12053 1593 12087
rect 1627 12053 1639 12087
rect 1854 12084 1860 12096
rect 1815 12056 1860 12084
rect 1581 12047 1639 12053
rect 1854 12044 1860 12056
rect 1912 12044 1918 12096
rect 1946 12044 1952 12096
rect 2004 12084 2010 12096
rect 2004 12056 2049 12084
rect 2004 12044 2010 12056
rect 2314 12044 2320 12096
rect 2372 12084 2378 12096
rect 2590 12084 2596 12096
rect 2372 12056 2596 12084
rect 2372 12044 2378 12056
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 2958 12044 2964 12096
rect 3016 12084 3022 12096
rect 3789 12087 3847 12093
rect 3789 12084 3801 12087
rect 3016 12056 3801 12084
rect 3016 12044 3022 12056
rect 3789 12053 3801 12056
rect 3835 12053 3847 12087
rect 3789 12047 3847 12053
rect 4062 12044 4068 12096
rect 4120 12044 4126 12096
rect 4706 12044 4712 12096
rect 4764 12084 4770 12096
rect 7116 12084 7144 12192
rect 8662 12180 8668 12232
rect 8720 12220 8726 12232
rect 8941 12223 8999 12229
rect 8941 12220 8953 12223
rect 8720 12192 8953 12220
rect 8720 12180 8726 12192
rect 8941 12189 8953 12192
rect 8987 12189 8999 12223
rect 11054 12220 11060 12232
rect 8941 12183 8999 12189
rect 9416 12192 11060 12220
rect 8021 12155 8079 12161
rect 8021 12121 8033 12155
rect 8067 12152 8079 12155
rect 8386 12152 8392 12164
rect 8067 12124 8392 12152
rect 8067 12121 8079 12124
rect 8021 12115 8079 12121
rect 8386 12112 8392 12124
rect 8444 12112 8450 12164
rect 9416 12152 9444 12192
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 11330 12180 11336 12232
rect 11388 12220 11394 12232
rect 11885 12223 11943 12229
rect 11885 12220 11897 12223
rect 11388 12192 11897 12220
rect 11388 12180 11394 12192
rect 11885 12189 11897 12192
rect 11931 12220 11943 12223
rect 14277 12223 14335 12229
rect 14277 12220 14289 12223
rect 11931 12192 14289 12220
rect 11931 12189 11943 12192
rect 11885 12183 11943 12189
rect 14277 12189 14289 12192
rect 14323 12220 14335 12223
rect 14323 12192 14872 12220
rect 14323 12189 14335 12192
rect 14277 12183 14335 12189
rect 8496 12124 9444 12152
rect 7282 12084 7288 12096
rect 4764 12056 7144 12084
rect 7243 12056 7288 12084
rect 4764 12044 4770 12056
rect 7282 12044 7288 12056
rect 7340 12044 7346 12096
rect 8110 12084 8116 12096
rect 8071 12056 8116 12084
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 8496 12093 8524 12124
rect 9490 12112 9496 12164
rect 9548 12152 9554 12164
rect 10137 12155 10195 12161
rect 10137 12152 10149 12155
rect 9548 12124 10149 12152
rect 9548 12112 9554 12124
rect 10137 12121 10149 12124
rect 10183 12121 10195 12155
rect 10137 12115 10195 12121
rect 10594 12112 10600 12164
rect 10652 12152 10658 12164
rect 11618 12155 11676 12161
rect 11618 12152 11630 12155
rect 10652 12124 11630 12152
rect 10652 12112 10658 12124
rect 11618 12121 11630 12124
rect 11664 12121 11676 12155
rect 11618 12115 11676 12121
rect 13173 12155 13231 12161
rect 13173 12121 13185 12155
rect 13219 12152 13231 12155
rect 13538 12152 13544 12164
rect 13219 12124 13544 12152
rect 13219 12121 13231 12124
rect 13173 12115 13231 12121
rect 13538 12112 13544 12124
rect 13596 12112 13602 12164
rect 14544 12155 14602 12161
rect 14544 12121 14556 12155
rect 14590 12152 14602 12155
rect 14734 12152 14740 12164
rect 14590 12124 14740 12152
rect 14590 12121 14602 12124
rect 14544 12115 14602 12121
rect 14734 12112 14740 12124
rect 14792 12112 14798 12164
rect 14844 12152 14872 12192
rect 14918 12180 14924 12232
rect 14976 12220 14982 12232
rect 15749 12223 15807 12229
rect 15749 12220 15761 12223
rect 14976 12192 15761 12220
rect 14976 12180 14982 12192
rect 15749 12189 15761 12192
rect 15795 12189 15807 12223
rect 15749 12183 15807 12189
rect 16942 12152 16948 12164
rect 14844 12124 16948 12152
rect 16942 12112 16948 12124
rect 17000 12112 17006 12164
rect 8481 12087 8539 12093
rect 8481 12053 8493 12087
rect 8527 12053 8539 12087
rect 10042 12084 10048 12096
rect 10003 12056 10048 12084
rect 8481 12047 8539 12053
rect 10042 12044 10048 12056
rect 10100 12044 10106 12096
rect 11238 12044 11244 12096
rect 11296 12084 11302 12096
rect 12253 12087 12311 12093
rect 12253 12084 12265 12087
rect 11296 12056 12265 12084
rect 11296 12044 11302 12056
rect 12253 12053 12265 12056
rect 12299 12053 12311 12087
rect 12253 12047 12311 12053
rect 12345 12087 12403 12093
rect 12345 12053 12357 12087
rect 12391 12084 12403 12087
rect 12805 12087 12863 12093
rect 12805 12084 12817 12087
rect 12391 12056 12817 12084
rect 12391 12053 12403 12056
rect 12345 12047 12403 12053
rect 12805 12053 12817 12056
rect 12851 12053 12863 12087
rect 13262 12084 13268 12096
rect 13223 12056 13268 12084
rect 12805 12047 12863 12053
rect 13262 12044 13268 12056
rect 13320 12044 13326 12096
rect 15562 12044 15568 12096
rect 15620 12084 15626 12096
rect 15657 12087 15715 12093
rect 15657 12084 15669 12087
rect 15620 12056 15669 12084
rect 15620 12044 15626 12056
rect 15657 12053 15669 12056
rect 15703 12053 15715 12087
rect 16390 12084 16396 12096
rect 16351 12056 16396 12084
rect 15657 12047 15715 12053
rect 16390 12044 16396 12056
rect 16448 12044 16454 12096
rect 1104 11994 21896 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21896 11994
rect 1104 11920 21896 11942
rect 1489 11883 1547 11889
rect 1489 11849 1501 11883
rect 1535 11880 1547 11883
rect 2314 11880 2320 11892
rect 1535 11852 2320 11880
rect 1535 11849 1547 11852
rect 1489 11843 1547 11849
rect 2314 11840 2320 11852
rect 2372 11880 2378 11892
rect 2372 11852 3004 11880
rect 2372 11840 2378 11852
rect 1946 11772 1952 11824
rect 2004 11812 2010 11824
rect 2222 11812 2228 11824
rect 2004 11784 2228 11812
rect 2004 11772 2010 11784
rect 2222 11772 2228 11784
rect 2280 11812 2286 11824
rect 2602 11815 2660 11821
rect 2602 11812 2614 11815
rect 2280 11784 2614 11812
rect 2280 11772 2286 11784
rect 2602 11781 2614 11784
rect 2648 11781 2660 11815
rect 2602 11775 2660 11781
rect 2976 11753 3004 11852
rect 3142 11840 3148 11892
rect 3200 11880 3206 11892
rect 3697 11883 3755 11889
rect 3697 11880 3709 11883
rect 3200 11852 3709 11880
rect 3200 11840 3206 11852
rect 3697 11849 3709 11852
rect 3743 11849 3755 11883
rect 3697 11843 3755 11849
rect 4157 11883 4215 11889
rect 4157 11849 4169 11883
rect 4203 11880 4215 11883
rect 4706 11880 4712 11892
rect 4203 11852 4712 11880
rect 4203 11849 4215 11852
rect 4157 11843 4215 11849
rect 4706 11840 4712 11852
rect 4764 11840 4770 11892
rect 4801 11883 4859 11889
rect 4801 11849 4813 11883
rect 4847 11880 4859 11883
rect 5166 11880 5172 11892
rect 4847 11852 5172 11880
rect 4847 11849 4859 11852
rect 4801 11843 4859 11849
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11713 2927 11747
rect 2869 11707 2927 11713
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11713 3019 11747
rect 2961 11707 3019 11713
rect 4065 11747 4123 11753
rect 4065 11713 4077 11747
rect 4111 11744 4123 11747
rect 4816 11744 4844 11843
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 5813 11883 5871 11889
rect 5813 11849 5825 11883
rect 5859 11849 5871 11883
rect 5813 11843 5871 11849
rect 6825 11883 6883 11889
rect 6825 11849 6837 11883
rect 6871 11880 6883 11883
rect 7098 11880 7104 11892
rect 6871 11852 7104 11880
rect 6871 11849 6883 11852
rect 6825 11843 6883 11849
rect 5626 11812 5632 11824
rect 4111 11716 4844 11744
rect 5184 11784 5632 11812
rect 4111 11713 4123 11716
rect 4065 11707 4123 11713
rect 2884 11676 2912 11707
rect 3326 11676 3332 11688
rect 2884 11648 3332 11676
rect 3326 11636 3332 11648
rect 3384 11636 3390 11688
rect 4249 11679 4307 11685
rect 4249 11676 4261 11679
rect 4080 11648 4261 11676
rect 4080 11620 4108 11648
rect 4249 11645 4261 11648
rect 4295 11645 4307 11679
rect 4249 11639 4307 11645
rect 3050 11608 3056 11620
rect 2884 11580 3056 11608
rect 1854 11500 1860 11552
rect 1912 11540 1918 11552
rect 2884 11540 2912 11580
rect 3050 11568 3056 11580
rect 3108 11608 3114 11620
rect 4062 11608 4068 11620
rect 3108 11580 4068 11608
rect 3108 11568 3114 11580
rect 4062 11568 4068 11580
rect 4120 11568 4126 11620
rect 1912 11512 2912 11540
rect 1912 11500 1918 11512
rect 2958 11500 2964 11552
rect 3016 11540 3022 11552
rect 3605 11543 3663 11549
rect 3605 11540 3617 11543
rect 3016 11512 3617 11540
rect 3016 11500 3022 11512
rect 3605 11509 3617 11512
rect 3651 11509 3663 11543
rect 3605 11503 3663 11509
rect 4246 11500 4252 11552
rect 4304 11540 4310 11552
rect 4356 11540 4384 11716
rect 5184 11685 5212 11784
rect 5626 11772 5632 11784
rect 5684 11772 5690 11824
rect 5828 11812 5856 11843
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 7285 11883 7343 11889
rect 7285 11849 7297 11883
rect 7331 11849 7343 11883
rect 7285 11843 7343 11849
rect 6917 11815 6975 11821
rect 6917 11812 6929 11815
rect 5828 11784 6929 11812
rect 6917 11781 6929 11784
rect 6963 11781 6975 11815
rect 7300 11812 7328 11843
rect 7558 11840 7564 11892
rect 7616 11880 7622 11892
rect 8205 11883 8263 11889
rect 8205 11880 8217 11883
rect 7616 11852 8217 11880
rect 7616 11840 7622 11852
rect 8205 11849 8217 11852
rect 8251 11849 8263 11883
rect 8205 11843 8263 11849
rect 8297 11883 8355 11889
rect 8297 11849 8309 11883
rect 8343 11880 8355 11883
rect 8570 11880 8576 11892
rect 8343 11852 8576 11880
rect 8343 11849 8355 11852
rect 8297 11843 8355 11849
rect 8570 11840 8576 11852
rect 8628 11840 8634 11892
rect 9030 11880 9036 11892
rect 8991 11852 9036 11880
rect 9030 11840 9036 11852
rect 9088 11840 9094 11892
rect 9122 11840 9128 11892
rect 9180 11880 9186 11892
rect 9490 11880 9496 11892
rect 9180 11852 9225 11880
rect 9451 11852 9496 11880
rect 9180 11840 9186 11852
rect 9490 11840 9496 11852
rect 9548 11840 9554 11892
rect 10045 11883 10103 11889
rect 10045 11849 10057 11883
rect 10091 11880 10103 11883
rect 10410 11880 10416 11892
rect 10091 11852 10416 11880
rect 10091 11849 10103 11852
rect 10045 11843 10103 11849
rect 10410 11840 10416 11852
rect 10468 11840 10474 11892
rect 11885 11883 11943 11889
rect 11885 11849 11897 11883
rect 11931 11880 11943 11883
rect 13173 11883 13231 11889
rect 13173 11880 13185 11883
rect 11931 11852 13185 11880
rect 11931 11849 11943 11852
rect 11885 11843 11943 11849
rect 13173 11849 13185 11852
rect 13219 11849 13231 11883
rect 13538 11880 13544 11892
rect 13499 11852 13544 11880
rect 13173 11843 13231 11849
rect 13538 11840 13544 11852
rect 13596 11840 13602 11892
rect 14277 11883 14335 11889
rect 14277 11849 14289 11883
rect 14323 11880 14335 11883
rect 14458 11880 14464 11892
rect 14323 11852 14464 11880
rect 14323 11849 14335 11852
rect 14277 11843 14335 11849
rect 14458 11840 14464 11852
rect 14516 11880 14522 11892
rect 14918 11880 14924 11892
rect 14516 11852 14924 11880
rect 14516 11840 14522 11852
rect 14918 11840 14924 11852
rect 14976 11840 14982 11892
rect 15746 11880 15752 11892
rect 15707 11852 15752 11880
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 10226 11812 10232 11824
rect 7300 11784 10232 11812
rect 6917 11775 6975 11781
rect 10226 11772 10232 11784
rect 10284 11772 10290 11824
rect 11333 11815 11391 11821
rect 11333 11781 11345 11815
rect 11379 11812 11391 11815
rect 12158 11812 12164 11824
rect 11379 11784 12164 11812
rect 11379 11781 11391 11784
rect 11333 11775 11391 11781
rect 12158 11772 12164 11784
rect 12216 11772 12222 11824
rect 13725 11815 13783 11821
rect 13725 11781 13737 11815
rect 13771 11812 13783 11815
rect 13814 11812 13820 11824
rect 13771 11784 13820 11812
rect 13771 11781 13783 11784
rect 13725 11775 13783 11781
rect 13814 11772 13820 11784
rect 13872 11812 13878 11824
rect 14366 11812 14372 11824
rect 13872 11784 14372 11812
rect 13872 11772 13878 11784
rect 14366 11772 14372 11784
rect 14424 11772 14430 11824
rect 16942 11812 16948 11824
rect 15672 11784 16948 11812
rect 5442 11744 5448 11756
rect 5403 11716 5448 11744
rect 5442 11704 5448 11716
rect 5500 11704 5506 11756
rect 5534 11704 5540 11756
rect 5592 11744 5598 11756
rect 7006 11744 7012 11756
rect 5592 11716 7012 11744
rect 5592 11704 5598 11716
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 8662 11704 8668 11756
rect 8720 11744 8726 11756
rect 11790 11744 11796 11756
rect 8720 11716 8892 11744
rect 8720 11704 8726 11716
rect 5169 11679 5227 11685
rect 5169 11645 5181 11679
rect 5215 11645 5227 11679
rect 5350 11676 5356 11688
rect 5311 11648 5356 11676
rect 5169 11639 5227 11645
rect 5350 11636 5356 11648
rect 5408 11636 5414 11688
rect 5902 11676 5908 11688
rect 5863 11648 5908 11676
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 6733 11679 6791 11685
rect 6733 11645 6745 11679
rect 6779 11676 6791 11679
rect 7282 11676 7288 11688
rect 6779 11648 7288 11676
rect 6779 11645 6791 11648
rect 6733 11639 6791 11645
rect 7282 11636 7288 11648
rect 7340 11636 7346 11688
rect 7377 11679 7435 11685
rect 7377 11645 7389 11679
rect 7423 11645 7435 11679
rect 7377 11639 7435 11645
rect 8113 11679 8171 11685
rect 8113 11645 8125 11679
rect 8159 11676 8171 11679
rect 8202 11676 8208 11688
rect 8159 11648 8208 11676
rect 8159 11645 8171 11648
rect 8113 11639 8171 11645
rect 5810 11568 5816 11620
rect 5868 11608 5874 11620
rect 7392 11608 7420 11639
rect 8202 11636 8208 11648
rect 8260 11636 8266 11688
rect 8864 11685 8892 11716
rect 10520 11716 11796 11744
rect 8849 11679 8907 11685
rect 8849 11645 8861 11679
rect 8895 11645 8907 11679
rect 8849 11639 8907 11645
rect 9030 11636 9036 11688
rect 9088 11676 9094 11688
rect 10520 11676 10548 11716
rect 11790 11704 11796 11716
rect 11848 11704 11854 11756
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 12342 11744 12348 11756
rect 11940 11716 12204 11744
rect 12303 11716 12348 11744
rect 11940 11704 11946 11716
rect 9088 11648 10548 11676
rect 9088 11636 9094 11648
rect 10594 11636 10600 11688
rect 10652 11676 10658 11688
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 10652 11648 12081 11676
rect 10652 11636 10658 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 12176 11676 12204 11716
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 15401 11747 15459 11753
rect 12544 11716 12940 11744
rect 12250 11676 12256 11688
rect 12176 11648 12256 11676
rect 12069 11639 12127 11645
rect 5868 11580 7420 11608
rect 5868 11568 5874 11580
rect 7558 11568 7564 11620
rect 7616 11608 7622 11620
rect 12084 11608 12112 11639
rect 12250 11636 12256 11648
rect 12308 11676 12314 11688
rect 12308 11648 12401 11676
rect 12308 11636 12314 11648
rect 12544 11608 12572 11716
rect 12912 11685 12940 11716
rect 15401 11713 15413 11747
rect 15447 11744 15459 11747
rect 15562 11744 15568 11756
rect 15447 11716 15568 11744
rect 15447 11713 15459 11716
rect 15401 11707 15459 11713
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 15672 11753 15700 11784
rect 16942 11772 16948 11784
rect 17000 11772 17006 11824
rect 15657 11747 15715 11753
rect 15657 11713 15669 11747
rect 15703 11713 15715 11747
rect 16114 11744 16120 11756
rect 16075 11716 16120 11744
rect 15657 11707 15715 11713
rect 16114 11704 16120 11716
rect 16172 11704 16178 11756
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11645 12955 11679
rect 12897 11639 12955 11645
rect 13081 11679 13139 11685
rect 13081 11645 13093 11679
rect 13127 11676 13139 11679
rect 13354 11676 13360 11688
rect 13127 11648 13360 11676
rect 13127 11645 13139 11648
rect 13081 11639 13139 11645
rect 13354 11636 13360 11648
rect 13412 11636 13418 11688
rect 15580 11676 15608 11704
rect 16206 11676 16212 11688
rect 15580 11648 15700 11676
rect 16167 11648 16212 11676
rect 13538 11608 13544 11620
rect 7616 11580 12020 11608
rect 12084 11580 12572 11608
rect 12636 11580 13544 11608
rect 7616 11568 7622 11580
rect 4304 11512 4384 11540
rect 4617 11543 4675 11549
rect 4304 11500 4310 11512
rect 4617 11509 4629 11543
rect 4663 11540 4675 11543
rect 4706 11540 4712 11552
rect 4663 11512 4712 11540
rect 4663 11509 4675 11512
rect 4617 11503 4675 11509
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 4893 11543 4951 11549
rect 4893 11540 4905 11543
rect 4856 11512 4905 11540
rect 4856 11500 4862 11512
rect 4893 11509 4905 11512
rect 4939 11509 4951 11543
rect 4893 11503 4951 11509
rect 5626 11500 5632 11552
rect 5684 11540 5690 11552
rect 6365 11543 6423 11549
rect 6365 11540 6377 11543
rect 5684 11512 6377 11540
rect 5684 11500 5690 11512
rect 6365 11509 6377 11512
rect 6411 11540 6423 11543
rect 7374 11540 7380 11552
rect 6411 11512 7380 11540
rect 6411 11509 6423 11512
rect 6365 11503 6423 11509
rect 7374 11500 7380 11512
rect 7432 11500 7438 11552
rect 8662 11540 8668 11552
rect 8623 11512 8668 11540
rect 8662 11500 8668 11512
rect 8720 11500 8726 11552
rect 11514 11540 11520 11552
rect 11475 11512 11520 11540
rect 11514 11500 11520 11512
rect 11572 11540 11578 11552
rect 11882 11540 11888 11552
rect 11572 11512 11888 11540
rect 11572 11500 11578 11512
rect 11882 11500 11888 11512
rect 11940 11500 11946 11552
rect 11992 11540 12020 11580
rect 12636 11540 12664 11580
rect 13538 11568 13544 11580
rect 13596 11568 13602 11620
rect 15672 11608 15700 11648
rect 16206 11636 16212 11648
rect 16264 11636 16270 11688
rect 16301 11679 16359 11685
rect 16301 11645 16313 11679
rect 16347 11645 16359 11679
rect 16301 11639 16359 11645
rect 16316 11608 16344 11639
rect 15672 11580 16344 11608
rect 11992 11512 12664 11540
rect 12713 11543 12771 11549
rect 12713 11509 12725 11543
rect 12759 11540 12771 11543
rect 13262 11540 13268 11552
rect 12759 11512 13268 11540
rect 12759 11509 12771 11512
rect 12713 11503 12771 11509
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 13722 11500 13728 11552
rect 13780 11540 13786 11552
rect 18506 11540 18512 11552
rect 13780 11512 18512 11540
rect 13780 11500 13786 11512
rect 18506 11500 18512 11512
rect 18564 11500 18570 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 1394 11336 1400 11348
rect 1355 11308 1400 11336
rect 1394 11296 1400 11308
rect 1452 11296 1458 11348
rect 2314 11336 2320 11348
rect 2275 11308 2320 11336
rect 2314 11296 2320 11308
rect 2372 11296 2378 11348
rect 3881 11339 3939 11345
rect 3881 11336 3893 11339
rect 2424 11308 3893 11336
rect 1765 11203 1823 11209
rect 1765 11169 1777 11203
rect 1811 11200 1823 11203
rect 1854 11200 1860 11212
rect 1811 11172 1860 11200
rect 1811 11169 1823 11172
rect 1765 11163 1823 11169
rect 1854 11160 1860 11172
rect 1912 11160 1918 11212
rect 2424 11200 2452 11308
rect 3881 11305 3893 11308
rect 3927 11336 3939 11339
rect 5074 11336 5080 11348
rect 3927 11308 5080 11336
rect 3927 11305 3939 11308
rect 3881 11299 3939 11305
rect 5074 11296 5080 11308
rect 5132 11296 5138 11348
rect 5353 11339 5411 11345
rect 5353 11305 5365 11339
rect 5399 11336 5411 11339
rect 5442 11336 5448 11348
rect 5399 11308 5448 11336
rect 5399 11305 5411 11308
rect 5353 11299 5411 11305
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 6086 11296 6092 11348
rect 6144 11336 6150 11348
rect 6914 11336 6920 11348
rect 6144 11308 6920 11336
rect 6144 11296 6150 11308
rect 6914 11296 6920 11308
rect 6972 11296 6978 11348
rect 7009 11339 7067 11345
rect 7009 11305 7021 11339
rect 7055 11336 7067 11339
rect 8110 11336 8116 11348
rect 7055 11308 8116 11336
rect 7055 11305 7067 11308
rect 7009 11299 7067 11305
rect 8110 11296 8116 11308
rect 8168 11296 8174 11348
rect 8478 11296 8484 11348
rect 8536 11336 8542 11348
rect 8573 11339 8631 11345
rect 8573 11336 8585 11339
rect 8536 11308 8585 11336
rect 8536 11296 8542 11308
rect 8573 11305 8585 11308
rect 8619 11305 8631 11339
rect 8573 11299 8631 11305
rect 9950 11296 9956 11348
rect 10008 11336 10014 11348
rect 10505 11339 10563 11345
rect 10505 11336 10517 11339
rect 10008 11308 10517 11336
rect 10008 11296 10014 11308
rect 10505 11305 10517 11308
rect 10551 11305 10563 11339
rect 14185 11339 14243 11345
rect 10505 11299 10563 11305
rect 11624 11308 13676 11336
rect 3418 11228 3424 11280
rect 3476 11268 3482 11280
rect 4430 11268 4436 11280
rect 3476 11240 4436 11268
rect 3476 11228 3482 11240
rect 4430 11228 4436 11240
rect 4488 11228 4494 11280
rect 6181 11271 6239 11277
rect 6181 11237 6193 11271
rect 6227 11268 6239 11271
rect 6227 11240 6684 11268
rect 6227 11237 6239 11240
rect 6181 11231 6239 11237
rect 1964 11172 2452 11200
rect 1964 11132 1992 11172
rect 2590 11160 2596 11212
rect 2648 11200 2654 11212
rect 2774 11200 2780 11212
rect 2648 11172 2780 11200
rect 2648 11160 2654 11172
rect 2774 11160 2780 11172
rect 2832 11200 2838 11212
rect 2869 11203 2927 11209
rect 2869 11200 2881 11203
rect 2832 11172 2881 11200
rect 2832 11160 2838 11172
rect 2869 11169 2881 11172
rect 2915 11169 2927 11203
rect 3050 11200 3056 11212
rect 3011 11172 3056 11200
rect 2869 11163 2927 11169
rect 3050 11160 3056 11172
rect 3108 11160 3114 11212
rect 3602 11200 3608 11212
rect 3515 11172 3608 11200
rect 3602 11160 3608 11172
rect 3660 11200 3666 11212
rect 3970 11200 3976 11212
rect 3660 11172 3976 11200
rect 3660 11160 3666 11172
rect 3970 11160 3976 11172
rect 4028 11160 4034 11212
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11200 4859 11203
rect 4890 11200 4896 11212
rect 4847 11172 4896 11200
rect 4847 11169 4859 11172
rect 4801 11163 4859 11169
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 5629 11203 5687 11209
rect 5629 11169 5641 11203
rect 5675 11200 5687 11203
rect 5718 11200 5724 11212
rect 5675 11172 5724 11200
rect 5675 11169 5687 11172
rect 5629 11163 5687 11169
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 6457 11203 6515 11209
rect 6457 11169 6469 11203
rect 6503 11169 6515 11203
rect 6457 11163 6515 11169
rect 1872 11104 1992 11132
rect 1872 11073 1900 11104
rect 2038 11092 2044 11144
rect 2096 11132 2102 11144
rect 4985 11135 5043 11141
rect 2096 11104 4752 11132
rect 2096 11092 2102 11104
rect 4724 11076 4752 11104
rect 4985 11101 4997 11135
rect 5031 11132 5043 11135
rect 5902 11132 5908 11144
rect 5031 11104 5908 11132
rect 5031 11101 5043 11104
rect 4985 11095 5043 11101
rect 5902 11092 5908 11104
rect 5960 11092 5966 11144
rect 1857 11067 1915 11073
rect 1857 11033 1869 11067
rect 1903 11033 1915 11067
rect 1857 11027 1915 11033
rect 1949 11067 2007 11073
rect 1949 11033 1961 11067
rect 1995 11064 2007 11067
rect 3237 11067 3295 11073
rect 3237 11064 3249 11067
rect 1995 11036 3249 11064
rect 1995 11033 2007 11036
rect 1949 11027 2007 11033
rect 3237 11033 3249 11036
rect 3283 11033 3295 11067
rect 3237 11027 3295 11033
rect 1578 10956 1584 11008
rect 1636 10996 1642 11008
rect 1872 10996 1900 11027
rect 3326 11024 3332 11076
rect 3384 11064 3390 11076
rect 3973 11067 4031 11073
rect 3973 11064 3985 11067
rect 3384 11036 3985 11064
rect 3384 11024 3390 11036
rect 3973 11033 3985 11036
rect 4019 11033 4031 11067
rect 4249 11067 4307 11073
rect 4249 11064 4261 11067
rect 3973 11027 4031 11033
rect 4080 11036 4261 11064
rect 1636 10968 1900 10996
rect 2409 10999 2467 11005
rect 1636 10956 1642 10968
rect 2409 10965 2421 10999
rect 2455 10996 2467 10999
rect 2498 10996 2504 11008
rect 2455 10968 2504 10996
rect 2455 10965 2467 10968
rect 2409 10959 2467 10965
rect 2498 10956 2504 10968
rect 2556 10956 2562 11008
rect 2777 10999 2835 11005
rect 2777 10965 2789 10999
rect 2823 10996 2835 10999
rect 3602 10996 3608 11008
rect 2823 10968 3608 10996
rect 2823 10965 2835 10968
rect 2777 10959 2835 10965
rect 3602 10956 3608 10968
rect 3660 10956 3666 11008
rect 3786 10956 3792 11008
rect 3844 10996 3850 11008
rect 4080 10996 4108 11036
rect 4249 11033 4261 11036
rect 4295 11064 4307 11067
rect 4295 11036 4660 11064
rect 4295 11033 4307 11036
rect 4249 11027 4307 11033
rect 3844 10968 4108 10996
rect 4632 10996 4660 11036
rect 4706 11024 4712 11076
rect 4764 11064 4770 11076
rect 4893 11067 4951 11073
rect 4893 11064 4905 11067
rect 4764 11036 4905 11064
rect 4764 11024 4770 11036
rect 4893 11033 4905 11036
rect 4939 11033 4951 11067
rect 5534 11064 5540 11076
rect 4893 11027 4951 11033
rect 5000 11036 5540 11064
rect 5000 10996 5028 11036
rect 5534 11024 5540 11036
rect 5592 11024 5598 11076
rect 5810 11064 5816 11076
rect 5771 11036 5816 11064
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 6472 11064 6500 11163
rect 6656 11141 6684 11240
rect 6822 11160 6828 11212
rect 6880 11200 6886 11212
rect 6880 11172 7328 11200
rect 6880 11160 6886 11172
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 6730 11092 6736 11144
rect 6788 11132 6794 11144
rect 7193 11135 7251 11141
rect 7193 11132 7205 11135
rect 6788 11104 7205 11132
rect 6788 11092 6794 11104
rect 7193 11101 7205 11104
rect 7239 11101 7251 11135
rect 7300 11132 7328 11172
rect 10594 11160 10600 11212
rect 10652 11200 10658 11212
rect 11057 11203 11115 11209
rect 11057 11200 11069 11203
rect 10652 11172 11069 11200
rect 10652 11160 10658 11172
rect 11057 11169 11069 11172
rect 11103 11169 11115 11203
rect 11057 11163 11115 11169
rect 11146 11160 11152 11212
rect 11204 11200 11210 11212
rect 11517 11203 11575 11209
rect 11517 11200 11529 11203
rect 11204 11172 11529 11200
rect 11204 11160 11210 11172
rect 11517 11169 11529 11172
rect 11563 11200 11575 11203
rect 11624 11200 11652 11308
rect 12069 11271 12127 11277
rect 12069 11237 12081 11271
rect 12115 11268 12127 11271
rect 13081 11271 13139 11277
rect 13081 11268 13093 11271
rect 12115 11240 12434 11268
rect 12115 11237 12127 11240
rect 12069 11231 12127 11237
rect 11563 11172 11652 11200
rect 11563 11169 11575 11172
rect 11517 11163 11575 11169
rect 8941 11135 8999 11141
rect 8941 11132 8953 11135
rect 7300 11104 8953 11132
rect 7193 11095 7251 11101
rect 8941 11101 8953 11104
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 10965 11135 11023 11141
rect 10965 11132 10977 11135
rect 9732 11104 10977 11132
rect 9732 11092 9738 11104
rect 10965 11101 10977 11104
rect 11011 11101 11023 11135
rect 10965 11095 11023 11101
rect 11609 11135 11667 11141
rect 11609 11101 11621 11135
rect 11655 11132 11667 11135
rect 11790 11132 11796 11144
rect 11655 11104 11796 11132
rect 11655 11101 11667 11104
rect 11609 11095 11667 11101
rect 11790 11092 11796 11104
rect 11848 11092 11854 11144
rect 12406 11132 12434 11240
rect 12636 11240 13093 11268
rect 12636 11141 12664 11240
rect 13081 11237 13093 11240
rect 13127 11237 13139 11271
rect 13081 11231 13139 11237
rect 13648 11268 13676 11308
rect 14185 11305 14197 11339
rect 14231 11336 14243 11339
rect 17218 11336 17224 11348
rect 14231 11308 17224 11336
rect 14231 11305 14243 11308
rect 14185 11299 14243 11305
rect 14737 11271 14795 11277
rect 14737 11268 14749 11271
rect 13648 11240 14749 11268
rect 12802 11200 12808 11212
rect 12763 11172 12808 11200
rect 12802 11160 12808 11172
rect 12860 11160 12866 11212
rect 13648 11209 13676 11240
rect 14737 11237 14749 11240
rect 14783 11237 14795 11271
rect 14737 11231 14795 11237
rect 13633 11203 13691 11209
rect 13633 11169 13645 11203
rect 13679 11169 13691 11203
rect 14844 11200 14872 11308
rect 17218 11296 17224 11308
rect 17276 11296 17282 11348
rect 13633 11163 13691 11169
rect 14292 11172 14872 11200
rect 12621 11135 12679 11141
rect 12406 11104 12572 11132
rect 7460 11067 7518 11073
rect 7460 11064 7472 11067
rect 6472 11036 7472 11064
rect 7460 11033 7472 11036
rect 7506 11064 7518 11067
rect 7834 11064 7840 11076
rect 7506 11036 7840 11064
rect 7506 11033 7518 11036
rect 7460 11027 7518 11033
rect 7834 11024 7840 11036
rect 7892 11024 7898 11076
rect 9208 11067 9266 11073
rect 9208 11033 9220 11067
rect 9254 11064 9266 11067
rect 9582 11064 9588 11076
rect 9254 11036 9588 11064
rect 9254 11033 9266 11036
rect 9208 11027 9266 11033
rect 9582 11024 9588 11036
rect 9640 11024 9646 11076
rect 10042 11024 10048 11076
rect 10100 11064 10106 11076
rect 11701 11067 11759 11073
rect 11701 11064 11713 11067
rect 10100 11036 11713 11064
rect 10100 11024 10106 11036
rect 11701 11033 11713 11036
rect 11747 11033 11759 11067
rect 11701 11027 11759 11033
rect 11974 11024 11980 11076
rect 12032 11064 12038 11076
rect 12544 11064 12572 11104
rect 12621 11101 12633 11135
rect 12667 11101 12679 11135
rect 12621 11095 12679 11101
rect 13449 11135 13507 11141
rect 13449 11101 13461 11135
rect 13495 11132 13507 11135
rect 13814 11132 13820 11144
rect 13495 11104 13820 11132
rect 13495 11101 13507 11104
rect 13449 11095 13507 11101
rect 12713 11067 12771 11073
rect 12713 11064 12725 11067
rect 12032 11036 12480 11064
rect 12544 11036 12725 11064
rect 12032 11024 12038 11036
rect 4632 10968 5028 10996
rect 3844 10956 3850 10968
rect 5074 10956 5080 11008
rect 5132 10996 5138 11008
rect 5721 10999 5779 11005
rect 5721 10996 5733 10999
rect 5132 10968 5733 10996
rect 5132 10956 5138 10968
rect 5721 10965 5733 10968
rect 5767 10996 5779 10999
rect 5994 10996 6000 11008
rect 5767 10968 6000 10996
rect 5767 10965 5779 10968
rect 5721 10959 5779 10965
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 6546 10996 6552 11008
rect 6507 10968 6552 10996
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 6638 10956 6644 11008
rect 6696 10996 6702 11008
rect 8110 10996 8116 11008
rect 6696 10968 8116 10996
rect 6696 10956 6702 10968
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 10318 10996 10324 11008
rect 10279 10968 10324 10996
rect 10318 10956 10324 10968
rect 10376 10956 10382 11008
rect 10594 10956 10600 11008
rect 10652 10996 10658 11008
rect 10873 10999 10931 11005
rect 10873 10996 10885 10999
rect 10652 10968 10885 10996
rect 10652 10956 10658 10968
rect 10873 10965 10885 10968
rect 10919 10996 10931 10999
rect 10962 10996 10968 11008
rect 10919 10968 10968 10996
rect 10919 10965 10931 10968
rect 10873 10959 10931 10965
rect 10962 10956 10968 10968
rect 11020 10956 11026 11008
rect 12250 10996 12256 11008
rect 12211 10968 12256 10996
rect 12250 10956 12256 10968
rect 12308 10956 12314 11008
rect 12452 10996 12480 11036
rect 12713 11033 12725 11036
rect 12759 11033 12771 11067
rect 13464 11064 13492 11095
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 12713 11027 12771 11033
rect 12820 11036 13492 11064
rect 12820 10996 12848 11036
rect 13538 11024 13544 11076
rect 13596 11064 13602 11076
rect 14292 11064 14320 11172
rect 14458 11092 14464 11144
rect 14516 11132 14522 11144
rect 16117 11135 16175 11141
rect 16117 11132 16129 11135
rect 14516 11104 16129 11132
rect 14516 11092 14522 11104
rect 16117 11101 16129 11104
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 13596 11036 14320 11064
rect 15872 11067 15930 11073
rect 13596 11024 13602 11036
rect 15872 11033 15884 11067
rect 15918 11064 15930 11067
rect 16390 11064 16396 11076
rect 15918 11036 16396 11064
rect 15918 11033 15930 11036
rect 15872 11027 15930 11033
rect 16390 11024 16396 11036
rect 16448 11024 16454 11076
rect 14642 10996 14648 11008
rect 12452 10968 12848 10996
rect 14603 10968 14648 10996
rect 14642 10956 14648 10968
rect 14700 10956 14706 11008
rect 1104 10906 21896 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21896 10906
rect 1104 10832 21896 10854
rect 4065 10795 4123 10801
rect 4065 10792 4077 10795
rect 1688 10764 4077 10792
rect 1688 10668 1716 10764
rect 4065 10761 4077 10764
rect 4111 10761 4123 10795
rect 4065 10755 4123 10761
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 4617 10795 4675 10801
rect 4617 10792 4629 10795
rect 4396 10764 4629 10792
rect 4396 10752 4402 10764
rect 4617 10761 4629 10764
rect 4663 10761 4675 10795
rect 4617 10755 4675 10761
rect 4985 10795 5043 10801
rect 4985 10761 4997 10795
rect 5031 10792 5043 10795
rect 5350 10792 5356 10804
rect 5031 10764 5356 10792
rect 5031 10761 5043 10764
rect 4985 10755 5043 10761
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 7466 10792 7472 10804
rect 5460 10764 7472 10792
rect 3881 10727 3939 10733
rect 3881 10724 3893 10727
rect 1964 10696 3893 10724
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 1670 10656 1676 10668
rect 1631 10628 1676 10656
rect 1670 10616 1676 10628
rect 1728 10616 1734 10668
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 1964 10665 1992 10696
rect 3881 10693 3893 10696
rect 3927 10693 3939 10727
rect 4890 10724 4896 10736
rect 3881 10687 3939 10693
rect 4448 10696 4896 10724
rect 1949 10659 2007 10665
rect 1949 10656 1961 10659
rect 1912 10628 1961 10656
rect 1912 10616 1918 10628
rect 1949 10625 1961 10628
rect 1995 10625 2007 10659
rect 1949 10619 2007 10625
rect 2314 10616 2320 10668
rect 2372 10656 2378 10668
rect 2665 10659 2723 10665
rect 2665 10656 2677 10659
rect 2372 10628 2677 10656
rect 2372 10616 2378 10628
rect 2665 10625 2677 10628
rect 2711 10625 2723 10659
rect 2665 10619 2723 10625
rect 3234 10616 3240 10668
rect 3292 10656 3298 10668
rect 3786 10656 3792 10668
rect 3292 10628 3792 10656
rect 3292 10616 3298 10628
rect 3786 10616 3792 10628
rect 3844 10616 3850 10668
rect 1412 10588 1440 10616
rect 2406 10588 2412 10600
rect 1412 10560 2268 10588
rect 2367 10560 2412 10588
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10520 1639 10523
rect 1946 10520 1952 10532
rect 1627 10492 1952 10520
rect 1627 10489 1639 10492
rect 1581 10483 1639 10489
rect 1946 10480 1952 10492
rect 2004 10480 2010 10532
rect 2130 10520 2136 10532
rect 2091 10492 2136 10520
rect 2130 10480 2136 10492
rect 2188 10480 2194 10532
rect 2240 10520 2268 10560
rect 2406 10548 2412 10560
rect 2464 10548 2470 10600
rect 4448 10597 4476 10696
rect 4890 10684 4896 10696
rect 4948 10684 4954 10736
rect 5258 10684 5264 10736
rect 5316 10724 5322 10736
rect 5460 10724 5488 10764
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 7745 10795 7803 10801
rect 7745 10761 7757 10795
rect 7791 10792 7803 10795
rect 7834 10792 7840 10804
rect 7791 10764 7840 10792
rect 7791 10761 7803 10764
rect 7745 10755 7803 10761
rect 7834 10752 7840 10764
rect 7892 10752 7898 10804
rect 8386 10752 8392 10804
rect 8444 10792 8450 10804
rect 8481 10795 8539 10801
rect 8481 10792 8493 10795
rect 8444 10764 8493 10792
rect 8444 10752 8450 10764
rect 8481 10761 8493 10764
rect 8527 10761 8539 10795
rect 8481 10755 8539 10761
rect 8662 10752 8668 10804
rect 8720 10792 8726 10804
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8720 10764 8953 10792
rect 8720 10752 8726 10764
rect 8941 10761 8953 10764
rect 8987 10761 8999 10795
rect 8941 10755 8999 10761
rect 9122 10752 9128 10804
rect 9180 10792 9186 10804
rect 9769 10795 9827 10801
rect 9769 10792 9781 10795
rect 9180 10764 9781 10792
rect 9180 10752 9186 10764
rect 9769 10761 9781 10764
rect 9815 10761 9827 10795
rect 9769 10755 9827 10761
rect 10229 10795 10287 10801
rect 10229 10761 10241 10795
rect 10275 10761 10287 10795
rect 10229 10755 10287 10761
rect 11241 10795 11299 10801
rect 11241 10761 11253 10795
rect 11287 10792 11299 10795
rect 11790 10792 11796 10804
rect 11287 10764 11796 10792
rect 11287 10761 11299 10764
rect 11241 10755 11299 10761
rect 6730 10724 6736 10736
rect 5316 10696 5488 10724
rect 6380 10696 6736 10724
rect 5316 10684 5322 10696
rect 4982 10616 4988 10668
rect 5040 10656 5046 10668
rect 5445 10659 5503 10665
rect 5445 10656 5457 10659
rect 5040 10628 5457 10656
rect 5040 10616 5046 10628
rect 5445 10625 5457 10628
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 5718 10616 5724 10668
rect 5776 10656 5782 10668
rect 6380 10665 6408 10696
rect 6730 10684 6736 10696
rect 6788 10684 6794 10736
rect 6822 10684 6828 10736
rect 6880 10684 6886 10736
rect 8849 10727 8907 10733
rect 8849 10693 8861 10727
rect 8895 10724 8907 10727
rect 10244 10724 10272 10755
rect 11790 10752 11796 10764
rect 11848 10752 11854 10804
rect 12250 10752 12256 10804
rect 12308 10792 12314 10804
rect 12529 10795 12587 10801
rect 12529 10792 12541 10795
rect 12308 10764 12541 10792
rect 12308 10752 12314 10764
rect 12529 10761 12541 10764
rect 12575 10761 12587 10795
rect 12529 10755 12587 10761
rect 12989 10795 13047 10801
rect 12989 10761 13001 10795
rect 13035 10792 13047 10795
rect 14550 10792 14556 10804
rect 13035 10764 14556 10792
rect 13035 10761 13047 10764
rect 12989 10755 13047 10761
rect 14550 10752 14556 10764
rect 14608 10752 14614 10804
rect 14642 10752 14648 10804
rect 14700 10792 14706 10804
rect 14921 10795 14979 10801
rect 14921 10792 14933 10795
rect 14700 10764 14933 10792
rect 14700 10752 14706 10764
rect 14921 10761 14933 10764
rect 14967 10761 14979 10795
rect 14921 10755 14979 10761
rect 15289 10795 15347 10801
rect 15289 10761 15301 10795
rect 15335 10792 15347 10795
rect 16114 10792 16120 10804
rect 15335 10764 16120 10792
rect 15335 10761 15347 10764
rect 15289 10755 15347 10761
rect 16114 10752 16120 10764
rect 16172 10752 16178 10804
rect 14829 10727 14887 10733
rect 14829 10724 14841 10727
rect 8895 10696 10272 10724
rect 10336 10696 14841 10724
rect 8895 10693 8907 10696
rect 8849 10687 8907 10693
rect 6638 10665 6644 10668
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 5776 10628 6377 10656
rect 5776 10616 5782 10628
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6632 10656 6644 10665
rect 6599 10628 6644 10656
rect 6365 10619 6423 10625
rect 6632 10619 6644 10628
rect 6638 10616 6644 10619
rect 6696 10616 6702 10668
rect 6840 10656 6868 10684
rect 9674 10656 9680 10668
rect 6840 10628 9168 10656
rect 9635 10628 9680 10656
rect 4433 10591 4491 10597
rect 4433 10557 4445 10591
rect 4479 10557 4491 10591
rect 4433 10551 4491 10557
rect 4525 10591 4583 10597
rect 4525 10557 4537 10591
rect 4571 10557 4583 10591
rect 5534 10588 5540 10600
rect 5495 10560 5540 10588
rect 4525 10551 4583 10557
rect 3789 10523 3847 10529
rect 2240 10492 2360 10520
rect 1857 10455 1915 10461
rect 1857 10421 1869 10455
rect 1903 10452 1915 10455
rect 2038 10452 2044 10464
rect 1903 10424 2044 10452
rect 1903 10421 1915 10424
rect 1857 10415 1915 10421
rect 2038 10412 2044 10424
rect 2096 10412 2102 10464
rect 2222 10452 2228 10464
rect 2183 10424 2228 10452
rect 2222 10412 2228 10424
rect 2280 10412 2286 10464
rect 2332 10452 2360 10492
rect 3789 10489 3801 10523
rect 3835 10520 3847 10523
rect 3970 10520 3976 10532
rect 3835 10492 3976 10520
rect 3835 10489 3847 10492
rect 3789 10483 3847 10489
rect 3970 10480 3976 10492
rect 4028 10480 4034 10532
rect 4062 10480 4068 10532
rect 4120 10520 4126 10532
rect 4540 10520 4568 10551
rect 5534 10548 5540 10560
rect 5592 10548 5598 10600
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 4120 10492 4568 10520
rect 4120 10480 4126 10492
rect 4614 10480 4620 10532
rect 4672 10520 4678 10532
rect 5077 10523 5135 10529
rect 5077 10520 5089 10523
rect 4672 10492 5089 10520
rect 4672 10480 4678 10492
rect 5077 10489 5089 10492
rect 5123 10489 5135 10523
rect 5644 10520 5672 10551
rect 7834 10548 7840 10600
rect 7892 10588 7898 10600
rect 9033 10591 9091 10597
rect 9033 10588 9045 10591
rect 7892 10560 9045 10588
rect 7892 10548 7898 10560
rect 9033 10557 9045 10560
rect 9079 10557 9091 10591
rect 9140 10588 9168 10628
rect 9674 10616 9680 10628
rect 9732 10616 9738 10668
rect 10336 10656 10364 10696
rect 14829 10693 14841 10696
rect 14875 10724 14887 10727
rect 15381 10727 15439 10733
rect 15381 10724 15393 10727
rect 14875 10696 15393 10724
rect 14875 10693 14887 10696
rect 14829 10687 14887 10693
rect 15381 10693 15393 10696
rect 15427 10724 15439 10727
rect 15470 10724 15476 10736
rect 15427 10696 15476 10724
rect 15427 10693 15439 10696
rect 15381 10687 15439 10693
rect 15470 10684 15476 10696
rect 15528 10684 15534 10736
rect 9784 10628 10364 10656
rect 10597 10659 10655 10665
rect 9784 10588 9812 10628
rect 10597 10625 10609 10659
rect 10643 10656 10655 10659
rect 11606 10656 11612 10668
rect 10643 10628 11612 10656
rect 10643 10625 10655 10628
rect 10597 10619 10655 10625
rect 11606 10616 11612 10628
rect 11664 10616 11670 10668
rect 12618 10656 12624 10668
rect 12579 10628 12624 10656
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 14182 10656 14188 10668
rect 14240 10665 14246 10668
rect 14152 10628 14188 10656
rect 14182 10616 14188 10628
rect 14240 10619 14252 10665
rect 14458 10656 14464 10668
rect 14419 10628 14464 10656
rect 14240 10616 14246 10619
rect 14458 10616 14464 10628
rect 14516 10616 14522 10668
rect 9950 10588 9956 10600
rect 9140 10560 9812 10588
rect 9863 10560 9956 10588
rect 9033 10551 9091 10557
rect 9950 10548 9956 10560
rect 10008 10588 10014 10600
rect 10318 10588 10324 10600
rect 10008 10560 10324 10588
rect 10008 10548 10014 10560
rect 10318 10548 10324 10560
rect 10376 10548 10382 10600
rect 10686 10588 10692 10600
rect 10647 10560 10692 10588
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 10873 10591 10931 10597
rect 10873 10557 10885 10591
rect 10919 10557 10931 10591
rect 11790 10588 11796 10600
rect 11751 10560 11796 10588
rect 10873 10551 10931 10557
rect 5077 10483 5135 10489
rect 5184 10492 5672 10520
rect 3326 10452 3332 10464
rect 2332 10424 3332 10452
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 3878 10412 3884 10464
rect 3936 10452 3942 10464
rect 5184 10452 5212 10492
rect 8202 10480 8208 10532
rect 8260 10520 8266 10532
rect 10888 10520 10916 10551
rect 11790 10548 11796 10560
rect 11848 10548 11854 10600
rect 12434 10548 12440 10600
rect 12492 10588 12498 10600
rect 14734 10588 14740 10600
rect 12492 10560 12537 10588
rect 14695 10560 14740 10588
rect 12492 10548 12498 10560
rect 14734 10548 14740 10560
rect 14792 10548 14798 10600
rect 13081 10523 13139 10529
rect 13081 10520 13093 10523
rect 8260 10492 13093 10520
rect 8260 10480 8266 10492
rect 13081 10489 13093 10492
rect 13127 10489 13139 10523
rect 13081 10483 13139 10489
rect 5902 10452 5908 10464
rect 3936 10424 5212 10452
rect 5863 10424 5908 10452
rect 3936 10412 3942 10424
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 5994 10412 6000 10464
rect 6052 10452 6058 10464
rect 6089 10455 6147 10461
rect 6089 10452 6101 10455
rect 6052 10424 6101 10452
rect 6052 10412 6058 10424
rect 6089 10421 6101 10424
rect 6135 10421 6147 10455
rect 6089 10415 6147 10421
rect 6638 10412 6644 10464
rect 6696 10452 6702 10464
rect 8220 10452 8248 10480
rect 9306 10452 9312 10464
rect 6696 10424 8248 10452
rect 9267 10424 9312 10452
rect 6696 10412 6702 10424
rect 9306 10412 9312 10424
rect 9364 10412 9370 10464
rect 11606 10452 11612 10464
rect 11519 10424 11612 10452
rect 11606 10412 11612 10424
rect 11664 10452 11670 10464
rect 12066 10452 12072 10464
rect 11664 10424 12072 10452
rect 11664 10412 11670 10424
rect 12066 10412 12072 10424
rect 12124 10452 12130 10464
rect 12250 10452 12256 10464
rect 12124 10424 12256 10452
rect 12124 10412 12130 10424
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 1486 10248 1492 10260
rect 1447 10220 1492 10248
rect 1486 10208 1492 10220
rect 1544 10208 1550 10260
rect 1762 10248 1768 10260
rect 1723 10220 1768 10248
rect 1762 10208 1768 10220
rect 1820 10208 1826 10260
rect 3789 10251 3847 10257
rect 3789 10217 3801 10251
rect 3835 10248 3847 10251
rect 3878 10248 3884 10260
rect 3835 10220 3884 10248
rect 3835 10217 3847 10220
rect 3789 10211 3847 10217
rect 3878 10208 3884 10220
rect 3936 10208 3942 10260
rect 3970 10208 3976 10260
rect 4028 10248 4034 10260
rect 5902 10248 5908 10260
rect 4028 10220 5908 10248
rect 4028 10208 4034 10220
rect 5902 10208 5908 10220
rect 5960 10208 5966 10260
rect 6546 10248 6552 10260
rect 6507 10220 6552 10248
rect 6546 10208 6552 10220
rect 6604 10208 6610 10260
rect 9582 10248 9588 10260
rect 9543 10220 9588 10248
rect 9582 10208 9588 10220
rect 9640 10208 9646 10260
rect 12434 10208 12440 10260
rect 12492 10248 12498 10260
rect 13538 10248 13544 10260
rect 12492 10220 13544 10248
rect 12492 10208 12498 10220
rect 13538 10208 13544 10220
rect 13596 10208 13602 10260
rect 15013 10251 15071 10257
rect 15013 10217 15025 10251
rect 15059 10248 15071 10251
rect 16206 10248 16212 10260
rect 15059 10220 16212 10248
rect 15059 10217 15071 10220
rect 15013 10211 15071 10217
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 5534 10140 5540 10192
rect 5592 10180 5598 10192
rect 7377 10183 7435 10189
rect 7377 10180 7389 10183
rect 5592 10152 7389 10180
rect 5592 10140 5598 10152
rect 7377 10149 7389 10152
rect 7423 10149 7435 10183
rect 7377 10143 7435 10149
rect 7466 10140 7472 10192
rect 7524 10180 7530 10192
rect 10502 10180 10508 10192
rect 7524 10152 10508 10180
rect 7524 10140 7530 10152
rect 10502 10140 10508 10152
rect 10560 10140 10566 10192
rect 3421 10115 3479 10121
rect 3421 10081 3433 10115
rect 3467 10112 3479 10115
rect 3602 10112 3608 10124
rect 3467 10084 3608 10112
rect 3467 10081 3479 10084
rect 3421 10075 3479 10081
rect 3602 10072 3608 10084
rect 3660 10072 3666 10124
rect 5169 10115 5227 10121
rect 5169 10081 5181 10115
rect 5215 10112 5227 10115
rect 5718 10112 5724 10124
rect 5215 10084 5724 10112
rect 5215 10081 5227 10084
rect 5169 10075 5227 10081
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 2406 10004 2412 10056
rect 2464 10044 2470 10056
rect 3237 10047 3295 10053
rect 3237 10044 3249 10047
rect 2464 10016 3249 10044
rect 2464 10004 2470 10016
rect 3237 10013 3249 10016
rect 3283 10044 3295 10047
rect 5184 10044 5212 10075
rect 5718 10072 5724 10084
rect 5776 10072 5782 10124
rect 5810 10072 5816 10124
rect 5868 10112 5874 10124
rect 5997 10115 6055 10121
rect 5997 10112 6009 10115
rect 5868 10084 6009 10112
rect 5868 10072 5874 10084
rect 5997 10081 6009 10084
rect 6043 10112 6055 10115
rect 6546 10112 6552 10124
rect 6043 10084 6552 10112
rect 6043 10081 6055 10084
rect 5997 10075 6055 10081
rect 6546 10072 6552 10084
rect 6604 10072 6610 10124
rect 6914 10072 6920 10124
rect 6972 10112 6978 10124
rect 7098 10112 7104 10124
rect 6972 10084 7104 10112
rect 6972 10072 6978 10084
rect 7098 10072 7104 10084
rect 7156 10112 7162 10124
rect 7929 10115 7987 10121
rect 7929 10112 7941 10115
rect 7156 10084 7941 10112
rect 7156 10072 7162 10084
rect 7929 10081 7941 10084
rect 7975 10081 7987 10115
rect 10321 10115 10379 10121
rect 10321 10112 10333 10115
rect 7929 10075 7987 10081
rect 8220 10084 10333 10112
rect 3283 10016 5212 10044
rect 3283 10013 3295 10016
rect 3237 10007 3295 10013
rect 5258 10004 5264 10056
rect 5316 10044 5322 10056
rect 5316 10016 5361 10044
rect 5316 10004 5322 10016
rect 5442 10004 5448 10056
rect 5500 10044 5506 10056
rect 6181 10047 6239 10053
rect 6181 10044 6193 10047
rect 5500 10016 6193 10044
rect 5500 10004 5506 10016
rect 6181 10013 6193 10016
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10013 6699 10047
rect 6641 10007 6699 10013
rect 2222 9936 2228 9988
rect 2280 9976 2286 9988
rect 2590 9976 2596 9988
rect 2280 9948 2596 9976
rect 2280 9936 2286 9948
rect 2590 9936 2596 9948
rect 2648 9936 2654 9988
rect 2958 9936 2964 9988
rect 3016 9985 3022 9988
rect 3016 9976 3028 9985
rect 4924 9979 4982 9985
rect 3016 9948 3061 9976
rect 3016 9939 3028 9948
rect 4924 9945 4936 9979
rect 4970 9976 4982 9979
rect 5074 9976 5080 9988
rect 4970 9948 5080 9976
rect 4970 9945 4982 9948
rect 4924 9939 4982 9945
rect 3016 9936 3022 9939
rect 5074 9936 5080 9948
rect 5132 9936 5138 9988
rect 5902 9936 5908 9988
rect 5960 9976 5966 9988
rect 6656 9976 6684 10007
rect 7006 10004 7012 10056
rect 7064 10044 7070 10056
rect 8220 10044 8248 10084
rect 10321 10081 10333 10084
rect 10367 10112 10379 10115
rect 10594 10112 10600 10124
rect 10367 10084 10600 10112
rect 10367 10081 10379 10084
rect 10321 10075 10379 10081
rect 10594 10072 10600 10084
rect 10652 10072 10658 10124
rect 14461 10115 14519 10121
rect 14461 10081 14473 10115
rect 14507 10112 14519 10115
rect 14734 10112 14740 10124
rect 14507 10084 14740 10112
rect 14507 10081 14519 10084
rect 14461 10075 14519 10081
rect 14734 10072 14740 10084
rect 14792 10072 14798 10124
rect 7064 10016 8248 10044
rect 7064 10004 7070 10016
rect 8478 10004 8484 10056
rect 8536 10044 8542 10056
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8536 10016 8953 10044
rect 8536 10004 8542 10016
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 8941 10007 8999 10013
rect 10689 10047 10747 10053
rect 10689 10013 10701 10047
rect 10735 10044 10747 10047
rect 12158 10044 12164 10056
rect 10735 10016 12164 10044
rect 10735 10013 10747 10016
rect 10689 10007 10747 10013
rect 11072 9988 11100 10016
rect 12158 10004 12164 10016
rect 12216 10004 12222 10056
rect 12428 10047 12486 10053
rect 12428 10044 12440 10047
rect 12406 10013 12440 10044
rect 12474 10044 12486 10047
rect 12802 10044 12808 10056
rect 12474 10016 12808 10044
rect 12474 10013 12486 10016
rect 12406 10007 12486 10013
rect 5960 9948 6684 9976
rect 7745 9979 7803 9985
rect 5960 9936 5966 9948
rect 7745 9945 7757 9979
rect 7791 9976 7803 9979
rect 8386 9976 8392 9988
rect 7791 9948 8392 9976
rect 7791 9945 7803 9948
rect 7745 9939 7803 9945
rect 8386 9936 8392 9948
rect 8444 9936 8450 9988
rect 10956 9979 11014 9985
rect 10956 9945 10968 9979
rect 11002 9945 11014 9979
rect 10956 9939 11014 9945
rect 1854 9908 1860 9920
rect 1815 9880 1860 9908
rect 1854 9868 1860 9880
rect 1912 9868 1918 9920
rect 3605 9911 3663 9917
rect 3605 9877 3617 9911
rect 3651 9908 3663 9911
rect 3786 9908 3792 9920
rect 3651 9880 3792 9908
rect 3651 9877 3663 9880
rect 3605 9871 3663 9877
rect 3786 9868 3792 9880
rect 3844 9868 3850 9920
rect 5534 9908 5540 9920
rect 5495 9880 5540 9908
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 5626 9868 5632 9920
rect 5684 9908 5690 9920
rect 6089 9911 6147 9917
rect 6089 9908 6101 9911
rect 5684 9880 6101 9908
rect 5684 9868 5690 9880
rect 6089 9877 6101 9880
rect 6135 9877 6147 9911
rect 6089 9871 6147 9877
rect 6638 9868 6644 9920
rect 6696 9908 6702 9920
rect 7285 9911 7343 9917
rect 7285 9908 7297 9911
rect 6696 9880 7297 9908
rect 6696 9868 6702 9880
rect 7285 9877 7297 9880
rect 7331 9877 7343 9911
rect 7285 9871 7343 9877
rect 7834 9868 7840 9920
rect 7892 9908 7898 9920
rect 7892 9880 7937 9908
rect 7892 9868 7898 9880
rect 9674 9868 9680 9920
rect 9732 9908 9738 9920
rect 10045 9911 10103 9917
rect 10045 9908 10057 9911
rect 9732 9880 10057 9908
rect 9732 9868 9738 9880
rect 10045 9877 10057 9880
rect 10091 9908 10103 9911
rect 10226 9908 10232 9920
rect 10091 9880 10232 9908
rect 10091 9877 10103 9880
rect 10045 9871 10103 9877
rect 10226 9868 10232 9880
rect 10284 9908 10290 9920
rect 10686 9908 10692 9920
rect 10284 9880 10692 9908
rect 10284 9868 10290 9880
rect 10686 9868 10692 9880
rect 10744 9868 10750 9920
rect 10980 9908 11008 9939
rect 11054 9936 11060 9988
rect 11112 9936 11118 9988
rect 11146 9908 11152 9920
rect 10980 9880 11152 9908
rect 11146 9868 11152 9880
rect 11204 9868 11210 9920
rect 11698 9868 11704 9920
rect 11756 9908 11762 9920
rect 12069 9911 12127 9917
rect 12069 9908 12081 9911
rect 11756 9880 12081 9908
rect 11756 9868 11762 9880
rect 12069 9877 12081 9880
rect 12115 9908 12127 9911
rect 12406 9908 12434 10007
rect 12802 10004 12808 10016
rect 12860 10004 12866 10056
rect 14185 10047 14243 10053
rect 14185 10013 14197 10047
rect 14231 10044 14243 10047
rect 14553 10047 14611 10053
rect 14553 10044 14565 10047
rect 14231 10016 14565 10044
rect 14231 10013 14243 10016
rect 14185 10007 14243 10013
rect 14553 10013 14565 10016
rect 14599 10044 14611 10047
rect 14642 10044 14648 10056
rect 14599 10016 14648 10044
rect 14599 10013 14611 10016
rect 14553 10007 14611 10013
rect 14642 10004 14648 10016
rect 14700 10004 14706 10056
rect 12115 9880 12434 9908
rect 14645 9911 14703 9917
rect 12115 9877 12127 9880
rect 12069 9871 12127 9877
rect 14645 9877 14657 9911
rect 14691 9908 14703 9911
rect 15286 9908 15292 9920
rect 14691 9880 15292 9908
rect 14691 9877 14703 9880
rect 14645 9871 14703 9877
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 1104 9818 21896 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21896 9818
rect 1104 9744 21896 9766
rect 1854 9664 1860 9716
rect 1912 9704 1918 9716
rect 3050 9704 3056 9716
rect 1912 9676 3056 9704
rect 1912 9664 1918 9676
rect 3050 9664 3056 9676
rect 3108 9664 3114 9716
rect 4617 9707 4675 9713
rect 4617 9673 4629 9707
rect 4663 9704 4675 9707
rect 5258 9704 5264 9716
rect 4663 9676 5264 9704
rect 4663 9673 4675 9676
rect 4617 9667 4675 9673
rect 5258 9664 5264 9676
rect 5316 9664 5322 9716
rect 6917 9707 6975 9713
rect 6917 9673 6929 9707
rect 6963 9704 6975 9707
rect 7098 9704 7104 9716
rect 6963 9676 7104 9704
rect 6963 9673 6975 9676
rect 6917 9667 6975 9673
rect 7098 9664 7104 9676
rect 7156 9664 7162 9716
rect 9122 9664 9128 9716
rect 9180 9704 9186 9716
rect 9490 9704 9496 9716
rect 9180 9676 9496 9704
rect 9180 9664 9186 9676
rect 9490 9664 9496 9676
rect 9548 9664 9554 9716
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 13262 9704 13268 9716
rect 10560 9676 13268 9704
rect 10560 9664 10566 9676
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 14185 9707 14243 9713
rect 14185 9673 14197 9707
rect 14231 9704 14243 9707
rect 14274 9704 14280 9716
rect 14231 9676 14280 9704
rect 14231 9673 14243 9676
rect 14185 9667 14243 9673
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 1762 9596 1768 9648
rect 1820 9636 1826 9648
rect 4154 9636 4160 9648
rect 1820 9608 4016 9636
rect 4115 9608 4160 9636
rect 1820 9596 1826 9608
rect 1486 9568 1492 9580
rect 1447 9540 1492 9568
rect 1486 9528 1492 9540
rect 1544 9528 1550 9580
rect 2866 9568 2872 9580
rect 2827 9540 2872 9568
rect 2866 9528 2872 9540
rect 2924 9528 2930 9580
rect 3142 9568 3148 9580
rect 3103 9540 3148 9568
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9568 3571 9571
rect 3878 9568 3884 9580
rect 3559 9540 3884 9568
rect 3559 9537 3571 9540
rect 3513 9531 3571 9537
rect 3878 9528 3884 9540
rect 3936 9528 3942 9580
rect 3988 9568 4016 9608
rect 4154 9596 4160 9608
rect 4212 9596 4218 9648
rect 4430 9596 4436 9648
rect 4488 9636 4494 9648
rect 4525 9639 4583 9645
rect 4525 9636 4537 9639
rect 4488 9608 4537 9636
rect 4488 9596 4494 9608
rect 4525 9605 4537 9608
rect 4571 9605 4583 9639
rect 4525 9599 4583 9605
rect 5074 9596 5080 9648
rect 5132 9636 5138 9648
rect 5132 9608 6500 9636
rect 5132 9596 5138 9608
rect 4798 9568 4804 9580
rect 3988 9540 4804 9568
rect 4798 9528 4804 9540
rect 4856 9528 4862 9580
rect 2406 9460 2412 9512
rect 2464 9500 2470 9512
rect 3237 9503 3295 9509
rect 3237 9500 3249 9503
rect 2464 9472 3249 9500
rect 2464 9460 2470 9472
rect 3237 9469 3249 9472
rect 3283 9469 3295 9503
rect 3237 9463 3295 9469
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9500 4491 9503
rect 5092 9500 5120 9596
rect 5442 9528 5448 9580
rect 5500 9568 5506 9580
rect 5721 9571 5779 9577
rect 5721 9568 5733 9571
rect 5500 9540 5733 9568
rect 5500 9528 5506 9540
rect 5721 9537 5733 9540
rect 5767 9537 5779 9571
rect 5721 9531 5779 9537
rect 5810 9528 5816 9580
rect 5868 9568 5874 9580
rect 5868 9540 5913 9568
rect 5868 9528 5874 9540
rect 5902 9500 5908 9512
rect 4479 9472 5120 9500
rect 5863 9472 5908 9500
rect 4479 9469 4491 9472
rect 4433 9463 4491 9469
rect 5902 9460 5908 9472
rect 5960 9460 5966 9512
rect 5994 9460 6000 9512
rect 6052 9500 6058 9512
rect 6365 9503 6423 9509
rect 6365 9500 6377 9503
rect 6052 9472 6377 9500
rect 6052 9460 6058 9472
rect 6365 9469 6377 9472
rect 6411 9469 6423 9503
rect 6472 9500 6500 9608
rect 6730 9596 6736 9648
rect 6788 9636 6794 9648
rect 6788 9608 8340 9636
rect 6788 9596 6794 9608
rect 8018 9528 8024 9580
rect 8076 9577 8082 9580
rect 8076 9568 8088 9577
rect 8076 9540 8121 9568
rect 8076 9531 8088 9540
rect 8076 9528 8082 9531
rect 8202 9528 8208 9580
rect 8260 9528 8266 9580
rect 8312 9577 8340 9608
rect 8478 9596 8484 9648
rect 8536 9636 8542 9648
rect 9674 9636 9680 9648
rect 8536 9608 9680 9636
rect 8536 9596 8542 9608
rect 9674 9596 9680 9608
rect 9732 9596 9738 9648
rect 9800 9639 9858 9645
rect 9800 9605 9812 9639
rect 9846 9636 9858 9639
rect 9950 9636 9956 9648
rect 9846 9608 9956 9636
rect 9846 9605 9858 9608
rect 9800 9599 9858 9605
rect 9950 9596 9956 9608
rect 10008 9596 10014 9648
rect 11054 9636 11060 9648
rect 10060 9608 11060 9636
rect 10060 9577 10088 9608
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 14366 9596 14372 9648
rect 14424 9636 14430 9648
rect 14734 9636 14740 9648
rect 14424 9608 14740 9636
rect 14424 9596 14430 9608
rect 14734 9596 14740 9608
rect 14792 9596 14798 9648
rect 8297 9571 8355 9577
rect 8297 9537 8309 9571
rect 8343 9537 8355 9571
rect 10045 9571 10103 9577
rect 8297 9531 8355 9537
rect 9048 9540 9996 9568
rect 6914 9500 6920 9512
rect 6472 9472 6920 9500
rect 6365 9463 6423 9469
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 8220 9500 8248 9528
rect 9048 9500 9076 9540
rect 8220 9472 9076 9500
rect 9968 9500 9996 9540
rect 10045 9537 10057 9571
rect 10091 9537 10103 9571
rect 10502 9568 10508 9580
rect 10463 9540 10508 9568
rect 10045 9531 10103 9537
rect 10502 9528 10508 9540
rect 10560 9528 10566 9580
rect 11882 9568 11888 9580
rect 11843 9540 11888 9568
rect 11882 9528 11888 9540
rect 11940 9528 11946 9580
rect 13538 9568 13544 9580
rect 13499 9540 13544 9568
rect 13538 9528 13544 9540
rect 13596 9528 13602 9580
rect 10318 9500 10324 9512
rect 9968 9472 10324 9500
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 10597 9503 10655 9509
rect 10597 9469 10609 9503
rect 10643 9469 10655 9503
rect 10597 9463 10655 9469
rect 10689 9503 10747 9509
rect 10689 9469 10701 9503
rect 10735 9469 10747 9503
rect 11698 9500 11704 9512
rect 11659 9472 11704 9500
rect 10689 9463 10747 9469
rect 1578 9392 1584 9444
rect 1636 9432 1642 9444
rect 1636 9404 2452 9432
rect 1636 9392 1642 9404
rect 2130 9364 2136 9376
rect 2091 9336 2136 9364
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 2222 9324 2228 9376
rect 2280 9364 2286 9376
rect 2424 9364 2452 9404
rect 2682 9392 2688 9444
rect 2740 9432 2746 9444
rect 2961 9435 3019 9441
rect 2961 9432 2973 9435
rect 2740 9404 2973 9432
rect 2740 9392 2746 9404
rect 2961 9401 2973 9404
rect 3007 9401 3019 9435
rect 5353 9435 5411 9441
rect 5353 9432 5365 9435
rect 2961 9395 3019 9401
rect 4080 9404 5365 9432
rect 4080 9364 4108 9404
rect 5353 9401 5365 9404
rect 5399 9401 5411 9435
rect 5353 9395 5411 9401
rect 10042 9392 10048 9444
rect 10100 9432 10106 9444
rect 10612 9432 10640 9463
rect 10100 9404 10640 9432
rect 10100 9392 10106 9404
rect 4982 9364 4988 9376
rect 2280 9336 2325 9364
rect 2424 9336 4108 9364
rect 4943 9336 4988 9364
rect 2280 9324 2286 9336
rect 4982 9324 4988 9336
rect 5040 9324 5046 9376
rect 5169 9367 5227 9373
rect 5169 9333 5181 9367
rect 5215 9364 5227 9367
rect 5258 9364 5264 9376
rect 5215 9336 5264 9364
rect 5215 9333 5227 9336
rect 5169 9327 5227 9333
rect 5258 9324 5264 9336
rect 5316 9324 5322 9376
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 6641 9367 6699 9373
rect 6641 9364 6653 9367
rect 6604 9336 6653 9364
rect 6604 9324 6610 9336
rect 6641 9333 6653 9336
rect 6687 9333 6699 9367
rect 6641 9327 6699 9333
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 8389 9367 8447 9373
rect 8389 9364 8401 9367
rect 6788 9336 8401 9364
rect 6788 9324 6794 9336
rect 8389 9333 8401 9336
rect 8435 9333 8447 9367
rect 8389 9327 8447 9333
rect 8665 9367 8723 9373
rect 8665 9333 8677 9367
rect 8711 9364 8723 9367
rect 9122 9364 9128 9376
rect 8711 9336 9128 9364
rect 8711 9333 8723 9336
rect 8665 9327 8723 9333
rect 9122 9324 9128 9336
rect 9180 9324 9186 9376
rect 10134 9364 10140 9376
rect 10095 9336 10140 9364
rect 10134 9324 10140 9336
rect 10192 9324 10198 9376
rect 10226 9324 10232 9376
rect 10284 9364 10290 9376
rect 10704 9364 10732 9463
rect 11698 9460 11704 9472
rect 11756 9460 11762 9512
rect 11793 9503 11851 9509
rect 11793 9469 11805 9503
rect 11839 9500 11851 9503
rect 12066 9500 12072 9512
rect 11839 9472 12072 9500
rect 11839 9469 11851 9472
rect 11793 9463 11851 9469
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 14366 9460 14372 9512
rect 14424 9500 14430 9512
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 14424 9472 14473 9500
rect 14424 9460 14430 9472
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 14461 9463 14519 9469
rect 12253 9435 12311 9441
rect 12253 9401 12265 9435
rect 12299 9432 12311 9435
rect 12618 9432 12624 9444
rect 12299 9404 12624 9432
rect 12299 9401 12311 9404
rect 12253 9395 12311 9401
rect 12618 9392 12624 9404
rect 12676 9392 12682 9444
rect 10284 9336 10732 9364
rect 10284 9324 10290 9336
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 2774 9160 2780 9172
rect 1412 9132 2780 9160
rect 1412 8965 1440 9132
rect 2774 9120 2780 9132
rect 2832 9160 2838 9172
rect 3970 9160 3976 9172
rect 2832 9132 3976 9160
rect 2832 9120 2838 9132
rect 3970 9120 3976 9132
rect 4028 9120 4034 9172
rect 5258 9120 5264 9172
rect 5316 9160 5322 9172
rect 5316 9132 5580 9160
rect 5316 9120 5322 9132
rect 2866 9092 2872 9104
rect 1964 9064 2872 9092
rect 1964 9036 1992 9064
rect 2866 9052 2872 9064
rect 2924 9092 2930 9104
rect 5552 9092 5580 9132
rect 5902 9120 5908 9172
rect 5960 9160 5966 9172
rect 5997 9163 6055 9169
rect 5997 9160 6009 9163
rect 5960 9132 6009 9160
rect 5960 9120 5966 9132
rect 5997 9129 6009 9132
rect 6043 9129 6055 9163
rect 7653 9163 7711 9169
rect 5997 9123 6055 9129
rect 6104 9132 7604 9160
rect 6104 9092 6132 9132
rect 2924 9064 4384 9092
rect 5552 9064 6132 9092
rect 7576 9092 7604 9132
rect 7653 9129 7665 9163
rect 7699 9160 7711 9163
rect 7834 9160 7840 9172
rect 7699 9132 7840 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 7834 9120 7840 9132
rect 7892 9120 7898 9172
rect 8570 9120 8576 9172
rect 8628 9160 8634 9172
rect 8665 9163 8723 9169
rect 8665 9160 8677 9163
rect 8628 9132 8677 9160
rect 8628 9120 8634 9132
rect 8665 9129 8677 9132
rect 8711 9129 8723 9163
rect 10502 9160 10508 9172
rect 8665 9123 8723 9129
rect 9232 9132 10508 9160
rect 8294 9092 8300 9104
rect 7576 9064 8300 9092
rect 2924 9052 2930 9064
rect 1946 9024 1952 9036
rect 1859 8996 1952 9024
rect 1946 8984 1952 8996
rect 2004 8984 2010 9036
rect 3050 8984 3056 9036
rect 3108 9024 3114 9036
rect 4356 9033 4384 9064
rect 8294 9052 8300 9064
rect 8352 9052 8358 9104
rect 3145 9027 3203 9033
rect 3145 9024 3157 9027
rect 3108 8996 3157 9024
rect 3108 8984 3114 8996
rect 3145 8993 3157 8996
rect 3191 8993 3203 9027
rect 3145 8987 3203 8993
rect 4341 9027 4399 9033
rect 4341 8993 4353 9027
rect 4387 8993 4399 9027
rect 4341 8987 4399 8993
rect 5718 8984 5724 9036
rect 5776 9024 5782 9036
rect 6089 9027 6147 9033
rect 6089 9024 6101 9027
rect 5776 8996 6101 9024
rect 5776 8984 5782 8996
rect 6089 8993 6101 8996
rect 6135 8993 6147 9027
rect 8205 9027 8263 9033
rect 8205 9024 8217 9027
rect 6089 8987 6147 8993
rect 7760 8996 8217 9024
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 2133 8959 2191 8965
rect 2133 8925 2145 8959
rect 2179 8956 2191 8959
rect 2866 8956 2872 8968
rect 2179 8928 2872 8956
rect 2179 8925 2191 8928
rect 2133 8919 2191 8925
rect 2866 8916 2872 8928
rect 2924 8916 2930 8968
rect 2958 8916 2964 8968
rect 3016 8956 3022 8968
rect 3234 8956 3240 8968
rect 3016 8928 3240 8956
rect 3016 8916 3022 8928
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 3418 8916 3424 8968
rect 3476 8916 3482 8968
rect 3878 8916 3884 8968
rect 3936 8956 3942 8968
rect 4617 8959 4675 8965
rect 3936 8928 4568 8956
rect 3936 8916 3942 8928
rect 2041 8891 2099 8897
rect 2041 8857 2053 8891
rect 2087 8888 2099 8891
rect 3053 8891 3111 8897
rect 2087 8860 2636 8888
rect 2087 8857 2099 8860
rect 2041 8851 2099 8857
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 2498 8820 2504 8832
rect 2459 8792 2504 8820
rect 2498 8780 2504 8792
rect 2556 8780 2562 8832
rect 2608 8829 2636 8860
rect 3053 8857 3065 8891
rect 3099 8888 3111 8891
rect 3436 8888 3464 8916
rect 3099 8860 3464 8888
rect 3099 8857 3111 8860
rect 3053 8851 3111 8857
rect 3970 8848 3976 8900
rect 4028 8888 4034 8900
rect 4540 8888 4568 8928
rect 4617 8925 4629 8959
rect 4663 8956 4675 8959
rect 5736 8956 5764 8984
rect 4663 8928 5764 8956
rect 6356 8959 6414 8965
rect 4663 8925 4675 8928
rect 4617 8919 4675 8925
rect 6356 8925 6368 8959
rect 6402 8956 6414 8959
rect 6638 8956 6644 8968
rect 6402 8928 6644 8956
rect 6402 8925 6414 8928
rect 6356 8919 6414 8925
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 4706 8888 4712 8900
rect 4028 8860 4476 8888
rect 4540 8860 4712 8888
rect 4028 8848 4034 8860
rect 2593 8823 2651 8829
rect 2593 8789 2605 8823
rect 2639 8789 2651 8823
rect 2593 8783 2651 8789
rect 3234 8780 3240 8832
rect 3292 8820 3298 8832
rect 3421 8823 3479 8829
rect 3421 8820 3433 8823
rect 3292 8792 3433 8820
rect 3292 8780 3298 8792
rect 3421 8789 3433 8792
rect 3467 8789 3479 8823
rect 3421 8783 3479 8789
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8820 3847 8823
rect 3878 8820 3884 8832
rect 3835 8792 3884 8820
rect 3835 8789 3847 8792
rect 3789 8783 3847 8789
rect 3878 8780 3884 8792
rect 3936 8780 3942 8832
rect 4154 8820 4160 8832
rect 4115 8792 4160 8820
rect 4154 8780 4160 8792
rect 4212 8780 4218 8832
rect 4246 8780 4252 8832
rect 4304 8820 4310 8832
rect 4448 8820 4476 8860
rect 4706 8848 4712 8860
rect 4764 8848 4770 8900
rect 4884 8891 4942 8897
rect 4884 8857 4896 8891
rect 4930 8888 4942 8891
rect 5902 8888 5908 8900
rect 4930 8860 5908 8888
rect 4930 8857 4942 8860
rect 4884 8851 4942 8857
rect 5902 8848 5908 8860
rect 5960 8848 5966 8900
rect 6730 8820 6736 8832
rect 4304 8792 4349 8820
rect 4448 8792 6736 8820
rect 4304 8780 4310 8792
rect 6730 8780 6736 8792
rect 6788 8780 6794 8832
rect 7466 8820 7472 8832
rect 7379 8792 7472 8820
rect 7466 8780 7472 8792
rect 7524 8820 7530 8832
rect 7760 8820 7788 8996
rect 8205 8993 8217 8996
rect 8251 8993 8263 9027
rect 8205 8987 8263 8993
rect 9125 9027 9183 9033
rect 9125 8993 9137 9027
rect 9171 9024 9183 9027
rect 9232 9024 9260 9132
rect 10502 9120 10508 9132
rect 10560 9120 10566 9172
rect 11882 9120 11888 9172
rect 11940 9160 11946 9172
rect 12161 9163 12219 9169
rect 12161 9160 12173 9163
rect 11940 9132 12173 9160
rect 11940 9120 11946 9132
rect 12161 9129 12173 9132
rect 12207 9129 12219 9163
rect 12161 9123 12219 9129
rect 10594 9052 10600 9104
rect 10652 9092 10658 9104
rect 17770 9092 17776 9104
rect 10652 9064 17776 9092
rect 10652 9052 10658 9064
rect 17770 9052 17776 9064
rect 17828 9052 17834 9104
rect 11054 9024 11060 9036
rect 9171 8996 9260 9024
rect 10336 8996 11060 9024
rect 9171 8993 9183 8996
rect 9125 8987 9183 8993
rect 8113 8959 8171 8965
rect 8113 8925 8125 8959
rect 8159 8956 8171 8959
rect 8570 8956 8576 8968
rect 8159 8928 8576 8956
rect 8159 8925 8171 8928
rect 8113 8919 8171 8925
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 10336 8956 10364 8996
rect 11054 8984 11060 8996
rect 11112 8984 11118 9036
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 11517 9027 11575 9033
rect 11517 9024 11529 9027
rect 11204 8996 11529 9024
rect 11204 8984 11210 8996
rect 11517 8993 11529 8996
rect 11563 9024 11575 9027
rect 11698 9024 11704 9036
rect 11563 8996 11704 9024
rect 11563 8993 11575 8996
rect 11517 8987 11575 8993
rect 11698 8984 11704 8996
rect 11756 8984 11762 9036
rect 13265 9027 13323 9033
rect 13265 8993 13277 9027
rect 13311 9024 13323 9027
rect 13814 9024 13820 9036
rect 13311 8996 13820 9024
rect 13311 8993 13323 8996
rect 13265 8987 13323 8993
rect 13814 8984 13820 8996
rect 13872 9024 13878 9036
rect 14185 9027 14243 9033
rect 14185 9024 14197 9027
rect 13872 8996 14197 9024
rect 13872 8984 13878 8996
rect 14185 8993 14197 8996
rect 14231 8993 14243 9027
rect 14185 8987 14243 8993
rect 15105 9027 15163 9033
rect 15105 8993 15117 9027
rect 15151 9024 15163 9027
rect 15562 9024 15568 9036
rect 15151 8996 15568 9024
rect 15151 8993 15163 8996
rect 15105 8987 15163 8993
rect 15562 8984 15568 8996
rect 15620 9024 15626 9036
rect 15620 8996 15792 9024
rect 15620 8984 15626 8996
rect 10594 8956 10600 8968
rect 9263 8928 10364 8956
rect 10428 8928 10600 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 7524 8792 7788 8820
rect 8021 8823 8079 8829
rect 7524 8780 7530 8792
rect 8021 8789 8033 8823
rect 8067 8820 8079 8823
rect 8478 8820 8484 8832
rect 8067 8792 8484 8820
rect 8067 8789 8079 8792
rect 8021 8783 8079 8789
rect 8478 8780 8484 8792
rect 8536 8780 8542 8832
rect 8588 8820 8616 8916
rect 8754 8848 8760 8900
rect 8812 8888 8818 8900
rect 9122 8888 9128 8900
rect 8812 8860 9128 8888
rect 8812 8848 8818 8860
rect 9122 8848 9128 8860
rect 9180 8888 9186 8900
rect 9484 8891 9542 8897
rect 9484 8888 9496 8891
rect 9180 8860 9496 8888
rect 9180 8848 9186 8860
rect 9484 8857 9496 8860
rect 9530 8888 9542 8891
rect 10226 8888 10232 8900
rect 9530 8860 10232 8888
rect 9530 8857 9542 8860
rect 9484 8851 9542 8857
rect 10226 8848 10232 8860
rect 10284 8848 10290 8900
rect 10428 8820 10456 8928
rect 10594 8916 10600 8928
rect 10652 8916 10658 8968
rect 10689 8959 10747 8965
rect 10689 8925 10701 8959
rect 10735 8925 10747 8959
rect 11790 8956 11796 8968
rect 11751 8928 11796 8956
rect 10689 8919 10747 8925
rect 10704 8888 10732 8919
rect 11790 8916 11796 8928
rect 11848 8916 11854 8968
rect 13446 8956 13452 8968
rect 13407 8928 13452 8956
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 14366 8916 14372 8968
rect 14424 8956 14430 8968
rect 14461 8959 14519 8965
rect 14461 8956 14473 8959
rect 14424 8928 14473 8956
rect 14424 8916 14430 8928
rect 14461 8925 14473 8928
rect 14507 8925 14519 8959
rect 14461 8919 14519 8925
rect 14826 8916 14832 8968
rect 14884 8916 14890 8968
rect 15764 8965 15792 8996
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8925 15807 8959
rect 15749 8919 15807 8925
rect 10612 8860 10732 8888
rect 11333 8891 11391 8897
rect 10612 8832 10640 8860
rect 11333 8857 11345 8891
rect 11379 8888 11391 8891
rect 12802 8888 12808 8900
rect 11379 8860 12808 8888
rect 11379 8857 11391 8860
rect 11333 8851 11391 8857
rect 12802 8848 12808 8860
rect 12860 8848 12866 8900
rect 12986 8848 12992 8900
rect 13044 8888 13050 8900
rect 13357 8891 13415 8897
rect 13357 8888 13369 8891
rect 13044 8860 13369 8888
rect 13044 8848 13050 8860
rect 13357 8857 13369 8860
rect 13403 8888 13415 8891
rect 13630 8888 13636 8900
rect 13403 8860 13636 8888
rect 13403 8857 13415 8860
rect 13357 8851 13415 8857
rect 13630 8848 13636 8860
rect 13688 8848 13694 8900
rect 14844 8888 14872 8916
rect 14384 8860 14872 8888
rect 10594 8820 10600 8832
rect 8588 8792 10456 8820
rect 10555 8792 10600 8820
rect 10594 8780 10600 8792
rect 10652 8780 10658 8832
rect 10962 8780 10968 8832
rect 11020 8820 11026 8832
rect 11701 8823 11759 8829
rect 11701 8820 11713 8823
rect 11020 8792 11713 8820
rect 11020 8780 11026 8792
rect 11701 8789 11713 8792
rect 11747 8789 11759 8823
rect 11701 8783 11759 8789
rect 13817 8823 13875 8829
rect 13817 8789 13829 8823
rect 13863 8820 13875 8823
rect 14274 8820 14280 8832
rect 13863 8792 14280 8820
rect 13863 8789 13875 8792
rect 13817 8783 13875 8789
rect 14274 8780 14280 8792
rect 14332 8780 14338 8832
rect 14384 8829 14412 8860
rect 14918 8848 14924 8900
rect 14976 8888 14982 8900
rect 15289 8891 15347 8897
rect 15289 8888 15301 8891
rect 14976 8860 15301 8888
rect 14976 8848 14982 8860
rect 15289 8857 15301 8860
rect 15335 8857 15347 8891
rect 15289 8851 15347 8857
rect 14369 8823 14427 8829
rect 14369 8789 14381 8823
rect 14415 8789 14427 8823
rect 14369 8783 14427 8789
rect 14550 8780 14556 8832
rect 14608 8820 14614 8832
rect 14829 8823 14887 8829
rect 14829 8820 14841 8823
rect 14608 8792 14841 8820
rect 14608 8780 14614 8792
rect 14829 8789 14841 8792
rect 14875 8789 14887 8823
rect 14829 8783 14887 8789
rect 15010 8780 15016 8832
rect 15068 8820 15074 8832
rect 15197 8823 15255 8829
rect 15197 8820 15209 8823
rect 15068 8792 15209 8820
rect 15068 8780 15074 8792
rect 15197 8789 15209 8792
rect 15243 8789 15255 8823
rect 15197 8783 15255 8789
rect 15378 8780 15384 8832
rect 15436 8820 15442 8832
rect 15657 8823 15715 8829
rect 15657 8820 15669 8823
rect 15436 8792 15669 8820
rect 15436 8780 15442 8792
rect 15657 8789 15669 8792
rect 15703 8789 15715 8823
rect 16390 8820 16396 8832
rect 16351 8792 16396 8820
rect 15657 8783 15715 8789
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 1104 8730 21896 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21896 8730
rect 1104 8656 21896 8678
rect 1946 8576 1952 8628
rect 2004 8616 2010 8628
rect 2133 8619 2191 8625
rect 2133 8616 2145 8619
rect 2004 8588 2145 8616
rect 2004 8576 2010 8588
rect 2133 8585 2145 8588
rect 2179 8585 2191 8619
rect 2133 8579 2191 8585
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 4212 8588 4445 8616
rect 4212 8576 4218 8588
rect 4433 8585 4445 8588
rect 4479 8585 4491 8619
rect 4433 8579 4491 8585
rect 4709 8619 4767 8625
rect 4709 8585 4721 8619
rect 4755 8616 4767 8619
rect 4982 8616 4988 8628
rect 4755 8588 4988 8616
rect 4755 8585 4767 8588
rect 4709 8579 4767 8585
rect 4982 8576 4988 8588
rect 5040 8616 5046 8628
rect 5626 8616 5632 8628
rect 5040 8588 5632 8616
rect 5040 8576 5046 8588
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 6365 8619 6423 8625
rect 6365 8616 6377 8619
rect 5868 8588 6377 8616
rect 5868 8576 5874 8588
rect 6365 8585 6377 8588
rect 6411 8585 6423 8619
rect 6365 8579 6423 8585
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 7285 8619 7343 8625
rect 7285 8616 7297 8619
rect 6779 8588 7297 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 7285 8585 7297 8588
rect 7331 8616 7343 8619
rect 7558 8616 7564 8628
rect 7331 8588 7564 8616
rect 7331 8585 7343 8588
rect 7285 8579 7343 8585
rect 7558 8576 7564 8588
rect 7616 8616 7622 8628
rect 7834 8616 7840 8628
rect 7616 8588 7840 8616
rect 7616 8576 7622 8588
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8018 8576 8024 8628
rect 8076 8616 8082 8628
rect 8113 8619 8171 8625
rect 8113 8616 8125 8619
rect 8076 8588 8125 8616
rect 8076 8576 8082 8588
rect 8113 8585 8125 8588
rect 8159 8585 8171 8619
rect 8113 8579 8171 8585
rect 8294 8576 8300 8628
rect 8352 8616 8358 8628
rect 8481 8619 8539 8625
rect 8481 8616 8493 8619
rect 8352 8588 8493 8616
rect 8352 8576 8358 8588
rect 8481 8585 8493 8588
rect 8527 8585 8539 8619
rect 8481 8579 8539 8585
rect 9033 8619 9091 8625
rect 9033 8585 9045 8619
rect 9079 8616 9091 8619
rect 9306 8616 9312 8628
rect 9079 8588 9312 8616
rect 9079 8585 9091 8588
rect 9033 8579 9091 8585
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 9493 8619 9551 8625
rect 9493 8585 9505 8619
rect 9539 8616 9551 8619
rect 9861 8619 9919 8625
rect 9861 8616 9873 8619
rect 9539 8588 9873 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 9861 8585 9873 8588
rect 9907 8585 9919 8619
rect 9861 8579 9919 8585
rect 9953 8619 10011 8625
rect 9953 8585 9965 8619
rect 9999 8616 10011 8619
rect 10134 8616 10140 8628
rect 9999 8588 10140 8616
rect 9999 8585 10011 8588
rect 9953 8579 10011 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 10318 8576 10324 8628
rect 10376 8616 10382 8628
rect 10962 8616 10968 8628
rect 10376 8588 10968 8616
rect 10376 8576 10382 8588
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11054 8576 11060 8628
rect 11112 8616 11118 8628
rect 11885 8619 11943 8625
rect 11885 8616 11897 8619
rect 11112 8588 11897 8616
rect 11112 8576 11118 8588
rect 11885 8585 11897 8588
rect 11931 8585 11943 8619
rect 11885 8579 11943 8585
rect 12066 8576 12072 8628
rect 12124 8616 12130 8628
rect 12253 8619 12311 8625
rect 12253 8616 12265 8619
rect 12124 8588 12265 8616
rect 12124 8576 12130 8588
rect 12253 8585 12265 8588
rect 12299 8585 12311 8619
rect 12253 8579 12311 8585
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 13722 8616 13728 8628
rect 12768 8588 13728 8616
rect 12768 8576 12774 8588
rect 13722 8576 13728 8588
rect 13780 8576 13786 8628
rect 14458 8576 14464 8628
rect 14516 8576 14522 8628
rect 15562 8616 15568 8628
rect 15523 8588 15568 8616
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 1397 8551 1455 8557
rect 1397 8517 1409 8551
rect 1443 8548 1455 8551
rect 2314 8548 2320 8560
rect 1443 8520 2320 8548
rect 1443 8517 1455 8520
rect 1397 8511 1455 8517
rect 2314 8508 2320 8520
rect 2372 8508 2378 8560
rect 3050 8508 3056 8560
rect 3108 8548 3114 8560
rect 3246 8551 3304 8557
rect 3246 8548 3258 8551
rect 3108 8520 3258 8548
rect 3108 8508 3114 8520
rect 3246 8517 3258 8520
rect 3292 8548 3304 8551
rect 5718 8548 5724 8560
rect 3292 8520 3464 8548
rect 3292 8517 3304 8520
rect 3246 8511 3304 8517
rect 3436 8492 3464 8520
rect 3528 8520 5724 8548
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 2958 8480 2964 8492
rect 2087 8452 2964 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2958 8440 2964 8452
rect 3016 8440 3022 8492
rect 3418 8480 3424 8492
rect 3331 8452 3424 8480
rect 3418 8440 3424 8452
rect 3476 8440 3482 8492
rect 3528 8489 3556 8520
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8449 3571 8483
rect 3513 8443 3571 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8480 4123 8483
rect 4154 8480 4160 8492
rect 4111 8452 4160 8480
rect 4111 8449 4123 8452
rect 4065 8443 4123 8449
rect 4154 8440 4160 8452
rect 4212 8480 4218 8492
rect 4430 8480 4436 8492
rect 4212 8452 4436 8480
rect 4212 8440 4218 8452
rect 4430 8440 4436 8452
rect 4488 8440 4494 8492
rect 4525 8483 4583 8489
rect 4525 8449 4537 8483
rect 4571 8480 4583 8483
rect 4614 8480 4620 8492
rect 4571 8452 4620 8480
rect 4571 8449 4583 8452
rect 4525 8443 4583 8449
rect 4614 8440 4620 8452
rect 4672 8440 4678 8492
rect 4816 8489 4844 8520
rect 5718 8508 5724 8520
rect 5776 8508 5782 8560
rect 6638 8508 6644 8560
rect 6696 8548 6702 8560
rect 8205 8551 8263 8557
rect 8205 8548 8217 8551
rect 6696 8520 8217 8548
rect 6696 8508 6702 8520
rect 8205 8517 8217 8520
rect 8251 8517 8263 8551
rect 8205 8511 8263 8517
rect 9214 8508 9220 8560
rect 9272 8548 9278 8560
rect 9272 8520 11192 8548
rect 9272 8508 9278 8520
rect 4801 8483 4859 8489
rect 4801 8449 4813 8483
rect 4847 8449 4859 8483
rect 4801 8443 4859 8449
rect 4890 8440 4896 8492
rect 4948 8480 4954 8492
rect 5057 8483 5115 8489
rect 5057 8480 5069 8483
rect 4948 8452 5069 8480
rect 4948 8440 4954 8452
rect 5057 8449 5069 8452
rect 5103 8449 5115 8483
rect 5057 8443 5115 8449
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 7098 8480 7104 8492
rect 6871 8452 7104 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 7098 8440 7104 8452
rect 7156 8440 7162 8492
rect 7466 8480 7472 8492
rect 7427 8452 7472 8480
rect 7466 8440 7472 8452
rect 7524 8440 7530 8492
rect 9122 8480 9128 8492
rect 9083 8452 9128 8480
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 11054 8480 11060 8492
rect 9232 8452 11060 8480
rect 3436 8412 3464 8440
rect 3789 8415 3847 8421
rect 3789 8412 3801 8415
rect 3436 8384 3801 8412
rect 3789 8381 3801 8384
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 3973 8415 4031 8421
rect 3973 8381 3985 8415
rect 4019 8412 4031 8415
rect 4706 8412 4712 8424
rect 4019 8384 4712 8412
rect 4019 8381 4031 8384
rect 3973 8375 4031 8381
rect 4706 8372 4712 8384
rect 4764 8372 4770 8424
rect 6917 8415 6975 8421
rect 6917 8412 6929 8415
rect 6196 8384 6929 8412
rect 1854 8304 1860 8356
rect 1912 8344 1918 8356
rect 1912 8316 2636 8344
rect 1912 8304 1918 8316
rect 2608 8276 2636 8316
rect 3528 8316 4844 8344
rect 3528 8276 3556 8316
rect 2608 8248 3556 8276
rect 4816 8276 4844 8316
rect 5902 8304 5908 8356
rect 5960 8344 5966 8356
rect 6196 8353 6224 8384
rect 6917 8381 6929 8384
rect 6963 8381 6975 8415
rect 6917 8375 6975 8381
rect 8754 8372 8760 8424
rect 8812 8412 8818 8424
rect 8849 8415 8907 8421
rect 8849 8412 8861 8415
rect 8812 8384 8861 8412
rect 8812 8372 8818 8384
rect 8849 8381 8861 8384
rect 8895 8381 8907 8415
rect 9232 8412 9260 8452
rect 11054 8440 11060 8452
rect 11112 8440 11118 8492
rect 8849 8375 8907 8381
rect 8956 8384 9260 8412
rect 9769 8415 9827 8421
rect 6181 8347 6239 8353
rect 6181 8344 6193 8347
rect 5960 8316 6193 8344
rect 5960 8304 5966 8316
rect 6181 8313 6193 8316
rect 6227 8313 6239 8347
rect 8956 8344 8984 8384
rect 9769 8381 9781 8415
rect 9815 8412 9827 8415
rect 10594 8412 10600 8424
rect 9815 8384 10600 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 10594 8372 10600 8384
rect 10652 8372 10658 8424
rect 11164 8421 11192 8520
rect 12158 8508 12164 8560
rect 12216 8548 12222 8560
rect 14476 8548 14504 8576
rect 12216 8520 14504 8548
rect 12216 8508 12222 8520
rect 12728 8489 12756 8520
rect 12713 8483 12771 8489
rect 12713 8449 12725 8483
rect 12759 8449 12771 8483
rect 12713 8443 12771 8449
rect 12980 8483 13038 8489
rect 12980 8449 12992 8483
rect 13026 8480 13038 8483
rect 13814 8480 13820 8492
rect 13026 8452 13820 8480
rect 13026 8449 13038 8452
rect 12980 8443 13038 8449
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 11698 8412 11704 8424
rect 11659 8384 11704 8412
rect 11149 8375 11207 8381
rect 11698 8372 11704 8384
rect 11756 8372 11762 8424
rect 11790 8372 11796 8424
rect 11848 8412 11854 8424
rect 11848 8384 11893 8412
rect 11848 8372 11854 8384
rect 6181 8307 6239 8313
rect 6288 8316 8984 8344
rect 10321 8347 10379 8353
rect 6288 8276 6316 8316
rect 10321 8313 10333 8347
rect 10367 8344 10379 8347
rect 12710 8344 12716 8356
rect 10367 8316 12716 8344
rect 10367 8313 10379 8316
rect 10321 8307 10379 8313
rect 12710 8304 12716 8316
rect 12768 8304 12774 8356
rect 10594 8276 10600 8288
rect 4816 8248 6316 8276
rect 10555 8248 10600 8276
rect 10594 8236 10600 8248
rect 10652 8236 10658 8288
rect 13740 8276 13768 8452
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 14200 8489 14228 8520
rect 14185 8483 14243 8489
rect 14185 8449 14197 8483
rect 14231 8449 14243 8483
rect 14441 8483 14499 8489
rect 14441 8480 14453 8483
rect 14185 8443 14243 8449
rect 14292 8452 14453 8480
rect 14292 8412 14320 8452
rect 14441 8449 14453 8452
rect 14487 8449 14499 8483
rect 14441 8443 14499 8449
rect 14108 8384 14320 8412
rect 13814 8304 13820 8356
rect 13872 8344 13878 8356
rect 14108 8353 14136 8384
rect 14093 8347 14151 8353
rect 14093 8344 14105 8347
rect 13872 8316 14105 8344
rect 13872 8304 13878 8316
rect 14093 8313 14105 8316
rect 14139 8313 14151 8347
rect 14093 8307 14151 8313
rect 14366 8276 14372 8288
rect 13740 8248 14372 8276
rect 14366 8236 14372 8248
rect 14424 8236 14430 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 1397 8075 1455 8081
rect 1397 8041 1409 8075
rect 1443 8072 1455 8075
rect 1486 8072 1492 8084
rect 1443 8044 1492 8072
rect 1443 8041 1455 8044
rect 1397 8035 1455 8041
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 2866 8072 2872 8084
rect 2827 8044 2872 8072
rect 2866 8032 2872 8044
rect 2924 8032 2930 8084
rect 3789 8075 3847 8081
rect 3789 8041 3801 8075
rect 3835 8072 3847 8075
rect 4246 8072 4252 8084
rect 3835 8044 4252 8072
rect 3835 8041 3847 8044
rect 3789 8035 3847 8041
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 5166 8072 5172 8084
rect 5127 8044 5172 8072
rect 5166 8032 5172 8044
rect 5224 8032 5230 8084
rect 5718 8072 5724 8084
rect 5679 8044 5724 8072
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 5810 8032 5816 8084
rect 5868 8072 5874 8084
rect 7098 8072 7104 8084
rect 5868 8044 6960 8072
rect 7059 8044 7104 8072
rect 5868 8032 5874 8044
rect 6546 8004 6552 8016
rect 2884 7976 6552 8004
rect 2884 7948 2912 7976
rect 2866 7896 2872 7948
rect 2924 7896 2930 7948
rect 3418 7936 3424 7948
rect 3379 7908 3424 7936
rect 3418 7896 3424 7908
rect 3476 7936 3482 7948
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 3476 7908 4353 7936
rect 3476 7896 3482 7908
rect 4341 7905 4353 7908
rect 4387 7905 4399 7939
rect 4939 7936 4967 7976
rect 6546 7964 6552 7976
rect 6604 7964 6610 8016
rect 6932 8004 6960 8044
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 9122 8032 9128 8084
rect 9180 8072 9186 8084
rect 9217 8075 9275 8081
rect 9217 8072 9229 8075
rect 9180 8044 9229 8072
rect 9180 8032 9186 8044
rect 9217 8041 9229 8044
rect 9263 8041 9275 8075
rect 9217 8035 9275 8041
rect 12894 8032 12900 8084
rect 12952 8072 12958 8084
rect 14829 8075 14887 8081
rect 12952 8044 14780 8072
rect 12952 8032 12958 8044
rect 8662 8004 8668 8016
rect 6932 7976 8668 8004
rect 8662 7964 8668 7976
rect 8720 7964 8726 8016
rect 14752 8004 14780 8044
rect 14829 8041 14841 8075
rect 14875 8072 14887 8075
rect 14918 8072 14924 8084
rect 14875 8044 14924 8072
rect 14875 8041 14887 8044
rect 14829 8035 14887 8041
rect 14918 8032 14924 8044
rect 14976 8032 14982 8084
rect 15013 8007 15071 8013
rect 15013 8004 15025 8007
rect 14752 7976 15025 8004
rect 15013 7973 15025 7976
rect 15059 8004 15071 8007
rect 15194 8004 15200 8016
rect 15059 7976 15200 8004
rect 15059 7973 15071 7976
rect 15013 7967 15071 7973
rect 15194 7964 15200 7976
rect 15252 7964 15258 8016
rect 4939 7908 5028 7936
rect 4341 7899 4399 7905
rect 2222 7828 2228 7880
rect 2280 7868 2286 7880
rect 2510 7871 2568 7877
rect 2510 7868 2522 7871
rect 2280 7840 2522 7868
rect 2280 7828 2286 7840
rect 2510 7837 2522 7840
rect 2556 7837 2568 7871
rect 2774 7868 2780 7880
rect 2735 7840 2780 7868
rect 2510 7831 2568 7837
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 3234 7868 3240 7880
rect 3195 7840 3240 7868
rect 3234 7828 3240 7840
rect 3292 7828 3298 7880
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 5000 7877 5028 7908
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 7653 7939 7711 7945
rect 7653 7936 7665 7939
rect 5684 7908 7665 7936
rect 5684 7896 5690 7908
rect 7653 7905 7665 7908
rect 7699 7905 7711 7939
rect 7653 7899 7711 7905
rect 9122 7896 9128 7948
rect 9180 7936 9186 7948
rect 9398 7936 9404 7948
rect 9180 7908 9404 7936
rect 9180 7896 9186 7908
rect 9398 7896 9404 7908
rect 9456 7936 9462 7948
rect 9677 7939 9735 7945
rect 9677 7936 9689 7939
rect 9456 7908 9689 7936
rect 9456 7896 9462 7908
rect 9677 7905 9689 7908
rect 9723 7905 9735 7939
rect 9677 7899 9735 7905
rect 9861 7939 9919 7945
rect 9861 7905 9873 7939
rect 9907 7936 9919 7939
rect 9950 7936 9956 7948
rect 9907 7908 9956 7936
rect 9907 7905 9919 7908
rect 9861 7899 9919 7905
rect 9950 7896 9956 7908
rect 10008 7896 10014 7948
rect 10244 7908 12434 7936
rect 4157 7871 4215 7877
rect 3384 7840 3429 7868
rect 3384 7828 3390 7840
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 4893 7871 4951 7877
rect 4203 7840 4844 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 2222 7692 2228 7744
rect 2280 7732 2286 7744
rect 3326 7732 3332 7744
rect 2280 7704 3332 7732
rect 2280 7692 2286 7704
rect 3326 7692 3332 7704
rect 3384 7692 3390 7744
rect 4246 7732 4252 7744
rect 4207 7704 4252 7732
rect 4246 7692 4252 7704
rect 4304 7692 4310 7744
rect 4706 7732 4712 7744
rect 4667 7704 4712 7732
rect 4706 7692 4712 7704
rect 4764 7692 4770 7744
rect 4816 7732 4844 7840
rect 4893 7837 4905 7871
rect 4939 7837 4951 7871
rect 4893 7831 4951 7837
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7837 5043 7871
rect 4985 7831 5043 7837
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7868 7527 7871
rect 7558 7868 7564 7880
rect 7515 7840 7564 7868
rect 7515 7837 7527 7840
rect 7469 7831 7527 7837
rect 4908 7800 4936 7831
rect 7558 7828 7564 7840
rect 7616 7828 7622 7880
rect 7926 7868 7932 7880
rect 7887 7840 7932 7868
rect 7926 7828 7932 7840
rect 7984 7828 7990 7880
rect 10244 7868 10272 7908
rect 10410 7868 10416 7880
rect 8680 7840 10272 7868
rect 10371 7840 10416 7868
rect 5074 7800 5080 7812
rect 4908 7772 5080 7800
rect 5074 7760 5080 7772
rect 5132 7800 5138 7812
rect 5534 7800 5540 7812
rect 5132 7772 5540 7800
rect 5132 7760 5138 7772
rect 5534 7760 5540 7772
rect 5592 7760 5598 7812
rect 7006 7800 7012 7812
rect 6967 7772 7012 7800
rect 7006 7760 7012 7772
rect 7064 7760 7070 7812
rect 8680 7809 8708 7840
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 8665 7803 8723 7809
rect 8665 7800 8677 7803
rect 7576 7772 8677 7800
rect 6546 7732 6552 7744
rect 4816 7704 6552 7732
rect 6546 7692 6552 7704
rect 6604 7692 6610 7744
rect 6822 7692 6828 7744
rect 6880 7732 6886 7744
rect 7576 7741 7604 7772
rect 8665 7769 8677 7772
rect 8711 7769 8723 7803
rect 12158 7800 12164 7812
rect 12119 7772 12164 7800
rect 8665 7763 8723 7769
rect 12158 7760 12164 7772
rect 12216 7760 12222 7812
rect 12406 7800 12434 7908
rect 13814 7896 13820 7948
rect 13872 7936 13878 7948
rect 14185 7939 14243 7945
rect 14185 7936 14197 7939
rect 13872 7908 14197 7936
rect 13872 7896 13878 7908
rect 14185 7905 14197 7908
rect 14231 7905 14243 7939
rect 14185 7899 14243 7905
rect 14274 7896 14280 7948
rect 14332 7936 14338 7948
rect 14369 7939 14427 7945
rect 14369 7936 14381 7939
rect 14332 7908 14381 7936
rect 14332 7896 14338 7908
rect 14369 7905 14381 7908
rect 14415 7905 14427 7939
rect 14369 7899 14427 7905
rect 14458 7896 14464 7948
rect 14516 7936 14522 7948
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 14516 7908 15301 7936
rect 14516 7896 14522 7908
rect 15289 7905 15301 7908
rect 15335 7905 15347 7939
rect 15289 7899 15347 7905
rect 12802 7828 12808 7880
rect 12860 7868 12866 7880
rect 13366 7871 13424 7877
rect 13366 7868 13378 7871
rect 12860 7840 13378 7868
rect 12860 7828 12866 7840
rect 13366 7837 13378 7840
rect 13412 7837 13424 7871
rect 13630 7868 13636 7880
rect 13591 7840 13636 7868
rect 13366 7831 13424 7837
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 15556 7871 15614 7877
rect 15556 7837 15568 7871
rect 15602 7868 15614 7871
rect 16390 7868 16396 7880
rect 15602 7840 16396 7868
rect 15602 7837 15614 7840
rect 15556 7831 15614 7837
rect 16390 7828 16396 7840
rect 16448 7828 16454 7880
rect 13722 7800 13728 7812
rect 12406 7772 13728 7800
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 14461 7803 14519 7809
rect 14461 7769 14473 7803
rect 14507 7800 14519 7803
rect 14550 7800 14556 7812
rect 14507 7772 14556 7800
rect 14507 7769 14519 7772
rect 14461 7763 14519 7769
rect 14550 7760 14556 7772
rect 14608 7760 14614 7812
rect 14844 7772 16712 7800
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 6880 7704 7573 7732
rect 6880 7692 6886 7704
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 8570 7732 8576 7744
rect 8531 7704 8576 7732
rect 7561 7695 7619 7701
rect 8570 7692 8576 7704
rect 8628 7692 8634 7744
rect 9122 7732 9128 7744
rect 9083 7704 9128 7732
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 9582 7732 9588 7744
rect 9543 7704 9588 7732
rect 9582 7692 9588 7704
rect 9640 7692 9646 7744
rect 10226 7732 10232 7744
rect 10187 7704 10232 7732
rect 10226 7692 10232 7704
rect 10284 7692 10290 7744
rect 10962 7692 10968 7744
rect 11020 7732 11026 7744
rect 12253 7735 12311 7741
rect 12253 7732 12265 7735
rect 11020 7704 12265 7732
rect 11020 7692 11026 7704
rect 12253 7701 12265 7704
rect 12299 7732 12311 7735
rect 12618 7732 12624 7744
rect 12299 7704 12624 7732
rect 12299 7701 12311 7704
rect 12253 7695 12311 7701
rect 12618 7692 12624 7704
rect 12676 7692 12682 7744
rect 13078 7692 13084 7744
rect 13136 7732 13142 7744
rect 14844 7732 14872 7772
rect 16684 7741 16712 7772
rect 13136 7704 14872 7732
rect 16669 7735 16727 7741
rect 13136 7692 13142 7704
rect 16669 7701 16681 7735
rect 16715 7732 16727 7735
rect 16942 7732 16948 7744
rect 16715 7704 16948 7732
rect 16715 7701 16727 7704
rect 16669 7695 16727 7701
rect 16942 7692 16948 7704
rect 17000 7692 17006 7744
rect 1104 7642 21896 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21896 7642
rect 1104 7568 21896 7590
rect 2317 7531 2375 7537
rect 2317 7497 2329 7531
rect 2363 7528 2375 7531
rect 2498 7528 2504 7540
rect 2363 7500 2504 7528
rect 2363 7497 2375 7500
rect 2317 7491 2375 7497
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 2685 7531 2743 7537
rect 2685 7497 2697 7531
rect 2731 7528 2743 7531
rect 3050 7528 3056 7540
rect 2731 7500 3056 7528
rect 2731 7497 2743 7500
rect 2685 7491 2743 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 3234 7528 3240 7540
rect 3191 7500 3240 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 3510 7528 3516 7540
rect 3471 7500 3516 7528
rect 3510 7488 3516 7500
rect 3568 7488 3574 7540
rect 4341 7531 4399 7537
rect 4341 7497 4353 7531
rect 4387 7497 4399 7531
rect 4341 7491 4399 7497
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 4982 7528 4988 7540
rect 4939 7500 4988 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 2225 7463 2283 7469
rect 2225 7429 2237 7463
rect 2271 7460 2283 7463
rect 3878 7460 3884 7472
rect 2271 7432 3884 7460
rect 2271 7429 2283 7432
rect 2225 7423 2283 7429
rect 3878 7420 3884 7432
rect 3936 7420 3942 7472
rect 4356 7460 4384 7491
rect 4982 7488 4988 7500
rect 5040 7488 5046 7540
rect 5442 7528 5448 7540
rect 5403 7500 5448 7528
rect 5442 7488 5448 7500
rect 5500 7488 5506 7540
rect 5813 7531 5871 7537
rect 5813 7497 5825 7531
rect 5859 7528 5871 7531
rect 5994 7528 6000 7540
rect 5859 7500 6000 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 5994 7488 6000 7500
rect 6052 7488 6058 7540
rect 8202 7488 8208 7540
rect 8260 7528 8266 7540
rect 8478 7528 8484 7540
rect 8260 7500 8484 7528
rect 8260 7488 8266 7500
rect 8478 7488 8484 7500
rect 8536 7488 8542 7540
rect 8665 7531 8723 7537
rect 8665 7497 8677 7531
rect 8711 7497 8723 7531
rect 8665 7491 8723 7497
rect 6914 7460 6920 7472
rect 4356 7432 6920 7460
rect 6914 7420 6920 7432
rect 6972 7420 6978 7472
rect 7552 7463 7610 7469
rect 7552 7429 7564 7463
rect 7598 7460 7610 7463
rect 8570 7460 8576 7472
rect 7598 7432 8576 7460
rect 7598 7429 7610 7432
rect 7552 7423 7610 7429
rect 8570 7420 8576 7432
rect 8628 7420 8634 7472
rect 8680 7460 8708 7491
rect 9490 7488 9496 7540
rect 9548 7528 9554 7540
rect 9585 7531 9643 7537
rect 9585 7528 9597 7531
rect 9548 7500 9597 7528
rect 9548 7488 9554 7500
rect 9585 7497 9597 7500
rect 9631 7528 9643 7531
rect 9858 7528 9864 7540
rect 9631 7500 9864 7528
rect 9631 7497 9643 7500
rect 9585 7491 9643 7497
rect 9858 7488 9864 7500
rect 9916 7488 9922 7540
rect 9953 7531 10011 7537
rect 9953 7497 9965 7531
rect 9999 7528 10011 7531
rect 10042 7528 10048 7540
rect 9999 7500 10048 7528
rect 9999 7497 10011 7500
rect 9953 7491 10011 7497
rect 10042 7488 10048 7500
rect 10100 7488 10106 7540
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 10413 7531 10471 7537
rect 10413 7528 10425 7531
rect 10284 7500 10425 7528
rect 10284 7488 10290 7500
rect 10413 7497 10425 7500
rect 10459 7497 10471 7531
rect 10413 7491 10471 7497
rect 10870 7488 10876 7540
rect 10928 7528 10934 7540
rect 12434 7528 12440 7540
rect 10928 7500 12440 7528
rect 10928 7488 10934 7500
rect 12434 7488 12440 7500
rect 12492 7488 12498 7540
rect 12526 7488 12532 7540
rect 12584 7528 12590 7540
rect 13265 7531 13323 7537
rect 13265 7528 13277 7531
rect 12584 7500 13277 7528
rect 12584 7488 12590 7500
rect 13265 7497 13277 7500
rect 13311 7497 13323 7531
rect 13265 7491 13323 7497
rect 13354 7488 13360 7540
rect 13412 7528 13418 7540
rect 13412 7500 13457 7528
rect 13412 7488 13418 7500
rect 13722 7488 13728 7540
rect 13780 7528 13786 7540
rect 13817 7531 13875 7537
rect 13817 7528 13829 7531
rect 13780 7500 13829 7528
rect 13780 7488 13786 7500
rect 13817 7497 13829 7500
rect 13863 7497 13875 7531
rect 13817 7491 13875 7497
rect 14277 7531 14335 7537
rect 14277 7497 14289 7531
rect 14323 7528 14335 7531
rect 14829 7531 14887 7537
rect 14829 7528 14841 7531
rect 14323 7500 14841 7528
rect 14323 7497 14335 7500
rect 14277 7491 14335 7497
rect 14829 7497 14841 7500
rect 14875 7497 14887 7531
rect 15194 7528 15200 7540
rect 15155 7500 15200 7528
rect 14829 7491 14887 7497
rect 8941 7463 8999 7469
rect 8941 7460 8953 7463
rect 8680 7432 8953 7460
rect 8941 7429 8953 7432
rect 8987 7460 8999 7463
rect 9214 7460 9220 7472
rect 8987 7432 9220 7460
rect 8987 7429 8999 7432
rect 8941 7423 8999 7429
rect 9214 7420 9220 7432
rect 9272 7420 9278 7472
rect 11241 7463 11299 7469
rect 11241 7460 11253 7463
rect 9324 7432 11253 7460
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 1670 7392 1676 7404
rect 1631 7364 1676 7392
rect 1670 7352 1676 7364
rect 1728 7392 1734 7404
rect 3053 7395 3111 7401
rect 1728 7364 2774 7392
rect 1728 7352 1734 7364
rect 1486 7284 1492 7336
rect 1544 7324 1550 7336
rect 2041 7327 2099 7333
rect 2041 7324 2053 7327
rect 1544 7296 2053 7324
rect 1544 7284 1550 7296
rect 2041 7293 2053 7296
rect 2087 7293 2099 7327
rect 2041 7287 2099 7293
rect 2314 7284 2320 7336
rect 2372 7324 2378 7336
rect 2590 7324 2596 7336
rect 2372 7296 2596 7324
rect 2372 7284 2378 7296
rect 2590 7284 2596 7296
rect 2648 7284 2654 7336
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 2498 7256 2504 7268
rect 1627 7228 2504 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 2498 7216 2504 7228
rect 2556 7216 2562 7268
rect 2746 7256 2774 7364
rect 3053 7361 3065 7395
rect 3099 7392 3111 7395
rect 3970 7392 3976 7404
rect 3099 7364 3188 7392
rect 3931 7364 3976 7392
rect 3099 7361 3111 7364
rect 3053 7355 3111 7361
rect 2958 7324 2964 7336
rect 2919 7296 2964 7324
rect 2958 7284 2964 7296
rect 3016 7284 3022 7336
rect 3160 7324 3188 7364
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 4246 7352 4252 7404
rect 4304 7392 4310 7404
rect 4985 7395 5043 7401
rect 4985 7392 4997 7395
rect 4304 7364 4997 7392
rect 4304 7352 4310 7364
rect 4985 7361 4997 7364
rect 5031 7392 5043 7395
rect 5350 7392 5356 7404
rect 5031 7364 5356 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 5350 7352 5356 7364
rect 5408 7352 5414 7404
rect 6086 7352 6092 7404
rect 6144 7392 6150 7404
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 6144 7364 6745 7392
rect 6144 7352 6150 7364
rect 6733 7361 6745 7364
rect 6779 7361 6791 7395
rect 9324 7392 9352 7432
rect 11241 7429 11253 7432
rect 11287 7429 11299 7463
rect 11241 7423 11299 7429
rect 12158 7420 12164 7472
rect 12216 7460 12222 7472
rect 13832 7460 13860 7491
rect 15194 7488 15200 7500
rect 15252 7528 15258 7540
rect 15930 7528 15936 7540
rect 15252 7500 15936 7528
rect 15252 7488 15258 7500
rect 15930 7488 15936 7500
rect 15988 7488 15994 7540
rect 15289 7463 15347 7469
rect 15289 7460 15301 7463
rect 12216 7432 12940 7460
rect 13832 7432 15301 7460
rect 12216 7420 12222 7432
rect 6733 7355 6791 7361
rect 6840 7364 9352 7392
rect 3326 7324 3332 7336
rect 3160 7296 3332 7324
rect 3326 7284 3332 7296
rect 3384 7284 3390 7336
rect 3418 7284 3424 7336
rect 3476 7324 3482 7336
rect 3697 7327 3755 7333
rect 3697 7324 3709 7327
rect 3476 7296 3709 7324
rect 3476 7284 3482 7296
rect 3697 7293 3709 7296
rect 3743 7293 3755 7327
rect 3878 7324 3884 7336
rect 3839 7296 3884 7324
rect 3697 7287 3755 7293
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 4801 7327 4859 7333
rect 4801 7293 4813 7327
rect 4847 7324 4859 7327
rect 5442 7324 5448 7336
rect 4847 7296 5448 7324
rect 4847 7293 4859 7296
rect 4801 7287 4859 7293
rect 5442 7284 5448 7296
rect 5500 7284 5506 7336
rect 5718 7284 5724 7336
rect 5776 7324 5782 7336
rect 5905 7327 5963 7333
rect 5905 7324 5917 7327
rect 5776 7296 5917 7324
rect 5776 7284 5782 7296
rect 5905 7293 5917 7296
rect 5951 7293 5963 7327
rect 5905 7287 5963 7293
rect 5994 7284 6000 7336
rect 6052 7324 6058 7336
rect 6546 7324 6552 7336
rect 6052 7296 6097 7324
rect 6507 7296 6552 7324
rect 6052 7284 6058 7296
rect 6546 7284 6552 7296
rect 6604 7284 6610 7336
rect 6641 7327 6699 7333
rect 6641 7293 6653 7327
rect 6687 7293 6699 7327
rect 6641 7287 6699 7293
rect 5353 7259 5411 7265
rect 2746 7228 4568 7256
rect 1857 7191 1915 7197
rect 1857 7157 1869 7191
rect 1903 7188 1915 7191
rect 4246 7188 4252 7200
rect 1903 7160 4252 7188
rect 1903 7157 1915 7160
rect 1857 7151 1915 7157
rect 4246 7148 4252 7160
rect 4304 7148 4310 7200
rect 4430 7188 4436 7200
rect 4391 7160 4436 7188
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 4540 7188 4568 7228
rect 5353 7225 5365 7259
rect 5399 7256 5411 7259
rect 6656 7256 6684 7287
rect 5399 7228 6684 7256
rect 5399 7225 5411 7228
rect 5353 7219 5411 7225
rect 6840 7188 6868 7364
rect 9858 7352 9864 7404
rect 9916 7392 9922 7404
rect 10321 7395 10379 7401
rect 10321 7392 10333 7395
rect 9916 7364 10333 7392
rect 9916 7352 9922 7364
rect 10321 7361 10333 7364
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 12618 7352 12624 7404
rect 12676 7401 12682 7404
rect 12912 7401 12940 7432
rect 15289 7429 15301 7432
rect 15335 7460 15347 7463
rect 16298 7460 16304 7472
rect 15335 7432 16304 7460
rect 15335 7429 15347 7432
rect 15289 7423 15347 7429
rect 16298 7420 16304 7432
rect 16356 7420 16362 7472
rect 12676 7392 12688 7401
rect 12897 7395 12955 7401
rect 12676 7364 12721 7392
rect 12676 7355 12688 7364
rect 12897 7361 12909 7395
rect 12943 7361 12955 7395
rect 12897 7355 12955 7361
rect 12676 7352 12682 7355
rect 13446 7352 13452 7404
rect 13504 7392 13510 7404
rect 14369 7395 14427 7401
rect 14369 7392 14381 7395
rect 13504 7364 14381 7392
rect 13504 7352 13510 7364
rect 14369 7361 14381 7364
rect 14415 7361 14427 7395
rect 14369 7355 14427 7361
rect 7282 7324 7288 7336
rect 7243 7296 7288 7324
rect 7282 7284 7288 7296
rect 7340 7284 7346 7336
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7293 9459 7327
rect 9401 7287 9459 7293
rect 9416 7256 9444 7287
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 10134 7324 10140 7336
rect 9548 7296 9593 7324
rect 10095 7296 10140 7324
rect 9548 7284 9554 7296
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 11057 7327 11115 7333
rect 11057 7324 11069 7327
rect 10336 7296 11069 7324
rect 9950 7256 9956 7268
rect 8220 7228 9352 7256
rect 9416 7228 9956 7256
rect 7098 7188 7104 7200
rect 4540 7160 6868 7188
rect 7059 7160 7104 7188
rect 7098 7148 7104 7160
rect 7156 7148 7162 7200
rect 7190 7148 7196 7200
rect 7248 7188 7254 7200
rect 8220 7188 8248 7228
rect 7248 7160 8248 7188
rect 8849 7191 8907 7197
rect 7248 7148 7254 7160
rect 8849 7157 8861 7191
rect 8895 7188 8907 7191
rect 9214 7188 9220 7200
rect 8895 7160 9220 7188
rect 8895 7157 8907 7160
rect 8849 7151 8907 7157
rect 9214 7148 9220 7160
rect 9272 7148 9278 7200
rect 9324 7188 9352 7228
rect 9950 7216 9956 7228
rect 10008 7216 10014 7268
rect 10336 7188 10364 7296
rect 11057 7293 11069 7296
rect 11103 7293 11115 7327
rect 13078 7324 13084 7336
rect 13039 7296 13084 7324
rect 11057 7287 11115 7293
rect 13078 7284 13084 7296
rect 13136 7284 13142 7336
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 14093 7327 14151 7333
rect 14093 7324 14105 7327
rect 13872 7296 14105 7324
rect 13872 7284 13878 7296
rect 14093 7293 14105 7296
rect 14139 7293 14151 7327
rect 14093 7287 14151 7293
rect 14458 7284 14464 7336
rect 14516 7324 14522 7336
rect 15381 7327 15439 7333
rect 14516 7296 15240 7324
rect 14516 7284 14522 7296
rect 10686 7216 10692 7268
rect 10744 7256 10750 7268
rect 11517 7259 11575 7265
rect 11517 7256 11529 7259
rect 10744 7228 11529 7256
rect 10744 7216 10750 7228
rect 11517 7225 11529 7228
rect 11563 7225 11575 7259
rect 11517 7219 11575 7225
rect 13725 7259 13783 7265
rect 13725 7225 13737 7259
rect 13771 7256 13783 7259
rect 14737 7259 14795 7265
rect 13771 7228 14688 7256
rect 13771 7225 13783 7228
rect 13725 7219 13783 7225
rect 10778 7188 10784 7200
rect 9324 7160 10364 7188
rect 10739 7160 10784 7188
rect 10778 7148 10784 7160
rect 10836 7148 10842 7200
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 14660 7188 14688 7228
rect 14737 7225 14749 7259
rect 14783 7256 14795 7259
rect 15010 7256 15016 7268
rect 14783 7228 15016 7256
rect 14783 7225 14795 7228
rect 14737 7219 14795 7225
rect 15010 7216 15016 7228
rect 15068 7216 15074 7268
rect 15212 7256 15240 7296
rect 15381 7293 15393 7327
rect 15427 7293 15439 7327
rect 15381 7287 15439 7293
rect 15396 7256 15424 7287
rect 15212 7228 15424 7256
rect 16390 7188 16396 7200
rect 10928 7160 10973 7188
rect 14660 7160 16396 7188
rect 10928 7148 10934 7160
rect 16390 7148 16396 7160
rect 16448 7148 16454 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 2869 6987 2927 6993
rect 2869 6953 2881 6987
rect 2915 6984 2927 6987
rect 3326 6984 3332 6996
rect 2915 6956 3332 6984
rect 2915 6953 2927 6956
rect 2869 6947 2927 6953
rect 3326 6944 3332 6956
rect 3384 6944 3390 6996
rect 4154 6944 4160 6996
rect 4212 6984 4218 6996
rect 4430 6984 4436 6996
rect 4212 6956 4436 6984
rect 4212 6944 4218 6956
rect 4430 6944 4436 6956
rect 4488 6984 4494 6996
rect 5166 6984 5172 6996
rect 4488 6956 5172 6984
rect 4488 6944 4494 6956
rect 5166 6944 5172 6956
rect 5224 6984 5230 6996
rect 5718 6984 5724 6996
rect 5224 6956 5724 6984
rect 5224 6944 5230 6956
rect 5718 6944 5724 6956
rect 5776 6944 5782 6996
rect 6086 6984 6092 6996
rect 6047 6956 6092 6984
rect 6086 6944 6092 6956
rect 6144 6944 6150 6996
rect 7190 6984 7196 6996
rect 6196 6956 7196 6984
rect 2777 6919 2835 6925
rect 2777 6885 2789 6919
rect 2823 6916 2835 6919
rect 3970 6916 3976 6928
rect 2823 6888 3976 6916
rect 2823 6885 2835 6888
rect 2777 6879 2835 6885
rect 3970 6876 3976 6888
rect 4028 6876 4034 6928
rect 4982 6916 4988 6928
rect 4448 6888 4988 6916
rect 1762 6848 1768 6860
rect 1412 6820 1768 6848
rect 1412 6792 1440 6820
rect 1762 6808 1768 6820
rect 1820 6808 1826 6860
rect 2225 6851 2283 6857
rect 2225 6817 2237 6851
rect 2271 6848 2283 6851
rect 2498 6848 2504 6860
rect 2271 6820 2504 6848
rect 2271 6817 2283 6820
rect 2225 6811 2283 6817
rect 2498 6808 2504 6820
rect 2556 6808 2562 6860
rect 3418 6848 3424 6860
rect 3379 6820 3424 6848
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6848 4307 6851
rect 4338 6848 4344 6860
rect 4295 6820 4344 6848
rect 4295 6817 4307 6820
rect 4249 6811 4307 6817
rect 1394 6780 1400 6792
rect 1355 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6740 1458 6792
rect 1670 6780 1676 6792
rect 1631 6752 1676 6780
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6780 2375 6783
rect 3694 6780 3700 6792
rect 2363 6752 3700 6780
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 3694 6740 3700 6752
rect 3752 6740 3758 6792
rect 4264 6712 4292 6811
rect 4338 6808 4344 6820
rect 4396 6808 4402 6860
rect 4448 6857 4476 6888
rect 4982 6876 4988 6888
rect 5040 6876 5046 6928
rect 5350 6876 5356 6928
rect 5408 6916 5414 6928
rect 6196 6916 6224 6956
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 7374 6944 7380 6996
rect 7432 6984 7438 6996
rect 7561 6987 7619 6993
rect 7561 6984 7573 6987
rect 7432 6956 7573 6984
rect 7432 6944 7438 6956
rect 7561 6953 7573 6956
rect 7607 6984 7619 6987
rect 7926 6984 7932 6996
rect 7607 6956 7932 6984
rect 7607 6953 7619 6956
rect 7561 6947 7619 6953
rect 7926 6944 7932 6956
rect 7984 6944 7990 6996
rect 9122 6984 9128 6996
rect 8036 6956 9128 6984
rect 8036 6916 8064 6956
rect 9122 6944 9128 6956
rect 9180 6944 9186 6996
rect 10042 6944 10048 6996
rect 10100 6984 10106 6996
rect 10870 6984 10876 6996
rect 10100 6956 10876 6984
rect 10100 6944 10106 6956
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 12713 6987 12771 6993
rect 12713 6953 12725 6987
rect 12759 6984 12771 6987
rect 13446 6984 13452 6996
rect 12759 6956 13452 6984
rect 12759 6953 12771 6956
rect 12713 6947 12771 6953
rect 13446 6944 13452 6956
rect 13504 6944 13510 6996
rect 15654 6984 15660 6996
rect 14476 6956 15660 6984
rect 5408 6888 6224 6916
rect 7668 6888 8064 6916
rect 8128 6888 8340 6916
rect 5408 6876 5414 6888
rect 4433 6851 4491 6857
rect 4433 6817 4445 6851
rect 4479 6817 4491 6851
rect 4433 6811 4491 6817
rect 4617 6851 4675 6857
rect 4617 6817 4629 6851
rect 4663 6848 4675 6851
rect 4890 6848 4896 6860
rect 4663 6820 4896 6848
rect 4663 6817 4675 6820
rect 4617 6811 4675 6817
rect 4890 6808 4896 6820
rect 4948 6808 4954 6860
rect 5442 6848 5448 6860
rect 5403 6820 5448 6848
rect 5442 6808 5448 6820
rect 5500 6808 5506 6860
rect 7466 6808 7472 6860
rect 7524 6848 7530 6860
rect 7668 6848 7696 6888
rect 7524 6820 7696 6848
rect 7524 6808 7530 6820
rect 7742 6808 7748 6860
rect 7800 6848 7806 6860
rect 8128 6848 8156 6888
rect 7800 6820 8156 6848
rect 8205 6851 8263 6857
rect 7800 6808 7806 6820
rect 8205 6817 8217 6851
rect 8251 6817 8263 6851
rect 8312 6848 8340 6888
rect 8478 6876 8484 6928
rect 8536 6916 8542 6928
rect 8938 6916 8944 6928
rect 8536 6888 8944 6916
rect 8536 6876 8542 6888
rect 8938 6876 8944 6888
rect 8996 6876 9002 6928
rect 10318 6876 10324 6928
rect 10376 6916 10382 6928
rect 10965 6919 11023 6925
rect 10965 6916 10977 6919
rect 10376 6888 10977 6916
rect 10376 6876 10382 6888
rect 10965 6885 10977 6888
rect 11011 6885 11023 6919
rect 14093 6919 14151 6925
rect 14093 6916 14105 6919
rect 10965 6879 11023 6885
rect 12176 6888 14105 6916
rect 8665 6851 8723 6857
rect 8665 6848 8677 6851
rect 8312 6820 8677 6848
rect 8205 6811 8263 6817
rect 8665 6817 8677 6820
rect 8711 6817 8723 6851
rect 8665 6811 8723 6817
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6780 5319 6783
rect 5626 6780 5632 6792
rect 5307 6752 5632 6780
rect 5307 6749 5319 6752
rect 5261 6743 5319 6749
rect 5626 6740 5632 6752
rect 5684 6740 5690 6792
rect 5994 6740 6000 6792
rect 6052 6780 6058 6792
rect 6181 6783 6239 6789
rect 6181 6780 6193 6783
rect 6052 6752 6193 6780
rect 6052 6740 6058 6752
rect 6181 6749 6193 6752
rect 6227 6780 6239 6783
rect 7282 6780 7288 6792
rect 6227 6752 7288 6780
rect 6227 6749 6239 6752
rect 6181 6743 6239 6749
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 8220 6780 8248 6811
rect 8754 6808 8760 6860
rect 8812 6848 8818 6860
rect 9125 6851 9183 6857
rect 9125 6848 9137 6851
rect 8812 6820 9137 6848
rect 8812 6808 8818 6820
rect 9125 6817 9137 6820
rect 9171 6817 9183 6851
rect 9125 6811 9183 6817
rect 9493 6851 9551 6857
rect 9493 6817 9505 6851
rect 9539 6848 9551 6851
rect 9858 6848 9864 6860
rect 9539 6820 9864 6848
rect 9539 6817 9551 6820
rect 9493 6811 9551 6817
rect 9858 6808 9864 6820
rect 9916 6848 9922 6860
rect 10134 6848 10140 6860
rect 9916 6820 10140 6848
rect 9916 6808 9922 6820
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 10226 6808 10232 6860
rect 10284 6848 10290 6860
rect 12176 6857 12204 6888
rect 14093 6885 14105 6888
rect 14139 6916 14151 6919
rect 14366 6916 14372 6928
rect 14139 6888 14372 6916
rect 14139 6885 14151 6888
rect 14093 6879 14151 6885
rect 14366 6876 14372 6888
rect 14424 6876 14430 6928
rect 10689 6851 10747 6857
rect 10689 6848 10701 6851
rect 10284 6820 10701 6848
rect 10284 6808 10290 6820
rect 10689 6817 10701 6820
rect 10735 6848 10747 6851
rect 11517 6851 11575 6857
rect 11517 6848 11529 6851
rect 10735 6820 11529 6848
rect 10735 6817 10747 6820
rect 10689 6811 10747 6817
rect 11517 6817 11529 6820
rect 11563 6817 11575 6851
rect 11517 6811 11575 6817
rect 12161 6851 12219 6857
rect 12161 6817 12173 6851
rect 12207 6817 12219 6851
rect 12802 6848 12808 6860
rect 12763 6820 12808 6848
rect 12161 6811 12219 6817
rect 12802 6808 12808 6820
rect 12860 6808 12866 6860
rect 12894 6808 12900 6860
rect 12952 6848 12958 6860
rect 14476 6848 14504 6956
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 12952 6820 14504 6848
rect 15473 6851 15531 6857
rect 12952 6808 12958 6820
rect 15473 6817 15485 6851
rect 15519 6848 15531 6851
rect 15746 6848 15752 6860
rect 15519 6820 15752 6848
rect 15519 6817 15531 6820
rect 15473 6811 15531 6817
rect 7392 6752 8248 6780
rect 1872 6684 4292 6712
rect 6448 6715 6506 6721
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 1762 6644 1768 6656
rect 1627 6616 1768 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 1762 6604 1768 6616
rect 1820 6604 1826 6656
rect 1872 6653 1900 6684
rect 6448 6681 6460 6715
rect 6494 6712 6506 6715
rect 6546 6712 6552 6724
rect 6494 6684 6552 6712
rect 6494 6681 6506 6684
rect 6448 6675 6506 6681
rect 6546 6672 6552 6684
rect 6604 6712 6610 6724
rect 6604 6684 6868 6712
rect 6604 6672 6610 6684
rect 1857 6647 1915 6653
rect 1857 6613 1869 6647
rect 1903 6613 1915 6647
rect 1857 6607 1915 6613
rect 2409 6647 2467 6653
rect 2409 6613 2421 6647
rect 2455 6644 2467 6647
rect 2958 6644 2964 6656
rect 2455 6616 2964 6644
rect 2455 6613 2467 6616
rect 2409 6607 2467 6613
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 3234 6644 3240 6656
rect 3195 6616 3240 6644
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 3326 6604 3332 6656
rect 3384 6644 3390 6656
rect 3786 6644 3792 6656
rect 3384 6616 3429 6644
rect 3747 6616 3792 6644
rect 3384 6604 3390 6616
rect 3786 6604 3792 6616
rect 3844 6604 3850 6656
rect 4157 6647 4215 6653
rect 4157 6613 4169 6647
rect 4203 6644 4215 6647
rect 4522 6644 4528 6656
rect 4203 6616 4528 6644
rect 4203 6613 4215 6616
rect 4157 6607 4215 6613
rect 4522 6604 4528 6616
rect 4580 6604 4586 6656
rect 5534 6604 5540 6656
rect 5592 6644 5598 6656
rect 5629 6647 5687 6653
rect 5629 6644 5641 6647
rect 5592 6616 5641 6644
rect 5592 6604 5598 6616
rect 5629 6613 5641 6616
rect 5675 6613 5687 6647
rect 5629 6607 5687 6613
rect 5721 6647 5779 6653
rect 5721 6613 5733 6647
rect 5767 6644 5779 6647
rect 6638 6644 6644 6656
rect 5767 6616 6644 6644
rect 5767 6613 5779 6616
rect 5721 6607 5779 6613
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 6840 6644 6868 6684
rect 7392 6644 7420 6752
rect 8386 6740 8392 6792
rect 8444 6780 8450 6792
rect 9582 6780 9588 6792
rect 8444 6752 9588 6780
rect 8444 6740 8450 6752
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 10962 6740 10968 6792
rect 11020 6780 11026 6792
rect 12253 6783 12311 6789
rect 12253 6780 12265 6783
rect 11020 6752 12265 6780
rect 11020 6740 11026 6752
rect 12253 6749 12265 6752
rect 12299 6749 12311 6783
rect 12253 6743 12311 6749
rect 12342 6740 12348 6792
rect 12400 6780 12406 6792
rect 12400 6752 12445 6780
rect 12400 6740 12406 6752
rect 13354 6740 13360 6792
rect 13412 6780 13418 6792
rect 13630 6780 13636 6792
rect 13412 6752 13636 6780
rect 13412 6740 13418 6752
rect 13630 6740 13636 6752
rect 13688 6780 13694 6792
rect 15488 6780 15516 6811
rect 15746 6808 15752 6820
rect 15804 6808 15810 6860
rect 13688 6752 15516 6780
rect 15565 6783 15623 6789
rect 13688 6740 13694 6752
rect 15565 6749 15577 6783
rect 15611 6780 15623 6783
rect 15654 6780 15660 6792
rect 15611 6752 15660 6780
rect 15611 6749 15623 6752
rect 15565 6743 15623 6749
rect 15654 6740 15660 6752
rect 15712 6740 15718 6792
rect 7926 6672 7932 6724
rect 7984 6712 7990 6724
rect 8021 6715 8079 6721
rect 8021 6712 8033 6715
rect 7984 6684 8033 6712
rect 7984 6672 7990 6684
rect 8021 6681 8033 6684
rect 8067 6681 8079 6715
rect 8021 6675 8079 6681
rect 8202 6672 8208 6724
rect 8260 6712 8266 6724
rect 8481 6715 8539 6721
rect 8481 6712 8493 6715
rect 8260 6684 8493 6712
rect 8260 6672 8266 6684
rect 8481 6681 8493 6684
rect 8527 6681 8539 6715
rect 8481 6675 8539 6681
rect 8662 6672 8668 6724
rect 8720 6712 8726 6724
rect 9490 6712 9496 6724
rect 8720 6684 9496 6712
rect 8720 6672 8726 6684
rect 9490 6672 9496 6684
rect 9548 6712 9554 6724
rect 9677 6715 9735 6721
rect 9677 6712 9689 6715
rect 9548 6684 9689 6712
rect 9548 6672 9554 6684
rect 9677 6681 9689 6684
rect 9723 6681 9735 6715
rect 10505 6715 10563 6721
rect 9677 6675 9735 6681
rect 10060 6684 10456 6712
rect 6840 6616 7420 6644
rect 7650 6604 7656 6656
rect 7708 6644 7714 6656
rect 8110 6644 8116 6656
rect 7708 6616 7753 6644
rect 8071 6616 8116 6644
rect 7708 6604 7714 6616
rect 8110 6604 8116 6616
rect 8168 6604 8174 6656
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 9950 6644 9956 6656
rect 9364 6616 9956 6644
rect 9364 6604 9370 6616
rect 9950 6604 9956 6616
rect 10008 6604 10014 6656
rect 10060 6653 10088 6684
rect 10045 6647 10103 6653
rect 10045 6613 10057 6647
rect 10091 6613 10103 6647
rect 10045 6607 10103 6613
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 10428 6644 10456 6684
rect 10505 6681 10517 6715
rect 10551 6712 10563 6715
rect 15228 6715 15286 6721
rect 10551 6684 10732 6712
rect 10551 6681 10563 6684
rect 10505 6675 10563 6681
rect 10597 6647 10655 6653
rect 10597 6644 10609 6647
rect 10192 6616 10237 6644
rect 10428 6616 10609 6644
rect 10192 6604 10198 6616
rect 10597 6613 10609 6616
rect 10643 6613 10655 6647
rect 10704 6644 10732 6684
rect 15228 6681 15240 6715
rect 15274 6712 15286 6715
rect 15470 6712 15476 6724
rect 15274 6684 15476 6712
rect 15274 6681 15286 6684
rect 15228 6675 15286 6681
rect 15470 6672 15476 6684
rect 15528 6672 15534 6724
rect 16206 6712 16212 6724
rect 16167 6684 16212 6712
rect 16206 6672 16212 6684
rect 16264 6672 16270 6724
rect 10778 6644 10784 6656
rect 10704 6616 10784 6644
rect 10597 6607 10655 6613
rect 10778 6604 10784 6616
rect 10836 6604 10842 6656
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11333 6647 11391 6653
rect 11333 6644 11345 6647
rect 11296 6616 11345 6644
rect 11296 6604 11302 6616
rect 11333 6613 11345 6616
rect 11379 6613 11391 6647
rect 11333 6607 11391 6613
rect 11425 6647 11483 6653
rect 11425 6613 11437 6647
rect 11471 6644 11483 6647
rect 11698 6644 11704 6656
rect 11471 6616 11704 6644
rect 11471 6613 11483 6616
rect 11425 6607 11483 6613
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 13906 6644 13912 6656
rect 11848 6616 11893 6644
rect 13867 6616 13912 6644
rect 11848 6604 11854 6616
rect 13906 6604 13912 6616
rect 13964 6604 13970 6656
rect 14734 6604 14740 6656
rect 14792 6644 14798 6656
rect 15654 6644 15660 6656
rect 14792 6616 15660 6644
rect 14792 6604 14798 6616
rect 15654 6604 15660 6616
rect 15712 6604 15718 6656
rect 1104 6554 21896 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21896 6554
rect 1104 6480 21896 6502
rect 1765 6443 1823 6449
rect 1765 6409 1777 6443
rect 1811 6440 1823 6443
rect 2590 6440 2596 6452
rect 1811 6412 2596 6440
rect 1811 6409 1823 6412
rect 1765 6403 1823 6409
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 3142 6400 3148 6452
rect 3200 6440 3206 6452
rect 3329 6443 3387 6449
rect 3329 6440 3341 6443
rect 3200 6412 3341 6440
rect 3200 6400 3206 6412
rect 3329 6409 3341 6412
rect 3375 6409 3387 6443
rect 3786 6440 3792 6452
rect 3747 6412 3792 6440
rect 3329 6403 3387 6409
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 4338 6400 4344 6452
rect 4396 6440 4402 6452
rect 4798 6440 4804 6452
rect 4396 6412 4804 6440
rect 4396 6400 4402 6412
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 6181 6443 6239 6449
rect 6181 6409 6193 6443
rect 6227 6440 6239 6443
rect 6546 6440 6552 6452
rect 6227 6412 6552 6440
rect 6227 6409 6239 6412
rect 6181 6403 6239 6409
rect 6546 6400 6552 6412
rect 6604 6400 6610 6452
rect 7098 6440 7104 6452
rect 7059 6412 7104 6440
rect 7098 6400 7104 6412
rect 7156 6400 7162 6452
rect 7193 6443 7251 6449
rect 7193 6409 7205 6443
rect 7239 6440 7251 6443
rect 7650 6440 7656 6452
rect 7239 6412 7656 6440
rect 7239 6409 7251 6412
rect 7193 6403 7251 6409
rect 7650 6400 7656 6412
rect 7708 6400 7714 6452
rect 8297 6443 8355 6449
rect 8297 6409 8309 6443
rect 8343 6440 8355 6443
rect 8570 6440 8576 6452
rect 8343 6412 8576 6440
rect 8343 6409 8355 6412
rect 8297 6403 8355 6409
rect 8570 6400 8576 6412
rect 8628 6400 8634 6452
rect 8754 6400 8760 6452
rect 8812 6440 8818 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 8812 6412 9505 6440
rect 8812 6400 8818 6412
rect 9493 6409 9505 6412
rect 9539 6409 9551 6443
rect 9493 6403 9551 6409
rect 9582 6400 9588 6452
rect 9640 6440 9646 6452
rect 11241 6443 11299 6449
rect 11241 6440 11253 6443
rect 9640 6412 11253 6440
rect 9640 6400 9646 6412
rect 11241 6409 11253 6412
rect 11287 6409 11299 6443
rect 11241 6403 11299 6409
rect 11882 6400 11888 6452
rect 11940 6440 11946 6452
rect 12253 6443 12311 6449
rect 12253 6440 12265 6443
rect 11940 6412 12265 6440
rect 11940 6400 11946 6412
rect 12253 6409 12265 6412
rect 12299 6409 12311 6443
rect 12986 6440 12992 6452
rect 12947 6412 12992 6440
rect 12253 6403 12311 6409
rect 12986 6400 12992 6412
rect 13044 6400 13050 6452
rect 13906 6400 13912 6452
rect 13964 6440 13970 6452
rect 16025 6443 16083 6449
rect 16025 6440 16037 6443
rect 13964 6412 16037 6440
rect 13964 6400 13970 6412
rect 16025 6409 16037 6412
rect 16071 6409 16083 6443
rect 16025 6403 16083 6409
rect 16390 6400 16396 6452
rect 16448 6440 16454 6452
rect 17129 6443 17187 6449
rect 17129 6440 17141 6443
rect 16448 6412 17141 6440
rect 16448 6400 16454 6412
rect 17129 6409 17141 6412
rect 17175 6409 17187 6443
rect 21358 6440 21364 6452
rect 21319 6412 21364 6440
rect 17129 6403 17187 6409
rect 21358 6400 21364 6412
rect 21416 6400 21422 6452
rect 2682 6372 2688 6384
rect 1872 6344 2688 6372
rect 1397 6307 1455 6313
rect 1397 6273 1409 6307
rect 1443 6304 1455 6307
rect 1578 6304 1584 6316
rect 1443 6276 1584 6304
rect 1443 6273 1455 6276
rect 1397 6267 1455 6273
rect 1578 6264 1584 6276
rect 1636 6264 1642 6316
rect 1872 6313 1900 6344
rect 2682 6332 2688 6344
rect 2740 6332 2746 6384
rect 2774 6332 2780 6384
rect 2832 6372 2838 6384
rect 5068 6375 5126 6381
rect 2832 6344 3013 6372
rect 2832 6332 2838 6344
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6273 1915 6307
rect 1857 6267 1915 6273
rect 1946 6264 1952 6316
rect 2004 6304 2010 6316
rect 2113 6307 2171 6313
rect 2113 6304 2125 6307
rect 2004 6276 2125 6304
rect 2004 6264 2010 6276
rect 2113 6273 2125 6276
rect 2159 6304 2171 6307
rect 2985 6304 3013 6344
rect 3620 6344 5028 6372
rect 3620 6304 3648 6344
rect 2159 6276 2912 6304
rect 2985 6276 3648 6304
rect 3697 6307 3755 6313
rect 2159 6273 2171 6276
rect 2113 6267 2171 6273
rect 1581 6103 1639 6109
rect 1581 6069 1593 6103
rect 1627 6100 1639 6103
rect 2774 6100 2780 6112
rect 1627 6072 2780 6100
rect 1627 6069 1639 6072
rect 1581 6063 1639 6069
rect 2774 6060 2780 6072
rect 2832 6060 2838 6112
rect 2884 6100 2912 6276
rect 3697 6273 3709 6307
rect 3743 6304 3755 6307
rect 4157 6307 4215 6313
rect 4157 6304 4169 6307
rect 3743 6276 4169 6304
rect 3743 6273 3755 6276
rect 3697 6267 3755 6273
rect 4157 6273 4169 6276
rect 4203 6273 4215 6307
rect 4157 6267 4215 6273
rect 4433 6307 4491 6313
rect 4433 6273 4445 6307
rect 4479 6304 4491 6307
rect 4522 6304 4528 6316
rect 4479 6276 4528 6304
rect 4479 6273 4491 6276
rect 4433 6267 4491 6273
rect 4522 6264 4528 6276
rect 4580 6264 4586 6316
rect 5000 6304 5028 6344
rect 5068 6341 5080 6375
rect 5114 6372 5126 6375
rect 5442 6372 5448 6384
rect 5114 6344 5448 6372
rect 5114 6341 5126 6344
rect 5068 6335 5126 6341
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 5810 6332 5816 6384
rect 5868 6372 5874 6384
rect 11517 6375 11575 6381
rect 11517 6372 11529 6375
rect 5868 6344 6316 6372
rect 5868 6332 5874 6344
rect 6288 6304 6316 6344
rect 9499 6344 11529 6372
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 5000 6276 6224 6304
rect 6288 6276 6377 6304
rect 3418 6236 3424 6248
rect 3331 6208 3424 6236
rect 3050 6128 3056 6180
rect 3108 6168 3114 6180
rect 3237 6171 3295 6177
rect 3237 6168 3249 6171
rect 3108 6140 3249 6168
rect 3108 6128 3114 6140
rect 3237 6137 3249 6140
rect 3283 6137 3295 6171
rect 3237 6131 3295 6137
rect 3344 6100 3372 6208
rect 3418 6196 3424 6208
rect 3476 6236 3482 6248
rect 3881 6239 3939 6245
rect 3881 6236 3893 6239
rect 3476 6208 3893 6236
rect 3476 6196 3482 6208
rect 3881 6205 3893 6208
rect 3927 6205 3939 6239
rect 4798 6236 4804 6248
rect 4759 6208 4804 6236
rect 3881 6199 3939 6205
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 6196 6236 6224 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 7208 6276 7696 6304
rect 7208 6236 7236 6276
rect 7374 6236 7380 6248
rect 6196 6208 7236 6236
rect 7335 6208 7380 6236
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 7668 6236 7696 6276
rect 7742 6264 7748 6316
rect 7800 6304 7806 6316
rect 7800 6276 7845 6304
rect 7800 6264 7806 6276
rect 8202 6264 8208 6316
rect 8260 6308 8266 6316
rect 8389 6308 8447 6313
rect 8260 6307 8616 6308
rect 8260 6280 8401 6307
rect 8260 6264 8266 6280
rect 8389 6273 8401 6280
rect 8435 6304 8616 6307
rect 8849 6307 8907 6313
rect 8435 6280 8800 6304
rect 8435 6273 8447 6280
rect 8588 6276 8800 6280
rect 8389 6267 8447 6273
rect 8294 6236 8300 6248
rect 7668 6208 8300 6236
rect 8294 6196 8300 6208
rect 8352 6196 8358 6248
rect 8570 6196 8576 6248
rect 8628 6236 8634 6248
rect 8772 6236 8800 6276
rect 8849 6273 8861 6307
rect 8895 6304 8907 6307
rect 9122 6304 9128 6316
rect 8895 6276 9128 6304
rect 8895 6273 8907 6276
rect 8849 6267 8907 6273
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 8628 6208 8673 6236
rect 8772 6208 8984 6236
rect 8628 6196 8634 6208
rect 3694 6128 3700 6180
rect 3752 6168 3758 6180
rect 4430 6168 4436 6180
rect 3752 6140 4436 6168
rect 3752 6128 3758 6140
rect 4430 6128 4436 6140
rect 4488 6128 4494 6180
rect 6914 6128 6920 6180
rect 6972 6168 6978 6180
rect 8478 6168 8484 6180
rect 6972 6140 8484 6168
rect 6972 6128 6978 6140
rect 8478 6128 8484 6140
rect 8536 6128 8542 6180
rect 8846 6128 8852 6180
rect 8904 6128 8910 6180
rect 2884 6072 3372 6100
rect 4617 6103 4675 6109
rect 4617 6069 4629 6103
rect 4663 6100 4675 6103
rect 5166 6100 5172 6112
rect 4663 6072 5172 6100
rect 4663 6069 4675 6072
rect 4617 6063 4675 6069
rect 5166 6060 5172 6072
rect 5224 6060 5230 6112
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 6546 6100 6552 6112
rect 5592 6072 6552 6100
rect 5592 6060 5598 6072
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 6638 6060 6644 6112
rect 6696 6100 6702 6112
rect 6733 6103 6791 6109
rect 6733 6100 6745 6103
rect 6696 6072 6745 6100
rect 6696 6060 6702 6072
rect 6733 6069 6745 6072
rect 6779 6069 6791 6103
rect 6733 6063 6791 6069
rect 7098 6060 7104 6112
rect 7156 6100 7162 6112
rect 7561 6103 7619 6109
rect 7561 6100 7573 6103
rect 7156 6072 7573 6100
rect 7156 6060 7162 6072
rect 7561 6069 7573 6072
rect 7607 6069 7619 6103
rect 7926 6100 7932 6112
rect 7887 6072 7932 6100
rect 7561 6063 7619 6069
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 8864 6100 8892 6128
rect 8352 6072 8892 6100
rect 8956 6100 8984 6208
rect 9398 6196 9404 6248
rect 9456 6236 9462 6248
rect 9499 6236 9527 6344
rect 11517 6341 11529 6344
rect 11563 6341 11575 6375
rect 11517 6335 11575 6341
rect 11974 6332 11980 6384
rect 12032 6372 12038 6384
rect 12069 6375 12127 6381
rect 12069 6372 12081 6375
rect 12032 6344 12081 6372
rect 12032 6332 12038 6344
rect 12069 6341 12081 6344
rect 12115 6341 12127 6375
rect 12894 6372 12900 6384
rect 12855 6344 12900 6372
rect 12069 6335 12127 6341
rect 12894 6332 12900 6344
rect 12952 6332 12958 6384
rect 15197 6375 15255 6381
rect 15197 6341 15209 6375
rect 15243 6372 15255 6375
rect 15286 6372 15292 6384
rect 15243 6344 15292 6372
rect 15243 6341 15255 6344
rect 15197 6335 15255 6341
rect 15286 6332 15292 6344
rect 15344 6332 15350 6384
rect 15562 6332 15568 6384
rect 15620 6372 15626 6384
rect 16117 6375 16175 6381
rect 16117 6372 16129 6375
rect 15620 6344 16129 6372
rect 15620 6332 15626 6344
rect 16117 6341 16129 6344
rect 16163 6341 16175 6375
rect 16117 6335 16175 6341
rect 9585 6307 9643 6313
rect 9585 6273 9597 6307
rect 9631 6304 9643 6307
rect 9674 6304 9680 6316
rect 9631 6276 9680 6304
rect 9631 6273 9643 6276
rect 9585 6267 9643 6273
rect 9674 6264 9680 6276
rect 9732 6264 9738 6316
rect 9858 6313 9864 6316
rect 9852 6267 9864 6313
rect 9916 6304 9922 6316
rect 10686 6304 10692 6316
rect 9916 6276 10692 6304
rect 9858 6264 9864 6267
rect 9916 6264 9922 6276
rect 10686 6264 10692 6276
rect 10744 6264 10750 6316
rect 10778 6264 10784 6316
rect 10836 6304 10842 6316
rect 10836 6276 12434 6304
rect 10836 6264 10842 6276
rect 9456 6208 9527 6236
rect 12406 6236 12434 6276
rect 12526 6264 12532 6316
rect 12584 6304 12590 6316
rect 13354 6304 13360 6316
rect 12584 6276 13360 6304
rect 12584 6264 12590 6276
rect 13354 6264 13360 6276
rect 13412 6264 13418 6316
rect 13630 6313 13636 6316
rect 13624 6304 13636 6313
rect 13591 6276 13636 6304
rect 13624 6267 13636 6276
rect 13630 6264 13636 6267
rect 13688 6264 13694 6316
rect 15470 6308 15476 6316
rect 15396 6280 15476 6308
rect 12621 6239 12679 6245
rect 12621 6236 12633 6239
rect 12406 6208 12633 6236
rect 9456 6196 9462 6208
rect 12621 6205 12633 6208
rect 12667 6205 12679 6239
rect 12621 6199 12679 6205
rect 12894 6196 12900 6248
rect 12952 6236 12958 6248
rect 12952 6208 13400 6236
rect 12952 6196 12958 6208
rect 11054 6128 11060 6180
rect 11112 6168 11118 6180
rect 13262 6168 13268 6180
rect 11112 6140 13268 6168
rect 11112 6128 11118 6140
rect 13262 6128 13268 6140
rect 13320 6128 13326 6180
rect 9858 6100 9864 6112
rect 8956 6072 9864 6100
rect 8352 6060 8358 6072
rect 9858 6060 9864 6072
rect 9916 6060 9922 6112
rect 10226 6060 10232 6112
rect 10284 6100 10290 6112
rect 10965 6103 11023 6109
rect 10965 6100 10977 6103
rect 10284 6072 10977 6100
rect 10284 6060 10290 6072
rect 10965 6069 10977 6072
rect 11011 6069 11023 6103
rect 10965 6063 11023 6069
rect 11149 6103 11207 6109
rect 11149 6069 11161 6103
rect 11195 6100 11207 6103
rect 11330 6100 11336 6112
rect 11195 6072 11336 6100
rect 11195 6069 11207 6072
rect 11149 6063 11207 6069
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 11606 6060 11612 6112
rect 11664 6100 11670 6112
rect 11701 6103 11759 6109
rect 11701 6100 11713 6103
rect 11664 6072 11713 6100
rect 11664 6060 11670 6072
rect 11701 6069 11713 6072
rect 11747 6069 11759 6103
rect 11882 6100 11888 6112
rect 11843 6072 11888 6100
rect 11701 6063 11759 6069
rect 11882 6060 11888 6072
rect 11940 6060 11946 6112
rect 12342 6060 12348 6112
rect 12400 6100 12406 6112
rect 12437 6103 12495 6109
rect 12437 6100 12449 6103
rect 12400 6072 12449 6100
rect 12400 6060 12406 6072
rect 12437 6069 12449 6072
rect 12483 6069 12495 6103
rect 13170 6100 13176 6112
rect 13131 6072 13176 6100
rect 12437 6063 12495 6069
rect 13170 6060 13176 6072
rect 13228 6060 13234 6112
rect 13372 6100 13400 6208
rect 14642 6196 14648 6248
rect 14700 6236 14706 6248
rect 15396 6245 15424 6280
rect 15470 6264 15476 6280
rect 15528 6304 15534 6316
rect 17037 6307 17095 6313
rect 15528 6276 16252 6304
rect 15528 6264 15534 6276
rect 16224 6245 16252 6276
rect 17037 6273 17049 6307
rect 17083 6304 17095 6307
rect 17497 6307 17555 6313
rect 17497 6304 17509 6307
rect 17083 6276 17509 6304
rect 17083 6273 17095 6276
rect 17037 6267 17095 6273
rect 17497 6273 17509 6276
rect 17543 6273 17555 6307
rect 18046 6304 18052 6316
rect 18007 6276 18052 6304
rect 17497 6267 17555 6273
rect 18046 6264 18052 6276
rect 18104 6264 18110 6316
rect 21269 6307 21327 6313
rect 21269 6273 21281 6307
rect 21315 6304 21327 6307
rect 21542 6304 21548 6316
rect 21315 6276 21548 6304
rect 21315 6273 21327 6276
rect 21269 6267 21327 6273
rect 21542 6264 21548 6276
rect 21600 6264 21606 6316
rect 15289 6239 15347 6245
rect 15289 6236 15301 6239
rect 14700 6208 15301 6236
rect 14700 6196 14706 6208
rect 15289 6205 15301 6208
rect 15335 6205 15347 6239
rect 15289 6199 15347 6205
rect 15381 6239 15439 6245
rect 15381 6205 15393 6239
rect 15427 6205 15439 6239
rect 15381 6199 15439 6205
rect 16209 6239 16267 6245
rect 16209 6205 16221 6239
rect 16255 6205 16267 6239
rect 16209 6199 16267 6205
rect 17218 6196 17224 6248
rect 17276 6236 17282 6248
rect 17276 6208 17321 6236
rect 17276 6196 17282 6208
rect 18230 6168 18236 6180
rect 14568 6140 18236 6168
rect 14568 6100 14596 6140
rect 18230 6128 18236 6140
rect 18288 6128 18294 6180
rect 14734 6100 14740 6112
rect 13372 6072 14596 6100
rect 14695 6072 14740 6100
rect 14734 6060 14740 6072
rect 14792 6060 14798 6112
rect 14826 6060 14832 6112
rect 14884 6100 14890 6112
rect 15654 6100 15660 6112
rect 14884 6072 14929 6100
rect 15615 6072 15660 6100
rect 14884 6060 14890 6072
rect 15654 6060 15660 6072
rect 15712 6060 15718 6112
rect 16669 6103 16727 6109
rect 16669 6069 16681 6103
rect 16715 6100 16727 6103
rect 16942 6100 16948 6112
rect 16715 6072 16948 6100
rect 16715 6069 16727 6072
rect 16669 6063 16727 6069
rect 16942 6060 16948 6072
rect 17000 6060 17006 6112
rect 18690 6100 18696 6112
rect 18651 6072 18696 6100
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 1857 5899 1915 5905
rect 1857 5865 1869 5899
rect 1903 5896 1915 5899
rect 1946 5896 1952 5908
rect 1903 5868 1952 5896
rect 1903 5865 1915 5868
rect 1857 5859 1915 5865
rect 1946 5856 1952 5868
rect 2004 5856 2010 5908
rect 2590 5856 2596 5908
rect 2648 5896 2654 5908
rect 3973 5899 4031 5905
rect 2648 5868 3280 5896
rect 2648 5856 2654 5868
rect 1673 5831 1731 5837
rect 1673 5797 1685 5831
rect 1719 5828 1731 5831
rect 2222 5828 2228 5840
rect 1719 5800 2228 5828
rect 1719 5797 1731 5800
rect 1673 5791 1731 5797
rect 2222 5788 2228 5800
rect 2280 5788 2286 5840
rect 3252 5828 3280 5868
rect 3973 5865 3985 5899
rect 4019 5896 4031 5899
rect 4062 5896 4068 5908
rect 4019 5868 4068 5896
rect 4019 5865 4031 5868
rect 3973 5859 4031 5865
rect 4062 5856 4068 5868
rect 4120 5856 4126 5908
rect 4430 5896 4436 5908
rect 4391 5868 4436 5896
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 4540 5868 5100 5896
rect 3510 5828 3516 5840
rect 3252 5800 3516 5828
rect 3252 5769 3280 5800
rect 3510 5788 3516 5800
rect 3568 5788 3574 5840
rect 3237 5763 3295 5769
rect 3237 5729 3249 5763
rect 3283 5729 3295 5763
rect 3602 5760 3608 5772
rect 3237 5723 3295 5729
rect 3344 5732 3608 5760
rect 3344 5701 3372 5732
rect 3602 5720 3608 5732
rect 3660 5720 3666 5772
rect 4540 5760 4568 5868
rect 5072 5828 5100 5868
rect 5442 5856 5448 5908
rect 5500 5896 5506 5908
rect 5902 5896 5908 5908
rect 5500 5868 5908 5896
rect 5500 5856 5506 5868
rect 5902 5856 5908 5868
rect 5960 5896 5966 5908
rect 6914 5896 6920 5908
rect 5960 5868 6920 5896
rect 5960 5856 5966 5868
rect 6914 5856 6920 5868
rect 6972 5896 6978 5908
rect 7101 5899 7159 5905
rect 7101 5896 7113 5899
rect 6972 5868 7113 5896
rect 6972 5856 6978 5868
rect 7101 5865 7113 5868
rect 7147 5865 7159 5899
rect 7101 5859 7159 5865
rect 7282 5856 7288 5908
rect 7340 5896 7346 5908
rect 12253 5899 12311 5905
rect 12253 5896 12265 5899
rect 7340 5868 8524 5896
rect 7340 5856 7346 5868
rect 7466 5828 7472 5840
rect 3804 5732 4568 5760
rect 4632 5800 5028 5828
rect 5072 5800 7472 5828
rect 3804 5701 3832 5732
rect 2970 5695 3028 5701
rect 2970 5661 2982 5695
rect 3016 5692 3028 5695
rect 3329 5695 3387 5701
rect 3016 5664 3096 5692
rect 3016 5661 3028 5664
rect 2970 5655 3028 5661
rect 3068 5636 3096 5664
rect 3329 5661 3341 5695
rect 3375 5661 3387 5695
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 3329 5655 3387 5661
rect 3436 5664 3801 5692
rect 1486 5624 1492 5636
rect 1447 5596 1492 5624
rect 1486 5584 1492 5596
rect 1544 5584 1550 5636
rect 3050 5584 3056 5636
rect 3108 5584 3114 5636
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 3436 5556 3464 5664
rect 3789 5661 3801 5664
rect 3835 5661 3847 5695
rect 3789 5655 3847 5661
rect 4065 5695 4123 5701
rect 4065 5661 4077 5695
rect 4111 5692 4123 5695
rect 4246 5692 4252 5704
rect 4111 5664 4252 5692
rect 4111 5661 4123 5664
rect 4065 5655 4123 5661
rect 4246 5652 4252 5664
rect 4304 5652 4310 5704
rect 4430 5652 4436 5704
rect 4488 5692 4494 5704
rect 4632 5692 4660 5800
rect 4890 5760 4896 5772
rect 4851 5732 4896 5760
rect 4890 5720 4896 5732
rect 4948 5720 4954 5772
rect 5000 5769 5028 5800
rect 7466 5788 7472 5800
rect 7524 5788 7530 5840
rect 8496 5769 8524 5868
rect 8956 5868 12265 5896
rect 8956 5840 8984 5868
rect 12253 5865 12265 5868
rect 12299 5865 12311 5899
rect 12894 5896 12900 5908
rect 12253 5859 12311 5865
rect 12406 5868 12900 5896
rect 8573 5831 8631 5837
rect 8573 5797 8585 5831
rect 8619 5797 8631 5831
rect 8573 5791 8631 5797
rect 4985 5763 5043 5769
rect 4985 5729 4997 5763
rect 5031 5729 5043 5763
rect 4985 5723 5043 5729
rect 8481 5763 8539 5769
rect 8481 5729 8493 5763
rect 8527 5729 8539 5763
rect 8588 5760 8616 5791
rect 8938 5788 8944 5840
rect 8996 5788 9002 5840
rect 11054 5788 11060 5840
rect 11112 5828 11118 5840
rect 11606 5828 11612 5840
rect 11112 5800 11612 5828
rect 11112 5788 11118 5800
rect 11606 5788 11612 5800
rect 11664 5828 11670 5840
rect 12406 5828 12434 5868
rect 12894 5856 12900 5868
rect 12952 5856 12958 5908
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 13320 5868 19288 5896
rect 13320 5856 13326 5868
rect 14826 5828 14832 5840
rect 11664 5800 12434 5828
rect 14568 5800 14832 5828
rect 11664 5788 11670 5800
rect 9306 5760 9312 5772
rect 8588 5732 9312 5760
rect 8481 5723 8539 5729
rect 9306 5720 9312 5732
rect 9364 5720 9370 5772
rect 10502 5720 10508 5772
rect 10560 5760 10566 5772
rect 11330 5760 11336 5772
rect 10560 5732 11336 5760
rect 10560 5720 10566 5732
rect 11330 5720 11336 5732
rect 11388 5720 11394 5772
rect 12161 5763 12219 5769
rect 12161 5729 12173 5763
rect 12207 5760 12219 5763
rect 12526 5760 12532 5772
rect 12207 5732 12532 5760
rect 12207 5729 12219 5732
rect 12161 5723 12219 5729
rect 4488 5664 4660 5692
rect 4488 5652 4494 5664
rect 4798 5652 4804 5704
rect 4856 5692 4862 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 4856 5664 5457 5692
rect 4856 5652 4862 5664
rect 5445 5661 5457 5664
rect 5491 5692 5503 5695
rect 5994 5692 6000 5704
rect 5491 5664 6000 5692
rect 5491 5661 5503 5664
rect 5445 5655 5503 5661
rect 5994 5652 6000 5664
rect 6052 5652 6058 5704
rect 7006 5692 7012 5704
rect 6919 5664 7012 5692
rect 7006 5652 7012 5664
rect 7064 5692 7070 5704
rect 8754 5692 8760 5704
rect 7064 5664 8432 5692
rect 8715 5664 8760 5692
rect 7064 5652 7070 5664
rect 6822 5624 6828 5636
rect 3528 5596 6828 5624
rect 3528 5565 3556 5596
rect 6822 5584 6828 5596
rect 6880 5584 6886 5636
rect 8202 5624 8208 5636
rect 8260 5633 8266 5636
rect 8172 5596 8208 5624
rect 8202 5584 8208 5596
rect 8260 5587 8272 5633
rect 8404 5624 8432 5664
rect 8754 5652 8760 5664
rect 8812 5652 8818 5704
rect 9674 5652 9680 5704
rect 9732 5692 9738 5704
rect 10321 5695 10379 5701
rect 10321 5692 10333 5695
rect 9732 5664 10333 5692
rect 9732 5652 9738 5664
rect 9968 5636 9996 5664
rect 10321 5661 10333 5664
rect 10367 5692 10379 5695
rect 12176 5692 12204 5723
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 14568 5769 14596 5800
rect 14826 5788 14832 5800
rect 14884 5788 14890 5840
rect 15562 5828 15568 5840
rect 15523 5800 15568 5828
rect 15562 5788 15568 5800
rect 15620 5788 15626 5840
rect 17037 5831 17095 5837
rect 17037 5797 17049 5831
rect 17083 5828 17095 5831
rect 17126 5828 17132 5840
rect 17083 5800 17132 5828
rect 17083 5797 17095 5800
rect 17037 5791 17095 5797
rect 17126 5788 17132 5800
rect 17184 5788 17190 5840
rect 14553 5763 14611 5769
rect 14553 5729 14565 5763
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 14737 5763 14795 5769
rect 14737 5729 14749 5763
rect 14783 5729 14795 5763
rect 14737 5723 14795 5729
rect 12796 5695 12854 5701
rect 12796 5692 12808 5695
rect 10367 5664 12204 5692
rect 12728 5664 12808 5692
rect 10367 5661 10379 5664
rect 10321 5655 10379 5661
rect 12728 5636 12756 5664
rect 12796 5661 12808 5664
rect 12842 5661 12854 5695
rect 14458 5692 14464 5704
rect 14419 5664 14464 5692
rect 12796 5655 12854 5661
rect 14458 5652 14464 5664
rect 14516 5652 14522 5704
rect 8404 5596 9260 5624
rect 8260 5584 8266 5587
rect 2924 5528 3464 5556
rect 3513 5559 3571 5565
rect 2924 5516 2930 5528
rect 3513 5525 3525 5559
rect 3559 5525 3571 5559
rect 3513 5519 3571 5525
rect 3602 5516 3608 5568
rect 3660 5556 3666 5568
rect 3970 5556 3976 5568
rect 3660 5528 3976 5556
rect 3660 5516 3666 5528
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 4249 5559 4307 5565
rect 4249 5525 4261 5559
rect 4295 5556 4307 5559
rect 4338 5556 4344 5568
rect 4295 5528 4344 5556
rect 4295 5525 4307 5528
rect 4249 5519 4307 5525
rect 4338 5516 4344 5528
rect 4396 5516 4402 5568
rect 4801 5559 4859 5565
rect 4801 5525 4813 5559
rect 4847 5556 4859 5559
rect 5258 5556 5264 5568
rect 4847 5528 5264 5556
rect 4847 5525 4859 5528
rect 4801 5519 4859 5525
rect 5258 5516 5264 5528
rect 5316 5516 5322 5568
rect 5718 5516 5724 5568
rect 5776 5556 5782 5568
rect 7742 5556 7748 5568
rect 5776 5528 7748 5556
rect 5776 5516 5782 5528
rect 7742 5516 7748 5528
rect 7800 5516 7806 5568
rect 8478 5516 8484 5568
rect 8536 5556 8542 5568
rect 8754 5556 8760 5568
rect 8536 5528 8760 5556
rect 8536 5516 8542 5528
rect 8754 5516 8760 5528
rect 8812 5516 8818 5568
rect 8941 5559 8999 5565
rect 8941 5525 8953 5559
rect 8987 5556 8999 5559
rect 9122 5556 9128 5568
rect 8987 5528 9128 5556
rect 8987 5525 8999 5528
rect 8941 5519 8999 5525
rect 9122 5516 9128 5528
rect 9180 5516 9186 5568
rect 9232 5556 9260 5596
rect 9950 5584 9956 5636
rect 10008 5584 10014 5636
rect 10076 5627 10134 5633
rect 10076 5593 10088 5627
rect 10122 5624 10134 5627
rect 10226 5624 10232 5636
rect 10122 5596 10232 5624
rect 10122 5593 10134 5596
rect 10076 5587 10134 5593
rect 10226 5584 10232 5596
rect 10284 5584 10290 5636
rect 10410 5624 10416 5636
rect 10371 5596 10416 5624
rect 10410 5584 10416 5596
rect 10468 5584 10474 5636
rect 12710 5584 12716 5636
rect 12768 5584 12774 5636
rect 12894 5584 12900 5636
rect 12952 5624 12958 5636
rect 13262 5624 13268 5636
rect 12952 5596 13268 5624
rect 12952 5584 12958 5596
rect 13262 5584 13268 5596
rect 13320 5584 13326 5636
rect 14752 5624 14780 5723
rect 15657 5695 15715 5701
rect 15657 5661 15669 5695
rect 15703 5692 15715 5695
rect 15746 5692 15752 5704
rect 15703 5664 15752 5692
rect 15703 5661 15715 5664
rect 15657 5655 15715 5661
rect 15746 5652 15752 5664
rect 15804 5692 15810 5704
rect 17034 5692 17040 5704
rect 15804 5664 17040 5692
rect 15804 5652 15810 5664
rect 17034 5652 17040 5664
rect 17092 5692 17098 5704
rect 19260 5701 19288 5868
rect 18509 5695 18567 5701
rect 18509 5692 18521 5695
rect 17092 5664 18521 5692
rect 17092 5652 17098 5664
rect 18509 5661 18521 5664
rect 18555 5661 18567 5695
rect 18509 5655 18567 5661
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5661 19303 5695
rect 19245 5655 19303 5661
rect 13924 5596 14780 5624
rect 15924 5627 15982 5633
rect 10428 5556 10456 5584
rect 9232 5528 10456 5556
rect 11146 5516 11152 5568
rect 11204 5556 11210 5568
rect 11882 5556 11888 5568
rect 11204 5528 11888 5556
rect 11204 5516 11210 5528
rect 11882 5516 11888 5528
rect 11940 5516 11946 5568
rect 13078 5516 13084 5568
rect 13136 5556 13142 5568
rect 13630 5556 13636 5568
rect 13136 5528 13636 5556
rect 13136 5516 13142 5528
rect 13630 5516 13636 5528
rect 13688 5556 13694 5568
rect 13924 5565 13952 5596
rect 15924 5593 15936 5627
rect 15970 5624 15982 5627
rect 16850 5624 16856 5636
rect 15970 5596 16856 5624
rect 15970 5593 15982 5596
rect 15924 5587 15982 5593
rect 16850 5584 16856 5596
rect 16908 5624 16914 5636
rect 17862 5624 17868 5636
rect 16908 5596 17868 5624
rect 16908 5584 16914 5596
rect 17862 5584 17868 5596
rect 17920 5584 17926 5636
rect 18264 5627 18322 5633
rect 18264 5593 18276 5627
rect 18310 5624 18322 5627
rect 18690 5624 18696 5636
rect 18310 5596 18696 5624
rect 18310 5593 18322 5596
rect 18264 5587 18322 5593
rect 18690 5584 18696 5596
rect 18748 5584 18754 5636
rect 13909 5559 13967 5565
rect 13909 5556 13921 5559
rect 13688 5528 13921 5556
rect 13688 5516 13694 5528
rect 13909 5525 13921 5528
rect 13955 5525 13967 5559
rect 14090 5556 14096 5568
rect 14051 5528 14096 5556
rect 13909 5519 13967 5525
rect 14090 5516 14096 5528
rect 14148 5516 14154 5568
rect 14642 5516 14648 5568
rect 14700 5556 14706 5568
rect 14921 5559 14979 5565
rect 14921 5556 14933 5559
rect 14700 5528 14933 5556
rect 14700 5516 14706 5528
rect 14921 5525 14933 5528
rect 14967 5525 14979 5559
rect 14921 5519 14979 5525
rect 17129 5559 17187 5565
rect 17129 5525 17141 5559
rect 17175 5556 17187 5559
rect 17218 5556 17224 5568
rect 17175 5528 17224 5556
rect 17175 5525 17187 5528
rect 17129 5519 17187 5525
rect 17218 5516 17224 5528
rect 17276 5516 17282 5568
rect 19429 5559 19487 5565
rect 19429 5525 19441 5559
rect 19475 5556 19487 5559
rect 19978 5556 19984 5568
rect 19475 5528 19984 5556
rect 19475 5525 19487 5528
rect 19429 5519 19487 5525
rect 19978 5516 19984 5528
rect 20036 5516 20042 5568
rect 1104 5466 21896 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21896 5466
rect 1104 5392 21896 5414
rect 1578 5352 1584 5364
rect 1539 5324 1584 5352
rect 1578 5312 1584 5324
rect 1636 5352 1642 5364
rect 2682 5352 2688 5364
rect 1636 5324 2688 5352
rect 1636 5312 1642 5324
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 3326 5312 3332 5364
rect 3384 5352 3390 5364
rect 3973 5355 4031 5361
rect 3973 5352 3985 5355
rect 3384 5324 3985 5352
rect 3384 5312 3390 5324
rect 3973 5321 3985 5324
rect 4019 5321 4031 5355
rect 3973 5315 4031 5321
rect 4341 5355 4399 5361
rect 4341 5321 4353 5355
rect 4387 5352 4399 5355
rect 5534 5352 5540 5364
rect 4387 5324 5540 5352
rect 4387 5321 4399 5324
rect 4341 5315 4399 5321
rect 5534 5312 5540 5324
rect 5592 5312 5598 5364
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 6181 5355 6239 5361
rect 6181 5352 6193 5355
rect 5684 5324 6193 5352
rect 5684 5312 5690 5324
rect 6181 5321 6193 5324
rect 6227 5321 6239 5355
rect 7006 5352 7012 5364
rect 6181 5315 6239 5321
rect 6380 5324 7012 5352
rect 2130 5244 2136 5296
rect 2188 5293 2194 5296
rect 2188 5287 2252 5293
rect 2188 5253 2206 5287
rect 2240 5253 2252 5287
rect 2188 5247 2252 5253
rect 2746 5256 3740 5284
rect 2188 5244 2194 5247
rect 1489 5219 1547 5225
rect 1489 5185 1501 5219
rect 1535 5185 1547 5219
rect 1489 5179 1547 5185
rect 1504 5148 1532 5179
rect 2038 5176 2044 5228
rect 2096 5216 2102 5228
rect 2590 5216 2596 5228
rect 2096 5188 2596 5216
rect 2096 5176 2102 5188
rect 2590 5176 2596 5188
rect 2648 5216 2654 5228
rect 2746 5216 2774 5256
rect 2648 5188 2774 5216
rect 2648 5176 2654 5188
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 3712 5225 3740 5256
rect 3786 5244 3792 5296
rect 3844 5284 3850 5296
rect 6380 5284 6408 5324
rect 7006 5312 7012 5324
rect 7064 5312 7070 5364
rect 7101 5355 7159 5361
rect 7101 5321 7113 5355
rect 7147 5352 7159 5355
rect 7190 5352 7196 5364
rect 7147 5324 7196 5352
rect 7147 5321 7159 5324
rect 7101 5315 7159 5321
rect 7190 5312 7196 5324
rect 7248 5312 7254 5364
rect 7561 5355 7619 5361
rect 7561 5321 7573 5355
rect 7607 5352 7619 5355
rect 7926 5352 7932 5364
rect 7607 5324 7932 5352
rect 7607 5321 7619 5324
rect 7561 5315 7619 5321
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 8021 5355 8079 5361
rect 8021 5321 8033 5355
rect 8067 5352 8079 5355
rect 8110 5352 8116 5364
rect 8067 5324 8116 5352
rect 8067 5321 8079 5324
rect 8021 5315 8079 5321
rect 8110 5312 8116 5324
rect 8168 5312 8174 5364
rect 8570 5352 8576 5364
rect 8531 5324 8576 5352
rect 8570 5312 8576 5324
rect 8628 5312 8634 5364
rect 9766 5312 9772 5364
rect 9824 5352 9830 5364
rect 10045 5355 10103 5361
rect 10045 5352 10057 5355
rect 9824 5324 10057 5352
rect 9824 5312 9830 5324
rect 10045 5321 10057 5324
rect 10091 5321 10103 5355
rect 10410 5352 10416 5364
rect 10371 5324 10416 5352
rect 10045 5315 10103 5321
rect 10410 5312 10416 5324
rect 10468 5352 10474 5364
rect 11146 5352 11152 5364
rect 10468 5324 11152 5352
rect 10468 5312 10474 5324
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 11238 5312 11244 5364
rect 11296 5352 11302 5364
rect 11333 5355 11391 5361
rect 11333 5352 11345 5355
rect 11296 5324 11345 5352
rect 11296 5312 11302 5324
rect 11333 5321 11345 5324
rect 11379 5321 11391 5355
rect 11333 5315 11391 5321
rect 11793 5355 11851 5361
rect 11793 5321 11805 5355
rect 11839 5352 11851 5355
rect 11882 5352 11888 5364
rect 11839 5324 11888 5352
rect 11839 5321 11851 5324
rect 11793 5315 11851 5321
rect 11882 5312 11888 5324
rect 11940 5352 11946 5364
rect 12621 5355 12679 5361
rect 12621 5352 12633 5355
rect 11940 5324 12633 5352
rect 11940 5312 11946 5324
rect 12621 5321 12633 5324
rect 12667 5321 12679 5355
rect 14090 5352 14096 5364
rect 14051 5324 14096 5352
rect 12621 5315 12679 5321
rect 3844 5256 6408 5284
rect 3844 5244 3850 5256
rect 7282 5244 7288 5296
rect 7340 5284 7346 5296
rect 8294 5284 8300 5296
rect 7340 5256 8300 5284
rect 7340 5244 7346 5256
rect 8294 5244 8300 5256
rect 8352 5244 8358 5296
rect 8662 5244 8668 5296
rect 8720 5284 8726 5296
rect 9686 5287 9744 5293
rect 9686 5284 9698 5287
rect 8720 5256 9698 5284
rect 8720 5244 8726 5256
rect 9686 5253 9698 5256
rect 9732 5253 9744 5287
rect 9686 5247 9744 5253
rect 11054 5244 11060 5296
rect 11112 5284 11118 5296
rect 12636 5284 12664 5315
rect 14090 5312 14096 5324
rect 14148 5312 14154 5364
rect 15194 5352 15200 5364
rect 15155 5324 15200 5352
rect 15194 5312 15200 5324
rect 15252 5312 15258 5364
rect 16025 5355 16083 5361
rect 16025 5321 16037 5355
rect 16071 5352 16083 5355
rect 18141 5355 18199 5361
rect 18141 5352 18153 5355
rect 16071 5324 18153 5352
rect 16071 5321 16083 5324
rect 16025 5315 16083 5321
rect 18141 5321 18153 5324
rect 18187 5321 18199 5355
rect 18141 5315 18199 5321
rect 15286 5284 15292 5296
rect 11112 5256 12572 5284
rect 12636 5256 15292 5284
rect 11112 5244 11118 5256
rect 3421 5219 3479 5225
rect 3421 5216 3433 5219
rect 3384 5188 3433 5216
rect 3384 5176 3390 5188
rect 3421 5185 3433 5188
rect 3467 5185 3479 5219
rect 3421 5179 3479 5185
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5185 3755 5219
rect 4430 5216 4436 5228
rect 4391 5188 4436 5216
rect 3697 5179 3755 5185
rect 4430 5176 4436 5188
rect 4488 5176 4494 5228
rect 4798 5216 4804 5228
rect 4759 5188 4804 5216
rect 4798 5176 4804 5188
rect 4856 5176 4862 5228
rect 4890 5176 4896 5228
rect 4948 5176 4954 5228
rect 5068 5219 5126 5225
rect 5068 5185 5080 5219
rect 5114 5216 5126 5219
rect 5350 5216 5356 5228
rect 5114 5188 5356 5216
rect 5114 5185 5126 5188
rect 5068 5179 5126 5185
rect 5350 5176 5356 5188
rect 5408 5176 5414 5228
rect 6454 5176 6460 5228
rect 6512 5216 6518 5228
rect 6641 5219 6699 5225
rect 6641 5216 6653 5219
rect 6512 5188 6653 5216
rect 6512 5176 6518 5188
rect 6641 5185 6653 5188
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 6730 5176 6736 5228
rect 6788 5216 6794 5228
rect 7650 5216 7656 5228
rect 6788 5188 6833 5216
rect 7611 5188 7656 5216
rect 6788 5176 6794 5188
rect 7650 5176 7656 5188
rect 7708 5176 7714 5228
rect 8113 5219 8171 5225
rect 8113 5185 8125 5219
rect 8159 5185 8171 5219
rect 8113 5179 8171 5185
rect 1854 5148 1860 5160
rect 1504 5120 1860 5148
rect 1854 5108 1860 5120
rect 1912 5108 1918 5160
rect 1946 5108 1952 5160
rect 2004 5148 2010 5160
rect 3970 5148 3976 5160
rect 2004 5120 2049 5148
rect 3620 5120 3976 5148
rect 2004 5108 2010 5120
rect 3050 5040 3056 5092
rect 3108 5080 3114 5092
rect 3620 5089 3648 5120
rect 3970 5108 3976 5120
rect 4028 5108 4034 5160
rect 4617 5151 4675 5157
rect 4617 5117 4629 5151
rect 4663 5148 4675 5151
rect 4908 5148 4936 5176
rect 4663 5120 4936 5148
rect 4663 5117 4675 5120
rect 4617 5111 4675 5117
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 6549 5151 6607 5157
rect 6549 5148 6561 5151
rect 5960 5120 6561 5148
rect 5960 5108 5966 5120
rect 6549 5117 6561 5120
rect 6595 5117 6607 5151
rect 6549 5111 6607 5117
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 7377 5151 7435 5157
rect 7377 5148 7389 5151
rect 6972 5120 7389 5148
rect 6972 5108 6978 5120
rect 7377 5117 7389 5120
rect 7423 5117 7435 5151
rect 7377 5111 7435 5117
rect 3329 5083 3387 5089
rect 3329 5080 3341 5083
rect 3108 5052 3341 5080
rect 3108 5040 3114 5052
rect 3329 5049 3341 5052
rect 3375 5049 3387 5083
rect 3329 5043 3387 5049
rect 3605 5083 3663 5089
rect 3605 5049 3617 5083
rect 3651 5049 3663 5083
rect 3605 5043 3663 5049
rect 1762 5012 1768 5024
rect 1723 4984 1768 5012
rect 1762 4972 1768 4984
rect 1820 5012 1826 5024
rect 3234 5012 3240 5024
rect 1820 4984 3240 5012
rect 1820 4972 1826 4984
rect 3234 4972 3240 4984
rect 3292 4972 3298 5024
rect 3344 5012 3372 5043
rect 3786 5040 3792 5092
rect 3844 5080 3850 5092
rect 3881 5083 3939 5089
rect 3881 5080 3893 5083
rect 3844 5052 3893 5080
rect 3844 5040 3850 5052
rect 3881 5049 3893 5052
rect 3927 5049 3939 5083
rect 4338 5080 4344 5092
rect 3881 5043 3939 5049
rect 3988 5052 4344 5080
rect 3988 5012 4016 5052
rect 4338 5040 4344 5052
rect 4396 5040 4402 5092
rect 6822 5040 6828 5092
rect 6880 5080 6886 5092
rect 8128 5080 8156 5179
rect 8478 5176 8484 5228
rect 8536 5216 8542 5228
rect 9398 5216 9404 5228
rect 8536 5188 9404 5216
rect 8536 5176 8542 5188
rect 9398 5176 9404 5188
rect 9456 5176 9462 5228
rect 9950 5216 9956 5228
rect 9911 5188 9956 5216
rect 9950 5176 9956 5188
rect 10008 5176 10014 5228
rect 10042 5176 10048 5228
rect 10100 5216 10106 5228
rect 10229 5219 10287 5225
rect 10229 5216 10241 5219
rect 10100 5188 10241 5216
rect 10100 5176 10106 5188
rect 10229 5185 10241 5188
rect 10275 5185 10287 5219
rect 10229 5179 10287 5185
rect 10410 5176 10416 5228
rect 10468 5216 10474 5228
rect 10965 5219 11023 5225
rect 10965 5216 10977 5219
rect 10468 5188 10977 5216
rect 10468 5176 10474 5188
rect 10965 5185 10977 5188
rect 11011 5185 11023 5219
rect 10965 5179 11023 5185
rect 11146 5176 11152 5228
rect 11204 5216 11210 5228
rect 11885 5219 11943 5225
rect 11885 5216 11897 5219
rect 11204 5188 11897 5216
rect 11204 5176 11210 5188
rect 11885 5185 11897 5188
rect 11931 5185 11943 5219
rect 11885 5179 11943 5185
rect 8294 5108 8300 5160
rect 8352 5148 8358 5160
rect 8389 5151 8447 5157
rect 8389 5148 8401 5151
rect 8352 5120 8401 5148
rect 8352 5108 8358 5120
rect 8389 5117 8401 5120
rect 8435 5117 8447 5151
rect 10686 5148 10692 5160
rect 10647 5120 10692 5148
rect 8389 5111 8447 5117
rect 6880 5052 8156 5080
rect 6880 5040 6886 5052
rect 3344 4984 4016 5012
rect 4246 4972 4252 5024
rect 4304 5012 4310 5024
rect 6730 5012 6736 5024
rect 4304 4984 6736 5012
rect 4304 4972 4310 4984
rect 6730 4972 6736 4984
rect 6788 5012 6794 5024
rect 7466 5012 7472 5024
rect 6788 4984 7472 5012
rect 6788 4972 6794 4984
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 8294 5012 8300 5024
rect 8255 4984 8300 5012
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 8404 5012 8432 5111
rect 10686 5108 10692 5120
rect 10744 5108 10750 5160
rect 10873 5151 10931 5157
rect 10873 5117 10885 5151
rect 10919 5148 10931 5151
rect 11238 5148 11244 5160
rect 10919 5120 11244 5148
rect 10919 5117 10931 5120
rect 10873 5111 10931 5117
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 11514 5108 11520 5160
rect 11572 5148 11578 5160
rect 11609 5151 11667 5157
rect 11609 5148 11621 5151
rect 11572 5120 11621 5148
rect 11572 5108 11578 5120
rect 11609 5117 11621 5120
rect 11655 5117 11667 5151
rect 11900 5148 11928 5179
rect 12250 5176 12256 5228
rect 12308 5216 12314 5228
rect 12345 5219 12403 5225
rect 12345 5216 12357 5219
rect 12308 5188 12357 5216
rect 12308 5176 12314 5188
rect 12345 5185 12357 5188
rect 12391 5185 12403 5219
rect 12544 5216 12572 5256
rect 15286 5244 15292 5256
rect 15344 5244 15350 5296
rect 17034 5284 17040 5296
rect 16684 5256 17040 5284
rect 12618 5216 12624 5228
rect 12544 5188 12624 5216
rect 12345 5179 12403 5185
rect 12618 5176 12624 5188
rect 12676 5176 12682 5228
rect 13262 5216 13268 5228
rect 13223 5188 13268 5216
rect 13262 5176 13268 5188
rect 13320 5176 13326 5228
rect 14734 5216 14740 5228
rect 13924 5188 14740 5216
rect 12802 5148 12808 5160
rect 11900 5120 12808 5148
rect 11609 5111 11667 5117
rect 12802 5108 12808 5120
rect 12860 5108 12866 5160
rect 13078 5148 13084 5160
rect 13039 5120 13084 5148
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13173 5151 13231 5157
rect 13173 5117 13185 5151
rect 13219 5148 13231 5151
rect 13722 5148 13728 5160
rect 13219 5120 13728 5148
rect 13219 5117 13231 5120
rect 13173 5111 13231 5117
rect 13722 5108 13728 5120
rect 13780 5108 13786 5160
rect 13924 5157 13952 5188
rect 14734 5176 14740 5188
rect 14792 5176 14798 5228
rect 15194 5176 15200 5228
rect 15252 5216 15258 5228
rect 16684 5225 16712 5256
rect 17034 5244 17040 5256
rect 17092 5244 17098 5296
rect 17126 5244 17132 5296
rect 17184 5244 17190 5296
rect 17954 5244 17960 5296
rect 18012 5284 18018 5296
rect 18509 5287 18567 5293
rect 18509 5284 18521 5287
rect 18012 5256 18521 5284
rect 18012 5244 18018 5256
rect 18509 5253 18521 5256
rect 18555 5253 18567 5287
rect 18509 5247 18567 5253
rect 16117 5219 16175 5225
rect 16117 5216 16129 5219
rect 15252 5188 16129 5216
rect 15252 5176 15258 5188
rect 16117 5185 16129 5188
rect 16163 5185 16175 5219
rect 16117 5179 16175 5185
rect 16669 5219 16727 5225
rect 16669 5185 16681 5219
rect 16715 5185 16727 5219
rect 16925 5219 16983 5225
rect 16925 5216 16937 5219
rect 16669 5179 16727 5185
rect 16776 5188 16937 5216
rect 13909 5151 13967 5157
rect 13909 5117 13921 5151
rect 13955 5117 13967 5151
rect 13909 5111 13967 5117
rect 14001 5151 14059 5157
rect 14001 5117 14013 5151
rect 14047 5117 14059 5151
rect 14553 5151 14611 5157
rect 14553 5148 14565 5151
rect 14001 5111 14059 5117
rect 14108 5120 14565 5148
rect 12529 5083 12587 5089
rect 9968 5052 12480 5080
rect 9968 5024 9996 5052
rect 9950 5012 9956 5024
rect 8404 4984 9956 5012
rect 9950 4972 9956 4984
rect 10008 4972 10014 5024
rect 10226 4972 10232 5024
rect 10284 5012 10290 5024
rect 10778 5012 10784 5024
rect 10284 4984 10784 5012
rect 10284 4972 10290 4984
rect 10778 4972 10784 4984
rect 10836 4972 10842 5024
rect 10870 4972 10876 5024
rect 10928 5012 10934 5024
rect 11514 5012 11520 5024
rect 10928 4984 11520 5012
rect 10928 4972 10934 4984
rect 11514 4972 11520 4984
rect 11572 4972 11578 5024
rect 12253 5015 12311 5021
rect 12253 4981 12265 5015
rect 12299 5012 12311 5015
rect 12342 5012 12348 5024
rect 12299 4984 12348 5012
rect 12299 4981 12311 4984
rect 12253 4975 12311 4981
rect 12342 4972 12348 4984
rect 12400 4972 12406 5024
rect 12452 5012 12480 5052
rect 12529 5049 12541 5083
rect 12575 5080 12587 5083
rect 12894 5080 12900 5092
rect 12575 5052 12900 5080
rect 12575 5049 12587 5052
rect 12529 5043 12587 5049
rect 12894 5040 12900 5052
rect 12952 5040 12958 5092
rect 13633 5083 13691 5089
rect 13633 5049 13645 5083
rect 13679 5080 13691 5083
rect 14016 5080 14044 5111
rect 13679 5052 14044 5080
rect 13679 5049 13691 5052
rect 13633 5043 13691 5049
rect 14108 5012 14136 5120
rect 14553 5117 14565 5120
rect 14599 5148 14611 5151
rect 15746 5148 15752 5160
rect 14599 5120 15752 5148
rect 14599 5117 14611 5120
rect 14553 5111 14611 5117
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 15933 5151 15991 5157
rect 15933 5117 15945 5151
rect 15979 5148 15991 5151
rect 16776 5148 16804 5188
rect 16925 5185 16937 5188
rect 16971 5216 16983 5219
rect 17144 5216 17172 5244
rect 16971 5188 17172 5216
rect 16971 5185 16983 5188
rect 16925 5179 16983 5185
rect 17862 5176 17868 5228
rect 17920 5216 17926 5228
rect 19978 5216 19984 5228
rect 17920 5188 18736 5216
rect 19939 5188 19984 5216
rect 17920 5176 17926 5188
rect 15979 5120 16804 5148
rect 15979 5117 15991 5120
rect 15933 5111 15991 5117
rect 17770 5108 17776 5160
rect 17828 5148 17834 5160
rect 18708 5157 18736 5188
rect 19978 5176 19984 5188
rect 20036 5176 20042 5228
rect 18601 5151 18659 5157
rect 18601 5148 18613 5151
rect 17828 5120 18613 5148
rect 17828 5108 17834 5120
rect 18601 5117 18613 5120
rect 18647 5117 18659 5151
rect 18601 5111 18659 5117
rect 18693 5151 18751 5157
rect 18693 5117 18705 5151
rect 18739 5117 18751 5151
rect 18693 5111 18751 5117
rect 14366 5040 14372 5092
rect 14424 5080 14430 5092
rect 14921 5083 14979 5089
rect 14921 5080 14933 5083
rect 14424 5052 14933 5080
rect 14424 5040 14430 5052
rect 14921 5049 14933 5052
rect 14967 5049 14979 5083
rect 14921 5043 14979 5049
rect 14458 5012 14464 5024
rect 12452 4984 14136 5012
rect 14419 4984 14464 5012
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 14826 5012 14832 5024
rect 14787 4984 14832 5012
rect 14826 4972 14832 4984
rect 14884 4972 14890 5024
rect 16485 5015 16543 5021
rect 16485 4981 16497 5015
rect 16531 5012 16543 5015
rect 16666 5012 16672 5024
rect 16531 4984 16672 5012
rect 16531 4981 16543 4984
rect 16485 4975 16543 4981
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 18046 5012 18052 5024
rect 18007 4984 18052 5012
rect 18046 4972 18052 4984
rect 18104 4972 18110 5024
rect 20165 5015 20223 5021
rect 20165 4981 20177 5015
rect 20211 5012 20223 5015
rect 20898 5012 20904 5024
rect 20211 4984 20904 5012
rect 20211 4981 20223 4984
rect 20165 4975 20223 4981
rect 20898 4972 20904 4984
rect 20956 4972 20962 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 1949 4811 2007 4817
rect 1949 4777 1961 4811
rect 1995 4808 2007 4811
rect 2038 4808 2044 4820
rect 1995 4780 2044 4808
rect 1995 4777 2007 4780
rect 1949 4771 2007 4777
rect 2038 4768 2044 4780
rect 2096 4768 2102 4820
rect 2314 4808 2320 4820
rect 2148 4780 2320 4808
rect 1673 4743 1731 4749
rect 1673 4709 1685 4743
rect 1719 4740 1731 4743
rect 2148 4740 2176 4780
rect 2314 4768 2320 4780
rect 2372 4768 2378 4820
rect 2777 4811 2835 4817
rect 2777 4777 2789 4811
rect 2823 4808 2835 4811
rect 2958 4808 2964 4820
rect 2823 4780 2964 4808
rect 2823 4777 2835 4780
rect 2777 4771 2835 4777
rect 2958 4768 2964 4780
rect 3016 4768 3022 4820
rect 3605 4811 3663 4817
rect 3605 4777 3617 4811
rect 3651 4808 3663 4811
rect 3878 4808 3884 4820
rect 3651 4780 3884 4808
rect 3651 4777 3663 4780
rect 3605 4771 3663 4777
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 4154 4768 4160 4820
rect 4212 4808 4218 4820
rect 4430 4808 4436 4820
rect 4212 4780 4436 4808
rect 4212 4768 4218 4780
rect 4430 4768 4436 4780
rect 4488 4768 4494 4820
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 5258 4808 5264 4820
rect 5040 4780 5264 4808
rect 5040 4768 5046 4780
rect 5258 4768 5264 4780
rect 5316 4768 5322 4820
rect 5810 4768 5816 4820
rect 5868 4808 5874 4820
rect 6822 4808 6828 4820
rect 5868 4780 6828 4808
rect 5868 4768 5874 4780
rect 6822 4768 6828 4780
rect 6880 4808 6886 4820
rect 7377 4811 7435 4817
rect 7377 4808 7389 4811
rect 6880 4780 7389 4808
rect 6880 4768 6886 4780
rect 7377 4777 7389 4780
rect 7423 4777 7435 4811
rect 7377 4771 7435 4777
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 7650 4808 7656 4820
rect 7607 4780 7656 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 8202 4768 8208 4820
rect 8260 4808 8266 4820
rect 9585 4811 9643 4817
rect 9585 4808 9597 4811
rect 8260 4780 9597 4808
rect 8260 4768 8266 4780
rect 9585 4777 9597 4780
rect 9631 4777 9643 4811
rect 9585 4771 9643 4777
rect 10686 4768 10692 4820
rect 10744 4808 10750 4820
rect 11422 4808 11428 4820
rect 10744 4780 11284 4808
rect 11383 4780 11428 4808
rect 10744 4768 10750 4780
rect 3050 4740 3056 4752
rect 1719 4712 2176 4740
rect 2240 4712 3056 4740
rect 1719 4709 1731 4712
rect 1673 4703 1731 4709
rect 2240 4681 2268 4712
rect 3050 4700 3056 4712
rect 3108 4700 3114 4752
rect 3142 4700 3148 4752
rect 3200 4740 3206 4752
rect 3789 4743 3847 4749
rect 3789 4740 3801 4743
rect 3200 4712 3801 4740
rect 3200 4700 3206 4712
rect 3789 4709 3801 4712
rect 3835 4709 3847 4743
rect 4706 4740 4712 4752
rect 3789 4703 3847 4709
rect 3896 4712 4712 4740
rect 2225 4675 2283 4681
rect 2225 4641 2237 4675
rect 2271 4641 2283 4675
rect 2225 4635 2283 4641
rect 2498 4632 2504 4684
rect 2556 4672 2562 4684
rect 2961 4675 3019 4681
rect 2961 4672 2973 4675
rect 2556 4644 2973 4672
rect 2556 4632 2562 4644
rect 2961 4641 2973 4644
rect 3007 4641 3019 4675
rect 3896 4672 3924 4712
rect 4706 4700 4712 4712
rect 4764 4700 4770 4752
rect 6546 4700 6552 4752
rect 6604 4740 6610 4752
rect 6730 4740 6736 4752
rect 6604 4712 6736 4740
rect 6604 4700 6610 4712
rect 6730 4700 6736 4712
rect 6788 4740 6794 4752
rect 6788 4712 7236 4740
rect 6788 4700 6794 4712
rect 2961 4635 3019 4641
rect 3068 4644 3924 4672
rect 4433 4675 4491 4681
rect 1489 4607 1547 4613
rect 1489 4573 1501 4607
rect 1535 4604 1547 4607
rect 1578 4604 1584 4616
rect 1535 4576 1584 4604
rect 1535 4573 1547 4576
rect 1489 4567 1547 4573
rect 1578 4564 1584 4576
rect 1636 4564 1642 4616
rect 1670 4564 1676 4616
rect 1728 4604 1734 4616
rect 1765 4607 1823 4613
rect 1765 4604 1777 4607
rect 1728 4576 1777 4604
rect 1728 4564 1734 4576
rect 1765 4573 1777 4576
rect 1811 4573 1823 4607
rect 2406 4604 2412 4616
rect 2367 4576 2412 4604
rect 1765 4567 1823 4573
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 2317 4539 2375 4545
rect 2317 4505 2329 4539
rect 2363 4536 2375 4539
rect 2682 4536 2688 4548
rect 2363 4508 2688 4536
rect 2363 4505 2375 4508
rect 2317 4499 2375 4505
rect 2682 4496 2688 4508
rect 2740 4496 2746 4548
rect 2866 4496 2872 4548
rect 2924 4536 2930 4548
rect 3068 4536 3096 4644
rect 4433 4641 4445 4675
rect 4479 4672 4491 4675
rect 4890 4672 4896 4684
rect 4479 4644 4896 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 4890 4632 4896 4644
rect 4948 4632 4954 4684
rect 6914 4672 6920 4684
rect 6875 4644 6920 4672
rect 6914 4632 6920 4644
rect 6972 4632 6978 4684
rect 3234 4564 3240 4616
rect 3292 4604 3298 4616
rect 3292 4576 6040 4604
rect 3292 4564 3298 4576
rect 2924 4508 3096 4536
rect 2924 4496 2930 4508
rect 4062 4496 4068 4548
rect 4120 4536 4126 4548
rect 4157 4539 4215 4545
rect 4157 4536 4169 4539
rect 4120 4508 4169 4536
rect 4120 4496 4126 4508
rect 4157 4505 4169 4508
rect 4203 4505 4215 4539
rect 4614 4536 4620 4548
rect 4575 4508 4620 4536
rect 4157 4499 4215 4505
rect 4614 4496 4620 4508
rect 4672 4496 4678 4548
rect 4706 4496 4712 4548
rect 4764 4536 4770 4548
rect 5914 4539 5972 4545
rect 5914 4536 5926 4539
rect 4764 4508 5926 4536
rect 4764 4496 4770 4508
rect 5914 4505 5926 4508
rect 5960 4505 5972 4539
rect 6012 4536 6040 4576
rect 6086 4564 6092 4616
rect 6144 4604 6150 4616
rect 6181 4607 6239 4613
rect 6181 4604 6193 4607
rect 6144 4576 6193 4604
rect 6144 4564 6150 4576
rect 6181 4573 6193 4576
rect 6227 4573 6239 4607
rect 6181 4567 6239 4573
rect 6270 4564 6276 4616
rect 6328 4604 6334 4616
rect 6641 4607 6699 4613
rect 6641 4604 6653 4607
rect 6328 4576 6653 4604
rect 6328 4564 6334 4576
rect 6641 4573 6653 4576
rect 6687 4573 6699 4607
rect 6641 4567 6699 4573
rect 7101 4607 7159 4613
rect 7101 4573 7113 4607
rect 7147 4573 7159 4607
rect 7208 4604 7236 4712
rect 8110 4700 8116 4752
rect 8168 4740 8174 4752
rect 11256 4740 11284 4780
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 11517 4811 11575 4817
rect 11517 4777 11529 4811
rect 11563 4808 11575 4811
rect 11698 4808 11704 4820
rect 11563 4780 11704 4808
rect 11563 4777 11575 4780
rect 11517 4771 11575 4777
rect 11698 4768 11704 4780
rect 11756 4768 11762 4820
rect 13262 4768 13268 4820
rect 13320 4808 13326 4820
rect 13357 4811 13415 4817
rect 13357 4808 13369 4811
rect 13320 4780 13369 4808
rect 13320 4768 13326 4780
rect 13357 4777 13369 4780
rect 13403 4777 13415 4811
rect 13357 4771 13415 4777
rect 13722 4768 13728 4820
rect 13780 4808 13786 4820
rect 14093 4811 14151 4817
rect 14093 4808 14105 4811
rect 13780 4780 14105 4808
rect 13780 4768 13786 4780
rect 14093 4777 14105 4780
rect 14139 4777 14151 4811
rect 18046 4808 18052 4820
rect 14093 4771 14151 4777
rect 16592 4780 18052 4808
rect 13449 4743 13507 4749
rect 13449 4740 13461 4743
rect 8168 4712 11192 4740
rect 11256 4712 12112 4740
rect 8168 4700 8174 4712
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 7834 4672 7840 4684
rect 7432 4644 7840 4672
rect 7432 4632 7438 4644
rect 7834 4632 7840 4644
rect 7892 4632 7898 4684
rect 8205 4675 8263 4681
rect 8205 4641 8217 4675
rect 8251 4672 8263 4675
rect 8570 4672 8576 4684
rect 8251 4644 8576 4672
rect 8251 4641 8263 4644
rect 8205 4635 8263 4641
rect 8570 4632 8576 4644
rect 8628 4672 8634 4684
rect 8628 4644 8984 4672
rect 8628 4632 8634 4644
rect 7929 4607 7987 4613
rect 7929 4604 7941 4607
rect 7208 4576 7941 4604
rect 7101 4567 7159 4573
rect 7929 4573 7941 4576
rect 7975 4573 7987 4607
rect 7929 4567 7987 4573
rect 7116 4536 7144 4567
rect 8018 4564 8024 4616
rect 8076 4604 8082 4616
rect 8386 4604 8392 4616
rect 8076 4576 8392 4604
rect 8076 4564 8082 4576
rect 8386 4564 8392 4576
rect 8444 4564 8450 4616
rect 8956 4613 8984 4644
rect 9122 4632 9128 4684
rect 9180 4672 9186 4684
rect 9953 4675 10011 4681
rect 9953 4672 9965 4675
rect 9180 4644 9965 4672
rect 9180 4632 9186 4644
rect 9953 4641 9965 4644
rect 9999 4641 10011 4675
rect 10870 4672 10876 4684
rect 10831 4644 10876 4672
rect 9953 4635 10011 4641
rect 10870 4632 10876 4644
rect 10928 4632 10934 4684
rect 10965 4675 11023 4681
rect 10965 4641 10977 4675
rect 11011 4672 11023 4675
rect 11054 4672 11060 4684
rect 11011 4644 11060 4672
rect 11011 4641 11023 4644
rect 10965 4635 11023 4641
rect 11054 4632 11060 4644
rect 11112 4632 11118 4684
rect 11164 4672 11192 4712
rect 12084 4681 12112 4712
rect 12268 4712 13461 4740
rect 12069 4675 12127 4681
rect 11164 4644 12020 4672
rect 8941 4607 8999 4613
rect 8941 4573 8953 4607
rect 8987 4573 8999 4607
rect 8941 4567 8999 4573
rect 10134 4564 10140 4616
rect 10192 4604 10198 4616
rect 10229 4607 10287 4613
rect 10229 4604 10241 4607
rect 10192 4576 10241 4604
rect 10192 4564 10198 4576
rect 10229 4573 10241 4576
rect 10275 4573 10287 4607
rect 11885 4607 11943 4613
rect 11885 4604 11897 4607
rect 10229 4567 10287 4573
rect 11808 4576 11897 4604
rect 6012 4508 7144 4536
rect 5914 4499 5972 4505
rect 8202 4496 8208 4548
rect 8260 4536 8266 4548
rect 8481 4539 8539 4545
rect 8481 4536 8493 4539
rect 8260 4508 8493 4536
rect 8260 4496 8266 4508
rect 8481 4505 8493 4508
rect 8527 4505 8539 4539
rect 8481 4499 8539 4505
rect 8665 4539 8723 4545
rect 8665 4505 8677 4539
rect 8711 4536 8723 4539
rect 8754 4536 8760 4548
rect 8711 4508 8760 4536
rect 8711 4505 8723 4508
rect 8665 4499 8723 4505
rect 8754 4496 8760 4508
rect 8812 4536 8818 4548
rect 9214 4536 9220 4548
rect 8812 4508 9220 4536
rect 8812 4496 8818 4508
rect 9214 4496 9220 4508
rect 9272 4536 9278 4548
rect 9490 4536 9496 4548
rect 9272 4508 9496 4536
rect 9272 4496 9278 4508
rect 9490 4496 9496 4508
rect 9548 4496 9554 4548
rect 11054 4536 11060 4548
rect 9600 4508 11060 4536
rect 3142 4468 3148 4480
rect 3103 4440 3148 4468
rect 3142 4428 3148 4440
rect 3200 4428 3206 4480
rect 3234 4428 3240 4480
rect 3292 4468 3298 4480
rect 3292 4440 3337 4468
rect 3292 4428 3298 4440
rect 3878 4428 3884 4480
rect 3936 4468 3942 4480
rect 4246 4468 4252 4480
rect 3936 4440 4252 4468
rect 3936 4428 3942 4440
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 4801 4471 4859 4477
rect 4801 4437 4813 4471
rect 4847 4468 4859 4471
rect 5442 4468 5448 4480
rect 4847 4440 5448 4468
rect 4847 4437 4859 4440
rect 4801 4431 4859 4437
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 5718 4428 5724 4480
rect 5776 4468 5782 4480
rect 6273 4471 6331 4477
rect 6273 4468 6285 4471
rect 5776 4440 6285 4468
rect 5776 4428 5782 4440
rect 6273 4437 6285 4440
rect 6319 4437 6331 4471
rect 6273 4431 6331 4437
rect 6546 4428 6552 4480
rect 6604 4468 6610 4480
rect 6733 4471 6791 4477
rect 6733 4468 6745 4471
rect 6604 4440 6745 4468
rect 6604 4428 6610 4440
rect 6733 4437 6745 4440
rect 6779 4437 6791 4471
rect 6733 4431 6791 4437
rect 7285 4471 7343 4477
rect 7285 4437 7297 4471
rect 7331 4468 7343 4471
rect 7742 4468 7748 4480
rect 7331 4440 7748 4468
rect 7331 4437 7343 4440
rect 7285 4431 7343 4437
rect 7742 4428 7748 4440
rect 7800 4428 7806 4480
rect 7834 4428 7840 4480
rect 7892 4468 7898 4480
rect 8021 4471 8079 4477
rect 8021 4468 8033 4471
rect 7892 4440 8033 4468
rect 7892 4428 7898 4440
rect 8021 4437 8033 4440
rect 8067 4437 8079 4471
rect 8021 4431 8079 4437
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 9600 4468 9628 4508
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 11422 4496 11428 4548
rect 11480 4536 11486 4548
rect 11808 4536 11836 4576
rect 11885 4573 11897 4576
rect 11931 4573 11943 4607
rect 11992 4604 12020 4644
rect 12069 4641 12081 4675
rect 12115 4641 12127 4675
rect 12069 4635 12127 4641
rect 12268 4604 12296 4712
rect 13449 4709 13461 4712
rect 13495 4709 13507 4743
rect 13449 4703 13507 4709
rect 13906 4700 13912 4752
rect 13964 4740 13970 4752
rect 15473 4743 15531 4749
rect 15473 4740 15485 4743
rect 13964 4712 15485 4740
rect 13964 4700 13970 4712
rect 15473 4709 15485 4712
rect 15519 4709 15531 4743
rect 15473 4703 15531 4709
rect 12710 4672 12716 4684
rect 12671 4644 12716 4672
rect 12710 4632 12716 4644
rect 12768 4632 12774 4684
rect 12802 4632 12808 4684
rect 12860 4672 12866 4684
rect 13817 4675 13875 4681
rect 13817 4672 13829 4675
rect 12860 4644 13829 4672
rect 12860 4632 12866 4644
rect 13817 4641 13829 4644
rect 13863 4641 13875 4675
rect 13817 4635 13875 4641
rect 14737 4675 14795 4681
rect 14737 4641 14749 4675
rect 14783 4641 14795 4675
rect 14737 4635 14795 4641
rect 11992 4576 12296 4604
rect 11885 4567 11943 4573
rect 12526 4564 12532 4616
rect 12584 4604 12590 4616
rect 13633 4607 13691 4613
rect 13633 4604 13645 4607
rect 12584 4576 13645 4604
rect 12584 4564 12590 4576
rect 13633 4573 13645 4576
rect 13679 4573 13691 4607
rect 14752 4604 14780 4635
rect 15654 4632 15660 4684
rect 15712 4672 15718 4684
rect 16592 4681 16620 4780
rect 18046 4768 18052 4780
rect 18104 4768 18110 4820
rect 17497 4743 17555 4749
rect 17497 4709 17509 4743
rect 17543 4740 17555 4743
rect 18138 4740 18144 4752
rect 17543 4712 18144 4740
rect 17543 4709 17555 4712
rect 17497 4703 17555 4709
rect 18138 4700 18144 4712
rect 18196 4700 18202 4752
rect 16577 4675 16635 4681
rect 15712 4644 15757 4672
rect 15712 4632 15718 4644
rect 16577 4641 16589 4675
rect 16623 4641 16635 4675
rect 16577 4635 16635 4641
rect 16666 4632 16672 4684
rect 16724 4672 16730 4684
rect 16761 4675 16819 4681
rect 16761 4672 16773 4675
rect 16724 4644 16773 4672
rect 16724 4632 16730 4644
rect 16761 4641 16773 4644
rect 16807 4641 16819 4675
rect 17954 4672 17960 4684
rect 17915 4644 17960 4672
rect 16761 4635 16819 4641
rect 17954 4632 17960 4644
rect 18012 4632 18018 4684
rect 15470 4604 15476 4616
rect 14752 4576 15476 4604
rect 13633 4567 13691 4573
rect 15470 4564 15476 4576
rect 15528 4564 15534 4616
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4604 16911 4607
rect 16942 4604 16948 4616
rect 16899 4576 16948 4604
rect 16899 4573 16911 4576
rect 16853 4567 16911 4573
rect 16942 4564 16948 4576
rect 17000 4564 17006 4616
rect 17313 4607 17371 4613
rect 17313 4604 17325 4607
rect 17236 4576 17325 4604
rect 12897 4539 12955 4545
rect 12897 4536 12909 4539
rect 11480 4508 11836 4536
rect 11900 4508 12909 4536
rect 11480 4496 11486 4508
rect 8352 4440 9628 4468
rect 8352 4428 8358 4440
rect 9674 4428 9680 4480
rect 9732 4468 9738 4480
rect 10042 4468 10048 4480
rect 9732 4440 10048 4468
rect 9732 4428 9738 4440
rect 10042 4428 10048 4440
rect 10100 4428 10106 4480
rect 10137 4471 10195 4477
rect 10137 4437 10149 4471
rect 10183 4468 10195 4471
rect 10318 4468 10324 4480
rect 10183 4440 10324 4468
rect 10183 4437 10195 4440
rect 10137 4431 10195 4437
rect 10318 4428 10324 4440
rect 10376 4428 10382 4480
rect 10597 4471 10655 4477
rect 10597 4437 10609 4471
rect 10643 4468 10655 4471
rect 10686 4468 10692 4480
rect 10643 4440 10692 4468
rect 10643 4437 10655 4440
rect 10597 4431 10655 4437
rect 10686 4428 10692 4440
rect 10744 4428 10750 4480
rect 10870 4428 10876 4480
rect 10928 4468 10934 4480
rect 11900 4468 11928 4508
rect 12897 4505 12909 4508
rect 12943 4505 12955 4539
rect 12897 4499 12955 4505
rect 12986 4496 12992 4548
rect 13044 4536 13050 4548
rect 13044 4508 13089 4536
rect 13044 4496 13050 4508
rect 13722 4496 13728 4548
rect 13780 4536 13786 4548
rect 15105 4539 15163 4545
rect 15105 4536 15117 4539
rect 13780 4508 15117 4536
rect 13780 4496 13786 4508
rect 15105 4505 15117 4508
rect 15151 4505 15163 4539
rect 15105 4499 15163 4505
rect 10928 4440 11928 4468
rect 11977 4471 12035 4477
rect 10928 4428 10934 4440
rect 11977 4437 11989 4471
rect 12023 4468 12035 4471
rect 12342 4468 12348 4480
rect 12023 4440 12348 4468
rect 12023 4437 12035 4440
rect 11977 4431 12035 4437
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 12492 4440 12537 4468
rect 12492 4428 12498 4440
rect 12618 4428 12624 4480
rect 12676 4468 12682 4480
rect 14182 4468 14188 4480
rect 12676 4440 14188 4468
rect 12676 4428 12682 4440
rect 14182 4428 14188 4440
rect 14240 4468 14246 4480
rect 14461 4471 14519 4477
rect 14461 4468 14473 4471
rect 14240 4440 14473 4468
rect 14240 4428 14246 4440
rect 14461 4437 14473 4440
rect 14507 4437 14519 4471
rect 14461 4431 14519 4437
rect 14550 4428 14556 4480
rect 14608 4468 14614 4480
rect 14918 4468 14924 4480
rect 14608 4440 14653 4468
rect 14879 4440 14924 4468
rect 14608 4428 14614 4440
rect 14918 4428 14924 4440
rect 14976 4428 14982 4480
rect 15381 4471 15439 4477
rect 15381 4437 15393 4471
rect 15427 4468 15439 4471
rect 15562 4468 15568 4480
rect 15427 4440 15568 4468
rect 15427 4437 15439 4440
rect 15381 4431 15439 4437
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 15838 4468 15844 4480
rect 15799 4440 15844 4468
rect 15838 4428 15844 4440
rect 15896 4428 15902 4480
rect 17236 4477 17264 4576
rect 17313 4573 17325 4576
rect 17359 4573 17371 4607
rect 17313 4567 17371 4573
rect 17770 4536 17776 4548
rect 17731 4508 17776 4536
rect 17770 4496 17776 4508
rect 17828 4496 17834 4548
rect 17221 4471 17279 4477
rect 17221 4437 17233 4471
rect 17267 4437 17279 4471
rect 17221 4431 17279 4437
rect 1104 4378 21896 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21896 4378
rect 1104 4304 21896 4326
rect 2406 4264 2412 4276
rect 2367 4236 2412 4264
rect 2406 4224 2412 4236
rect 2464 4224 2470 4276
rect 2501 4267 2559 4273
rect 2501 4233 2513 4267
rect 2547 4264 2559 4267
rect 2866 4264 2872 4276
rect 2547 4236 2872 4264
rect 2547 4233 2559 4236
rect 2501 4227 2559 4233
rect 2866 4224 2872 4236
rect 2924 4224 2930 4276
rect 2961 4267 3019 4273
rect 2961 4233 2973 4267
rect 3007 4264 3019 4267
rect 3142 4264 3148 4276
rect 3007 4236 3148 4264
rect 3007 4233 3019 4236
rect 2961 4227 3019 4233
rect 3142 4224 3148 4236
rect 3200 4224 3206 4276
rect 3234 4224 3240 4276
rect 3292 4264 3298 4276
rect 3789 4267 3847 4273
rect 3789 4264 3801 4267
rect 3292 4236 3801 4264
rect 3292 4224 3298 4236
rect 3789 4233 3801 4236
rect 3835 4233 3847 4267
rect 7098 4264 7104 4276
rect 3789 4227 3847 4233
rect 4080 4236 7104 4264
rect 3329 4199 3387 4205
rect 1964 4168 2728 4196
rect 658 4088 664 4140
rect 716 4128 722 4140
rect 1964 4128 1992 4168
rect 716 4100 1992 4128
rect 716 4088 722 4100
rect 2038 4088 2044 4140
rect 2096 4128 2102 4140
rect 2700 4128 2728 4168
rect 3329 4165 3341 4199
rect 3375 4196 3387 4199
rect 4080 4196 4108 4236
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 7466 4224 7472 4276
rect 7524 4264 7530 4276
rect 7653 4267 7711 4273
rect 7653 4264 7665 4267
rect 7524 4236 7665 4264
rect 7524 4224 7530 4236
rect 7653 4233 7665 4236
rect 7699 4233 7711 4267
rect 7653 4227 7711 4233
rect 7742 4224 7748 4276
rect 7800 4264 7806 4276
rect 10870 4264 10876 4276
rect 7800 4236 10876 4264
rect 7800 4224 7806 4236
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 12161 4267 12219 4273
rect 12161 4264 12173 4267
rect 10980 4236 12173 4264
rect 4430 4196 4436 4208
rect 3375 4168 4108 4196
rect 4172 4168 4436 4196
rect 3375 4165 3387 4168
rect 3329 4159 3387 4165
rect 3142 4128 3148 4140
rect 2096 4100 2141 4128
rect 2700 4100 3148 4128
rect 2096 4088 2102 4100
rect 3142 4088 3148 4100
rect 3200 4088 3206 4140
rect 4062 4128 4068 4140
rect 3436 4100 4068 4128
rect 2317 4063 2375 4069
rect 2317 4029 2329 4063
rect 2363 4060 2375 4063
rect 3234 4060 3240 4072
rect 2363 4032 3240 4060
rect 2363 4029 2375 4032
rect 2317 4023 2375 4029
rect 3234 4020 3240 4032
rect 3292 4020 3298 4072
rect 3436 4069 3464 4100
rect 4062 4088 4068 4100
rect 4120 4088 4126 4140
rect 4172 4137 4200 4168
rect 4430 4156 4436 4168
rect 4488 4196 4494 4208
rect 4890 4196 4896 4208
rect 4488 4168 4896 4196
rect 4488 4156 4494 4168
rect 4890 4156 4896 4168
rect 4948 4156 4954 4208
rect 5258 4156 5264 4208
rect 5316 4156 5322 4208
rect 6181 4199 6239 4205
rect 6181 4165 6193 4199
rect 6227 4196 6239 4199
rect 6733 4199 6791 4205
rect 6733 4196 6745 4199
rect 6227 4168 6745 4196
rect 6227 4165 6239 4168
rect 6181 4159 6239 4165
rect 6733 4165 6745 4168
rect 6779 4165 6791 4199
rect 6733 4159 6791 4165
rect 7006 4156 7012 4208
rect 7064 4196 7070 4208
rect 10980 4205 11008 4236
rect 12161 4233 12173 4236
rect 12207 4233 12219 4267
rect 12161 4227 12219 4233
rect 12710 4224 12716 4276
rect 12768 4264 12774 4276
rect 15381 4267 15439 4273
rect 15381 4264 15393 4267
rect 12768 4236 15393 4264
rect 12768 4224 12774 4236
rect 15381 4233 15393 4236
rect 15427 4264 15439 4267
rect 15470 4264 15476 4276
rect 15427 4236 15476 4264
rect 15427 4233 15439 4236
rect 15381 4227 15439 4233
rect 15470 4224 15476 4236
rect 15528 4224 15534 4276
rect 7561 4199 7619 4205
rect 7561 4196 7573 4199
rect 7064 4168 7573 4196
rect 7064 4156 7070 4168
rect 7561 4165 7573 4168
rect 7607 4196 7619 4199
rect 10965 4199 11023 4205
rect 10965 4196 10977 4199
rect 7607 4168 10977 4196
rect 7607 4165 7619 4168
rect 7561 4159 7619 4165
rect 10965 4165 10977 4168
rect 11011 4165 11023 4199
rect 10965 4159 11023 4165
rect 11054 4156 11060 4208
rect 11112 4196 11118 4208
rect 12069 4199 12127 4205
rect 12069 4196 12081 4199
rect 11112 4168 12081 4196
rect 11112 4156 11118 4168
rect 12069 4165 12081 4168
rect 12115 4165 12127 4199
rect 12069 4159 12127 4165
rect 14182 4156 14188 4208
rect 14240 4196 14246 4208
rect 17954 4196 17960 4208
rect 14240 4168 17960 4196
rect 14240 4156 14246 4168
rect 17954 4156 17960 4168
rect 18012 4156 18018 4208
rect 4157 4131 4215 4137
rect 4157 4097 4169 4131
rect 4203 4097 4215 4131
rect 5166 4128 5172 4140
rect 5127 4100 5172 4128
rect 4157 4091 4215 4097
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 5276 4128 5304 4156
rect 5721 4131 5779 4137
rect 5276 4100 5580 4128
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4029 3479 4063
rect 3421 4023 3479 4029
rect 3513 4063 3571 4069
rect 3513 4029 3525 4063
rect 3559 4029 3571 4063
rect 4246 4060 4252 4072
rect 4207 4032 4252 4060
rect 3513 4023 3571 4029
rect 1302 3952 1308 4004
rect 1360 3992 1366 4004
rect 2222 3992 2228 4004
rect 1360 3964 2228 3992
rect 1360 3952 1366 3964
rect 2222 3952 2228 3964
rect 2280 3952 2286 4004
rect 3050 3952 3056 4004
rect 3108 3992 3114 4004
rect 3528 3992 3556 4023
rect 4246 4020 4252 4032
rect 4304 4020 4310 4072
rect 4338 4020 4344 4072
rect 4396 4060 4402 4072
rect 5258 4060 5264 4072
rect 4396 4032 4441 4060
rect 5219 4032 5264 4060
rect 4396 4020 4402 4032
rect 5258 4020 5264 4032
rect 5316 4020 5322 4072
rect 5442 4060 5448 4072
rect 5403 4032 5448 4060
rect 5442 4020 5448 4032
rect 5500 4020 5506 4072
rect 5552 4060 5580 4100
rect 5721 4097 5733 4131
rect 5767 4128 5779 4131
rect 6638 4128 6644 4140
rect 5767 4100 6644 4128
rect 5767 4097 5779 4100
rect 5721 4091 5779 4097
rect 6638 4088 6644 4100
rect 6696 4088 6702 4140
rect 8294 4128 8300 4140
rect 7392 4100 8300 4128
rect 6825 4063 6883 4069
rect 6825 4060 6837 4063
rect 5552 4032 6837 4060
rect 6825 4029 6837 4032
rect 6871 4029 6883 4063
rect 6825 4023 6883 4029
rect 6914 4020 6920 4072
rect 6972 4060 6978 4072
rect 6972 4032 7017 4060
rect 6972 4020 6978 4032
rect 3108 3964 3556 3992
rect 3108 3952 3114 3964
rect 4430 3952 4436 4004
rect 4488 3992 4494 4004
rect 6365 3995 6423 4001
rect 6365 3992 6377 3995
rect 4488 3964 6377 3992
rect 4488 3952 4494 3964
rect 6365 3961 6377 3964
rect 6411 3961 6423 3995
rect 6365 3955 6423 3961
rect 6638 3952 6644 4004
rect 6696 3992 6702 4004
rect 7392 3992 7420 4100
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8478 4128 8484 4140
rect 8439 4100 8484 4128
rect 8478 4088 8484 4100
rect 8536 4088 8542 4140
rect 9306 4128 9312 4140
rect 9267 4100 9312 4128
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9950 4088 9956 4140
rect 10008 4128 10014 4140
rect 10045 4131 10103 4137
rect 10045 4128 10057 4131
rect 10008 4100 10057 4128
rect 10008 4088 10014 4100
rect 10045 4097 10057 4100
rect 10091 4097 10103 4131
rect 10045 4091 10103 4097
rect 10137 4131 10195 4137
rect 10137 4097 10149 4131
rect 10183 4128 10195 4131
rect 12434 4128 12440 4140
rect 10183 4100 12440 4128
rect 10183 4097 10195 4100
rect 10137 4091 10195 4097
rect 12434 4088 12440 4100
rect 12492 4088 12498 4140
rect 12526 4088 12532 4140
rect 12584 4128 12590 4140
rect 12621 4131 12679 4137
rect 12621 4128 12633 4131
rect 12584 4100 12633 4128
rect 12584 4088 12590 4100
rect 12621 4097 12633 4100
rect 12667 4097 12679 4131
rect 12621 4091 12679 4097
rect 13541 4131 13599 4137
rect 13541 4097 13553 4131
rect 13587 4128 13599 4131
rect 13630 4128 13636 4140
rect 13587 4100 13636 4128
rect 13587 4097 13599 4100
rect 13541 4091 13599 4097
rect 13630 4088 13636 4100
rect 13688 4088 13694 4140
rect 14274 4137 14280 4140
rect 14268 4091 14280 4137
rect 14332 4128 14338 4140
rect 14332 4100 14368 4128
rect 14274 4088 14280 4091
rect 14332 4088 14338 4100
rect 14734 4088 14740 4140
rect 14792 4128 14798 4140
rect 20254 4128 20260 4140
rect 14792 4100 20260 4128
rect 14792 4088 14798 4100
rect 20254 4088 20260 4100
rect 20312 4088 20318 4140
rect 7469 4063 7527 4069
rect 7469 4029 7481 4063
rect 7515 4029 7527 4063
rect 7469 4023 7527 4029
rect 6696 3964 7420 3992
rect 7484 3992 7512 4023
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 8573 4063 8631 4069
rect 8573 4060 8585 4063
rect 7708 4032 8585 4060
rect 7708 4020 7714 4032
rect 8573 4029 8585 4032
rect 8619 4029 8631 4063
rect 8754 4060 8760 4072
rect 8715 4032 8760 4060
rect 8573 4023 8631 4029
rect 8202 3992 8208 4004
rect 7484 3964 8208 3992
rect 6696 3952 6702 3964
rect 8202 3952 8208 3964
rect 8260 3992 8266 4004
rect 8478 3992 8484 4004
rect 8260 3964 8484 3992
rect 8260 3952 8266 3964
rect 8478 3952 8484 3964
rect 8536 3952 8542 4004
rect 1397 3927 1455 3933
rect 1397 3893 1409 3927
rect 1443 3924 1455 3927
rect 2038 3924 2044 3936
rect 1443 3896 2044 3924
rect 1443 3893 1455 3896
rect 1397 3887 1455 3893
rect 2038 3884 2044 3896
rect 2096 3884 2102 3936
rect 2869 3927 2927 3933
rect 2869 3893 2881 3927
rect 2915 3924 2927 3927
rect 4062 3924 4068 3936
rect 2915 3896 4068 3924
rect 2915 3893 2927 3896
rect 2869 3887 2927 3893
rect 4062 3884 4068 3896
rect 4120 3884 4126 3936
rect 4614 3924 4620 3936
rect 4575 3896 4620 3924
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4798 3924 4804 3936
rect 4759 3896 4804 3924
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 5810 3884 5816 3936
rect 5868 3924 5874 3936
rect 5905 3927 5963 3933
rect 5905 3924 5917 3927
rect 5868 3896 5917 3924
rect 5868 3884 5874 3896
rect 5905 3893 5917 3896
rect 5951 3893 5963 3927
rect 5905 3887 5963 3893
rect 7098 3884 7104 3936
rect 7156 3924 7162 3936
rect 7374 3924 7380 3936
rect 7156 3896 7380 3924
rect 7156 3884 7162 3896
rect 7374 3884 7380 3896
rect 7432 3884 7438 3936
rect 8018 3924 8024 3936
rect 7979 3896 8024 3924
rect 8018 3884 8024 3896
rect 8076 3884 8082 3936
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 8294 3924 8300 3936
rect 8159 3896 8300 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 8294 3884 8300 3896
rect 8352 3884 8358 3936
rect 8588 3924 8616 4023
rect 8754 4020 8760 4032
rect 8812 4020 8818 4072
rect 9033 4063 9091 4069
rect 9033 4029 9045 4063
rect 9079 4029 9091 4063
rect 9214 4060 9220 4072
rect 9175 4032 9220 4060
rect 9033 4023 9091 4029
rect 9048 3992 9076 4023
rect 9214 4020 9220 4032
rect 9272 4020 9278 4072
rect 9398 4020 9404 4072
rect 9456 4060 9462 4072
rect 9861 4063 9919 4069
rect 9861 4060 9873 4063
rect 9456 4032 9873 4060
rect 9456 4020 9462 4032
rect 9861 4029 9873 4032
rect 9907 4029 9919 4063
rect 10686 4060 10692 4072
rect 10647 4032 10692 4060
rect 9861 4023 9919 4029
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 11514 4060 11520 4072
rect 11475 4032 11520 4060
rect 11514 4020 11520 4032
rect 11572 4020 11578 4072
rect 11977 4063 12035 4069
rect 11977 4029 11989 4063
rect 12023 4029 12035 4063
rect 13078 4060 13084 4072
rect 11977 4023 12035 4029
rect 12406 4032 13084 4060
rect 9122 3992 9128 4004
rect 9048 3964 9128 3992
rect 9122 3952 9128 3964
rect 9180 3952 9186 4004
rect 9677 3995 9735 4001
rect 9677 3961 9689 3995
rect 9723 3992 9735 3995
rect 11992 3992 12020 4023
rect 12406 3992 12434 4032
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 13354 4020 13360 4072
rect 13412 4060 13418 4072
rect 14001 4063 14059 4069
rect 14001 4060 14013 4063
rect 13412 4032 14013 4060
rect 13412 4020 13418 4032
rect 14001 4029 14013 4032
rect 14047 4029 14059 4063
rect 14001 4023 14059 4029
rect 15010 4020 15016 4072
rect 15068 4060 15074 4072
rect 15841 4063 15899 4069
rect 15841 4060 15853 4063
rect 15068 4032 15853 4060
rect 15068 4020 15074 4032
rect 15841 4029 15853 4032
rect 15887 4029 15899 4063
rect 15841 4023 15899 4029
rect 16298 4020 16304 4072
rect 16356 4060 16362 4072
rect 16482 4060 16488 4072
rect 16356 4032 16488 4060
rect 16356 4020 16362 4032
rect 16482 4020 16488 4032
rect 16540 4020 16546 4072
rect 9723 3964 11928 3992
rect 11992 3964 12434 3992
rect 12529 3995 12587 4001
rect 9723 3961 9735 3964
rect 9677 3955 9735 3961
rect 10410 3924 10416 3936
rect 8588 3896 10416 3924
rect 10410 3884 10416 3896
rect 10468 3884 10474 3936
rect 10505 3927 10563 3933
rect 10505 3893 10517 3927
rect 10551 3924 10563 3927
rect 10686 3924 10692 3936
rect 10551 3896 10692 3924
rect 10551 3893 10563 3896
rect 10505 3887 10563 3893
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 11333 3927 11391 3933
rect 11333 3924 11345 3927
rect 11296 3896 11345 3924
rect 11296 3884 11302 3896
rect 11333 3893 11345 3896
rect 11379 3893 11391 3927
rect 11900 3924 11928 3964
rect 12529 3961 12541 3995
rect 12575 3992 12587 3995
rect 12575 3964 14044 3992
rect 12575 3961 12587 3964
rect 12529 3955 12587 3961
rect 12342 3924 12348 3936
rect 11900 3896 12348 3924
rect 11333 3887 11391 3893
rect 12342 3884 12348 3896
rect 12400 3884 12406 3936
rect 13262 3924 13268 3936
rect 13223 3896 13268 3924
rect 13262 3884 13268 3896
rect 13320 3884 13326 3936
rect 13357 3927 13415 3933
rect 13357 3893 13369 3927
rect 13403 3924 13415 3927
rect 13446 3924 13452 3936
rect 13403 3896 13452 3924
rect 13403 3893 13415 3896
rect 13357 3887 13415 3893
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 13630 3924 13636 3936
rect 13591 3896 13636 3924
rect 13630 3884 13636 3896
rect 13688 3884 13694 3936
rect 13814 3924 13820 3936
rect 13775 3896 13820 3924
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 14016 3924 14044 3964
rect 15286 3952 15292 4004
rect 15344 3992 15350 4004
rect 15473 3995 15531 4001
rect 15473 3992 15485 3995
rect 15344 3964 15485 3992
rect 15344 3952 15350 3964
rect 15473 3961 15485 3964
rect 15519 3961 15531 3995
rect 15473 3955 15531 3961
rect 15930 3952 15936 4004
rect 15988 3992 15994 4004
rect 16393 3995 16451 4001
rect 16393 3992 16405 3995
rect 15988 3964 16405 3992
rect 15988 3952 15994 3964
rect 16393 3961 16405 3964
rect 16439 3961 16451 3995
rect 16393 3955 16451 3961
rect 15194 3924 15200 3936
rect 14016 3896 15200 3924
rect 15194 3884 15200 3896
rect 15252 3884 15258 3936
rect 15654 3924 15660 3936
rect 15615 3896 15660 3924
rect 15654 3884 15660 3896
rect 15712 3884 15718 3936
rect 16022 3924 16028 3936
rect 15983 3896 16028 3924
rect 16022 3884 16028 3896
rect 16080 3884 16086 3936
rect 16298 3924 16304 3936
rect 16259 3896 16304 3924
rect 16298 3884 16304 3896
rect 16356 3884 16362 3936
rect 16666 3924 16672 3936
rect 16627 3896 16672 3924
rect 16666 3884 16672 3896
rect 16724 3884 16730 3936
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 1302 3680 1308 3732
rect 1360 3720 1366 3732
rect 1397 3723 1455 3729
rect 1397 3720 1409 3723
rect 1360 3692 1409 3720
rect 1360 3680 1366 3692
rect 1397 3689 1409 3692
rect 1443 3689 1455 3723
rect 1397 3683 1455 3689
rect 1670 3680 1676 3732
rect 1728 3720 1734 3732
rect 1765 3723 1823 3729
rect 1765 3720 1777 3723
rect 1728 3692 1777 3720
rect 1728 3680 1734 3692
rect 1765 3689 1777 3692
rect 1811 3689 1823 3723
rect 1765 3683 1823 3689
rect 2130 3680 2136 3732
rect 2188 3720 2194 3732
rect 3329 3723 3387 3729
rect 2188 3692 2912 3720
rect 2188 3680 2194 3692
rect 2884 3652 2912 3692
rect 3329 3689 3341 3723
rect 3375 3720 3387 3723
rect 3418 3720 3424 3732
rect 3375 3692 3424 3720
rect 3375 3689 3387 3692
rect 3329 3683 3387 3689
rect 3418 3680 3424 3692
rect 3476 3680 3482 3732
rect 3605 3723 3663 3729
rect 3605 3689 3617 3723
rect 3651 3720 3663 3723
rect 3878 3720 3884 3732
rect 3651 3692 3884 3720
rect 3651 3689 3663 3692
rect 3605 3683 3663 3689
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 4617 3723 4675 3729
rect 4617 3689 4629 3723
rect 4663 3720 4675 3723
rect 5166 3720 5172 3732
rect 4663 3692 5172 3720
rect 4663 3689 4675 3692
rect 4617 3683 4675 3689
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 6362 3720 6368 3732
rect 6323 3692 6368 3720
rect 6362 3680 6368 3692
rect 6420 3680 6426 3732
rect 7650 3720 7656 3732
rect 7392 3692 7656 3720
rect 4522 3652 4528 3664
rect 2884 3624 4528 3652
rect 4522 3612 4528 3624
rect 4580 3612 4586 3664
rect 4706 3652 4712 3664
rect 4667 3624 4712 3652
rect 4706 3612 4712 3624
rect 4764 3612 4770 3664
rect 7392 3652 7420 3692
rect 7650 3680 7656 3692
rect 7708 3680 7714 3732
rect 8386 3680 8392 3732
rect 8444 3720 8450 3732
rect 8941 3723 8999 3729
rect 8941 3720 8953 3723
rect 8444 3692 8953 3720
rect 8444 3680 8450 3692
rect 8941 3689 8953 3692
rect 8987 3689 8999 3723
rect 8941 3683 8999 3689
rect 9122 3680 9128 3732
rect 9180 3720 9186 3732
rect 10597 3723 10655 3729
rect 10597 3720 10609 3723
rect 9180 3692 10609 3720
rect 9180 3680 9186 3692
rect 10597 3689 10609 3692
rect 10643 3689 10655 3723
rect 10778 3720 10784 3732
rect 10739 3692 10784 3720
rect 10597 3683 10655 3689
rect 6656 3624 7420 3652
rect 10612 3652 10640 3683
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 13630 3720 13636 3732
rect 11020 3692 13636 3720
rect 11020 3680 11026 3692
rect 13630 3680 13636 3692
rect 13688 3680 13694 3732
rect 13909 3723 13967 3729
rect 13909 3689 13921 3723
rect 13955 3720 13967 3723
rect 14277 3723 14335 3729
rect 13955 3692 14228 3720
rect 13955 3689 13967 3692
rect 13909 3683 13967 3689
rect 12437 3655 12495 3661
rect 10612 3624 10999 3652
rect 1670 3544 1676 3596
rect 1728 3544 1734 3596
rect 1946 3584 1952 3596
rect 1907 3556 1952 3584
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 4065 3587 4123 3593
rect 4065 3553 4077 3587
rect 4111 3584 4123 3587
rect 4338 3584 4344 3596
rect 4111 3556 4344 3584
rect 4111 3553 4123 3556
rect 4065 3547 4123 3553
rect 4338 3544 4344 3556
rect 4396 3584 4402 3596
rect 4724 3584 4752 3612
rect 6656 3584 6684 3624
rect 4396 3556 4752 3584
rect 6012 3556 6684 3584
rect 6733 3587 6791 3593
rect 4396 3544 4402 3556
rect 1688 3516 1716 3544
rect 2216 3519 2274 3525
rect 2216 3516 2228 3519
rect 1688 3488 2228 3516
rect 2216 3485 2228 3488
rect 2262 3516 2274 3519
rect 2498 3516 2504 3528
rect 2262 3488 2504 3516
rect 2262 3485 2274 3488
rect 2216 3479 2274 3485
rect 2498 3476 2504 3488
rect 2556 3476 2562 3528
rect 2958 3476 2964 3528
rect 3016 3516 3022 3528
rect 3421 3519 3479 3525
rect 3421 3516 3433 3519
rect 3016 3488 3433 3516
rect 3016 3476 3022 3488
rect 3421 3485 3433 3488
rect 3467 3485 3479 3519
rect 3421 3479 3479 3485
rect 3878 3476 3884 3528
rect 3936 3516 3942 3528
rect 4154 3516 4160 3528
rect 3936 3488 4160 3516
rect 3936 3476 3942 3488
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4249 3519 4307 3525
rect 4249 3485 4261 3519
rect 4295 3516 4307 3519
rect 4430 3516 4436 3528
rect 4295 3488 4436 3516
rect 4295 3485 4307 3488
rect 4249 3479 4307 3485
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 6012 3516 6040 3556
rect 6733 3553 6745 3587
rect 6779 3584 6791 3587
rect 6779 3556 7512 3584
rect 6779 3553 6791 3556
rect 6733 3547 6791 3553
rect 5092 3488 6040 3516
rect 6089 3519 6147 3525
rect 1673 3451 1731 3457
rect 1673 3417 1685 3451
rect 1719 3448 1731 3451
rect 1719 3420 2176 3448
rect 1719 3417 1731 3420
rect 1673 3411 1731 3417
rect 2148 3380 2176 3420
rect 3970 3408 3976 3460
rect 4028 3448 4034 3460
rect 5092 3448 5120 3488
rect 6089 3485 6101 3519
rect 6135 3516 6147 3519
rect 7377 3519 7435 3525
rect 7377 3516 7389 3519
rect 6135 3488 7389 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 7377 3485 7389 3488
rect 7423 3485 7435 3519
rect 7484 3516 7512 3556
rect 7650 3525 7656 3528
rect 7644 3516 7656 3525
rect 7484 3488 7656 3516
rect 7377 3479 7435 3485
rect 7644 3479 7656 3488
rect 7708 3516 7714 3528
rect 8478 3516 8484 3528
rect 7708 3488 8484 3516
rect 4028 3420 5120 3448
rect 4028 3408 4034 3420
rect 5166 3408 5172 3460
rect 5224 3448 5230 3460
rect 5626 3448 5632 3460
rect 5224 3420 5632 3448
rect 5224 3408 5230 3420
rect 5626 3408 5632 3420
rect 5684 3448 5690 3460
rect 5822 3451 5880 3457
rect 5822 3448 5834 3451
rect 5684 3420 5834 3448
rect 5684 3408 5690 3420
rect 5822 3417 5834 3420
rect 5868 3417 5880 3451
rect 5822 3411 5880 3417
rect 5994 3408 6000 3460
rect 6052 3448 6058 3460
rect 6104 3448 6132 3479
rect 7650 3476 7656 3479
rect 7708 3476 7714 3488
rect 8478 3476 8484 3488
rect 8536 3476 8542 3528
rect 9030 3516 9036 3528
rect 8588 3488 9036 3516
rect 6270 3448 6276 3460
rect 6052 3420 6132 3448
rect 6231 3420 6276 3448
rect 6052 3408 6058 3420
rect 6270 3408 6276 3420
rect 6328 3408 6334 3460
rect 8588 3448 8616 3488
rect 9030 3476 9036 3488
rect 9088 3516 9094 3528
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 9088 3488 9137 3516
rect 9088 3476 9094 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9217 3519 9275 3525
rect 9217 3485 9229 3519
rect 9263 3516 9275 3519
rect 9766 3516 9772 3528
rect 9263 3488 9772 3516
rect 9263 3485 9275 3488
rect 9217 3479 9275 3485
rect 9766 3476 9772 3488
rect 9824 3476 9830 3528
rect 10871 3519 10929 3525
rect 10871 3516 10883 3519
rect 10704 3488 10883 3516
rect 6564 3420 8616 3448
rect 9484 3451 9542 3457
rect 2866 3380 2872 3392
rect 2148 3352 2872 3380
rect 2866 3340 2872 3352
rect 2924 3340 2930 3392
rect 4154 3380 4160 3392
rect 4115 3352 4160 3380
rect 4154 3340 4160 3352
rect 4212 3340 4218 3392
rect 4614 3340 4620 3392
rect 4672 3380 4678 3392
rect 6564 3380 6592 3420
rect 9484 3417 9496 3451
rect 9530 3448 9542 3451
rect 10410 3448 10416 3460
rect 9530 3420 10416 3448
rect 9530 3417 9542 3420
rect 9484 3411 9542 3417
rect 4672 3352 6592 3380
rect 4672 3340 4678 3352
rect 6638 3340 6644 3392
rect 6696 3380 6702 3392
rect 6825 3383 6883 3389
rect 6825 3380 6837 3383
rect 6696 3352 6837 3380
rect 6696 3340 6702 3352
rect 6825 3349 6837 3352
rect 6871 3349 6883 3383
rect 6825 3343 6883 3349
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7285 3383 7343 3389
rect 6972 3352 7017 3380
rect 6972 3340 6978 3352
rect 7285 3349 7297 3383
rect 7331 3380 7343 3383
rect 7374 3380 7380 3392
rect 7331 3352 7380 3380
rect 7331 3349 7343 3352
rect 7285 3343 7343 3349
rect 7374 3340 7380 3352
rect 7432 3340 7438 3392
rect 8386 3340 8392 3392
rect 8444 3380 8450 3392
rect 8757 3383 8815 3389
rect 8757 3380 8769 3383
rect 8444 3352 8769 3380
rect 8444 3340 8450 3352
rect 8757 3349 8769 3352
rect 8803 3380 8815 3383
rect 9499 3380 9527 3411
rect 10410 3408 10416 3420
rect 10468 3408 10474 3460
rect 10704 3448 10732 3488
rect 10871 3485 10883 3488
rect 10917 3485 10929 3519
rect 10871 3479 10929 3485
rect 10971 3448 10999 3624
rect 12437 3621 12449 3655
rect 12483 3652 12495 3655
rect 12526 3652 12532 3664
rect 12483 3624 12532 3652
rect 12483 3621 12495 3624
rect 12437 3615 12495 3621
rect 12526 3612 12532 3624
rect 12584 3612 12590 3664
rect 13998 3612 14004 3664
rect 14056 3652 14062 3664
rect 14200 3652 14228 3692
rect 14277 3689 14289 3723
rect 14323 3720 14335 3723
rect 14550 3720 14556 3732
rect 14323 3692 14556 3720
rect 14323 3689 14335 3692
rect 14277 3683 14335 3689
rect 14550 3680 14556 3692
rect 14608 3680 14614 3732
rect 14734 3680 14740 3732
rect 14792 3720 14798 3732
rect 15010 3720 15016 3732
rect 14792 3692 15016 3720
rect 14792 3680 14798 3692
rect 15010 3680 15016 3692
rect 15068 3720 15074 3732
rect 15105 3723 15163 3729
rect 15105 3720 15117 3723
rect 15068 3692 15117 3720
rect 15068 3680 15074 3692
rect 15105 3689 15117 3692
rect 15151 3689 15163 3723
rect 15105 3683 15163 3689
rect 15746 3680 15752 3732
rect 15804 3720 15810 3732
rect 16114 3720 16120 3732
rect 15804 3692 16120 3720
rect 15804 3680 15810 3692
rect 16114 3680 16120 3692
rect 16172 3720 16178 3732
rect 16209 3723 16267 3729
rect 16209 3720 16221 3723
rect 16172 3692 16221 3720
rect 16172 3680 16178 3692
rect 16209 3689 16221 3692
rect 16255 3689 16267 3723
rect 16209 3683 16267 3689
rect 16390 3680 16396 3732
rect 16448 3680 16454 3732
rect 16574 3680 16580 3732
rect 16632 3720 16638 3732
rect 17037 3723 17095 3729
rect 17037 3720 17049 3723
rect 16632 3692 17049 3720
rect 16632 3680 16638 3692
rect 17037 3689 17049 3692
rect 17083 3720 17095 3723
rect 17218 3720 17224 3732
rect 17083 3692 17224 3720
rect 17083 3689 17095 3692
rect 17037 3683 17095 3689
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 17405 3723 17463 3729
rect 17405 3689 17417 3723
rect 17451 3720 17463 3723
rect 17494 3720 17500 3732
rect 17451 3692 17500 3720
rect 17451 3689 17463 3692
rect 17405 3683 17463 3689
rect 17494 3680 17500 3692
rect 17552 3720 17558 3732
rect 17770 3720 17776 3732
rect 17552 3692 17776 3720
rect 17552 3680 17558 3692
rect 17770 3680 17776 3692
rect 17828 3680 17834 3732
rect 17954 3680 17960 3732
rect 18012 3720 18018 3732
rect 21361 3723 21419 3729
rect 21361 3720 21373 3723
rect 18012 3692 21373 3720
rect 18012 3680 18018 3692
rect 21361 3689 21373 3692
rect 21407 3689 21419 3723
rect 21361 3683 21419 3689
rect 14056 3624 14872 3652
rect 14056 3612 14062 3624
rect 14844 3593 14872 3624
rect 15470 3612 15476 3664
rect 15528 3652 15534 3664
rect 15841 3655 15899 3661
rect 15841 3652 15853 3655
rect 15528 3624 15853 3652
rect 15528 3612 15534 3624
rect 15841 3621 15853 3624
rect 15887 3621 15899 3655
rect 15841 3615 15899 3621
rect 16025 3655 16083 3661
rect 16025 3621 16037 3655
rect 16071 3652 16083 3655
rect 16408 3652 16436 3680
rect 16071 3624 16436 3652
rect 16071 3621 16083 3624
rect 16025 3615 16083 3621
rect 14829 3587 14887 3593
rect 14829 3553 14841 3587
rect 14875 3553 14887 3587
rect 15562 3584 15568 3596
rect 14829 3547 14887 3553
rect 15212 3556 15568 3584
rect 11057 3519 11115 3525
rect 11057 3485 11069 3519
rect 11103 3516 11115 3519
rect 12529 3519 12587 3525
rect 12529 3516 12541 3519
rect 11103 3488 12541 3516
rect 11103 3485 11115 3488
rect 11057 3479 11115 3485
rect 12529 3485 12541 3488
rect 12575 3516 12587 3519
rect 13354 3516 13360 3528
rect 12575 3488 13360 3516
rect 12575 3485 12587 3488
rect 12529 3479 12587 3485
rect 13354 3476 13360 3488
rect 13412 3476 13418 3528
rect 15212 3516 15240 3556
rect 15562 3544 15568 3556
rect 15620 3584 15626 3596
rect 16390 3584 16396 3596
rect 15620 3556 16396 3584
rect 15620 3544 15626 3556
rect 16390 3544 16396 3556
rect 16448 3584 16454 3596
rect 16577 3587 16635 3593
rect 16577 3584 16589 3587
rect 16448 3556 16589 3584
rect 16448 3544 16454 3556
rect 16577 3553 16589 3556
rect 16623 3553 16635 3587
rect 16577 3547 16635 3553
rect 17957 3587 18015 3593
rect 17957 3553 17969 3587
rect 18003 3584 18015 3587
rect 18230 3584 18236 3596
rect 18003 3556 18236 3584
rect 18003 3553 18015 3556
rect 17957 3547 18015 3553
rect 18230 3544 18236 3556
rect 18288 3544 18294 3596
rect 15378 3516 15384 3528
rect 14752 3488 15240 3516
rect 15339 3488 15384 3516
rect 11302 3451 11360 3457
rect 11302 3448 11314 3451
rect 10704 3420 10824 3448
rect 10971 3420 11314 3448
rect 10796 3392 10824 3420
rect 11302 3417 11314 3420
rect 11348 3417 11360 3451
rect 11302 3411 11360 3417
rect 12796 3451 12854 3457
rect 12796 3417 12808 3451
rect 12842 3448 12854 3451
rect 13262 3448 13268 3460
rect 12842 3420 13268 3448
rect 12842 3417 12854 3420
rect 12796 3411 12854 3417
rect 13262 3408 13268 3420
rect 13320 3408 13326 3460
rect 14752 3457 14780 3488
rect 15378 3476 15384 3488
rect 15436 3476 15442 3528
rect 15838 3476 15844 3528
rect 15896 3516 15902 3528
rect 16482 3516 16488 3528
rect 15896 3488 16488 3516
rect 15896 3476 15902 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 18138 3516 18144 3528
rect 18099 3488 18144 3516
rect 18138 3476 18144 3488
rect 18196 3476 18202 3528
rect 21269 3519 21327 3525
rect 21269 3485 21281 3519
rect 21315 3516 21327 3519
rect 21545 3519 21603 3525
rect 21545 3516 21557 3519
rect 21315 3488 21557 3516
rect 21315 3485 21327 3488
rect 21269 3479 21327 3485
rect 21545 3485 21557 3488
rect 21591 3516 21603 3519
rect 22646 3516 22652 3528
rect 21591 3488 22652 3516
rect 21591 3485 21603 3488
rect 21545 3479 21603 3485
rect 22646 3476 22652 3488
rect 22704 3476 22710 3528
rect 14737 3451 14795 3457
rect 14737 3448 14749 3451
rect 14200 3420 14749 3448
rect 14200 3392 14228 3420
rect 14737 3417 14749 3420
rect 14783 3417 14795 3451
rect 14737 3411 14795 3417
rect 15194 3408 15200 3460
rect 15252 3448 15258 3460
rect 15657 3451 15715 3457
rect 15657 3448 15669 3451
rect 15252 3420 15669 3448
rect 15252 3408 15258 3420
rect 15657 3417 15669 3420
rect 15703 3417 15715 3451
rect 15657 3411 15715 3417
rect 16206 3408 16212 3460
rect 16264 3448 16270 3460
rect 19518 3448 19524 3460
rect 16264 3420 19524 3448
rect 16264 3408 16270 3420
rect 19518 3408 19524 3420
rect 19576 3408 19582 3460
rect 8803 3352 9527 3380
rect 8803 3349 8815 3352
rect 8757 3343 8815 3349
rect 10318 3340 10324 3392
rect 10376 3380 10382 3392
rect 10594 3380 10600 3392
rect 10376 3352 10600 3380
rect 10376 3340 10382 3352
rect 10594 3340 10600 3352
rect 10652 3340 10658 3392
rect 10778 3340 10784 3392
rect 10836 3380 10842 3392
rect 13814 3380 13820 3392
rect 10836 3352 13820 3380
rect 10836 3340 10842 3352
rect 13814 3340 13820 3352
rect 13872 3340 13878 3392
rect 14182 3380 14188 3392
rect 14143 3352 14188 3380
rect 14182 3340 14188 3352
rect 14240 3340 14246 3392
rect 14645 3383 14703 3389
rect 14645 3349 14657 3383
rect 14691 3380 14703 3383
rect 15010 3380 15016 3392
rect 14691 3352 15016 3380
rect 14691 3349 14703 3352
rect 14645 3343 14703 3349
rect 15010 3340 15016 3352
rect 15068 3340 15074 3392
rect 15562 3380 15568 3392
rect 15523 3352 15568 3380
rect 15562 3340 15568 3352
rect 15620 3340 15626 3392
rect 15746 3340 15752 3392
rect 15804 3380 15810 3392
rect 16393 3383 16451 3389
rect 16393 3380 16405 3383
rect 15804 3352 16405 3380
rect 15804 3340 15810 3352
rect 16393 3349 16405 3352
rect 16439 3349 16451 3383
rect 16393 3343 16451 3349
rect 16853 3383 16911 3389
rect 16853 3349 16865 3383
rect 16899 3380 16911 3383
rect 16942 3380 16948 3392
rect 16899 3352 16948 3380
rect 16899 3349 16911 3352
rect 16853 3343 16911 3349
rect 16942 3340 16948 3352
rect 17000 3340 17006 3392
rect 18325 3383 18383 3389
rect 18325 3349 18337 3383
rect 18371 3380 18383 3383
rect 19058 3380 19064 3392
rect 18371 3352 19064 3380
rect 18371 3349 18383 3352
rect 18325 3343 18383 3349
rect 19058 3340 19064 3352
rect 19116 3340 19122 3392
rect 1104 3290 21896 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21896 3290
rect 1104 3216 21896 3238
rect 1670 3176 1676 3188
rect 1631 3148 1676 3176
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 2038 3136 2044 3188
rect 2096 3176 2102 3188
rect 2096 3148 3188 3176
rect 2096 3136 2102 3148
rect 1946 3068 1952 3120
rect 2004 3108 2010 3120
rect 3160 3108 3188 3148
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 4617 3179 4675 3185
rect 4617 3176 4629 3179
rect 3292 3148 4629 3176
rect 3292 3136 3298 3148
rect 4617 3145 4629 3148
rect 4663 3176 4675 3179
rect 5166 3176 5172 3188
rect 4663 3148 5172 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5350 3176 5356 3188
rect 5311 3148 5356 3176
rect 5350 3136 5356 3148
rect 5408 3136 5414 3188
rect 5445 3179 5503 3185
rect 5445 3145 5457 3179
rect 5491 3145 5503 3179
rect 5902 3176 5908 3188
rect 5863 3148 5908 3176
rect 5445 3139 5503 3145
rect 3482 3111 3540 3117
rect 3482 3108 3494 3111
rect 2004 3080 3096 3108
rect 3160 3080 3494 3108
rect 2004 3068 2010 3080
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 3068 3049 3096 3080
rect 3482 3077 3494 3080
rect 3528 3077 3540 3111
rect 3482 3071 3540 3077
rect 4154 3068 4160 3120
rect 4212 3108 4218 3120
rect 5460 3108 5488 3139
rect 5902 3136 5908 3148
rect 5960 3136 5966 3188
rect 6822 3176 6828 3188
rect 6783 3148 6828 3176
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7377 3179 7435 3185
rect 7377 3145 7389 3179
rect 7423 3176 7435 3179
rect 7742 3176 7748 3188
rect 7423 3148 7748 3176
rect 7423 3145 7435 3148
rect 7377 3139 7435 3145
rect 7742 3136 7748 3148
rect 7800 3136 7806 3188
rect 8294 3176 8300 3188
rect 8255 3148 8300 3176
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 8665 3179 8723 3185
rect 8665 3145 8677 3179
rect 8711 3176 8723 3179
rect 9214 3176 9220 3188
rect 8711 3148 9220 3176
rect 8711 3145 8723 3148
rect 8665 3139 8723 3145
rect 9214 3136 9220 3148
rect 9272 3136 9278 3188
rect 9306 3136 9312 3188
rect 9364 3176 9370 3188
rect 9769 3179 9827 3185
rect 9769 3176 9781 3179
rect 9364 3148 9781 3176
rect 9364 3136 9370 3148
rect 9769 3145 9781 3148
rect 9815 3145 9827 3179
rect 10134 3176 10140 3188
rect 10095 3148 10140 3176
rect 9769 3139 9827 3145
rect 10134 3136 10140 3148
rect 10192 3136 10198 3188
rect 10594 3136 10600 3188
rect 10652 3176 10658 3188
rect 10652 3148 10697 3176
rect 10652 3136 10658 3148
rect 14274 3136 14280 3188
rect 14332 3176 14338 3188
rect 14553 3179 14611 3185
rect 14553 3176 14565 3179
rect 14332 3148 14565 3176
rect 14332 3136 14338 3148
rect 14553 3145 14565 3148
rect 14599 3145 14611 3179
rect 14553 3139 14611 3145
rect 14829 3179 14887 3185
rect 14829 3145 14841 3179
rect 14875 3145 14887 3179
rect 14829 3139 14887 3145
rect 14921 3179 14979 3185
rect 14921 3145 14933 3179
rect 14967 3176 14979 3179
rect 15102 3176 15108 3188
rect 14967 3148 15108 3176
rect 14967 3145 14979 3148
rect 14921 3139 14979 3145
rect 4212 3080 5488 3108
rect 4212 3068 4218 3080
rect 5994 3068 6000 3120
rect 6052 3108 6058 3120
rect 6365 3111 6423 3117
rect 6365 3108 6377 3111
rect 6052 3080 6377 3108
rect 6052 3068 6058 3080
rect 6365 3077 6377 3080
rect 6411 3077 6423 3111
rect 6365 3071 6423 3077
rect 6917 3111 6975 3117
rect 6917 3077 6929 3111
rect 6963 3108 6975 3111
rect 7006 3108 7012 3120
rect 6963 3080 7012 3108
rect 6963 3077 6975 3080
rect 6917 3071 6975 3077
rect 7006 3068 7012 3080
rect 7064 3068 7070 3120
rect 7282 3068 7288 3120
rect 7340 3108 7346 3120
rect 7469 3111 7527 3117
rect 7469 3108 7481 3111
rect 7340 3080 7481 3108
rect 7340 3068 7346 3080
rect 7469 3077 7481 3080
rect 7515 3077 7527 3111
rect 7469 3071 7527 3077
rect 8018 3068 8024 3120
rect 8076 3108 8082 3120
rect 8205 3111 8263 3117
rect 8205 3108 8217 3111
rect 8076 3080 8217 3108
rect 8076 3068 8082 3080
rect 8205 3077 8217 3080
rect 8251 3077 8263 3111
rect 8205 3071 8263 3077
rect 8849 3111 8907 3117
rect 8849 3077 8861 3111
rect 8895 3108 8907 3111
rect 10229 3111 10287 3117
rect 8895 3080 10180 3108
rect 8895 3077 8907 3080
rect 8849 3071 8907 3077
rect 2797 3043 2855 3049
rect 2797 3009 2809 3043
rect 2843 3040 2855 3043
rect 3053 3043 3111 3049
rect 2843 3012 3004 3040
rect 2843 3009 2855 3012
rect 2797 3003 2855 3009
rect 2976 2972 3004 3012
rect 3053 3009 3065 3043
rect 3099 3040 3111 3043
rect 4709 3043 4767 3049
rect 3099 3012 3280 3040
rect 3099 3009 3111 3012
rect 3053 3003 3111 3009
rect 3252 2984 3280 3012
rect 4709 3009 4721 3043
rect 4755 3040 4767 3043
rect 5442 3040 5448 3052
rect 4755 3012 5448 3040
rect 4755 3009 4767 3012
rect 4709 3003 4767 3009
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 5626 3000 5632 3052
rect 5684 3040 5690 3052
rect 5813 3043 5871 3049
rect 5813 3040 5825 3043
rect 5684 3012 5825 3040
rect 5684 3000 5690 3012
rect 5813 3009 5825 3012
rect 5859 3040 5871 3043
rect 6086 3040 6092 3052
rect 5859 3012 6092 3040
rect 5859 3009 5871 3012
rect 5813 3003 5871 3009
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 6546 3040 6552 3052
rect 6507 3012 6552 3040
rect 6546 3000 6552 3012
rect 6604 3000 6610 3052
rect 6656 3012 7420 3040
rect 3234 2972 3240 2984
rect 2976 2944 3096 2972
rect 3195 2944 3240 2972
rect 3068 2916 3096 2944
rect 3234 2932 3240 2944
rect 3292 2932 3298 2984
rect 4430 2932 4436 2984
rect 4488 2972 4494 2984
rect 5534 2972 5540 2984
rect 4488 2944 5540 2972
rect 4488 2932 4494 2944
rect 5534 2932 5540 2944
rect 5592 2932 5598 2984
rect 5997 2975 6055 2981
rect 5997 2972 6009 2975
rect 5644 2944 6009 2972
rect 3050 2864 3056 2916
rect 3108 2864 3114 2916
rect 4246 2864 4252 2916
rect 4304 2904 4310 2916
rect 5442 2904 5448 2916
rect 4304 2876 5448 2904
rect 4304 2864 4310 2876
rect 5442 2864 5448 2876
rect 5500 2864 5506 2916
rect 1578 2836 1584 2848
rect 1539 2808 1584 2836
rect 1578 2796 1584 2808
rect 1636 2796 1642 2848
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 5644 2836 5672 2944
rect 5997 2941 6009 2944
rect 6043 2941 6055 2975
rect 5997 2935 6055 2941
rect 6178 2932 6184 2984
rect 6236 2972 6242 2984
rect 6656 2972 6684 3012
rect 6236 2944 6684 2972
rect 7285 2975 7343 2981
rect 6236 2932 6242 2944
rect 7285 2941 7297 2975
rect 7331 2941 7343 2975
rect 7392 2972 7420 3012
rect 7926 3000 7932 3052
rect 7984 3040 7990 3052
rect 9309 3043 9367 3049
rect 9309 3040 9321 3043
rect 7984 3012 9321 3040
rect 7984 3000 7990 3012
rect 9309 3009 9321 3012
rect 9355 3009 9367 3043
rect 9309 3003 9367 3009
rect 9398 3000 9404 3052
rect 9456 3040 9462 3052
rect 10042 3040 10048 3052
rect 9456 3012 10048 3040
rect 9456 3000 9462 3012
rect 10042 3000 10048 3012
rect 10100 3000 10106 3052
rect 10152 3040 10180 3080
rect 10229 3077 10241 3111
rect 10275 3108 10287 3111
rect 10318 3108 10324 3120
rect 10275 3080 10324 3108
rect 10275 3077 10287 3080
rect 10229 3071 10287 3077
rect 10318 3068 10324 3080
rect 10376 3068 10382 3120
rect 11238 3108 11244 3120
rect 10796 3080 11244 3108
rect 10152 3012 10548 3040
rect 8113 2975 8171 2981
rect 7392 2944 7972 2972
rect 7285 2935 7343 2941
rect 7300 2904 7328 2935
rect 7650 2904 7656 2916
rect 7300 2876 7656 2904
rect 7650 2864 7656 2876
rect 7708 2864 7714 2916
rect 5224 2808 5672 2836
rect 5224 2796 5230 2808
rect 7742 2796 7748 2848
rect 7800 2836 7806 2848
rect 7837 2839 7895 2845
rect 7837 2836 7849 2839
rect 7800 2808 7849 2836
rect 7800 2796 7806 2808
rect 7837 2805 7849 2808
rect 7883 2805 7895 2839
rect 7944 2836 7972 2944
rect 8113 2941 8125 2975
rect 8159 2972 8171 2975
rect 8386 2972 8392 2984
rect 8159 2944 8392 2972
rect 8159 2941 8171 2944
rect 8113 2935 8171 2941
rect 8386 2932 8392 2944
rect 8444 2932 8450 2984
rect 8938 2932 8944 2984
rect 8996 2972 9002 2984
rect 9033 2975 9091 2981
rect 9033 2972 9045 2975
rect 8996 2944 9045 2972
rect 8996 2932 9002 2944
rect 9033 2941 9045 2944
rect 9079 2941 9091 2975
rect 9033 2935 9091 2941
rect 9217 2975 9275 2981
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 9582 2972 9588 2984
rect 9263 2944 9588 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 9582 2932 9588 2944
rect 9640 2932 9646 2984
rect 10410 2972 10416 2984
rect 10371 2944 10416 2972
rect 10410 2932 10416 2944
rect 10468 2932 10474 2984
rect 10520 2972 10548 3012
rect 10796 2972 10824 3080
rect 11238 3068 11244 3080
rect 11296 3108 11302 3120
rect 11609 3111 11667 3117
rect 11609 3108 11621 3111
rect 11296 3080 11621 3108
rect 11296 3068 11302 3080
rect 11609 3077 11621 3080
rect 11655 3077 11667 3111
rect 11609 3071 11667 3077
rect 11793 3111 11851 3117
rect 11793 3077 11805 3111
rect 11839 3108 11851 3111
rect 11882 3108 11888 3120
rect 11839 3080 11888 3108
rect 11839 3077 11851 3080
rect 11793 3071 11851 3077
rect 11882 3068 11888 3080
rect 11940 3068 11946 3120
rect 12526 3108 12532 3120
rect 12268 3080 12532 3108
rect 10870 3000 10876 3052
rect 10928 3040 10934 3052
rect 10965 3043 11023 3049
rect 10965 3040 10977 3043
rect 10928 3012 10977 3040
rect 10928 3000 10934 3012
rect 10965 3009 10977 3012
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11112 3012 11157 3040
rect 11112 3000 11118 3012
rect 10520 2944 10824 2972
rect 11241 2975 11299 2981
rect 11241 2941 11253 2975
rect 11287 2972 11299 2975
rect 11330 2972 11336 2984
rect 11287 2944 11336 2972
rect 11287 2941 11299 2944
rect 11241 2935 11299 2941
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 12268 2981 12296 3080
rect 12526 3068 12532 3080
rect 12584 3068 12590 3120
rect 14844 3108 14872 3139
rect 15102 3136 15108 3148
rect 15160 3136 15166 3188
rect 17957 3179 18015 3185
rect 17957 3145 17969 3179
rect 18003 3145 18015 3179
rect 17957 3139 18015 3145
rect 14844 3080 15516 3108
rect 12434 3000 12440 3052
rect 12492 3040 12498 3052
rect 12894 3040 12900 3052
rect 12492 3012 12537 3040
rect 12855 3012 12900 3040
rect 12492 3000 12498 3012
rect 12894 3000 12900 3012
rect 12952 3000 12958 3052
rect 13173 3043 13231 3049
rect 13173 3009 13185 3043
rect 13219 3009 13231 3043
rect 13446 3040 13452 3052
rect 13407 3012 13452 3040
rect 13173 3003 13231 3009
rect 12253 2975 12311 2981
rect 12253 2941 12265 2975
rect 12299 2941 12311 2975
rect 12253 2935 12311 2941
rect 12345 2975 12403 2981
rect 12345 2941 12357 2975
rect 12391 2941 12403 2975
rect 13188 2972 13216 3003
rect 13446 3000 13452 3012
rect 13504 3000 13510 3052
rect 13909 3043 13967 3049
rect 13909 3009 13921 3043
rect 13955 3040 13967 3043
rect 13998 3040 14004 3052
rect 13955 3012 14004 3040
rect 13955 3009 13967 3012
rect 13909 3003 13967 3009
rect 13998 3000 14004 3012
rect 14056 3000 14062 3052
rect 14458 3000 14464 3052
rect 14516 3040 14522 3052
rect 14645 3043 14703 3049
rect 14645 3040 14657 3043
rect 14516 3012 14657 3040
rect 14516 3000 14522 3012
rect 14645 3009 14657 3012
rect 14691 3009 14703 3043
rect 15102 3040 15108 3052
rect 15063 3012 15108 3040
rect 14645 3003 14703 3009
rect 15102 3000 15108 3012
rect 15160 3000 15166 3052
rect 15378 3040 15384 3052
rect 15339 3012 15384 3040
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 15488 3049 15516 3080
rect 15746 3068 15752 3120
rect 15804 3108 15810 3120
rect 17972 3108 18000 3139
rect 18046 3136 18052 3188
rect 18104 3176 18110 3188
rect 18325 3179 18383 3185
rect 18325 3176 18337 3179
rect 18104 3148 18337 3176
rect 18104 3136 18110 3148
rect 18325 3145 18337 3148
rect 18371 3145 18383 3179
rect 18325 3139 18383 3145
rect 18598 3136 18604 3188
rect 18656 3176 18662 3188
rect 18877 3179 18935 3185
rect 18877 3176 18889 3179
rect 18656 3148 18889 3176
rect 18656 3136 18662 3148
rect 18877 3145 18889 3148
rect 18923 3145 18935 3179
rect 18877 3139 18935 3145
rect 19245 3179 19303 3185
rect 19245 3145 19257 3179
rect 19291 3176 19303 3179
rect 19978 3176 19984 3188
rect 19291 3148 19984 3176
rect 19291 3145 19303 3148
rect 19245 3139 19303 3145
rect 19978 3136 19984 3148
rect 20036 3136 20042 3188
rect 20254 3176 20260 3188
rect 20215 3148 20260 3176
rect 20254 3136 20260 3148
rect 20312 3136 20318 3188
rect 15804 3080 16344 3108
rect 17972 3080 20944 3108
rect 15804 3068 15810 3080
rect 15473 3043 15531 3049
rect 15473 3009 15485 3043
rect 15519 3009 15531 3043
rect 15473 3003 15531 3009
rect 15838 3000 15844 3052
rect 15896 3024 15902 3052
rect 16025 3044 16083 3049
rect 16114 3044 16120 3052
rect 16025 3043 16120 3044
rect 15933 3027 15991 3033
rect 15933 3024 15945 3027
rect 15896 3000 15945 3024
rect 15856 2996 15945 3000
rect 15933 2993 15945 2996
rect 15979 2993 15991 3027
rect 16025 3009 16037 3043
rect 16071 3016 16120 3043
rect 16071 3009 16083 3016
rect 16025 3003 16083 3009
rect 16114 3000 16120 3016
rect 16172 3000 16178 3052
rect 16316 3049 16344 3080
rect 16301 3043 16359 3049
rect 16301 3009 16313 3043
rect 16347 3009 16359 3043
rect 16301 3003 16359 3009
rect 16390 3000 16396 3052
rect 16448 3040 16454 3052
rect 16853 3043 16911 3049
rect 16853 3040 16865 3043
rect 16448 3012 16865 3040
rect 16448 3000 16454 3012
rect 16853 3009 16865 3012
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3040 17003 3043
rect 17034 3040 17040 3052
rect 16991 3012 17040 3040
rect 16991 3009 17003 3012
rect 16945 3003 17003 3009
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 17218 3040 17224 3052
rect 17179 3012 17224 3040
rect 17218 3000 17224 3012
rect 17276 3000 17282 3052
rect 17494 3040 17500 3052
rect 17455 3012 17500 3040
rect 17494 3000 17500 3012
rect 17552 3000 17558 3052
rect 17773 3043 17831 3049
rect 17773 3009 17785 3043
rect 17819 3040 17831 3043
rect 17954 3040 17960 3052
rect 17819 3012 17960 3040
rect 17819 3009 17831 3012
rect 17773 3003 17831 3009
rect 17954 3000 17960 3012
rect 18012 3000 18018 3052
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3040 18107 3043
rect 18230 3040 18236 3052
rect 18095 3012 18236 3040
rect 18095 3009 18107 3012
rect 18049 3003 18107 3009
rect 18230 3000 18236 3012
rect 18288 3000 18294 3052
rect 18598 3040 18604 3052
rect 18559 3012 18604 3040
rect 18598 3000 18604 3012
rect 18656 3000 18662 3052
rect 18782 3000 18788 3052
rect 18840 3040 18846 3052
rect 19061 3043 19119 3049
rect 19061 3040 19073 3043
rect 18840 3012 19073 3040
rect 18840 3000 18846 3012
rect 19061 3009 19073 3012
rect 19107 3040 19119 3043
rect 19337 3043 19395 3049
rect 19337 3040 19349 3043
rect 19107 3012 19349 3040
rect 19107 3009 19119 3012
rect 19061 3003 19119 3009
rect 19337 3009 19349 3012
rect 19383 3009 19395 3043
rect 19518 3040 19524 3052
rect 19479 3012 19524 3040
rect 19337 3003 19395 3009
rect 19518 3000 19524 3012
rect 19576 3040 19582 3052
rect 19797 3043 19855 3049
rect 19797 3040 19809 3043
rect 19576 3012 19809 3040
rect 19576 3000 19582 3012
rect 19797 3009 19809 3012
rect 19843 3009 19855 3043
rect 19797 3003 19855 3009
rect 20254 3000 20260 3052
rect 20312 3040 20318 3052
rect 20916 3049 20944 3080
rect 20441 3043 20499 3049
rect 20441 3040 20453 3043
rect 20312 3012 20453 3040
rect 20312 3000 20318 3012
rect 20441 3009 20453 3012
rect 20487 3009 20499 3043
rect 20441 3003 20499 3009
rect 20901 3043 20959 3049
rect 20901 3009 20913 3043
rect 20947 3009 20959 3043
rect 20901 3003 20959 3009
rect 21269 3043 21327 3049
rect 21269 3009 21281 3043
rect 21315 3009 21327 3043
rect 21269 3003 21327 3009
rect 15933 2987 15991 2993
rect 12345 2935 12403 2941
rect 12820 2944 13216 2972
rect 9677 2907 9735 2913
rect 9677 2873 9689 2907
rect 9723 2904 9735 2907
rect 12360 2904 12388 2935
rect 12820 2913 12848 2944
rect 13262 2932 13268 2984
rect 13320 2972 13326 2984
rect 13725 2975 13783 2981
rect 13725 2972 13737 2975
rect 13320 2944 13737 2972
rect 13320 2932 13326 2944
rect 13725 2941 13737 2944
rect 13771 2941 13783 2975
rect 21284 2972 21312 3003
rect 13725 2935 13783 2941
rect 16500 2944 21312 2972
rect 9723 2876 12388 2904
rect 12805 2907 12863 2913
rect 9723 2873 9735 2876
rect 9677 2867 9735 2873
rect 12805 2873 12817 2907
rect 12851 2873 12863 2907
rect 12805 2867 12863 2873
rect 13633 2907 13691 2913
rect 13633 2873 13645 2907
rect 13679 2904 13691 2907
rect 13814 2904 13820 2916
rect 13679 2876 13820 2904
rect 13679 2873 13691 2876
rect 13633 2867 13691 2873
rect 13814 2864 13820 2876
rect 13872 2864 13878 2916
rect 16500 2913 16528 2944
rect 16485 2907 16543 2913
rect 16485 2873 16497 2907
rect 16531 2873 16543 2907
rect 16485 2867 16543 2873
rect 17405 2907 17463 2913
rect 17405 2873 17417 2907
rect 17451 2904 17463 2907
rect 17494 2904 17500 2916
rect 17451 2876 17500 2904
rect 17451 2873 17463 2876
rect 17405 2867 17463 2873
rect 17494 2864 17500 2876
rect 17552 2864 17558 2916
rect 18785 2907 18843 2913
rect 18785 2873 18797 2907
rect 18831 2904 18843 2907
rect 19610 2904 19616 2916
rect 18831 2876 19616 2904
rect 18831 2873 18843 2876
rect 18785 2867 18843 2873
rect 19610 2864 19616 2876
rect 19668 2864 19674 2916
rect 19705 2907 19763 2913
rect 19705 2873 19717 2907
rect 19751 2904 19763 2907
rect 20438 2904 20444 2916
rect 19751 2876 20444 2904
rect 19751 2873 19763 2876
rect 19705 2867 19763 2873
rect 20438 2864 20444 2876
rect 20496 2864 20502 2916
rect 21085 2907 21143 2913
rect 21085 2873 21097 2907
rect 21131 2904 21143 2907
rect 22186 2904 22192 2916
rect 21131 2876 22192 2904
rect 21131 2873 21143 2876
rect 21085 2867 21143 2873
rect 22186 2864 22192 2876
rect 22244 2864 22250 2916
rect 10226 2836 10232 2848
rect 7944 2808 10232 2836
rect 7837 2799 7895 2805
rect 10226 2796 10232 2808
rect 10284 2796 10290 2848
rect 11882 2836 11888 2848
rect 11843 2808 11888 2836
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 13078 2836 13084 2848
rect 13039 2808 13084 2836
rect 13078 2796 13084 2808
rect 13136 2796 13142 2848
rect 13354 2836 13360 2848
rect 13315 2808 13360 2836
rect 13354 2796 13360 2808
rect 13412 2796 13418 2848
rect 15194 2836 15200 2848
rect 15155 2808 15200 2836
rect 15194 2796 15200 2808
rect 15252 2796 15258 2848
rect 15562 2796 15568 2848
rect 15620 2836 15626 2848
rect 15657 2839 15715 2845
rect 15657 2836 15669 2839
rect 15620 2808 15669 2836
rect 15620 2796 15626 2808
rect 15657 2805 15669 2808
rect 15703 2805 15715 2839
rect 15657 2799 15715 2805
rect 15746 2796 15752 2848
rect 15804 2836 15810 2848
rect 16206 2836 16212 2848
rect 15804 2808 15849 2836
rect 16167 2808 16212 2836
rect 15804 2796 15810 2808
rect 16206 2796 16212 2808
rect 16264 2796 16270 2848
rect 16669 2839 16727 2845
rect 16669 2805 16681 2839
rect 16715 2836 16727 2839
rect 16758 2836 16764 2848
rect 16715 2808 16764 2836
rect 16715 2805 16727 2808
rect 16669 2799 16727 2805
rect 16758 2796 16764 2808
rect 16816 2796 16822 2848
rect 17126 2836 17132 2848
rect 17087 2808 17132 2836
rect 17126 2796 17132 2808
rect 17184 2796 17190 2848
rect 17681 2839 17739 2845
rect 17681 2805 17693 2839
rect 17727 2836 17739 2839
rect 17770 2836 17776 2848
rect 17727 2808 17776 2836
rect 17727 2805 17739 2808
rect 17681 2799 17739 2805
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 18230 2836 18236 2848
rect 18191 2808 18236 2836
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 20625 2839 20683 2845
rect 20625 2805 20637 2839
rect 20671 2836 20683 2839
rect 20990 2836 20996 2848
rect 20671 2808 20996 2836
rect 20671 2805 20683 2808
rect 20625 2799 20683 2805
rect 20990 2796 20996 2808
rect 21048 2796 21054 2848
rect 21453 2839 21511 2845
rect 21453 2805 21465 2839
rect 21499 2836 21511 2839
rect 21726 2836 21732 2848
rect 21499 2808 21732 2836
rect 21499 2805 21511 2808
rect 21453 2799 21511 2805
rect 21726 2796 21732 2808
rect 21784 2796 21790 2848
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 3513 2635 3571 2641
rect 3513 2601 3525 2635
rect 3559 2632 3571 2635
rect 3970 2632 3976 2644
rect 3559 2604 3976 2632
rect 3559 2601 3571 2604
rect 3513 2595 3571 2601
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 4617 2635 4675 2641
rect 4617 2601 4629 2635
rect 4663 2632 4675 2635
rect 5258 2632 5264 2644
rect 4663 2604 5264 2632
rect 4663 2601 4675 2604
rect 4617 2595 4675 2601
rect 5258 2592 5264 2604
rect 5316 2592 5322 2644
rect 5442 2592 5448 2644
rect 5500 2632 5506 2644
rect 6178 2632 6184 2644
rect 5500 2604 6184 2632
rect 5500 2592 5506 2604
rect 6178 2592 6184 2604
rect 6236 2592 6242 2644
rect 6454 2632 6460 2644
rect 6415 2604 6460 2632
rect 6454 2592 6460 2604
rect 6512 2592 6518 2644
rect 6546 2592 6552 2644
rect 6604 2632 6610 2644
rect 6730 2632 6736 2644
rect 6604 2604 6736 2632
rect 6604 2592 6610 2604
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 6825 2635 6883 2641
rect 6825 2601 6837 2635
rect 6871 2632 6883 2635
rect 7190 2632 7196 2644
rect 6871 2604 7196 2632
rect 6871 2601 6883 2604
rect 6825 2595 6883 2601
rect 7190 2592 7196 2604
rect 7248 2592 7254 2644
rect 7282 2592 7288 2644
rect 7340 2632 7346 2644
rect 7558 2632 7564 2644
rect 7340 2604 7564 2632
rect 7340 2592 7346 2604
rect 7558 2592 7564 2604
rect 7616 2592 7622 2644
rect 7837 2635 7895 2641
rect 7837 2601 7849 2635
rect 7883 2632 7895 2635
rect 7926 2632 7932 2644
rect 7883 2604 7932 2632
rect 7883 2601 7895 2604
rect 7837 2595 7895 2601
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 9033 2635 9091 2641
rect 9033 2601 9045 2635
rect 9079 2632 9091 2635
rect 9214 2632 9220 2644
rect 9079 2604 9220 2632
rect 9079 2601 9091 2604
rect 9033 2595 9091 2601
rect 9214 2592 9220 2604
rect 9272 2592 9278 2644
rect 9398 2632 9404 2644
rect 9359 2604 9404 2632
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 9582 2592 9588 2644
rect 9640 2632 9646 2644
rect 10597 2635 10655 2641
rect 10597 2632 10609 2635
rect 9640 2604 10609 2632
rect 9640 2592 9646 2604
rect 10597 2601 10609 2604
rect 10643 2601 10655 2635
rect 10597 2595 10655 2601
rect 12802 2592 12808 2644
rect 12860 2632 12866 2644
rect 15102 2632 15108 2644
rect 12860 2604 15108 2632
rect 12860 2592 12866 2604
rect 15102 2592 15108 2604
rect 15160 2592 15166 2644
rect 4338 2564 4344 2576
rect 3988 2536 4344 2564
rect 2222 2496 2228 2508
rect 2183 2468 2228 2496
rect 2222 2456 2228 2468
rect 2280 2456 2286 2508
rect 3988 2505 4016 2536
rect 4338 2524 4344 2536
rect 4396 2524 4402 2576
rect 4893 2567 4951 2573
rect 4893 2533 4905 2567
rect 4939 2564 4951 2567
rect 7006 2564 7012 2576
rect 4939 2536 7012 2564
rect 4939 2533 4951 2536
rect 4893 2527 4951 2533
rect 7006 2524 7012 2536
rect 7064 2524 7070 2576
rect 8294 2564 8300 2576
rect 7300 2536 8300 2564
rect 2869 2499 2927 2505
rect 2869 2465 2881 2499
rect 2915 2496 2927 2499
rect 3973 2499 4031 2505
rect 2915 2468 3924 2496
rect 2915 2465 2927 2468
rect 2869 2459 2927 2465
rect 1946 2428 1952 2440
rect 1907 2400 1952 2428
rect 1946 2388 1952 2400
rect 2004 2388 2010 2440
rect 3142 2428 3148 2440
rect 3103 2400 3148 2428
rect 3142 2388 3148 2400
rect 3200 2388 3206 2440
rect 3896 2428 3924 2468
rect 3973 2465 3985 2499
rect 4019 2465 4031 2499
rect 3973 2459 4031 2465
rect 4062 2456 4068 2508
rect 4120 2496 4126 2508
rect 4157 2499 4215 2505
rect 4157 2496 4169 2499
rect 4120 2468 4169 2496
rect 4120 2456 4126 2468
rect 4157 2465 4169 2468
rect 4203 2465 4215 2499
rect 5534 2496 5540 2508
rect 5495 2468 5540 2496
rect 4157 2459 4215 2465
rect 5534 2456 5540 2468
rect 5592 2456 5598 2508
rect 7193 2499 7251 2505
rect 5736 2468 7144 2496
rect 4614 2428 4620 2440
rect 3896 2400 4620 2428
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2428 4767 2431
rect 5736 2428 5764 2468
rect 7116 2440 7144 2468
rect 7193 2465 7205 2499
rect 7239 2496 7251 2499
rect 7300 2496 7328 2536
rect 8294 2524 8300 2536
rect 8352 2524 8358 2576
rect 10410 2524 10416 2576
rect 10468 2564 10474 2576
rect 10468 2536 11192 2564
rect 10468 2524 10474 2536
rect 8478 2496 8484 2508
rect 7239 2468 7328 2496
rect 8439 2468 8484 2496
rect 7239 2465 7251 2468
rect 7193 2459 7251 2465
rect 8478 2456 8484 2468
rect 8536 2456 8542 2508
rect 8570 2456 8576 2508
rect 8628 2456 8634 2508
rect 9490 2456 9496 2508
rect 9548 2456 9554 2508
rect 10226 2496 10232 2508
rect 10187 2468 10232 2496
rect 10226 2456 10232 2468
rect 10284 2456 10290 2508
rect 10686 2456 10692 2508
rect 10744 2496 10750 2508
rect 11164 2505 11192 2536
rect 13354 2524 13360 2576
rect 13412 2564 13418 2576
rect 13412 2536 13584 2564
rect 13412 2524 13418 2536
rect 11057 2499 11115 2505
rect 11057 2496 11069 2499
rect 10744 2468 11069 2496
rect 10744 2456 10750 2468
rect 11057 2465 11069 2468
rect 11103 2465 11115 2499
rect 11057 2459 11115 2465
rect 11149 2499 11207 2505
rect 11149 2465 11161 2499
rect 11195 2465 11207 2499
rect 12066 2496 12072 2508
rect 12027 2468 12072 2496
rect 11149 2459 11207 2465
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 12158 2456 12164 2508
rect 12216 2496 12222 2508
rect 12216 2468 12434 2496
rect 12216 2456 12222 2468
rect 4755 2400 5764 2428
rect 5813 2431 5871 2437
rect 4755 2397 4767 2400
rect 4709 2391 4767 2397
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 6730 2428 6736 2440
rect 5859 2400 6736 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 3418 2360 3424 2372
rect 3379 2332 3424 2360
rect 3418 2320 3424 2332
rect 3476 2320 3482 2372
rect 4249 2363 4307 2369
rect 4249 2329 4261 2363
rect 4295 2360 4307 2363
rect 5718 2360 5724 2372
rect 4295 2332 5724 2360
rect 4295 2329 4307 2332
rect 4249 2323 4307 2329
rect 5718 2320 5724 2332
rect 5776 2320 5782 2372
rect 4890 2252 4896 2304
rect 4948 2292 4954 2304
rect 5828 2292 5856 2391
rect 6730 2388 6736 2400
rect 6788 2388 6794 2440
rect 7098 2388 7104 2440
rect 7156 2388 7162 2440
rect 7374 2428 7380 2440
rect 7335 2400 7380 2428
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 7742 2428 7748 2440
rect 7515 2400 7748 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7742 2388 7748 2400
rect 7800 2388 7806 2440
rect 8110 2388 8116 2440
rect 8168 2428 8174 2440
rect 8588 2428 8616 2456
rect 8757 2431 8815 2437
rect 8757 2428 8769 2431
rect 8168 2400 8769 2428
rect 8168 2388 8174 2400
rect 8757 2397 8769 2400
rect 8803 2397 8815 2431
rect 9508 2428 9536 2456
rect 10505 2431 10563 2437
rect 10505 2428 10517 2431
rect 9508 2400 10517 2428
rect 8757 2391 8815 2397
rect 10505 2397 10517 2400
rect 10551 2397 10563 2431
rect 10505 2391 10563 2397
rect 10594 2388 10600 2440
rect 10652 2428 10658 2440
rect 10965 2431 11023 2437
rect 10965 2428 10977 2431
rect 10652 2400 10977 2428
rect 10652 2388 10658 2400
rect 10965 2397 10977 2400
rect 11011 2397 11023 2431
rect 10965 2391 11023 2397
rect 11882 2388 11888 2440
rect 11940 2428 11946 2440
rect 12299 2431 12357 2437
rect 12299 2428 12311 2431
rect 11940 2400 12311 2428
rect 11940 2388 11946 2400
rect 12299 2397 12311 2400
rect 12345 2397 12357 2431
rect 12406 2428 12434 2468
rect 13078 2456 13084 2508
rect 13136 2496 13142 2508
rect 13136 2468 13400 2496
rect 13136 2456 13142 2468
rect 12989 2431 13047 2437
rect 12989 2428 13001 2431
rect 12406 2400 13001 2428
rect 12299 2391 12357 2397
rect 12989 2397 13001 2400
rect 13035 2397 13047 2431
rect 13262 2428 13268 2440
rect 13175 2400 13268 2428
rect 12989 2391 13047 2397
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 13372 2437 13400 2468
rect 13357 2431 13415 2437
rect 13357 2397 13369 2431
rect 13403 2397 13415 2431
rect 13556 2428 13584 2536
rect 13722 2524 13728 2576
rect 13780 2564 13786 2576
rect 14277 2567 14335 2573
rect 14277 2564 14289 2567
rect 13780 2536 14289 2564
rect 13780 2524 13786 2536
rect 14277 2533 14289 2536
rect 14323 2533 14335 2567
rect 14277 2527 14335 2533
rect 13725 2431 13783 2437
rect 13725 2428 13737 2431
rect 13556 2400 13737 2428
rect 13357 2391 13415 2397
rect 13725 2397 13737 2400
rect 13771 2397 13783 2431
rect 13725 2391 13783 2397
rect 13814 2388 13820 2440
rect 13872 2428 13878 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13872 2400 14105 2428
rect 13872 2388 13878 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 14461 2431 14519 2437
rect 14461 2397 14473 2431
rect 14507 2397 14519 2431
rect 14461 2391 14519 2397
rect 15105 2431 15163 2437
rect 15105 2397 15117 2431
rect 15151 2428 15163 2431
rect 15194 2428 15200 2440
rect 15151 2400 15200 2428
rect 15151 2397 15163 2400
rect 15105 2391 15163 2397
rect 6086 2360 6092 2372
rect 6047 2332 6092 2360
rect 6086 2320 6092 2332
rect 6144 2320 6150 2372
rect 6178 2320 6184 2372
rect 6236 2320 6242 2372
rect 6546 2360 6552 2372
rect 6507 2332 6552 2360
rect 6546 2320 6552 2332
rect 6604 2320 6610 2372
rect 6917 2363 6975 2369
rect 6917 2329 6929 2363
rect 6963 2360 6975 2363
rect 7650 2360 7656 2372
rect 6963 2332 7656 2360
rect 6963 2329 6975 2332
rect 6917 2323 6975 2329
rect 7650 2320 7656 2332
rect 7708 2320 7714 2372
rect 8662 2320 8668 2372
rect 8720 2360 8726 2372
rect 9125 2363 9183 2369
rect 9125 2360 9137 2363
rect 8720 2332 9137 2360
rect 8720 2320 8726 2332
rect 9125 2329 9137 2332
rect 9171 2329 9183 2363
rect 9125 2323 9183 2329
rect 9493 2363 9551 2369
rect 9493 2329 9505 2363
rect 9539 2360 9551 2363
rect 10410 2360 10416 2372
rect 9539 2332 10416 2360
rect 9539 2329 9551 2332
rect 9493 2323 9551 2329
rect 10410 2320 10416 2332
rect 10468 2320 10474 2372
rect 12434 2320 12440 2372
rect 12492 2360 12498 2372
rect 13280 2360 13308 2388
rect 14476 2360 14504 2391
rect 15194 2388 15200 2400
rect 15252 2388 15258 2440
rect 15562 2428 15568 2440
rect 15523 2400 15568 2428
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 15746 2428 15752 2440
rect 15707 2400 15752 2428
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 16206 2428 16212 2440
rect 16167 2400 16212 2428
rect 16206 2388 16212 2400
rect 16264 2388 16270 2440
rect 16666 2428 16672 2440
rect 16627 2400 16672 2428
rect 16666 2388 16672 2400
rect 16724 2388 16730 2440
rect 17126 2428 17132 2440
rect 17087 2400 17132 2428
rect 17126 2388 17132 2400
rect 17184 2388 17190 2440
rect 17586 2428 17592 2440
rect 17547 2400 17592 2428
rect 17586 2388 17592 2400
rect 17644 2388 17650 2440
rect 17678 2388 17684 2440
rect 17736 2428 17742 2440
rect 18049 2431 18107 2437
rect 18049 2428 18061 2431
rect 17736 2400 18061 2428
rect 17736 2388 17742 2400
rect 18049 2397 18061 2400
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 18230 2388 18236 2440
rect 18288 2428 18294 2440
rect 18509 2431 18567 2437
rect 18509 2428 18521 2431
rect 18288 2400 18521 2428
rect 18288 2388 18294 2400
rect 18509 2397 18521 2400
rect 18555 2397 18567 2431
rect 18509 2391 18567 2397
rect 19058 2388 19064 2440
rect 19116 2428 19122 2440
rect 19245 2431 19303 2437
rect 19245 2428 19257 2431
rect 19116 2400 19257 2428
rect 19116 2388 19122 2400
rect 19245 2397 19257 2400
rect 19291 2397 19303 2431
rect 19610 2428 19616 2440
rect 19571 2400 19616 2428
rect 19245 2391 19303 2397
rect 19610 2388 19616 2400
rect 19668 2388 19674 2440
rect 19978 2428 19984 2440
rect 19939 2400 19984 2428
rect 19978 2388 19984 2400
rect 20036 2388 20042 2440
rect 20438 2428 20444 2440
rect 20399 2400 20444 2428
rect 20438 2388 20444 2400
rect 20496 2388 20502 2440
rect 20898 2428 20904 2440
rect 20859 2400 20904 2428
rect 20898 2388 20904 2400
rect 20956 2388 20962 2440
rect 20990 2388 20996 2440
rect 21048 2428 21054 2440
rect 21269 2431 21327 2437
rect 21269 2428 21281 2431
rect 21048 2400 21281 2428
rect 21048 2388 21054 2400
rect 21269 2397 21281 2400
rect 21315 2397 21327 2431
rect 21269 2391 21327 2397
rect 12492 2332 13308 2360
rect 13924 2332 14504 2360
rect 12492 2320 12498 2332
rect 4948 2264 5856 2292
rect 5997 2295 6055 2301
rect 4948 2252 4954 2264
rect 5997 2261 6009 2295
rect 6043 2292 6055 2295
rect 6196 2292 6224 2320
rect 8294 2292 8300 2304
rect 6043 2264 8300 2292
rect 6043 2261 6055 2264
rect 5997 2255 6055 2261
rect 8294 2252 8300 2264
rect 8352 2252 8358 2304
rect 13262 2252 13268 2304
rect 13320 2292 13326 2304
rect 13924 2301 13952 2332
rect 13541 2295 13599 2301
rect 13541 2292 13553 2295
rect 13320 2264 13553 2292
rect 13320 2252 13326 2264
rect 13541 2261 13553 2264
rect 13587 2261 13599 2295
rect 13541 2255 13599 2261
rect 13909 2295 13967 2301
rect 13909 2261 13921 2295
rect 13955 2261 13967 2295
rect 13909 2255 13967 2261
rect 14366 2252 14372 2304
rect 14424 2292 14430 2304
rect 14645 2295 14703 2301
rect 14645 2292 14657 2295
rect 14424 2264 14657 2292
rect 14424 2252 14430 2264
rect 14645 2261 14657 2264
rect 14691 2261 14703 2295
rect 14645 2255 14703 2261
rect 14734 2252 14740 2304
rect 14792 2292 14798 2304
rect 14921 2295 14979 2301
rect 14921 2292 14933 2295
rect 14792 2264 14933 2292
rect 14792 2252 14798 2264
rect 14921 2261 14933 2264
rect 14967 2261 14979 2295
rect 14921 2255 14979 2261
rect 15194 2252 15200 2304
rect 15252 2292 15258 2304
rect 15381 2295 15439 2301
rect 15381 2292 15393 2295
rect 15252 2264 15393 2292
rect 15252 2252 15258 2264
rect 15381 2261 15393 2264
rect 15427 2261 15439 2295
rect 15381 2255 15439 2261
rect 15654 2252 15660 2304
rect 15712 2292 15718 2304
rect 15933 2295 15991 2301
rect 15933 2292 15945 2295
rect 15712 2264 15945 2292
rect 15712 2252 15718 2264
rect 15933 2261 15945 2264
rect 15979 2261 15991 2295
rect 15933 2255 15991 2261
rect 16114 2252 16120 2304
rect 16172 2292 16178 2304
rect 16393 2295 16451 2301
rect 16393 2292 16405 2295
rect 16172 2264 16405 2292
rect 16172 2252 16178 2264
rect 16393 2261 16405 2264
rect 16439 2261 16451 2295
rect 16393 2255 16451 2261
rect 16853 2295 16911 2301
rect 16853 2261 16865 2295
rect 16899 2292 16911 2295
rect 16942 2292 16948 2304
rect 16899 2264 16948 2292
rect 16899 2261 16911 2264
rect 16853 2255 16911 2261
rect 16942 2252 16948 2264
rect 17000 2252 17006 2304
rect 17034 2252 17040 2304
rect 17092 2292 17098 2304
rect 17313 2295 17371 2301
rect 17313 2292 17325 2295
rect 17092 2264 17325 2292
rect 17092 2252 17098 2264
rect 17313 2261 17325 2264
rect 17359 2261 17371 2295
rect 17313 2255 17371 2261
rect 17494 2252 17500 2304
rect 17552 2292 17558 2304
rect 17773 2295 17831 2301
rect 17773 2292 17785 2295
rect 17552 2264 17785 2292
rect 17552 2252 17558 2264
rect 17773 2261 17785 2264
rect 17819 2261 17831 2295
rect 17773 2255 17831 2261
rect 17954 2252 17960 2304
rect 18012 2292 18018 2304
rect 18233 2295 18291 2301
rect 18233 2292 18245 2295
rect 18012 2264 18245 2292
rect 18012 2252 18018 2264
rect 18233 2261 18245 2264
rect 18279 2261 18291 2295
rect 18233 2255 18291 2261
rect 18414 2252 18420 2304
rect 18472 2292 18478 2304
rect 18693 2295 18751 2301
rect 18693 2292 18705 2295
rect 18472 2264 18705 2292
rect 18472 2252 18478 2264
rect 18693 2261 18705 2264
rect 18739 2261 18751 2295
rect 18693 2255 18751 2261
rect 18966 2252 18972 2304
rect 19024 2292 19030 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 19024 2264 19441 2292
rect 19024 2252 19030 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 19429 2255 19487 2261
rect 19518 2252 19524 2304
rect 19576 2292 19582 2304
rect 19797 2295 19855 2301
rect 19797 2292 19809 2295
rect 19576 2264 19809 2292
rect 19576 2252 19582 2264
rect 19797 2261 19809 2264
rect 19843 2261 19855 2295
rect 19797 2255 19855 2261
rect 19886 2252 19892 2304
rect 19944 2292 19950 2304
rect 20165 2295 20223 2301
rect 20165 2292 20177 2295
rect 19944 2264 20177 2292
rect 19944 2252 19950 2264
rect 20165 2261 20177 2264
rect 20211 2261 20223 2295
rect 20165 2255 20223 2261
rect 20346 2252 20352 2304
rect 20404 2292 20410 2304
rect 20625 2295 20683 2301
rect 20625 2292 20637 2295
rect 20404 2264 20637 2292
rect 20404 2252 20410 2264
rect 20625 2261 20637 2264
rect 20671 2261 20683 2295
rect 20625 2255 20683 2261
rect 20806 2252 20812 2304
rect 20864 2292 20870 2304
rect 21085 2295 21143 2301
rect 21085 2292 21097 2295
rect 20864 2264 21097 2292
rect 20864 2252 20870 2264
rect 21085 2261 21097 2264
rect 21131 2261 21143 2295
rect 21085 2255 21143 2261
rect 21266 2252 21272 2304
rect 21324 2292 21330 2304
rect 21453 2295 21511 2301
rect 21453 2292 21465 2295
rect 21324 2264 21465 2292
rect 21324 2252 21330 2264
rect 21453 2261 21465 2264
rect 21499 2261 21511 2295
rect 21453 2255 21511 2261
rect 1104 2202 21896 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21896 2202
rect 1104 2128 21896 2150
rect 3234 2048 3240 2100
rect 3292 2088 3298 2100
rect 6638 2088 6644 2100
rect 3292 2060 6644 2088
rect 3292 2048 3298 2060
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 6730 2048 6736 2100
rect 6788 2088 6794 2100
rect 14826 2088 14832 2100
rect 6788 2060 14832 2088
rect 6788 2048 6794 2060
rect 14826 2048 14832 2060
rect 14884 2048 14890 2100
rect 1946 1980 1952 2032
rect 2004 2020 2010 2032
rect 7834 2020 7840 2032
rect 2004 1992 7840 2020
rect 2004 1980 2010 1992
rect 7834 1980 7840 1992
rect 7892 1980 7898 2032
rect 7650 1844 7656 1896
rect 7708 1884 7714 1896
rect 8202 1884 8208 1896
rect 7708 1856 8208 1884
rect 7708 1844 7714 1856
rect 8202 1844 8208 1856
rect 8260 1844 8266 1896
rect 8294 1844 8300 1896
rect 8352 1884 8358 1896
rect 12894 1884 12900 1896
rect 8352 1856 12900 1884
rect 8352 1844 8358 1856
rect 12894 1844 12900 1856
rect 12952 1844 12958 1896
rect 5902 1776 5908 1828
rect 5960 1816 5966 1828
rect 6822 1816 6828 1828
rect 5960 1788 6828 1816
rect 5960 1776 5966 1788
rect 6822 1776 6828 1788
rect 6880 1816 6886 1828
rect 15286 1816 15292 1828
rect 6880 1788 15292 1816
rect 6880 1776 6886 1788
rect 15286 1776 15292 1788
rect 15344 1776 15350 1828
rect 1578 1708 1584 1760
rect 1636 1748 1642 1760
rect 14642 1748 14648 1760
rect 1636 1720 14648 1748
rect 1636 1708 1642 1720
rect 14642 1708 14648 1720
rect 14700 1708 14706 1760
rect 6546 1640 6552 1692
rect 6604 1680 6610 1692
rect 6730 1680 6736 1692
rect 6604 1652 6736 1680
rect 6604 1640 6610 1652
rect 6730 1640 6736 1652
rect 6788 1680 6794 1692
rect 14918 1680 14924 1692
rect 6788 1652 14924 1680
rect 6788 1640 6794 1652
rect 14918 1640 14924 1652
rect 14976 1640 14982 1692
rect 3510 1572 3516 1624
rect 3568 1612 3574 1624
rect 14182 1612 14188 1624
rect 3568 1584 14188 1612
rect 3568 1572 3574 1584
rect 14182 1572 14188 1584
rect 14240 1572 14246 1624
rect 4062 1028 4068 1080
rect 4120 1068 4126 1080
rect 6914 1068 6920 1080
rect 4120 1040 6920 1068
rect 4120 1028 4126 1040
rect 6914 1028 6920 1040
rect 6972 1028 6978 1080
<< via1 >>
rect 10232 20748 10284 20800
rect 11244 20748 11296 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 3056 20544 3108 20596
rect 4620 20544 4672 20596
rect 4896 20544 4948 20596
rect 6644 20544 6696 20596
rect 7564 20544 7616 20596
rect 9312 20544 9364 20596
rect 5172 20476 5224 20528
rect 10232 20544 10284 20596
rect 12900 20544 12952 20596
rect 13084 20544 13136 20596
rect 13544 20544 13596 20596
rect 14004 20544 14056 20596
rect 14464 20544 14516 20596
rect 15200 20587 15252 20596
rect 15200 20553 15209 20587
rect 15209 20553 15243 20587
rect 15243 20553 15252 20587
rect 15200 20544 15252 20553
rect 15384 20544 15436 20596
rect 15844 20544 15896 20596
rect 16304 20544 16356 20596
rect 17224 20544 17276 20596
rect 17960 20587 18012 20596
rect 17960 20553 17969 20587
rect 17969 20553 18003 20587
rect 18003 20553 18012 20587
rect 17960 20544 18012 20553
rect 18144 20544 18196 20596
rect 18604 20544 18656 20596
rect 19340 20544 19392 20596
rect 19524 20544 19576 20596
rect 19984 20544 20036 20596
rect 20444 20544 20496 20596
rect 20904 20544 20956 20596
rect 11244 20476 11296 20528
rect 2044 20451 2096 20460
rect 2044 20417 2053 20451
rect 2053 20417 2087 20451
rect 2087 20417 2096 20451
rect 2044 20408 2096 20417
rect 2136 20408 2188 20460
rect 3516 20451 3568 20460
rect 3516 20417 3525 20451
rect 3525 20417 3559 20451
rect 3559 20417 3568 20451
rect 3516 20408 3568 20417
rect 2688 20383 2740 20392
rect 2688 20349 2697 20383
rect 2697 20349 2731 20383
rect 2731 20349 2740 20383
rect 2688 20340 2740 20349
rect 4160 20340 4212 20392
rect 4620 20383 4672 20392
rect 4620 20349 4629 20383
rect 4629 20349 4663 20383
rect 4663 20349 4672 20383
rect 4620 20340 4672 20349
rect 4896 20451 4948 20460
rect 4896 20417 4905 20451
rect 4905 20417 4939 20451
rect 4939 20417 4948 20451
rect 5448 20451 5500 20460
rect 4896 20408 4948 20417
rect 5448 20417 5457 20451
rect 5457 20417 5491 20451
rect 5491 20417 5500 20451
rect 5448 20408 5500 20417
rect 6368 20451 6420 20460
rect 5172 20340 5224 20392
rect 5540 20383 5592 20392
rect 5540 20349 5549 20383
rect 5549 20349 5583 20383
rect 5583 20349 5592 20383
rect 5540 20340 5592 20349
rect 5632 20383 5684 20392
rect 5632 20349 5641 20383
rect 5641 20349 5675 20383
rect 5675 20349 5684 20383
rect 6368 20417 6377 20451
rect 6377 20417 6411 20451
rect 6411 20417 6420 20451
rect 6368 20408 6420 20417
rect 7104 20408 7156 20460
rect 9404 20408 9456 20460
rect 10140 20408 10192 20460
rect 5632 20340 5684 20349
rect 7564 20340 7616 20392
rect 8300 20340 8352 20392
rect 1308 20204 1360 20256
rect 5908 20272 5960 20324
rect 8668 20272 8720 20324
rect 9312 20340 9364 20392
rect 10048 20340 10100 20392
rect 10416 20383 10468 20392
rect 10416 20349 10425 20383
rect 10425 20349 10459 20383
rect 10459 20349 10468 20383
rect 10416 20340 10468 20349
rect 10600 20340 10652 20392
rect 9680 20272 9732 20324
rect 10876 20272 10928 20324
rect 3976 20204 4028 20256
rect 4804 20247 4856 20256
rect 4804 20213 4813 20247
rect 4813 20213 4847 20247
rect 4847 20213 4856 20247
rect 4804 20204 4856 20213
rect 5816 20204 5868 20256
rect 7840 20247 7892 20256
rect 7840 20213 7849 20247
rect 7849 20213 7883 20247
rect 7883 20213 7892 20247
rect 7840 20204 7892 20213
rect 9312 20204 9364 20256
rect 9404 20204 9456 20256
rect 10048 20204 10100 20256
rect 11152 20340 11204 20392
rect 12440 20408 12492 20460
rect 13268 20408 13320 20460
rect 13544 20408 13596 20460
rect 13636 20451 13688 20460
rect 13636 20417 13645 20451
rect 13645 20417 13679 20451
rect 13679 20417 13688 20451
rect 13636 20408 13688 20417
rect 13820 20408 13872 20460
rect 14280 20408 14332 20460
rect 14832 20408 14884 20460
rect 15108 20408 15160 20460
rect 15936 20451 15988 20460
rect 15936 20417 15945 20451
rect 15945 20417 15979 20451
rect 15979 20417 15988 20451
rect 15936 20408 15988 20417
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 17040 20451 17092 20460
rect 17040 20417 17049 20451
rect 17049 20417 17083 20451
rect 17083 20417 17092 20451
rect 17040 20408 17092 20417
rect 17132 20408 17184 20460
rect 17684 20408 17736 20460
rect 17960 20408 18012 20460
rect 18328 20408 18380 20460
rect 18788 20408 18840 20460
rect 19708 20408 19760 20460
rect 20536 20451 20588 20460
rect 20536 20417 20545 20451
rect 20545 20417 20579 20451
rect 20579 20417 20588 20451
rect 20536 20408 20588 20417
rect 11060 20272 11112 20324
rect 12440 20272 12492 20324
rect 13452 20272 13504 20324
rect 14372 20272 14424 20324
rect 11888 20204 11940 20256
rect 16948 20272 17000 20324
rect 18420 20272 18472 20324
rect 21180 20408 21232 20460
rect 22744 20408 22796 20460
rect 20904 20204 20956 20256
rect 21364 20247 21416 20256
rect 21364 20213 21373 20247
rect 21373 20213 21407 20247
rect 21407 20213 21416 20247
rect 21364 20204 21416 20213
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 1124 19864 1176 19916
rect 1768 19864 1820 19916
rect 1952 19839 2004 19848
rect 1952 19805 1961 19839
rect 1961 19805 1995 19839
rect 1995 19805 2004 19839
rect 1952 19796 2004 19805
rect 3240 19796 3292 19848
rect 3516 19839 3568 19848
rect 3516 19805 3525 19839
rect 3525 19805 3559 19839
rect 3559 19805 3568 19839
rect 3516 19796 3568 19805
rect 5540 20000 5592 20052
rect 10140 20000 10192 20052
rect 10692 20000 10744 20052
rect 10416 19932 10468 19984
rect 11152 20000 11204 20052
rect 11704 20000 11756 20052
rect 13544 20043 13596 20052
rect 3700 19660 3752 19712
rect 3976 19660 4028 19712
rect 4160 19728 4212 19780
rect 4528 19728 4580 19780
rect 5356 19660 5408 19712
rect 6368 19864 6420 19916
rect 7104 19907 7156 19916
rect 7104 19873 7113 19907
rect 7113 19873 7147 19907
rect 7147 19873 7156 19907
rect 7104 19864 7156 19873
rect 6000 19796 6052 19848
rect 6828 19839 6880 19848
rect 6828 19805 6837 19839
rect 6837 19805 6871 19839
rect 6871 19805 6880 19839
rect 6828 19796 6880 19805
rect 8668 19796 8720 19848
rect 11060 19864 11112 19916
rect 13544 20009 13553 20043
rect 13553 20009 13587 20043
rect 13587 20009 13596 20043
rect 13544 20000 13596 20009
rect 14280 20043 14332 20052
rect 14280 20009 14289 20043
rect 14289 20009 14323 20043
rect 14323 20009 14332 20043
rect 14280 20000 14332 20009
rect 14832 20043 14884 20052
rect 14832 20009 14841 20043
rect 14841 20009 14875 20043
rect 14875 20009 14884 20043
rect 14832 20000 14884 20009
rect 15108 20043 15160 20052
rect 15108 20009 15117 20043
rect 15117 20009 15151 20043
rect 15151 20009 15160 20043
rect 15108 20000 15160 20009
rect 15936 20000 15988 20052
rect 17040 20000 17092 20052
rect 17684 20043 17736 20052
rect 17684 20009 17693 20043
rect 17693 20009 17727 20043
rect 17727 20009 17736 20043
rect 17684 20000 17736 20009
rect 17960 20043 18012 20052
rect 17960 20009 17969 20043
rect 17969 20009 18003 20043
rect 18003 20009 18012 20043
rect 17960 20000 18012 20009
rect 18328 20000 18380 20052
rect 18788 20000 18840 20052
rect 19708 20000 19760 20052
rect 20536 20000 20588 20052
rect 21180 20000 21232 20052
rect 21456 20043 21508 20052
rect 21456 20009 21465 20043
rect 21465 20009 21499 20043
rect 21499 20009 21508 20043
rect 21456 20000 21508 20009
rect 14372 19932 14424 19984
rect 16672 19932 16724 19984
rect 21824 19932 21876 19984
rect 12348 19839 12400 19848
rect 12348 19805 12357 19839
rect 12357 19805 12391 19839
rect 12391 19805 12400 19839
rect 12348 19796 12400 19805
rect 12532 19796 12584 19848
rect 13360 19839 13412 19848
rect 13360 19805 13369 19839
rect 13369 19805 13403 19839
rect 13403 19805 13412 19839
rect 13360 19796 13412 19805
rect 13728 19796 13780 19848
rect 14280 19796 14332 19848
rect 14372 19839 14424 19848
rect 14372 19805 14381 19839
rect 14381 19805 14415 19839
rect 14415 19805 14424 19839
rect 14372 19796 14424 19805
rect 14740 19796 14792 19848
rect 5540 19728 5592 19780
rect 9220 19728 9272 19780
rect 9864 19728 9916 19780
rect 10968 19728 11020 19780
rect 12624 19728 12676 19780
rect 13544 19728 13596 19780
rect 15292 19796 15344 19848
rect 15384 19796 15436 19848
rect 15936 19839 15988 19848
rect 15936 19805 15945 19839
rect 15945 19805 15979 19839
rect 15979 19805 15988 19839
rect 15936 19796 15988 19805
rect 17408 19839 17460 19848
rect 17408 19805 17417 19839
rect 17417 19805 17451 19839
rect 17451 19805 17460 19839
rect 17408 19796 17460 19805
rect 17500 19839 17552 19848
rect 17500 19805 17509 19839
rect 17509 19805 17543 19839
rect 17543 19805 17552 19839
rect 17776 19839 17828 19848
rect 17500 19796 17552 19805
rect 17776 19805 17785 19839
rect 17785 19805 17819 19839
rect 17819 19805 17828 19839
rect 17776 19796 17828 19805
rect 6828 19660 6880 19712
rect 7380 19660 7432 19712
rect 8116 19703 8168 19712
rect 8116 19669 8125 19703
rect 8125 19669 8159 19703
rect 8159 19669 8168 19703
rect 8116 19660 8168 19669
rect 9496 19660 9548 19712
rect 10140 19660 10192 19712
rect 16580 19771 16632 19780
rect 16580 19737 16589 19771
rect 16589 19737 16623 19771
rect 16623 19737 16632 19771
rect 16580 19728 16632 19737
rect 16948 19728 17000 19780
rect 19064 19796 19116 19848
rect 19616 19839 19668 19848
rect 19616 19805 19625 19839
rect 19625 19805 19659 19839
rect 19659 19805 19668 19839
rect 19616 19796 19668 19805
rect 20904 19839 20956 19848
rect 20904 19805 20913 19839
rect 20913 19805 20947 19839
rect 20947 19805 20956 19839
rect 20904 19796 20956 19805
rect 16304 19660 16356 19712
rect 18420 19660 18472 19712
rect 18604 19703 18656 19712
rect 18604 19669 18613 19703
rect 18613 19669 18647 19703
rect 18647 19669 18656 19703
rect 18604 19660 18656 19669
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 2412 19456 2464 19508
rect 1400 19388 1452 19440
rect 2504 19388 2556 19440
rect 2044 19320 2096 19372
rect 4160 19388 4212 19440
rect 4436 19456 4488 19508
rect 4528 19456 4580 19508
rect 5632 19456 5684 19508
rect 7104 19499 7156 19508
rect 204 19252 256 19304
rect 2228 19295 2280 19304
rect 2228 19261 2237 19295
rect 2237 19261 2271 19295
rect 2271 19261 2280 19295
rect 2228 19252 2280 19261
rect 4436 19320 4488 19372
rect 5540 19320 5592 19372
rect 5908 19363 5960 19372
rect 7104 19465 7113 19499
rect 7113 19465 7147 19499
rect 7147 19465 7156 19499
rect 7104 19456 7156 19465
rect 8668 19499 8720 19508
rect 8668 19465 8677 19499
rect 8677 19465 8711 19499
rect 8711 19465 8720 19499
rect 8668 19456 8720 19465
rect 9864 19456 9916 19508
rect 10508 19456 10560 19508
rect 8116 19388 8168 19440
rect 9312 19388 9364 19440
rect 10048 19388 10100 19440
rect 10324 19388 10376 19440
rect 12440 19388 12492 19440
rect 12900 19456 12952 19508
rect 13452 19456 13504 19508
rect 13636 19456 13688 19508
rect 14372 19499 14424 19508
rect 14372 19465 14381 19499
rect 14381 19465 14415 19499
rect 14415 19465 14424 19499
rect 14372 19456 14424 19465
rect 14740 19499 14792 19508
rect 14740 19465 14749 19499
rect 14749 19465 14783 19499
rect 14783 19465 14792 19499
rect 14740 19456 14792 19465
rect 15936 19456 15988 19508
rect 16304 19456 16356 19508
rect 16948 19456 17000 19508
rect 17132 19499 17184 19508
rect 17132 19465 17141 19499
rect 17141 19465 17175 19499
rect 17175 19465 17184 19499
rect 17132 19456 17184 19465
rect 19616 19456 19668 19508
rect 5908 19329 5926 19363
rect 5926 19329 5960 19363
rect 5908 19320 5960 19329
rect 6460 19320 6512 19372
rect 10508 19320 10560 19372
rect 12072 19363 12124 19372
rect 12072 19329 12081 19363
rect 12081 19329 12115 19363
rect 12115 19329 12124 19363
rect 12072 19320 12124 19329
rect 6552 19252 6604 19304
rect 8484 19295 8536 19304
rect 8484 19261 8493 19295
rect 8493 19261 8527 19295
rect 8527 19261 8536 19295
rect 8484 19252 8536 19261
rect 10324 19252 10376 19304
rect 10416 19252 10468 19304
rect 11060 19252 11112 19304
rect 11980 19252 12032 19304
rect 12256 19295 12308 19304
rect 12256 19261 12265 19295
rect 12265 19261 12299 19295
rect 12299 19261 12308 19295
rect 12256 19252 12308 19261
rect 3148 19184 3200 19236
rect 6184 19184 6236 19236
rect 2964 19116 3016 19168
rect 5448 19116 5500 19168
rect 5540 19116 5592 19168
rect 6828 19116 6880 19168
rect 10692 19116 10744 19168
rect 10876 19184 10928 19236
rect 12164 19184 12216 19236
rect 12716 19320 12768 19372
rect 12808 19320 12860 19372
rect 13084 19363 13136 19372
rect 13084 19329 13093 19363
rect 13093 19329 13127 19363
rect 13127 19329 13136 19363
rect 13084 19320 13136 19329
rect 14740 19320 14792 19372
rect 15016 19363 15068 19372
rect 15016 19329 15025 19363
rect 15025 19329 15059 19363
rect 15059 19329 15068 19363
rect 15016 19320 15068 19329
rect 17040 19388 17092 19440
rect 13728 19184 13780 19236
rect 11704 19116 11756 19168
rect 12440 19116 12492 19168
rect 12900 19116 12952 19168
rect 12992 19116 13044 19168
rect 15476 19227 15528 19236
rect 15476 19193 15485 19227
rect 15485 19193 15519 19227
rect 15519 19193 15528 19227
rect 15476 19184 15528 19193
rect 14280 19159 14332 19168
rect 14280 19125 14289 19159
rect 14289 19125 14323 19159
rect 14323 19125 14332 19159
rect 14280 19116 14332 19125
rect 15292 19159 15344 19168
rect 15292 19125 15301 19159
rect 15301 19125 15335 19159
rect 15335 19125 15344 19159
rect 15660 19159 15712 19168
rect 15292 19116 15344 19125
rect 15660 19125 15669 19159
rect 15669 19125 15703 19159
rect 15703 19125 15712 19159
rect 15660 19116 15712 19125
rect 15752 19116 15804 19168
rect 17224 19320 17276 19372
rect 18512 19320 18564 19372
rect 17408 19252 17460 19304
rect 22284 19252 22336 19304
rect 17224 19159 17276 19168
rect 17224 19125 17233 19159
rect 17233 19125 17267 19159
rect 17267 19125 17276 19159
rect 17408 19159 17460 19168
rect 17224 19116 17276 19125
rect 17408 19125 17417 19159
rect 17417 19125 17451 19159
rect 17451 19125 17460 19159
rect 17408 19116 17460 19125
rect 17776 19159 17828 19168
rect 17776 19125 17785 19159
rect 17785 19125 17819 19159
rect 17819 19125 17828 19159
rect 17776 19116 17828 19125
rect 18512 19159 18564 19168
rect 18512 19125 18521 19159
rect 18521 19125 18555 19159
rect 18555 19125 18564 19159
rect 18512 19116 18564 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 1492 18955 1544 18964
rect 1492 18921 1501 18955
rect 1501 18921 1535 18955
rect 1535 18921 1544 18955
rect 1492 18912 1544 18921
rect 3148 18912 3200 18964
rect 2780 18844 2832 18896
rect 6736 18912 6788 18964
rect 10232 18912 10284 18964
rect 10324 18912 10376 18964
rect 10508 18887 10560 18896
rect 3332 18819 3384 18828
rect 1584 18708 1636 18760
rect 3332 18785 3341 18819
rect 3341 18785 3375 18819
rect 3375 18785 3384 18819
rect 3332 18776 3384 18785
rect 2780 18751 2832 18760
rect 2780 18717 2789 18751
rect 2789 18717 2823 18751
rect 2823 18717 2832 18751
rect 2780 18708 2832 18717
rect 4988 18708 5040 18760
rect 2228 18640 2280 18692
rect 4712 18683 4764 18692
rect 3148 18572 3200 18624
rect 3332 18572 3384 18624
rect 4712 18649 4721 18683
rect 4721 18649 4755 18683
rect 4755 18649 4764 18683
rect 4712 18640 4764 18649
rect 4160 18615 4212 18624
rect 4160 18581 4169 18615
rect 4169 18581 4203 18615
rect 4203 18581 4212 18615
rect 4160 18572 4212 18581
rect 4436 18572 4488 18624
rect 5080 18572 5132 18624
rect 10508 18853 10517 18887
rect 10517 18853 10551 18887
rect 10551 18853 10560 18887
rect 10508 18844 10560 18853
rect 6552 18819 6604 18828
rect 6552 18785 6561 18819
rect 6561 18785 6595 18819
rect 6595 18785 6604 18819
rect 9404 18819 9456 18828
rect 6552 18776 6604 18785
rect 6460 18708 6512 18760
rect 6644 18708 6696 18760
rect 9404 18785 9413 18819
rect 9413 18785 9447 18819
rect 9447 18785 9456 18819
rect 9404 18776 9456 18785
rect 9496 18819 9548 18828
rect 9496 18785 9505 18819
rect 9505 18785 9539 18819
rect 9539 18785 9548 18819
rect 11244 18912 11296 18964
rect 12348 18912 12400 18964
rect 12624 18912 12676 18964
rect 13360 18912 13412 18964
rect 13636 18912 13688 18964
rect 14648 18955 14700 18964
rect 14648 18921 14657 18955
rect 14657 18921 14691 18955
rect 14691 18921 14700 18955
rect 14648 18912 14700 18921
rect 11980 18887 12032 18896
rect 11980 18853 11989 18887
rect 11989 18853 12023 18887
rect 12023 18853 12032 18887
rect 11980 18844 12032 18853
rect 12808 18844 12860 18896
rect 13268 18844 13320 18896
rect 13912 18844 13964 18896
rect 9496 18776 9548 18785
rect 8484 18708 8536 18760
rect 8576 18708 8628 18760
rect 6552 18640 6604 18692
rect 7012 18640 7064 18692
rect 7840 18640 7892 18692
rect 8116 18572 8168 18624
rect 9404 18640 9456 18692
rect 11612 18776 11664 18828
rect 11980 18708 12032 18760
rect 12164 18708 12216 18760
rect 12808 18751 12860 18760
rect 8944 18615 8996 18624
rect 8944 18581 8953 18615
rect 8953 18581 8987 18615
rect 8987 18581 8996 18615
rect 8944 18572 8996 18581
rect 9312 18615 9364 18624
rect 9312 18581 9321 18615
rect 9321 18581 9355 18615
rect 9355 18581 9364 18615
rect 9312 18572 9364 18581
rect 9956 18572 10008 18624
rect 11152 18572 11204 18624
rect 12256 18572 12308 18624
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 12900 18708 12952 18760
rect 12624 18640 12676 18692
rect 14832 18683 14884 18692
rect 14832 18649 14841 18683
rect 14841 18649 14875 18683
rect 14875 18649 14884 18683
rect 14832 18640 14884 18649
rect 17960 18640 18012 18692
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 2320 18368 2372 18420
rect 2780 18411 2832 18420
rect 2780 18377 2789 18411
rect 2789 18377 2823 18411
rect 2823 18377 2832 18411
rect 2780 18368 2832 18377
rect 2872 18300 2924 18352
rect 1952 18232 2004 18284
rect 2320 18232 2372 18284
rect 2688 18232 2740 18284
rect 2780 18232 2832 18284
rect 3792 18368 3844 18420
rect 4252 18368 4304 18420
rect 4436 18411 4488 18420
rect 4436 18377 4445 18411
rect 4445 18377 4479 18411
rect 4479 18377 4488 18411
rect 4436 18368 4488 18377
rect 6000 18368 6052 18420
rect 6828 18368 6880 18420
rect 8300 18368 8352 18420
rect 9312 18368 9364 18420
rect 9588 18368 9640 18420
rect 9680 18368 9732 18420
rect 11152 18411 11204 18420
rect 11152 18377 11161 18411
rect 11161 18377 11195 18411
rect 11195 18377 11204 18411
rect 11152 18368 11204 18377
rect 12164 18368 12216 18420
rect 11612 18300 11664 18352
rect 14464 18368 14516 18420
rect 12348 18300 12400 18352
rect 3424 18232 3476 18284
rect 4528 18232 4580 18284
rect 4804 18275 4856 18284
rect 4804 18241 4813 18275
rect 4813 18241 4847 18275
rect 4847 18241 4856 18275
rect 4804 18232 4856 18241
rect 6552 18275 6604 18284
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 2320 18028 2372 18080
rect 2504 18028 2556 18080
rect 2688 18071 2740 18080
rect 2688 18037 2697 18071
rect 2697 18037 2731 18071
rect 2731 18037 2740 18071
rect 2688 18028 2740 18037
rect 4896 18164 4948 18216
rect 5080 18207 5132 18216
rect 5080 18173 5089 18207
rect 5089 18173 5123 18207
rect 5123 18173 5132 18207
rect 5080 18164 5132 18173
rect 5632 18164 5684 18216
rect 6552 18241 6561 18275
rect 6561 18241 6595 18275
rect 6595 18241 6604 18275
rect 6552 18232 6604 18241
rect 6828 18232 6880 18284
rect 8116 18275 8168 18284
rect 8116 18241 8125 18275
rect 8125 18241 8159 18275
rect 8159 18241 8168 18275
rect 8116 18232 8168 18241
rect 8944 18232 8996 18284
rect 9128 18275 9180 18284
rect 9128 18241 9137 18275
rect 9137 18241 9171 18275
rect 9171 18241 9180 18275
rect 9128 18232 9180 18241
rect 9772 18275 9824 18284
rect 6920 18207 6972 18216
rect 6920 18173 6929 18207
rect 6929 18173 6963 18207
rect 6963 18173 6972 18207
rect 6920 18164 6972 18173
rect 9772 18241 9781 18275
rect 9781 18241 9815 18275
rect 9815 18241 9824 18275
rect 9772 18232 9824 18241
rect 10692 18275 10744 18284
rect 10692 18241 10701 18275
rect 10701 18241 10735 18275
rect 10735 18241 10744 18275
rect 10692 18232 10744 18241
rect 11704 18275 11756 18284
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 7012 18096 7064 18148
rect 4620 18028 4672 18080
rect 4896 18028 4948 18080
rect 9220 18139 9272 18148
rect 7196 18028 7248 18080
rect 9220 18105 9229 18139
rect 9229 18105 9263 18139
rect 9263 18105 9272 18139
rect 9220 18096 9272 18105
rect 10600 18164 10652 18216
rect 11060 18164 11112 18216
rect 12624 18232 12676 18284
rect 13084 18232 13136 18284
rect 13268 18300 13320 18352
rect 13452 18275 13504 18284
rect 13452 18241 13461 18275
rect 13461 18241 13495 18275
rect 13495 18241 13504 18275
rect 13452 18232 13504 18241
rect 10416 18071 10468 18080
rect 10416 18037 10425 18071
rect 10425 18037 10459 18071
rect 10459 18037 10468 18071
rect 10416 18028 10468 18037
rect 10508 18071 10560 18080
rect 10508 18037 10517 18071
rect 10517 18037 10551 18071
rect 10551 18037 10560 18071
rect 10508 18028 10560 18037
rect 10968 18028 11020 18080
rect 14832 18028 14884 18080
rect 17776 18028 17828 18080
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 1860 17867 1912 17876
rect 1860 17833 1869 17867
rect 1869 17833 1903 17867
rect 1903 17833 1912 17867
rect 1860 17824 1912 17833
rect 2228 17867 2280 17876
rect 2228 17833 2237 17867
rect 2237 17833 2271 17867
rect 2271 17833 2280 17867
rect 2228 17824 2280 17833
rect 2596 17867 2648 17876
rect 2596 17833 2605 17867
rect 2605 17833 2639 17867
rect 2639 17833 2648 17867
rect 2596 17824 2648 17833
rect 3056 17867 3108 17876
rect 3056 17833 3065 17867
rect 3065 17833 3099 17867
rect 3099 17833 3108 17867
rect 3056 17824 3108 17833
rect 3424 17867 3476 17876
rect 3424 17833 3433 17867
rect 3433 17833 3467 17867
rect 3467 17833 3476 17867
rect 3424 17824 3476 17833
rect 4068 17824 4120 17876
rect 10784 17824 10836 17876
rect 12992 17824 13044 17876
rect 13084 17824 13136 17876
rect 13820 17867 13872 17876
rect 13820 17833 13829 17867
rect 13829 17833 13863 17867
rect 13863 17833 13872 17867
rect 13820 17824 13872 17833
rect 4804 17756 4856 17808
rect 5540 17688 5592 17740
rect 6644 17688 6696 17740
rect 1676 17663 1728 17672
rect 1676 17629 1685 17663
rect 1685 17629 1719 17663
rect 1719 17629 1728 17663
rect 1676 17620 1728 17629
rect 2228 17620 2280 17672
rect 2596 17620 2648 17672
rect 2872 17663 2924 17672
rect 2872 17629 2881 17663
rect 2881 17629 2915 17663
rect 2915 17629 2924 17663
rect 3240 17663 3292 17672
rect 2872 17620 2924 17629
rect 3240 17629 3249 17663
rect 3249 17629 3283 17663
rect 3283 17629 3292 17663
rect 3240 17620 3292 17629
rect 4528 17620 4580 17672
rect 5264 17663 5316 17672
rect 5264 17629 5273 17663
rect 5273 17629 5307 17663
rect 5307 17629 5316 17663
rect 5264 17620 5316 17629
rect 7196 17663 7248 17672
rect 3056 17552 3108 17604
rect 3148 17552 3200 17604
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 7472 17731 7524 17740
rect 7472 17697 7481 17731
rect 7481 17697 7515 17731
rect 7515 17697 7524 17731
rect 7472 17688 7524 17697
rect 7564 17688 7616 17740
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 5080 17484 5132 17536
rect 5540 17484 5592 17536
rect 6644 17527 6696 17536
rect 6644 17493 6653 17527
rect 6653 17493 6687 17527
rect 6687 17493 6696 17527
rect 6644 17484 6696 17493
rect 6736 17484 6788 17536
rect 7012 17484 7064 17536
rect 7564 17484 7616 17536
rect 10048 17756 10100 17808
rect 10876 17756 10928 17808
rect 9036 17731 9088 17740
rect 9036 17697 9045 17731
rect 9045 17697 9079 17731
rect 9079 17697 9088 17731
rect 9036 17688 9088 17697
rect 9680 17688 9732 17740
rect 10784 17688 10836 17740
rect 10232 17663 10284 17672
rect 10232 17629 10241 17663
rect 10241 17629 10275 17663
rect 10275 17629 10284 17663
rect 10232 17620 10284 17629
rect 8484 17552 8536 17604
rect 11244 17620 11296 17672
rect 9404 17484 9456 17536
rect 10048 17527 10100 17536
rect 10048 17493 10057 17527
rect 10057 17493 10091 17527
rect 10091 17493 10100 17527
rect 10048 17484 10100 17493
rect 10784 17527 10836 17536
rect 10784 17493 10793 17527
rect 10793 17493 10827 17527
rect 10827 17493 10836 17527
rect 11704 17552 11756 17604
rect 10784 17484 10836 17493
rect 11152 17484 11204 17536
rect 13360 17620 13412 17672
rect 12624 17484 12676 17536
rect 21088 17527 21140 17536
rect 21088 17493 21097 17527
rect 21097 17493 21131 17527
rect 21131 17493 21140 17527
rect 21088 17484 21140 17493
rect 21456 17527 21508 17536
rect 21456 17493 21465 17527
rect 21465 17493 21499 17527
rect 21499 17493 21508 17527
rect 21456 17484 21508 17493
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 1768 17280 1820 17332
rect 3332 17280 3384 17332
rect 7104 17280 7156 17332
rect 1768 17144 1820 17196
rect 2044 17187 2096 17196
rect 2044 17153 2053 17187
rect 2053 17153 2087 17187
rect 2087 17153 2096 17187
rect 2044 17144 2096 17153
rect 2136 17144 2188 17196
rect 2780 17144 2832 17196
rect 1584 17076 1636 17128
rect 6644 17212 6696 17264
rect 3424 17187 3476 17196
rect 3424 17153 3433 17187
rect 3433 17153 3467 17187
rect 3467 17153 3476 17187
rect 3424 17144 3476 17153
rect 4160 17144 4212 17196
rect 4620 17144 4672 17196
rect 6184 17144 6236 17196
rect 6276 17144 6328 17196
rect 6828 17187 6880 17196
rect 6828 17153 6837 17187
rect 6837 17153 6871 17187
rect 6871 17153 6880 17187
rect 6828 17144 6880 17153
rect 4344 17119 4396 17128
rect 1216 17008 1268 17060
rect 2320 17008 2372 17060
rect 4344 17085 4353 17119
rect 4353 17085 4387 17119
rect 4387 17085 4396 17119
rect 4344 17076 4396 17085
rect 5080 17076 5132 17128
rect 6092 17119 6144 17128
rect 6092 17085 6101 17119
rect 6101 17085 6135 17119
rect 6135 17085 6144 17119
rect 6092 17076 6144 17085
rect 8300 17144 8352 17196
rect 9036 17144 9088 17196
rect 10324 17212 10376 17264
rect 10784 17280 10836 17332
rect 12532 17280 12584 17332
rect 13360 17323 13412 17332
rect 13360 17289 13369 17323
rect 13369 17289 13403 17323
rect 13403 17289 13412 17323
rect 13360 17280 13412 17289
rect 11796 17212 11848 17264
rect 10416 17144 10468 17196
rect 13176 17187 13228 17196
rect 13176 17153 13185 17187
rect 13185 17153 13219 17187
rect 13219 17153 13228 17187
rect 13176 17144 13228 17153
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 2964 16940 3016 16992
rect 4160 17008 4212 17060
rect 4804 17008 4856 17060
rect 5448 16940 5500 16992
rect 6184 16940 6236 16992
rect 7104 16940 7156 16992
rect 9772 17051 9824 17060
rect 9772 17017 9781 17051
rect 9781 17017 9815 17051
rect 9815 17017 9824 17051
rect 9772 17008 9824 17017
rect 11704 17008 11756 17060
rect 14372 17076 14424 17128
rect 10140 16940 10192 16992
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 1676 16736 1728 16788
rect 3240 16779 3292 16788
rect 3240 16745 3249 16779
rect 3249 16745 3283 16779
rect 3283 16745 3292 16779
rect 3240 16736 3292 16745
rect 4160 16736 4212 16788
rect 3424 16668 3476 16720
rect 3884 16668 3936 16720
rect 4528 16668 4580 16720
rect 6092 16736 6144 16788
rect 7472 16736 7524 16788
rect 1860 16532 1912 16584
rect 1308 16464 1360 16516
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 2412 16575 2464 16584
rect 2412 16541 2421 16575
rect 2421 16541 2455 16575
rect 2455 16541 2464 16575
rect 4804 16600 4856 16652
rect 2412 16532 2464 16541
rect 3056 16532 3108 16584
rect 3976 16532 4028 16584
rect 5080 16532 5132 16584
rect 5540 16532 5592 16584
rect 6092 16532 6144 16584
rect 7012 16532 7064 16584
rect 8576 16736 8628 16788
rect 9128 16736 9180 16788
rect 8392 16668 8444 16720
rect 8484 16600 8536 16652
rect 8760 16643 8812 16652
rect 8760 16609 8769 16643
rect 8769 16609 8803 16643
rect 8803 16609 8812 16643
rect 8760 16600 8812 16609
rect 10140 16643 10192 16652
rect 10140 16609 10149 16643
rect 10149 16609 10183 16643
rect 10183 16609 10192 16643
rect 10140 16600 10192 16609
rect 11152 16736 11204 16788
rect 11888 16736 11940 16788
rect 13176 16736 13228 16788
rect 14464 16668 14516 16720
rect 8300 16532 8352 16584
rect 11244 16600 11296 16652
rect 11704 16600 11756 16652
rect 13820 16600 13872 16652
rect 11060 16532 11112 16584
rect 2688 16396 2740 16448
rect 2780 16396 2832 16448
rect 3976 16396 4028 16448
rect 4436 16439 4488 16448
rect 4436 16405 4445 16439
rect 4445 16405 4479 16439
rect 4479 16405 4488 16439
rect 4436 16396 4488 16405
rect 6828 16464 6880 16516
rect 10140 16464 10192 16516
rect 12624 16464 12676 16516
rect 8208 16396 8260 16448
rect 9496 16396 9548 16448
rect 9956 16439 10008 16448
rect 9956 16405 9965 16439
rect 9965 16405 9999 16439
rect 9999 16405 10008 16439
rect 9956 16396 10008 16405
rect 10784 16439 10836 16448
rect 10784 16405 10793 16439
rect 10793 16405 10827 16439
rect 10827 16405 10836 16439
rect 11152 16439 11204 16448
rect 10784 16396 10836 16405
rect 11152 16405 11161 16439
rect 11161 16405 11195 16439
rect 11195 16405 11204 16439
rect 11152 16396 11204 16405
rect 11796 16396 11848 16448
rect 13084 16439 13136 16448
rect 13084 16405 13093 16439
rect 13093 16405 13127 16439
rect 13127 16405 13136 16439
rect 13084 16396 13136 16405
rect 13544 16396 13596 16448
rect 14740 16439 14792 16448
rect 14740 16405 14749 16439
rect 14749 16405 14783 16439
rect 14783 16405 14792 16439
rect 14740 16396 14792 16405
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 1860 16235 1912 16244
rect 1860 16201 1869 16235
rect 1869 16201 1903 16235
rect 1903 16201 1912 16235
rect 1860 16192 1912 16201
rect 2044 16192 2096 16244
rect 2872 16235 2924 16244
rect 2872 16201 2881 16235
rect 2881 16201 2915 16235
rect 2915 16201 2924 16235
rect 2872 16192 2924 16201
rect 4804 16192 4856 16244
rect 5264 16235 5316 16244
rect 5264 16201 5273 16235
rect 5273 16201 5307 16235
rect 5307 16201 5316 16235
rect 5264 16192 5316 16201
rect 8208 16235 8260 16244
rect 8208 16201 8217 16235
rect 8217 16201 8251 16235
rect 8251 16201 8260 16235
rect 8208 16192 8260 16201
rect 9496 16235 9548 16244
rect 9496 16201 9505 16235
rect 9505 16201 9539 16235
rect 9539 16201 9548 16235
rect 9496 16192 9548 16201
rect 1952 16124 2004 16176
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 2136 16056 2188 16108
rect 2320 16099 2372 16108
rect 2320 16065 2329 16099
rect 2329 16065 2363 16099
rect 2363 16065 2372 16099
rect 2320 16056 2372 16065
rect 2780 16124 2832 16176
rect 5632 16124 5684 16176
rect 6552 16124 6604 16176
rect 8300 16124 8352 16176
rect 9404 16167 9456 16176
rect 9404 16133 9413 16167
rect 9413 16133 9447 16167
rect 9447 16133 9456 16167
rect 9404 16124 9456 16133
rect 2688 16099 2740 16108
rect 2688 16065 2697 16099
rect 2697 16065 2731 16099
rect 2731 16065 2740 16099
rect 2688 16056 2740 16065
rect 2872 16056 2924 16108
rect 3424 16099 3476 16108
rect 3424 16065 3433 16099
rect 3433 16065 3467 16099
rect 3467 16065 3476 16099
rect 3424 16056 3476 16065
rect 3884 16099 3936 16108
rect 3884 16065 3893 16099
rect 3893 16065 3927 16099
rect 3927 16065 3936 16099
rect 3884 16056 3936 16065
rect 4160 16099 4212 16108
rect 4160 16065 4194 16099
rect 4194 16065 4212 16099
rect 4160 16056 4212 16065
rect 3332 15988 3384 16040
rect 5448 16099 5500 16108
rect 5448 16065 5457 16099
rect 5457 16065 5491 16099
rect 5491 16065 5500 16099
rect 6736 16099 6788 16108
rect 5448 16056 5500 16065
rect 6736 16065 6745 16099
rect 6745 16065 6779 16099
rect 6779 16065 6788 16099
rect 6736 16056 6788 16065
rect 7012 16056 7064 16108
rect 8208 16056 8260 16108
rect 8576 16099 8628 16108
rect 8576 16065 8585 16099
rect 8585 16065 8619 16099
rect 8619 16065 8628 16099
rect 8576 16056 8628 16065
rect 10048 16192 10100 16244
rect 10140 16235 10192 16244
rect 10140 16201 10149 16235
rect 10149 16201 10183 16235
rect 10183 16201 10192 16235
rect 10140 16192 10192 16201
rect 11152 16192 11204 16244
rect 13084 16192 13136 16244
rect 13820 16235 13872 16244
rect 13820 16201 13829 16235
rect 13829 16201 13863 16235
rect 13863 16201 13872 16235
rect 13820 16192 13872 16201
rect 10324 16124 10376 16176
rect 17408 16124 17460 16176
rect 11888 16099 11940 16108
rect 1492 15963 1544 15972
rect 1492 15929 1501 15963
rect 1501 15929 1535 15963
rect 1535 15929 1544 15963
rect 1492 15920 1544 15929
rect 1768 15920 1820 15972
rect 2228 15920 2280 15972
rect 3884 15920 3936 15972
rect 3148 15895 3200 15904
rect 3148 15861 3157 15895
rect 3157 15861 3191 15895
rect 3191 15861 3200 15895
rect 3148 15852 3200 15861
rect 3332 15852 3384 15904
rect 6552 15988 6604 16040
rect 7840 16031 7892 16040
rect 7840 15997 7849 16031
rect 7849 15997 7883 16031
rect 7883 15997 7892 16031
rect 7840 15988 7892 15997
rect 7932 16031 7984 16040
rect 7932 15997 7941 16031
rect 7941 15997 7975 16031
rect 7975 15997 7984 16031
rect 7932 15988 7984 15997
rect 8392 15988 8444 16040
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 8484 15920 8536 15972
rect 9772 15988 9824 16040
rect 10140 15988 10192 16040
rect 11152 15988 11204 16040
rect 9956 15920 10008 15972
rect 12992 16056 13044 16108
rect 5816 15852 5868 15904
rect 7472 15852 7524 15904
rect 12348 15920 12400 15972
rect 15752 15852 15804 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 2136 15691 2188 15700
rect 2136 15657 2145 15691
rect 2145 15657 2179 15691
rect 2179 15657 2188 15691
rect 2136 15648 2188 15657
rect 2320 15648 2372 15700
rect 3424 15691 3476 15700
rect 3424 15657 3433 15691
rect 3433 15657 3467 15691
rect 3467 15657 3476 15691
rect 3424 15648 3476 15657
rect 4252 15648 4304 15700
rect 4436 15648 4488 15700
rect 5080 15648 5132 15700
rect 5540 15691 5592 15700
rect 5540 15657 5549 15691
rect 5549 15657 5583 15691
rect 5583 15657 5592 15691
rect 5540 15648 5592 15657
rect 8484 15691 8536 15700
rect 1676 15580 1728 15632
rect 2596 15580 2648 15632
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 2044 15487 2096 15496
rect 2044 15453 2053 15487
rect 2053 15453 2087 15487
rect 2087 15453 2096 15487
rect 2044 15444 2096 15453
rect 2412 15444 2464 15496
rect 2596 15487 2648 15496
rect 2596 15453 2605 15487
rect 2605 15453 2639 15487
rect 2639 15453 2648 15487
rect 2596 15444 2648 15453
rect 3332 15512 3384 15564
rect 3516 15555 3568 15564
rect 3516 15521 3525 15555
rect 3525 15521 3559 15555
rect 3559 15521 3568 15555
rect 3516 15512 3568 15521
rect 4160 15555 4212 15564
rect 4160 15521 4169 15555
rect 4169 15521 4203 15555
rect 4203 15521 4212 15555
rect 4160 15512 4212 15521
rect 4344 15580 4396 15632
rect 4988 15580 5040 15632
rect 8484 15657 8493 15691
rect 8493 15657 8527 15691
rect 8527 15657 8536 15691
rect 8484 15648 8536 15657
rect 13544 15691 13596 15700
rect 13544 15657 13553 15691
rect 13553 15657 13587 15691
rect 13587 15657 13596 15691
rect 13544 15648 13596 15657
rect 3148 15487 3200 15496
rect 3148 15453 3157 15487
rect 3157 15453 3191 15487
rect 3191 15453 3200 15487
rect 3148 15444 3200 15453
rect 1400 15376 1452 15428
rect 3056 15376 3108 15428
rect 3884 15444 3936 15496
rect 5540 15512 5592 15564
rect 8300 15512 8352 15564
rect 12348 15512 12400 15564
rect 12992 15555 13044 15564
rect 12992 15521 13001 15555
rect 13001 15521 13035 15555
rect 13035 15521 13044 15555
rect 12992 15512 13044 15521
rect 7748 15444 7800 15496
rect 8208 15444 8260 15496
rect 11704 15444 11756 15496
rect 14740 15444 14792 15496
rect 16212 15487 16264 15496
rect 4068 15376 4120 15428
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 1860 15351 1912 15360
rect 1860 15317 1869 15351
rect 1869 15317 1903 15351
rect 1903 15317 1912 15351
rect 1860 15308 1912 15317
rect 3976 15308 4028 15360
rect 6828 15376 6880 15428
rect 7012 15419 7064 15428
rect 7012 15385 7021 15419
rect 7021 15385 7055 15419
rect 7055 15385 7064 15419
rect 7012 15376 7064 15385
rect 7104 15376 7156 15428
rect 10416 15419 10468 15428
rect 10416 15385 10425 15419
rect 10425 15385 10459 15419
rect 10459 15385 10468 15419
rect 10416 15376 10468 15385
rect 13820 15376 13872 15428
rect 4252 15351 4304 15360
rect 4252 15317 4261 15351
rect 4261 15317 4295 15351
rect 4295 15317 4304 15351
rect 4252 15308 4304 15317
rect 6000 15308 6052 15360
rect 7472 15308 7524 15360
rect 8576 15308 8628 15360
rect 12256 15308 12308 15360
rect 13176 15351 13228 15360
rect 13176 15317 13185 15351
rect 13185 15317 13219 15351
rect 13219 15317 13228 15351
rect 16212 15453 16221 15487
rect 16221 15453 16255 15487
rect 16255 15453 16264 15487
rect 16212 15444 16264 15453
rect 13176 15308 13228 15317
rect 15660 15308 15712 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 1676 15104 1728 15156
rect 2596 15104 2648 15156
rect 3148 15147 3200 15156
rect 3148 15113 3157 15147
rect 3157 15113 3191 15147
rect 3191 15113 3200 15147
rect 3148 15104 3200 15113
rect 2412 15036 2464 15088
rect 1860 14968 1912 15020
rect 1952 14968 2004 15020
rect 2228 14968 2280 15020
rect 6000 15104 6052 15156
rect 3424 15036 3476 15088
rect 1768 14900 1820 14952
rect 3976 14968 4028 15020
rect 6552 15104 6604 15156
rect 7840 15104 7892 15156
rect 9128 15104 9180 15156
rect 9312 15104 9364 15156
rect 9588 15104 9640 15156
rect 11060 15104 11112 15156
rect 11796 15104 11848 15156
rect 12900 15147 12952 15156
rect 12900 15113 12909 15147
rect 12909 15113 12943 15147
rect 12943 15113 12952 15147
rect 12900 15104 12952 15113
rect 13176 15104 13228 15156
rect 13820 15147 13872 15156
rect 13820 15113 13829 15147
rect 13829 15113 13863 15147
rect 13863 15113 13872 15147
rect 13820 15104 13872 15113
rect 7472 15011 7524 15020
rect 7472 14977 7490 15011
rect 7490 14977 7524 15011
rect 7472 14968 7524 14977
rect 7748 15011 7800 15020
rect 7748 14977 7757 15011
rect 7757 14977 7791 15011
rect 7791 14977 7800 15011
rect 7748 14968 7800 14977
rect 8576 14968 8628 15020
rect 9036 14968 9088 15020
rect 9496 14968 9548 15020
rect 10140 15011 10192 15020
rect 3332 14900 3384 14952
rect 3700 14943 3752 14952
rect 3700 14909 3709 14943
rect 3709 14909 3743 14943
rect 3743 14909 3752 14943
rect 3700 14900 3752 14909
rect 4068 14943 4120 14952
rect 2044 14832 2096 14884
rect 3516 14832 3568 14884
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 3240 14764 3292 14816
rect 4068 14909 4077 14943
rect 4077 14909 4111 14943
rect 4111 14909 4120 14943
rect 4068 14900 4120 14909
rect 8024 14900 8076 14952
rect 8760 14943 8812 14952
rect 8760 14909 8769 14943
rect 8769 14909 8803 14943
rect 8803 14909 8812 14943
rect 8760 14900 8812 14909
rect 10140 14977 10174 15011
rect 10174 14977 10192 15011
rect 10140 14968 10192 14977
rect 12348 15036 12400 15088
rect 11796 15011 11848 15020
rect 11796 14977 11830 15011
rect 11830 14977 11848 15011
rect 11796 14968 11848 14977
rect 5448 14875 5500 14884
rect 5448 14841 5457 14875
rect 5457 14841 5491 14875
rect 5491 14841 5500 14875
rect 5448 14832 5500 14841
rect 12624 14968 12676 15020
rect 13728 14968 13780 15020
rect 15292 14968 15344 15020
rect 15568 14968 15620 15020
rect 13452 14943 13504 14952
rect 13452 14909 13461 14943
rect 13461 14909 13495 14943
rect 13495 14909 13504 14943
rect 13452 14900 13504 14909
rect 15108 14943 15160 14952
rect 15108 14909 15117 14943
rect 15117 14909 15151 14943
rect 15151 14909 15160 14943
rect 15108 14900 15160 14909
rect 13820 14832 13872 14884
rect 7104 14764 7156 14816
rect 7472 14764 7524 14816
rect 9680 14764 9732 14816
rect 10600 14764 10652 14816
rect 15568 14807 15620 14816
rect 15568 14773 15577 14807
rect 15577 14773 15611 14807
rect 15611 14773 15620 14807
rect 15568 14764 15620 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 3332 14560 3384 14612
rect 3884 14560 3936 14612
rect 6644 14560 6696 14612
rect 1308 14424 1360 14476
rect 2044 14356 2096 14408
rect 4068 14424 4120 14476
rect 2228 14356 2280 14408
rect 1400 14288 1452 14340
rect 3332 14331 3384 14340
rect 3332 14297 3350 14331
rect 3350 14297 3384 14331
rect 4528 14356 4580 14408
rect 4988 14467 5040 14476
rect 4988 14433 4997 14467
rect 4997 14433 5031 14467
rect 5031 14433 5040 14467
rect 4988 14424 5040 14433
rect 5632 14356 5684 14408
rect 5816 14399 5868 14408
rect 5816 14365 5850 14399
rect 5850 14365 5868 14399
rect 5816 14356 5868 14365
rect 3332 14288 3384 14297
rect 4620 14288 4672 14340
rect 5448 14288 5500 14340
rect 7472 14560 7524 14612
rect 7564 14560 7616 14612
rect 7748 14560 7800 14612
rect 8024 14560 8076 14612
rect 9128 14603 9180 14612
rect 9128 14569 9137 14603
rect 9137 14569 9171 14603
rect 9171 14569 9180 14603
rect 9128 14560 9180 14569
rect 7196 14492 7248 14544
rect 7932 14492 7984 14544
rect 8576 14492 8628 14544
rect 9864 14560 9916 14612
rect 10784 14560 10836 14612
rect 11244 14560 11296 14612
rect 13728 14603 13780 14612
rect 13728 14569 13737 14603
rect 13737 14569 13771 14603
rect 13771 14569 13780 14603
rect 13728 14560 13780 14569
rect 8024 14424 8076 14476
rect 6828 14288 6880 14340
rect 10048 14492 10100 14544
rect 10968 14492 11020 14544
rect 10140 14424 10192 14476
rect 11152 14467 11204 14476
rect 9772 14399 9824 14408
rect 9772 14365 9781 14399
rect 9781 14365 9815 14399
rect 9815 14365 9824 14399
rect 11152 14433 11161 14467
rect 11161 14433 11195 14467
rect 11195 14433 11204 14467
rect 11152 14424 11204 14433
rect 12624 14467 12676 14476
rect 12624 14433 12633 14467
rect 12633 14433 12667 14467
rect 12667 14433 12676 14467
rect 12624 14424 12676 14433
rect 13268 14492 13320 14544
rect 19064 14560 19116 14612
rect 13820 14424 13872 14476
rect 16212 14424 16264 14476
rect 9772 14356 9824 14365
rect 12348 14356 12400 14408
rect 14280 14356 14332 14408
rect 15660 14399 15712 14408
rect 15660 14365 15678 14399
rect 15678 14365 15712 14399
rect 15660 14356 15712 14365
rect 16948 14356 17000 14408
rect 9680 14288 9732 14340
rect 16488 14331 16540 14340
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 2504 14220 2556 14272
rect 3240 14220 3292 14272
rect 3608 14220 3660 14272
rect 3884 14220 3936 14272
rect 4896 14263 4948 14272
rect 4896 14229 4905 14263
rect 4905 14229 4939 14263
rect 4939 14229 4948 14263
rect 5264 14263 5316 14272
rect 4896 14220 4948 14229
rect 5264 14229 5273 14263
rect 5273 14229 5307 14263
rect 5307 14229 5316 14263
rect 5264 14220 5316 14229
rect 5356 14220 5408 14272
rect 7472 14220 7524 14272
rect 7564 14220 7616 14272
rect 8116 14263 8168 14272
rect 8116 14229 8125 14263
rect 8125 14229 8159 14263
rect 8159 14229 8168 14263
rect 8116 14220 8168 14229
rect 8208 14263 8260 14272
rect 8208 14229 8217 14263
rect 8217 14229 8251 14263
rect 8251 14229 8260 14263
rect 8208 14220 8260 14229
rect 8392 14220 8444 14272
rect 8668 14220 8720 14272
rect 9864 14263 9916 14272
rect 9864 14229 9873 14263
rect 9873 14229 9907 14263
rect 9907 14229 9916 14263
rect 9864 14220 9916 14229
rect 10692 14220 10744 14272
rect 10968 14263 11020 14272
rect 10968 14229 10977 14263
rect 10977 14229 11011 14263
rect 11011 14229 11020 14263
rect 10968 14220 11020 14229
rect 11796 14220 11848 14272
rect 12072 14220 12124 14272
rect 12624 14220 12676 14272
rect 13268 14263 13320 14272
rect 13268 14229 13277 14263
rect 13277 14229 13311 14263
rect 13311 14229 13320 14263
rect 13268 14220 13320 14229
rect 13636 14220 13688 14272
rect 14740 14220 14792 14272
rect 14924 14220 14976 14272
rect 16488 14297 16497 14331
rect 16497 14297 16531 14331
rect 16531 14297 16540 14331
rect 16488 14288 16540 14297
rect 16396 14263 16448 14272
rect 16396 14229 16405 14263
rect 16405 14229 16439 14263
rect 16439 14229 16448 14263
rect 16396 14220 16448 14229
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 1860 14059 1912 14068
rect 1860 14025 1869 14059
rect 1869 14025 1903 14059
rect 1903 14025 1912 14059
rect 1860 14016 1912 14025
rect 2044 14016 2096 14068
rect 3424 14016 3476 14068
rect 3608 14059 3660 14068
rect 3608 14025 3617 14059
rect 3617 14025 3651 14059
rect 3651 14025 3660 14059
rect 3608 14016 3660 14025
rect 3976 14059 4028 14068
rect 3976 14025 3985 14059
rect 3985 14025 4019 14059
rect 4019 14025 4028 14059
rect 3976 14016 4028 14025
rect 4160 14016 4212 14068
rect 4988 14016 5040 14068
rect 7564 14059 7616 14068
rect 7564 14025 7573 14059
rect 7573 14025 7607 14059
rect 7607 14025 7616 14059
rect 7564 14016 7616 14025
rect 7656 14016 7708 14068
rect 8116 14016 8168 14068
rect 10692 14059 10744 14068
rect 10692 14025 10701 14059
rect 10701 14025 10735 14059
rect 10735 14025 10744 14059
rect 10692 14016 10744 14025
rect 11888 14016 11940 14068
rect 12348 14016 12400 14068
rect 13820 14059 13872 14068
rect 13820 14025 13829 14059
rect 13829 14025 13863 14059
rect 13863 14025 13872 14059
rect 13820 14016 13872 14025
rect 14924 14059 14976 14068
rect 14924 14025 14933 14059
rect 14933 14025 14967 14059
rect 14967 14025 14976 14059
rect 14924 14016 14976 14025
rect 16396 14016 16448 14068
rect 9312 13948 9364 14000
rect 9864 13948 9916 14000
rect 10600 13948 10652 14000
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 2044 13923 2096 13932
rect 2044 13889 2053 13923
rect 2053 13889 2087 13923
rect 2087 13889 2096 13923
rect 2044 13880 2096 13889
rect 2504 13923 2556 13932
rect 2504 13889 2513 13923
rect 2513 13889 2547 13923
rect 2547 13889 2556 13923
rect 2504 13880 2556 13889
rect 3332 13880 3384 13932
rect 2688 13812 2740 13864
rect 4160 13880 4212 13932
rect 3516 13855 3568 13864
rect 3516 13821 3525 13855
rect 3525 13821 3559 13855
rect 3559 13821 3568 13855
rect 5356 13880 5408 13932
rect 5540 13923 5592 13932
rect 5540 13889 5549 13923
rect 5549 13889 5583 13923
rect 5583 13889 5592 13923
rect 5540 13880 5592 13889
rect 7288 13880 7340 13932
rect 8024 13880 8076 13932
rect 8300 13880 8352 13932
rect 3516 13812 3568 13821
rect 5724 13812 5776 13864
rect 6552 13744 6604 13796
rect 9312 13855 9364 13864
rect 9312 13821 9321 13855
rect 9321 13821 9355 13855
rect 9355 13821 9364 13855
rect 9312 13812 9364 13821
rect 7472 13744 7524 13796
rect 7564 13744 7616 13796
rect 9496 13880 9548 13932
rect 10232 13880 10284 13932
rect 12808 13948 12860 14000
rect 15108 13948 15160 14000
rect 11152 13880 11204 13932
rect 12072 13880 12124 13932
rect 13728 13923 13780 13932
rect 9864 13855 9916 13864
rect 9864 13821 9873 13855
rect 9873 13821 9907 13855
rect 9907 13821 9916 13855
rect 9864 13812 9916 13821
rect 11060 13812 11112 13864
rect 11796 13812 11848 13864
rect 12808 13787 12860 13796
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 7104 13719 7156 13728
rect 7104 13685 7113 13719
rect 7113 13685 7147 13719
rect 7147 13685 7156 13719
rect 7932 13719 7984 13728
rect 7104 13676 7156 13685
rect 7932 13685 7941 13719
rect 7941 13685 7975 13719
rect 7975 13685 7984 13719
rect 7932 13676 7984 13685
rect 12808 13753 12817 13787
rect 12817 13753 12851 13787
rect 12851 13753 12860 13787
rect 12808 13744 12860 13753
rect 13728 13889 13737 13923
rect 13737 13889 13771 13923
rect 13771 13889 13780 13923
rect 13728 13880 13780 13889
rect 16304 13880 16356 13932
rect 21364 13880 21416 13932
rect 14740 13855 14792 13864
rect 14740 13821 14749 13855
rect 14749 13821 14783 13855
rect 14783 13821 14792 13855
rect 14740 13812 14792 13821
rect 16304 13744 16356 13796
rect 9772 13676 9824 13728
rect 11888 13676 11940 13728
rect 12348 13676 12400 13728
rect 15568 13676 15620 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 1676 13472 1728 13524
rect 2596 13472 2648 13524
rect 3424 13515 3476 13524
rect 3424 13481 3433 13515
rect 3433 13481 3467 13515
rect 3467 13481 3476 13515
rect 3424 13472 3476 13481
rect 4436 13472 4488 13524
rect 4896 13472 4948 13524
rect 8208 13472 8260 13524
rect 9128 13472 9180 13524
rect 9680 13472 9732 13524
rect 11704 13472 11756 13524
rect 15108 13472 15160 13524
rect 16304 13515 16356 13524
rect 16304 13481 16313 13515
rect 16313 13481 16347 13515
rect 16347 13481 16356 13515
rect 16304 13472 16356 13481
rect 16396 13472 16448 13524
rect 17040 13472 17092 13524
rect 2872 13404 2924 13456
rect 8024 13447 8076 13456
rect 8024 13413 8033 13447
rect 8033 13413 8067 13447
rect 8067 13413 8076 13447
rect 8024 13404 8076 13413
rect 8576 13404 8628 13456
rect 9496 13404 9548 13456
rect 15476 13404 15528 13456
rect 2228 13336 2280 13388
rect 2780 13336 2832 13388
rect 3424 13336 3476 13388
rect 5540 13336 5592 13388
rect 8208 13336 8260 13388
rect 8668 13379 8720 13388
rect 8668 13345 8677 13379
rect 8677 13345 8711 13379
rect 8711 13345 8720 13379
rect 8668 13336 8720 13345
rect 9036 13336 9088 13388
rect 9404 13336 9456 13388
rect 10508 13336 10560 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 1860 13268 1912 13320
rect 2964 13268 3016 13320
rect 1584 13175 1636 13184
rect 1584 13141 1593 13175
rect 1593 13141 1627 13175
rect 1627 13141 1636 13175
rect 1584 13132 1636 13141
rect 2136 13132 2188 13184
rect 2412 13175 2464 13184
rect 2412 13141 2421 13175
rect 2421 13141 2455 13175
rect 2455 13141 2464 13175
rect 2412 13132 2464 13141
rect 2504 13175 2556 13184
rect 2504 13141 2513 13175
rect 2513 13141 2547 13175
rect 2547 13141 2556 13175
rect 5448 13268 5500 13320
rect 6644 13268 6696 13320
rect 7012 13311 7064 13320
rect 7012 13277 7021 13311
rect 7021 13277 7055 13311
rect 7055 13277 7064 13311
rect 10416 13311 10468 13320
rect 7012 13268 7064 13277
rect 10416 13277 10425 13311
rect 10425 13277 10459 13311
rect 10459 13277 10468 13311
rect 10416 13268 10468 13277
rect 5632 13200 5684 13252
rect 7564 13243 7616 13252
rect 7564 13209 7573 13243
rect 7573 13209 7607 13243
rect 7607 13209 7616 13243
rect 7564 13200 7616 13209
rect 2504 13132 2556 13141
rect 5724 13175 5776 13184
rect 5724 13141 5733 13175
rect 5733 13141 5767 13175
rect 5767 13141 5776 13175
rect 5724 13132 5776 13141
rect 5816 13132 5868 13184
rect 7840 13132 7892 13184
rect 9128 13132 9180 13184
rect 9404 13132 9456 13184
rect 9864 13175 9916 13184
rect 9864 13141 9873 13175
rect 9873 13141 9907 13175
rect 9907 13141 9916 13175
rect 9864 13132 9916 13141
rect 9956 13175 10008 13184
rect 9956 13141 9965 13175
rect 9965 13141 9999 13175
rect 9999 13141 10008 13175
rect 9956 13132 10008 13141
rect 11244 13132 11296 13184
rect 11704 13175 11756 13184
rect 11704 13141 11713 13175
rect 11713 13141 11747 13175
rect 11747 13141 11756 13175
rect 11704 13132 11756 13141
rect 14740 13336 14792 13388
rect 12900 13268 12952 13320
rect 15752 13268 15804 13320
rect 16948 13268 17000 13320
rect 21364 13200 21416 13252
rect 12808 13132 12860 13184
rect 13176 13132 13228 13184
rect 13728 13175 13780 13184
rect 13728 13141 13737 13175
rect 13737 13141 13771 13175
rect 13771 13141 13780 13175
rect 13728 13132 13780 13141
rect 15200 13132 15252 13184
rect 15384 13175 15436 13184
rect 15384 13141 15393 13175
rect 15393 13141 15427 13175
rect 15427 13141 15436 13175
rect 15384 13132 15436 13141
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 1860 12971 1912 12980
rect 1860 12937 1869 12971
rect 1869 12937 1903 12971
rect 1903 12937 1912 12971
rect 1860 12928 1912 12937
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 2136 12928 2188 12980
rect 5816 12928 5868 12980
rect 6736 12928 6788 12980
rect 7748 12928 7800 12980
rect 7840 12928 7892 12980
rect 11152 12928 11204 12980
rect 2596 12860 2648 12912
rect 3148 12835 3200 12844
rect 3148 12801 3157 12835
rect 3157 12801 3191 12835
rect 3191 12801 3200 12835
rect 3148 12792 3200 12801
rect 5724 12860 5776 12912
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 2228 12656 2280 12708
rect 4896 12792 4948 12844
rect 7932 12860 7984 12912
rect 8668 12860 8720 12912
rect 11336 12860 11388 12912
rect 11704 12928 11756 12980
rect 12900 12971 12952 12980
rect 12900 12937 12909 12971
rect 12909 12937 12943 12971
rect 12943 12937 12952 12971
rect 12900 12928 12952 12937
rect 13360 12971 13412 12980
rect 13360 12937 13369 12971
rect 13369 12937 13403 12971
rect 13403 12937 13412 12971
rect 13360 12928 13412 12937
rect 13452 12928 13504 12980
rect 14648 12928 14700 12980
rect 15476 12971 15528 12980
rect 15476 12937 15485 12971
rect 15485 12937 15519 12971
rect 15519 12937 15528 12971
rect 15476 12928 15528 12937
rect 15568 12971 15620 12980
rect 15568 12937 15577 12971
rect 15577 12937 15611 12971
rect 15611 12937 15620 12971
rect 15568 12928 15620 12937
rect 7472 12792 7524 12844
rect 8208 12792 8260 12844
rect 8484 12792 8536 12844
rect 9312 12792 9364 12844
rect 9496 12835 9548 12844
rect 9496 12801 9530 12835
rect 9530 12801 9548 12835
rect 9496 12792 9548 12801
rect 7012 12767 7064 12776
rect 7012 12733 7021 12767
rect 7021 12733 7055 12767
rect 7055 12733 7064 12767
rect 7012 12724 7064 12733
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 4804 12656 4856 12708
rect 6552 12656 6604 12708
rect 6828 12656 6880 12708
rect 11060 12724 11112 12776
rect 16396 12860 16448 12912
rect 12072 12792 12124 12844
rect 15752 12792 15804 12844
rect 13176 12767 13228 12776
rect 13176 12733 13185 12767
rect 13185 12733 13219 12767
rect 13219 12733 13228 12767
rect 13176 12724 13228 12733
rect 13452 12724 13504 12776
rect 14464 12724 14516 12776
rect 15568 12724 15620 12776
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 4068 12588 4120 12640
rect 5080 12588 5132 12640
rect 6644 12588 6696 12640
rect 9220 12656 9272 12708
rect 8668 12588 8720 12640
rect 10600 12631 10652 12640
rect 10600 12597 10609 12631
rect 10609 12597 10643 12631
rect 10643 12597 10652 12631
rect 10600 12588 10652 12597
rect 11704 12588 11756 12640
rect 15200 12656 15252 12708
rect 13360 12588 13412 12640
rect 14832 12588 14884 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 2964 12384 3016 12436
rect 3332 12384 3384 12436
rect 5540 12384 5592 12436
rect 6644 12384 6696 12436
rect 7012 12384 7064 12436
rect 7380 12384 7432 12436
rect 7656 12384 7708 12436
rect 9496 12384 9548 12436
rect 9864 12384 9916 12436
rect 10508 12427 10560 12436
rect 10508 12393 10517 12427
rect 10517 12393 10551 12427
rect 10551 12393 10560 12427
rect 10508 12384 10560 12393
rect 12072 12384 12124 12436
rect 12716 12427 12768 12436
rect 12716 12393 12725 12427
rect 12725 12393 12759 12427
rect 12759 12393 12768 12427
rect 12716 12384 12768 12393
rect 14648 12384 14700 12436
rect 15016 12384 15068 12436
rect 8392 12316 8444 12368
rect 8760 12316 8812 12368
rect 9036 12316 9088 12368
rect 5540 12291 5592 12300
rect 1492 12180 1544 12232
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 5540 12257 5549 12291
rect 5549 12257 5583 12291
rect 5583 12257 5592 12291
rect 5540 12248 5592 12257
rect 8484 12248 8536 12300
rect 10784 12316 10836 12368
rect 3332 12223 3384 12232
rect 3332 12189 3341 12223
rect 3341 12189 3375 12223
rect 3375 12189 3384 12223
rect 3332 12180 3384 12189
rect 5724 12180 5776 12232
rect 10600 12248 10652 12300
rect 12900 12248 12952 12300
rect 4160 12112 4212 12164
rect 5632 12112 5684 12164
rect 6552 12112 6604 12164
rect 6828 12112 6880 12164
rect 1860 12087 1912 12096
rect 1860 12053 1869 12087
rect 1869 12053 1903 12087
rect 1903 12053 1912 12087
rect 1860 12044 1912 12053
rect 1952 12087 2004 12096
rect 1952 12053 1961 12087
rect 1961 12053 1995 12087
rect 1995 12053 2004 12087
rect 1952 12044 2004 12053
rect 2320 12044 2372 12096
rect 2596 12044 2648 12096
rect 2964 12044 3016 12096
rect 4068 12044 4120 12096
rect 4712 12044 4764 12096
rect 8668 12180 8720 12232
rect 8392 12112 8444 12164
rect 11060 12180 11112 12232
rect 11336 12180 11388 12232
rect 7288 12087 7340 12096
rect 7288 12053 7297 12087
rect 7297 12053 7331 12087
rect 7331 12053 7340 12087
rect 7288 12044 7340 12053
rect 8116 12087 8168 12096
rect 8116 12053 8125 12087
rect 8125 12053 8159 12087
rect 8159 12053 8168 12087
rect 8116 12044 8168 12053
rect 9496 12112 9548 12164
rect 10600 12112 10652 12164
rect 13544 12112 13596 12164
rect 14740 12112 14792 12164
rect 14924 12180 14976 12232
rect 16948 12112 17000 12164
rect 10048 12087 10100 12096
rect 10048 12053 10057 12087
rect 10057 12053 10091 12087
rect 10091 12053 10100 12087
rect 10048 12044 10100 12053
rect 11244 12044 11296 12096
rect 13268 12087 13320 12096
rect 13268 12053 13277 12087
rect 13277 12053 13311 12087
rect 13311 12053 13320 12087
rect 13268 12044 13320 12053
rect 15568 12044 15620 12096
rect 16396 12087 16448 12096
rect 16396 12053 16405 12087
rect 16405 12053 16439 12087
rect 16439 12053 16448 12087
rect 16396 12044 16448 12053
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 2320 11840 2372 11892
rect 1952 11772 2004 11824
rect 2228 11772 2280 11824
rect 3148 11840 3200 11892
rect 4712 11840 4764 11892
rect 5172 11840 5224 11892
rect 3332 11636 3384 11688
rect 1860 11500 1912 11552
rect 3056 11568 3108 11620
rect 4068 11568 4120 11620
rect 2964 11500 3016 11552
rect 4252 11500 4304 11552
rect 5632 11772 5684 11824
rect 7104 11840 7156 11892
rect 7564 11840 7616 11892
rect 8576 11840 8628 11892
rect 9036 11883 9088 11892
rect 9036 11849 9045 11883
rect 9045 11849 9079 11883
rect 9079 11849 9088 11883
rect 9036 11840 9088 11849
rect 9128 11883 9180 11892
rect 9128 11849 9137 11883
rect 9137 11849 9171 11883
rect 9171 11849 9180 11883
rect 9496 11883 9548 11892
rect 9128 11840 9180 11849
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 10416 11840 10468 11892
rect 13544 11883 13596 11892
rect 13544 11849 13553 11883
rect 13553 11849 13587 11883
rect 13587 11849 13596 11883
rect 13544 11840 13596 11849
rect 14464 11840 14516 11892
rect 14924 11840 14976 11892
rect 15752 11883 15804 11892
rect 15752 11849 15761 11883
rect 15761 11849 15795 11883
rect 15795 11849 15804 11883
rect 15752 11840 15804 11849
rect 10232 11772 10284 11824
rect 12164 11772 12216 11824
rect 13820 11772 13872 11824
rect 14372 11772 14424 11824
rect 5448 11747 5500 11756
rect 5448 11713 5457 11747
rect 5457 11713 5491 11747
rect 5491 11713 5500 11747
rect 5448 11704 5500 11713
rect 5540 11704 5592 11756
rect 7012 11704 7064 11756
rect 8668 11704 8720 11756
rect 5356 11679 5408 11688
rect 5356 11645 5365 11679
rect 5365 11645 5399 11679
rect 5399 11645 5408 11679
rect 5356 11636 5408 11645
rect 5908 11679 5960 11688
rect 5908 11645 5917 11679
rect 5917 11645 5951 11679
rect 5951 11645 5960 11679
rect 5908 11636 5960 11645
rect 7288 11636 7340 11688
rect 5816 11568 5868 11620
rect 8208 11636 8260 11688
rect 9036 11636 9088 11688
rect 11796 11704 11848 11756
rect 11888 11704 11940 11756
rect 12348 11747 12400 11756
rect 10600 11636 10652 11688
rect 12348 11713 12357 11747
rect 12357 11713 12391 11747
rect 12391 11713 12400 11747
rect 12348 11704 12400 11713
rect 12256 11679 12308 11688
rect 7564 11568 7616 11620
rect 12256 11645 12265 11679
rect 12265 11645 12299 11679
rect 12299 11645 12308 11679
rect 12256 11636 12308 11645
rect 15568 11704 15620 11756
rect 16948 11772 17000 11824
rect 16120 11747 16172 11756
rect 16120 11713 16129 11747
rect 16129 11713 16163 11747
rect 16163 11713 16172 11747
rect 16120 11704 16172 11713
rect 13360 11636 13412 11688
rect 16212 11679 16264 11688
rect 4712 11500 4764 11552
rect 4804 11500 4856 11552
rect 5632 11500 5684 11552
rect 7380 11500 7432 11552
rect 8668 11543 8720 11552
rect 8668 11509 8677 11543
rect 8677 11509 8711 11543
rect 8711 11509 8720 11543
rect 8668 11500 8720 11509
rect 11520 11543 11572 11552
rect 11520 11509 11529 11543
rect 11529 11509 11563 11543
rect 11563 11509 11572 11543
rect 11520 11500 11572 11509
rect 11888 11500 11940 11552
rect 13544 11568 13596 11620
rect 16212 11645 16221 11679
rect 16221 11645 16255 11679
rect 16255 11645 16264 11679
rect 16212 11636 16264 11645
rect 13268 11500 13320 11552
rect 13728 11500 13780 11552
rect 18512 11500 18564 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 1400 11339 1452 11348
rect 1400 11305 1409 11339
rect 1409 11305 1443 11339
rect 1443 11305 1452 11339
rect 1400 11296 1452 11305
rect 2320 11339 2372 11348
rect 2320 11305 2329 11339
rect 2329 11305 2363 11339
rect 2363 11305 2372 11339
rect 2320 11296 2372 11305
rect 1860 11160 1912 11212
rect 5080 11296 5132 11348
rect 5448 11296 5500 11348
rect 6092 11296 6144 11348
rect 6920 11296 6972 11348
rect 8116 11296 8168 11348
rect 8484 11296 8536 11348
rect 9956 11296 10008 11348
rect 3424 11228 3476 11280
rect 4436 11271 4488 11280
rect 4436 11237 4445 11271
rect 4445 11237 4479 11271
rect 4479 11237 4488 11271
rect 4436 11228 4488 11237
rect 2596 11160 2648 11212
rect 2780 11160 2832 11212
rect 3056 11203 3108 11212
rect 3056 11169 3065 11203
rect 3065 11169 3099 11203
rect 3099 11169 3108 11203
rect 3056 11160 3108 11169
rect 3608 11203 3660 11212
rect 3608 11169 3617 11203
rect 3617 11169 3651 11203
rect 3651 11169 3660 11203
rect 3608 11160 3660 11169
rect 3976 11160 4028 11212
rect 4896 11160 4948 11212
rect 5724 11160 5776 11212
rect 2044 11092 2096 11144
rect 5908 11092 5960 11144
rect 1584 10956 1636 11008
rect 3332 11024 3384 11076
rect 2504 10956 2556 11008
rect 3608 10956 3660 11008
rect 3792 10956 3844 11008
rect 4712 11024 4764 11076
rect 5540 11024 5592 11076
rect 5816 11067 5868 11076
rect 5816 11033 5825 11067
rect 5825 11033 5859 11067
rect 5859 11033 5868 11067
rect 5816 11024 5868 11033
rect 6828 11160 6880 11212
rect 6736 11092 6788 11144
rect 10600 11160 10652 11212
rect 11152 11160 11204 11212
rect 9680 11092 9732 11144
rect 11796 11092 11848 11144
rect 12808 11203 12860 11212
rect 12808 11169 12817 11203
rect 12817 11169 12851 11203
rect 12851 11169 12860 11203
rect 12808 11160 12860 11169
rect 17224 11296 17276 11348
rect 7840 11024 7892 11076
rect 9588 11024 9640 11076
rect 10048 11024 10100 11076
rect 11980 11024 12032 11076
rect 5080 10956 5132 11008
rect 6000 10956 6052 11008
rect 6552 10999 6604 11008
rect 6552 10965 6561 10999
rect 6561 10965 6595 10999
rect 6595 10965 6604 10999
rect 6552 10956 6604 10965
rect 6644 10956 6696 11008
rect 8116 10956 8168 11008
rect 10324 10999 10376 11008
rect 10324 10965 10333 10999
rect 10333 10965 10367 10999
rect 10367 10965 10376 10999
rect 10324 10956 10376 10965
rect 10600 10956 10652 11008
rect 10968 10956 11020 11008
rect 12256 10999 12308 11008
rect 12256 10965 12265 10999
rect 12265 10965 12299 10999
rect 12299 10965 12308 10999
rect 12256 10956 12308 10965
rect 13820 11092 13872 11144
rect 13544 11067 13596 11076
rect 13544 11033 13553 11067
rect 13553 11033 13587 11067
rect 13587 11033 13596 11067
rect 14464 11092 14516 11144
rect 13544 11024 13596 11033
rect 16396 11024 16448 11076
rect 14648 10999 14700 11008
rect 14648 10965 14657 10999
rect 14657 10965 14691 10999
rect 14691 10965 14700 10999
rect 14648 10956 14700 10965
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 4344 10752 4396 10804
rect 5356 10752 5408 10804
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 1860 10616 1912 10668
rect 2320 10616 2372 10668
rect 3240 10616 3292 10668
rect 3792 10616 3844 10668
rect 2412 10591 2464 10600
rect 1952 10480 2004 10532
rect 2136 10523 2188 10532
rect 2136 10489 2145 10523
rect 2145 10489 2179 10523
rect 2179 10489 2188 10523
rect 2136 10480 2188 10489
rect 2412 10557 2421 10591
rect 2421 10557 2455 10591
rect 2455 10557 2464 10591
rect 2412 10548 2464 10557
rect 4896 10684 4948 10736
rect 5264 10684 5316 10736
rect 7472 10752 7524 10804
rect 7840 10752 7892 10804
rect 8392 10752 8444 10804
rect 8668 10752 8720 10804
rect 9128 10752 9180 10804
rect 4988 10616 5040 10668
rect 5724 10616 5776 10668
rect 6736 10684 6788 10736
rect 6828 10684 6880 10736
rect 11796 10752 11848 10804
rect 12256 10752 12308 10804
rect 14556 10752 14608 10804
rect 14648 10752 14700 10804
rect 16120 10752 16172 10804
rect 6644 10659 6696 10668
rect 6644 10625 6678 10659
rect 6678 10625 6696 10659
rect 6644 10616 6696 10625
rect 9680 10659 9732 10668
rect 5540 10591 5592 10600
rect 2044 10412 2096 10464
rect 2228 10455 2280 10464
rect 2228 10421 2237 10455
rect 2237 10421 2271 10455
rect 2271 10421 2280 10455
rect 2228 10412 2280 10421
rect 3976 10480 4028 10532
rect 4068 10480 4120 10532
rect 5540 10557 5549 10591
rect 5549 10557 5583 10591
rect 5583 10557 5592 10591
rect 5540 10548 5592 10557
rect 4620 10480 4672 10532
rect 7840 10548 7892 10600
rect 9680 10625 9689 10659
rect 9689 10625 9723 10659
rect 9723 10625 9732 10659
rect 9680 10616 9732 10625
rect 15476 10684 15528 10736
rect 11612 10616 11664 10668
rect 12624 10659 12676 10668
rect 12624 10625 12633 10659
rect 12633 10625 12667 10659
rect 12667 10625 12676 10659
rect 12624 10616 12676 10625
rect 14188 10659 14240 10668
rect 14188 10625 14206 10659
rect 14206 10625 14240 10659
rect 14188 10616 14240 10625
rect 14464 10659 14516 10668
rect 14464 10625 14473 10659
rect 14473 10625 14507 10659
rect 14507 10625 14516 10659
rect 14464 10616 14516 10625
rect 9956 10591 10008 10600
rect 9956 10557 9965 10591
rect 9965 10557 9999 10591
rect 9999 10557 10008 10591
rect 9956 10548 10008 10557
rect 10324 10548 10376 10600
rect 10692 10591 10744 10600
rect 10692 10557 10701 10591
rect 10701 10557 10735 10591
rect 10735 10557 10744 10591
rect 10692 10548 10744 10557
rect 11796 10591 11848 10600
rect 3332 10412 3384 10464
rect 3884 10412 3936 10464
rect 8208 10480 8260 10532
rect 11796 10557 11805 10591
rect 11805 10557 11839 10591
rect 11839 10557 11848 10591
rect 11796 10548 11848 10557
rect 12440 10591 12492 10600
rect 12440 10557 12449 10591
rect 12449 10557 12483 10591
rect 12483 10557 12492 10591
rect 14740 10591 14792 10600
rect 12440 10548 12492 10557
rect 14740 10557 14749 10591
rect 14749 10557 14783 10591
rect 14783 10557 14792 10591
rect 14740 10548 14792 10557
rect 5908 10455 5960 10464
rect 5908 10421 5917 10455
rect 5917 10421 5951 10455
rect 5951 10421 5960 10455
rect 5908 10412 5960 10421
rect 6000 10412 6052 10464
rect 6644 10412 6696 10464
rect 9312 10455 9364 10464
rect 9312 10421 9321 10455
rect 9321 10421 9355 10455
rect 9355 10421 9364 10455
rect 9312 10412 9364 10421
rect 11612 10455 11664 10464
rect 11612 10421 11621 10455
rect 11621 10421 11655 10455
rect 11655 10421 11664 10455
rect 11612 10412 11664 10421
rect 12072 10412 12124 10464
rect 12256 10412 12308 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 1492 10251 1544 10260
rect 1492 10217 1501 10251
rect 1501 10217 1535 10251
rect 1535 10217 1544 10251
rect 1492 10208 1544 10217
rect 1768 10251 1820 10260
rect 1768 10217 1777 10251
rect 1777 10217 1811 10251
rect 1811 10217 1820 10251
rect 1768 10208 1820 10217
rect 3884 10208 3936 10260
rect 3976 10208 4028 10260
rect 5908 10208 5960 10260
rect 6552 10251 6604 10260
rect 6552 10217 6561 10251
rect 6561 10217 6595 10251
rect 6595 10217 6604 10251
rect 6552 10208 6604 10217
rect 9588 10251 9640 10260
rect 9588 10217 9597 10251
rect 9597 10217 9631 10251
rect 9631 10217 9640 10251
rect 9588 10208 9640 10217
rect 12440 10208 12492 10260
rect 13544 10251 13596 10260
rect 13544 10217 13553 10251
rect 13553 10217 13587 10251
rect 13587 10217 13596 10251
rect 13544 10208 13596 10217
rect 16212 10208 16264 10260
rect 5540 10140 5592 10192
rect 7472 10140 7524 10192
rect 10508 10140 10560 10192
rect 3608 10072 3660 10124
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 2412 10004 2464 10056
rect 5724 10072 5776 10124
rect 5816 10072 5868 10124
rect 6552 10072 6604 10124
rect 6920 10072 6972 10124
rect 7104 10072 7156 10124
rect 5264 10047 5316 10056
rect 5264 10013 5273 10047
rect 5273 10013 5307 10047
rect 5307 10013 5316 10047
rect 5264 10004 5316 10013
rect 5448 10004 5500 10056
rect 2228 9936 2280 9988
rect 2596 9936 2648 9988
rect 2964 9979 3016 9988
rect 2964 9945 2982 9979
rect 2982 9945 3016 9979
rect 2964 9936 3016 9945
rect 5080 9936 5132 9988
rect 5908 9936 5960 9988
rect 7012 10004 7064 10056
rect 10600 10072 10652 10124
rect 14740 10072 14792 10124
rect 8484 10004 8536 10056
rect 12164 10047 12216 10056
rect 12164 10013 12173 10047
rect 12173 10013 12207 10047
rect 12207 10013 12216 10047
rect 12164 10004 12216 10013
rect 8392 9936 8444 9988
rect 1860 9911 1912 9920
rect 1860 9877 1869 9911
rect 1869 9877 1903 9911
rect 1903 9877 1912 9911
rect 1860 9868 1912 9877
rect 3792 9868 3844 9920
rect 5540 9911 5592 9920
rect 5540 9877 5549 9911
rect 5549 9877 5583 9911
rect 5583 9877 5592 9911
rect 5540 9868 5592 9877
rect 5632 9868 5684 9920
rect 6644 9868 6696 9920
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 9680 9868 9732 9920
rect 10232 9868 10284 9920
rect 10692 9868 10744 9920
rect 11060 9936 11112 9988
rect 11152 9868 11204 9920
rect 11704 9868 11756 9920
rect 12808 10004 12860 10056
rect 14648 10004 14700 10056
rect 15292 9868 15344 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 1860 9664 1912 9716
rect 3056 9664 3108 9716
rect 5264 9664 5316 9716
rect 7104 9664 7156 9716
rect 9128 9664 9180 9716
rect 9496 9664 9548 9716
rect 10508 9664 10560 9716
rect 13268 9664 13320 9716
rect 14280 9664 14332 9716
rect 1768 9596 1820 9648
rect 4160 9639 4212 9648
rect 1492 9571 1544 9580
rect 1492 9537 1501 9571
rect 1501 9537 1535 9571
rect 1535 9537 1544 9571
rect 1492 9528 1544 9537
rect 2872 9571 2924 9580
rect 2872 9537 2881 9571
rect 2881 9537 2915 9571
rect 2915 9537 2924 9571
rect 2872 9528 2924 9537
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 3884 9528 3936 9580
rect 4160 9605 4169 9639
rect 4169 9605 4203 9639
rect 4203 9605 4212 9639
rect 4160 9596 4212 9605
rect 4436 9596 4488 9648
rect 5080 9596 5132 9648
rect 4804 9528 4856 9580
rect 2412 9460 2464 9512
rect 5448 9528 5500 9580
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 5908 9503 5960 9512
rect 5908 9469 5917 9503
rect 5917 9469 5951 9503
rect 5951 9469 5960 9503
rect 5908 9460 5960 9469
rect 6000 9460 6052 9512
rect 6736 9596 6788 9648
rect 8024 9571 8076 9580
rect 8024 9537 8042 9571
rect 8042 9537 8076 9571
rect 8024 9528 8076 9537
rect 8208 9528 8260 9580
rect 8484 9596 8536 9648
rect 9680 9596 9732 9648
rect 9956 9596 10008 9648
rect 11060 9596 11112 9648
rect 14372 9596 14424 9648
rect 14740 9596 14792 9648
rect 6920 9460 6972 9512
rect 10508 9571 10560 9580
rect 10508 9537 10517 9571
rect 10517 9537 10551 9571
rect 10551 9537 10560 9571
rect 10508 9528 10560 9537
rect 11888 9571 11940 9580
rect 11888 9537 11897 9571
rect 11897 9537 11931 9571
rect 11931 9537 11940 9571
rect 11888 9528 11940 9537
rect 13544 9571 13596 9580
rect 13544 9537 13553 9571
rect 13553 9537 13587 9571
rect 13587 9537 13596 9571
rect 13544 9528 13596 9537
rect 10324 9460 10376 9512
rect 11704 9503 11756 9512
rect 1584 9392 1636 9444
rect 2136 9367 2188 9376
rect 2136 9333 2145 9367
rect 2145 9333 2179 9367
rect 2179 9333 2188 9367
rect 2136 9324 2188 9333
rect 2228 9367 2280 9376
rect 2228 9333 2237 9367
rect 2237 9333 2271 9367
rect 2271 9333 2280 9367
rect 2688 9392 2740 9444
rect 10048 9392 10100 9444
rect 4988 9367 5040 9376
rect 2228 9324 2280 9333
rect 4988 9333 4997 9367
rect 4997 9333 5031 9367
rect 5031 9333 5040 9367
rect 4988 9324 5040 9333
rect 5264 9324 5316 9376
rect 6552 9324 6604 9376
rect 6736 9324 6788 9376
rect 9128 9324 9180 9376
rect 10140 9367 10192 9376
rect 10140 9333 10149 9367
rect 10149 9333 10183 9367
rect 10183 9333 10192 9367
rect 10140 9324 10192 9333
rect 10232 9324 10284 9376
rect 11704 9469 11713 9503
rect 11713 9469 11747 9503
rect 11747 9469 11756 9503
rect 11704 9460 11756 9469
rect 12072 9460 12124 9512
rect 14372 9460 14424 9512
rect 12624 9392 12676 9444
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 2780 9120 2832 9172
rect 3976 9120 4028 9172
rect 5264 9120 5316 9172
rect 2872 9052 2924 9104
rect 5908 9120 5960 9172
rect 7840 9120 7892 9172
rect 8576 9120 8628 9172
rect 1952 9027 2004 9036
rect 1952 8993 1961 9027
rect 1961 8993 1995 9027
rect 1995 8993 2004 9027
rect 1952 8984 2004 8993
rect 3056 8984 3108 9036
rect 8300 9052 8352 9104
rect 5724 8984 5776 9036
rect 2872 8916 2924 8968
rect 2964 8959 3016 8968
rect 2964 8925 2973 8959
rect 2973 8925 3007 8959
rect 3007 8925 3016 8959
rect 2964 8916 3016 8925
rect 3240 8916 3292 8968
rect 3424 8916 3476 8968
rect 3884 8916 3936 8968
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 2504 8823 2556 8832
rect 2504 8789 2513 8823
rect 2513 8789 2547 8823
rect 2547 8789 2556 8823
rect 2504 8780 2556 8789
rect 3976 8848 4028 8900
rect 6644 8916 6696 8968
rect 3240 8780 3292 8832
rect 3884 8780 3936 8832
rect 4160 8823 4212 8832
rect 4160 8789 4169 8823
rect 4169 8789 4203 8823
rect 4203 8789 4212 8823
rect 4160 8780 4212 8789
rect 4252 8823 4304 8832
rect 4252 8789 4261 8823
rect 4261 8789 4295 8823
rect 4295 8789 4304 8823
rect 4712 8848 4764 8900
rect 5908 8848 5960 8900
rect 4252 8780 4304 8789
rect 6736 8780 6788 8832
rect 7472 8823 7524 8832
rect 7472 8789 7481 8823
rect 7481 8789 7515 8823
rect 7515 8789 7524 8823
rect 10508 9120 10560 9172
rect 11888 9120 11940 9172
rect 10600 9052 10652 9104
rect 17776 9052 17828 9104
rect 8576 8916 8628 8968
rect 11060 8984 11112 9036
rect 11152 8984 11204 9036
rect 11704 8984 11756 9036
rect 13820 8984 13872 9036
rect 15568 8984 15620 9036
rect 7472 8780 7524 8789
rect 8484 8823 8536 8832
rect 8484 8789 8493 8823
rect 8493 8789 8527 8823
rect 8527 8789 8536 8823
rect 8484 8780 8536 8789
rect 8760 8848 8812 8900
rect 9128 8848 9180 8900
rect 10232 8848 10284 8900
rect 10600 8916 10652 8968
rect 11796 8959 11848 8968
rect 11796 8925 11805 8959
rect 11805 8925 11839 8959
rect 11839 8925 11848 8959
rect 11796 8916 11848 8925
rect 13452 8959 13504 8968
rect 13452 8925 13461 8959
rect 13461 8925 13495 8959
rect 13495 8925 13504 8959
rect 13452 8916 13504 8925
rect 14372 8916 14424 8968
rect 14832 8916 14884 8968
rect 12808 8848 12860 8900
rect 12992 8891 13044 8900
rect 12992 8857 13001 8891
rect 13001 8857 13035 8891
rect 13035 8857 13044 8891
rect 12992 8848 13044 8857
rect 13636 8848 13688 8900
rect 10600 8823 10652 8832
rect 10600 8789 10609 8823
rect 10609 8789 10643 8823
rect 10643 8789 10652 8823
rect 10600 8780 10652 8789
rect 10968 8780 11020 8832
rect 14280 8780 14332 8832
rect 14924 8848 14976 8900
rect 14556 8780 14608 8832
rect 15016 8780 15068 8832
rect 15384 8780 15436 8832
rect 16396 8823 16448 8832
rect 16396 8789 16405 8823
rect 16405 8789 16439 8823
rect 16439 8789 16448 8823
rect 16396 8780 16448 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 1952 8576 2004 8628
rect 4160 8576 4212 8628
rect 4988 8576 5040 8628
rect 5632 8576 5684 8628
rect 5816 8576 5868 8628
rect 7564 8576 7616 8628
rect 7840 8576 7892 8628
rect 8024 8576 8076 8628
rect 8300 8576 8352 8628
rect 9312 8576 9364 8628
rect 10140 8576 10192 8628
rect 10324 8576 10376 8628
rect 10968 8619 11020 8628
rect 10968 8585 10977 8619
rect 10977 8585 11011 8619
rect 11011 8585 11020 8619
rect 10968 8576 11020 8585
rect 11060 8576 11112 8628
rect 12072 8576 12124 8628
rect 12716 8576 12768 8628
rect 13728 8576 13780 8628
rect 14464 8576 14516 8628
rect 15568 8619 15620 8628
rect 15568 8585 15577 8619
rect 15577 8585 15611 8619
rect 15611 8585 15620 8619
rect 15568 8576 15620 8585
rect 2320 8508 2372 8560
rect 3056 8508 3108 8560
rect 2964 8440 3016 8492
rect 3424 8440 3476 8492
rect 4160 8440 4212 8492
rect 4436 8440 4488 8492
rect 4620 8440 4672 8492
rect 5724 8508 5776 8560
rect 6644 8508 6696 8560
rect 9220 8508 9272 8560
rect 4896 8440 4948 8492
rect 7104 8440 7156 8492
rect 7472 8483 7524 8492
rect 7472 8449 7481 8483
rect 7481 8449 7515 8483
rect 7515 8449 7524 8483
rect 7472 8440 7524 8449
rect 9128 8483 9180 8492
rect 9128 8449 9137 8483
rect 9137 8449 9171 8483
rect 9171 8449 9180 8483
rect 9128 8440 9180 8449
rect 11060 8483 11112 8492
rect 4712 8372 4764 8424
rect 1860 8304 1912 8356
rect 5908 8304 5960 8356
rect 8760 8372 8812 8424
rect 11060 8449 11069 8483
rect 11069 8449 11103 8483
rect 11103 8449 11112 8483
rect 11060 8440 11112 8449
rect 10600 8372 10652 8424
rect 12164 8508 12216 8560
rect 11704 8415 11756 8424
rect 11704 8381 11713 8415
rect 11713 8381 11747 8415
rect 11747 8381 11756 8415
rect 11704 8372 11756 8381
rect 11796 8415 11848 8424
rect 11796 8381 11805 8415
rect 11805 8381 11839 8415
rect 11839 8381 11848 8415
rect 11796 8372 11848 8381
rect 12716 8304 12768 8356
rect 10600 8279 10652 8288
rect 10600 8245 10609 8279
rect 10609 8245 10643 8279
rect 10643 8245 10652 8279
rect 10600 8236 10652 8245
rect 13820 8440 13872 8492
rect 13820 8304 13872 8356
rect 14372 8236 14424 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 1492 8032 1544 8084
rect 2872 8075 2924 8084
rect 2872 8041 2881 8075
rect 2881 8041 2915 8075
rect 2915 8041 2924 8075
rect 2872 8032 2924 8041
rect 4252 8032 4304 8084
rect 5172 8075 5224 8084
rect 5172 8041 5181 8075
rect 5181 8041 5215 8075
rect 5215 8041 5224 8075
rect 5172 8032 5224 8041
rect 5724 8075 5776 8084
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 5816 8032 5868 8084
rect 7104 8075 7156 8084
rect 2872 7896 2924 7948
rect 3424 7939 3476 7948
rect 3424 7905 3433 7939
rect 3433 7905 3467 7939
rect 3467 7905 3476 7939
rect 3424 7896 3476 7905
rect 6552 7964 6604 8016
rect 7104 8041 7113 8075
rect 7113 8041 7147 8075
rect 7147 8041 7156 8075
rect 7104 8032 7156 8041
rect 9128 8032 9180 8084
rect 12900 8032 12952 8084
rect 8668 7964 8720 8016
rect 14924 8032 14976 8084
rect 15200 7964 15252 8016
rect 2228 7828 2280 7880
rect 2780 7871 2832 7880
rect 2780 7837 2789 7871
rect 2789 7837 2823 7871
rect 2823 7837 2832 7871
rect 2780 7828 2832 7837
rect 3240 7871 3292 7880
rect 3240 7837 3249 7871
rect 3249 7837 3283 7871
rect 3283 7837 3292 7871
rect 3240 7828 3292 7837
rect 3332 7871 3384 7880
rect 3332 7837 3341 7871
rect 3341 7837 3375 7871
rect 3375 7837 3384 7871
rect 5632 7896 5684 7948
rect 9128 7896 9180 7948
rect 9404 7896 9456 7948
rect 9956 7896 10008 7948
rect 3332 7828 3384 7837
rect 2228 7692 2280 7744
rect 3332 7692 3384 7744
rect 4252 7735 4304 7744
rect 4252 7701 4261 7735
rect 4261 7701 4295 7735
rect 4295 7701 4304 7735
rect 4252 7692 4304 7701
rect 4712 7735 4764 7744
rect 4712 7701 4721 7735
rect 4721 7701 4755 7735
rect 4755 7701 4764 7735
rect 4712 7692 4764 7701
rect 7564 7828 7616 7880
rect 7932 7871 7984 7880
rect 7932 7837 7941 7871
rect 7941 7837 7975 7871
rect 7975 7837 7984 7871
rect 7932 7828 7984 7837
rect 10416 7871 10468 7880
rect 5080 7760 5132 7812
rect 5540 7760 5592 7812
rect 7012 7803 7064 7812
rect 7012 7769 7021 7803
rect 7021 7769 7055 7803
rect 7055 7769 7064 7803
rect 7012 7760 7064 7769
rect 10416 7837 10425 7871
rect 10425 7837 10459 7871
rect 10459 7837 10468 7871
rect 10416 7828 10468 7837
rect 6552 7692 6604 7744
rect 6828 7692 6880 7744
rect 12164 7803 12216 7812
rect 12164 7769 12173 7803
rect 12173 7769 12207 7803
rect 12207 7769 12216 7803
rect 12164 7760 12216 7769
rect 13820 7896 13872 7948
rect 14280 7896 14332 7948
rect 14464 7896 14516 7948
rect 12808 7828 12860 7880
rect 13636 7871 13688 7880
rect 13636 7837 13645 7871
rect 13645 7837 13679 7871
rect 13679 7837 13688 7871
rect 13636 7828 13688 7837
rect 16396 7828 16448 7880
rect 13728 7760 13780 7812
rect 14556 7760 14608 7812
rect 8576 7735 8628 7744
rect 8576 7701 8585 7735
rect 8585 7701 8619 7735
rect 8619 7701 8628 7735
rect 8576 7692 8628 7701
rect 9128 7735 9180 7744
rect 9128 7701 9137 7735
rect 9137 7701 9171 7735
rect 9171 7701 9180 7735
rect 9128 7692 9180 7701
rect 9588 7735 9640 7744
rect 9588 7701 9597 7735
rect 9597 7701 9631 7735
rect 9631 7701 9640 7735
rect 9588 7692 9640 7701
rect 10232 7735 10284 7744
rect 10232 7701 10241 7735
rect 10241 7701 10275 7735
rect 10275 7701 10284 7735
rect 10232 7692 10284 7701
rect 10968 7692 11020 7744
rect 12624 7692 12676 7744
rect 13084 7692 13136 7744
rect 16948 7692 17000 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 2504 7488 2556 7540
rect 3056 7488 3108 7540
rect 3240 7488 3292 7540
rect 3516 7531 3568 7540
rect 3516 7497 3525 7531
rect 3525 7497 3559 7531
rect 3559 7497 3568 7531
rect 3516 7488 3568 7497
rect 3884 7420 3936 7472
rect 4988 7488 5040 7540
rect 5448 7531 5500 7540
rect 5448 7497 5457 7531
rect 5457 7497 5491 7531
rect 5491 7497 5500 7531
rect 5448 7488 5500 7497
rect 6000 7488 6052 7540
rect 8208 7488 8260 7540
rect 8484 7488 8536 7540
rect 6920 7420 6972 7472
rect 8576 7420 8628 7472
rect 9496 7488 9548 7540
rect 9864 7488 9916 7540
rect 10048 7488 10100 7540
rect 10232 7488 10284 7540
rect 10876 7488 10928 7540
rect 12440 7488 12492 7540
rect 12532 7488 12584 7540
rect 13360 7531 13412 7540
rect 13360 7497 13369 7531
rect 13369 7497 13403 7531
rect 13403 7497 13412 7531
rect 13360 7488 13412 7497
rect 13728 7488 13780 7540
rect 15200 7531 15252 7540
rect 9220 7420 9272 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 1492 7284 1544 7336
rect 2320 7284 2372 7336
rect 2596 7284 2648 7336
rect 2504 7216 2556 7268
rect 3976 7395 4028 7404
rect 2964 7327 3016 7336
rect 2964 7293 2973 7327
rect 2973 7293 3007 7327
rect 3007 7293 3016 7327
rect 2964 7284 3016 7293
rect 3976 7361 3985 7395
rect 3985 7361 4019 7395
rect 4019 7361 4028 7395
rect 3976 7352 4028 7361
rect 4252 7352 4304 7404
rect 5356 7352 5408 7404
rect 6092 7352 6144 7404
rect 12164 7420 12216 7472
rect 15200 7497 15209 7531
rect 15209 7497 15243 7531
rect 15243 7497 15252 7531
rect 15200 7488 15252 7497
rect 15936 7488 15988 7540
rect 3332 7284 3384 7336
rect 3424 7284 3476 7336
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 5448 7284 5500 7336
rect 5724 7284 5776 7336
rect 6000 7327 6052 7336
rect 6000 7293 6009 7327
rect 6009 7293 6043 7327
rect 6043 7293 6052 7327
rect 6552 7327 6604 7336
rect 6000 7284 6052 7293
rect 6552 7293 6561 7327
rect 6561 7293 6595 7327
rect 6595 7293 6604 7327
rect 6552 7284 6604 7293
rect 4252 7148 4304 7200
rect 4436 7191 4488 7200
rect 4436 7157 4445 7191
rect 4445 7157 4479 7191
rect 4479 7157 4488 7191
rect 4436 7148 4488 7157
rect 9864 7352 9916 7404
rect 12624 7395 12676 7404
rect 16304 7420 16356 7472
rect 12624 7361 12642 7395
rect 12642 7361 12676 7395
rect 12624 7352 12676 7361
rect 13452 7352 13504 7404
rect 7288 7327 7340 7336
rect 7288 7293 7297 7327
rect 7297 7293 7331 7327
rect 7331 7293 7340 7327
rect 7288 7284 7340 7293
rect 9496 7327 9548 7336
rect 9496 7293 9505 7327
rect 9505 7293 9539 7327
rect 9539 7293 9548 7327
rect 10140 7327 10192 7336
rect 9496 7284 9548 7293
rect 10140 7293 10149 7327
rect 10149 7293 10183 7327
rect 10183 7293 10192 7327
rect 10140 7284 10192 7293
rect 7104 7191 7156 7200
rect 7104 7157 7113 7191
rect 7113 7157 7147 7191
rect 7147 7157 7156 7191
rect 7104 7148 7156 7157
rect 7196 7148 7248 7200
rect 9220 7148 9272 7200
rect 9956 7216 10008 7268
rect 13084 7327 13136 7336
rect 13084 7293 13093 7327
rect 13093 7293 13127 7327
rect 13127 7293 13136 7327
rect 13084 7284 13136 7293
rect 13820 7284 13872 7336
rect 14464 7284 14516 7336
rect 10692 7216 10744 7268
rect 10784 7191 10836 7200
rect 10784 7157 10793 7191
rect 10793 7157 10827 7191
rect 10827 7157 10836 7191
rect 10784 7148 10836 7157
rect 10876 7191 10928 7200
rect 10876 7157 10885 7191
rect 10885 7157 10919 7191
rect 10919 7157 10928 7191
rect 15016 7216 15068 7268
rect 10876 7148 10928 7157
rect 16396 7148 16448 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 3332 6944 3384 6996
rect 4160 6944 4212 6996
rect 4436 6944 4488 6996
rect 5172 6944 5224 6996
rect 5724 6944 5776 6996
rect 6092 6987 6144 6996
rect 6092 6953 6101 6987
rect 6101 6953 6135 6987
rect 6135 6953 6144 6987
rect 6092 6944 6144 6953
rect 3976 6876 4028 6928
rect 1768 6808 1820 6860
rect 2504 6808 2556 6860
rect 3424 6851 3476 6860
rect 3424 6817 3433 6851
rect 3433 6817 3467 6851
rect 3467 6817 3476 6851
rect 3424 6808 3476 6817
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 1676 6783 1728 6792
rect 1676 6749 1685 6783
rect 1685 6749 1719 6783
rect 1719 6749 1728 6783
rect 1676 6740 1728 6749
rect 3700 6740 3752 6792
rect 4344 6808 4396 6860
rect 4988 6876 5040 6928
rect 5356 6876 5408 6928
rect 7196 6944 7248 6996
rect 7380 6944 7432 6996
rect 7932 6944 7984 6996
rect 9128 6944 9180 6996
rect 10048 6944 10100 6996
rect 10876 6944 10928 6996
rect 13452 6944 13504 6996
rect 4896 6808 4948 6860
rect 5448 6851 5500 6860
rect 5448 6817 5457 6851
rect 5457 6817 5491 6851
rect 5491 6817 5500 6851
rect 5448 6808 5500 6817
rect 7472 6808 7524 6860
rect 7748 6808 7800 6860
rect 8484 6876 8536 6928
rect 8944 6919 8996 6928
rect 8944 6885 8953 6919
rect 8953 6885 8987 6919
rect 8987 6885 8996 6919
rect 8944 6876 8996 6885
rect 10324 6876 10376 6928
rect 5632 6740 5684 6792
rect 6000 6740 6052 6792
rect 7288 6740 7340 6792
rect 8760 6808 8812 6860
rect 9864 6808 9916 6860
rect 10140 6808 10192 6860
rect 10232 6808 10284 6860
rect 14372 6876 14424 6928
rect 12808 6851 12860 6860
rect 12808 6817 12817 6851
rect 12817 6817 12851 6851
rect 12851 6817 12860 6851
rect 12808 6808 12860 6817
rect 12900 6808 12952 6860
rect 15660 6944 15712 6996
rect 1768 6604 1820 6656
rect 6552 6672 6604 6724
rect 2964 6604 3016 6656
rect 3240 6647 3292 6656
rect 3240 6613 3249 6647
rect 3249 6613 3283 6647
rect 3283 6613 3292 6647
rect 3240 6604 3292 6613
rect 3332 6647 3384 6656
rect 3332 6613 3341 6647
rect 3341 6613 3375 6647
rect 3375 6613 3384 6647
rect 3792 6647 3844 6656
rect 3332 6604 3384 6613
rect 3792 6613 3801 6647
rect 3801 6613 3835 6647
rect 3835 6613 3844 6647
rect 3792 6604 3844 6613
rect 4528 6604 4580 6656
rect 5540 6604 5592 6656
rect 6644 6604 6696 6656
rect 8392 6740 8444 6792
rect 9588 6783 9640 6792
rect 9588 6749 9597 6783
rect 9597 6749 9631 6783
rect 9631 6749 9640 6783
rect 9588 6740 9640 6749
rect 10968 6740 11020 6792
rect 12348 6783 12400 6792
rect 12348 6749 12357 6783
rect 12357 6749 12391 6783
rect 12391 6749 12400 6783
rect 12348 6740 12400 6749
rect 13360 6740 13412 6792
rect 13636 6740 13688 6792
rect 15752 6808 15804 6860
rect 15660 6740 15712 6792
rect 7932 6672 7984 6724
rect 8208 6672 8260 6724
rect 8668 6672 8720 6724
rect 9496 6672 9548 6724
rect 7656 6647 7708 6656
rect 7656 6613 7665 6647
rect 7665 6613 7699 6647
rect 7699 6613 7708 6647
rect 8116 6647 8168 6656
rect 7656 6604 7708 6613
rect 8116 6613 8125 6647
rect 8125 6613 8159 6647
rect 8159 6613 8168 6647
rect 8116 6604 8168 6613
rect 9312 6604 9364 6656
rect 9956 6604 10008 6656
rect 10140 6647 10192 6656
rect 10140 6613 10149 6647
rect 10149 6613 10183 6647
rect 10183 6613 10192 6647
rect 10140 6604 10192 6613
rect 15476 6672 15528 6724
rect 16212 6715 16264 6724
rect 16212 6681 16221 6715
rect 16221 6681 16255 6715
rect 16255 6681 16264 6715
rect 16212 6672 16264 6681
rect 10784 6604 10836 6656
rect 11244 6604 11296 6656
rect 11704 6604 11756 6656
rect 11796 6647 11848 6656
rect 11796 6613 11805 6647
rect 11805 6613 11839 6647
rect 11839 6613 11848 6647
rect 13912 6647 13964 6656
rect 11796 6604 11848 6613
rect 13912 6613 13921 6647
rect 13921 6613 13955 6647
rect 13955 6613 13964 6647
rect 13912 6604 13964 6613
rect 14740 6604 14792 6656
rect 15660 6604 15712 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 2596 6400 2648 6452
rect 3148 6400 3200 6452
rect 3792 6443 3844 6452
rect 3792 6409 3801 6443
rect 3801 6409 3835 6443
rect 3835 6409 3844 6443
rect 3792 6400 3844 6409
rect 4344 6400 4396 6452
rect 4804 6400 4856 6452
rect 6552 6400 6604 6452
rect 7104 6443 7156 6452
rect 7104 6409 7113 6443
rect 7113 6409 7147 6443
rect 7147 6409 7156 6443
rect 7104 6400 7156 6409
rect 7656 6400 7708 6452
rect 8576 6400 8628 6452
rect 8760 6400 8812 6452
rect 9588 6400 9640 6452
rect 11888 6400 11940 6452
rect 12992 6443 13044 6452
rect 12992 6409 13001 6443
rect 13001 6409 13035 6443
rect 13035 6409 13044 6443
rect 12992 6400 13044 6409
rect 13912 6400 13964 6452
rect 16396 6400 16448 6452
rect 21364 6443 21416 6452
rect 21364 6409 21373 6443
rect 21373 6409 21407 6443
rect 21407 6409 21416 6443
rect 21364 6400 21416 6409
rect 1584 6264 1636 6316
rect 2688 6332 2740 6384
rect 2780 6332 2832 6384
rect 1952 6264 2004 6316
rect 2780 6060 2832 6112
rect 4528 6264 4580 6316
rect 5448 6332 5500 6384
rect 5816 6332 5868 6384
rect 3056 6128 3108 6180
rect 3424 6196 3476 6248
rect 4804 6239 4856 6248
rect 4804 6205 4813 6239
rect 4813 6205 4847 6239
rect 4847 6205 4856 6239
rect 4804 6196 4856 6205
rect 7380 6239 7432 6248
rect 7380 6205 7389 6239
rect 7389 6205 7423 6239
rect 7423 6205 7432 6239
rect 7380 6196 7432 6205
rect 7748 6307 7800 6316
rect 7748 6273 7757 6307
rect 7757 6273 7791 6307
rect 7791 6273 7800 6307
rect 7748 6264 7800 6273
rect 8208 6264 8260 6316
rect 8300 6196 8352 6248
rect 8576 6239 8628 6248
rect 8576 6205 8585 6239
rect 8585 6205 8619 6239
rect 8619 6205 8628 6239
rect 9128 6264 9180 6316
rect 8576 6196 8628 6205
rect 3700 6128 3752 6180
rect 4436 6128 4488 6180
rect 6920 6128 6972 6180
rect 8484 6128 8536 6180
rect 8852 6128 8904 6180
rect 5172 6060 5224 6112
rect 5540 6060 5592 6112
rect 6552 6103 6604 6112
rect 6552 6069 6561 6103
rect 6561 6069 6595 6103
rect 6595 6069 6604 6103
rect 6552 6060 6604 6069
rect 6644 6060 6696 6112
rect 7104 6060 7156 6112
rect 7932 6103 7984 6112
rect 7932 6069 7941 6103
rect 7941 6069 7975 6103
rect 7975 6069 7984 6103
rect 7932 6060 7984 6069
rect 8300 6060 8352 6112
rect 9404 6196 9456 6248
rect 11980 6332 12032 6384
rect 12900 6375 12952 6384
rect 12900 6341 12909 6375
rect 12909 6341 12943 6375
rect 12943 6341 12952 6375
rect 12900 6332 12952 6341
rect 15292 6332 15344 6384
rect 15568 6332 15620 6384
rect 9680 6264 9732 6316
rect 9864 6307 9916 6316
rect 9864 6273 9898 6307
rect 9898 6273 9916 6307
rect 9864 6264 9916 6273
rect 10692 6264 10744 6316
rect 10784 6264 10836 6316
rect 12532 6264 12584 6316
rect 13360 6307 13412 6316
rect 13360 6273 13369 6307
rect 13369 6273 13403 6307
rect 13403 6273 13412 6307
rect 13360 6264 13412 6273
rect 13636 6307 13688 6316
rect 13636 6273 13670 6307
rect 13670 6273 13688 6307
rect 13636 6264 13688 6273
rect 12900 6196 12952 6248
rect 11060 6128 11112 6180
rect 13268 6128 13320 6180
rect 9864 6060 9916 6112
rect 10232 6060 10284 6112
rect 11336 6060 11388 6112
rect 11612 6060 11664 6112
rect 11888 6103 11940 6112
rect 11888 6069 11897 6103
rect 11897 6069 11931 6103
rect 11931 6069 11940 6103
rect 11888 6060 11940 6069
rect 12348 6060 12400 6112
rect 13176 6103 13228 6112
rect 13176 6069 13185 6103
rect 13185 6069 13219 6103
rect 13219 6069 13228 6103
rect 13176 6060 13228 6069
rect 14648 6196 14700 6248
rect 15476 6264 15528 6316
rect 18052 6307 18104 6316
rect 18052 6273 18061 6307
rect 18061 6273 18095 6307
rect 18095 6273 18104 6307
rect 18052 6264 18104 6273
rect 21548 6307 21600 6316
rect 21548 6273 21557 6307
rect 21557 6273 21591 6307
rect 21591 6273 21600 6307
rect 21548 6264 21600 6273
rect 17224 6239 17276 6248
rect 17224 6205 17233 6239
rect 17233 6205 17267 6239
rect 17267 6205 17276 6239
rect 17224 6196 17276 6205
rect 18236 6128 18288 6180
rect 14740 6103 14792 6112
rect 14740 6069 14749 6103
rect 14749 6069 14783 6103
rect 14783 6069 14792 6103
rect 14740 6060 14792 6069
rect 14832 6103 14884 6112
rect 14832 6069 14841 6103
rect 14841 6069 14875 6103
rect 14875 6069 14884 6103
rect 15660 6103 15712 6112
rect 14832 6060 14884 6069
rect 15660 6069 15669 6103
rect 15669 6069 15703 6103
rect 15703 6069 15712 6103
rect 15660 6060 15712 6069
rect 16948 6060 17000 6112
rect 18696 6103 18748 6112
rect 18696 6069 18705 6103
rect 18705 6069 18739 6103
rect 18739 6069 18748 6103
rect 18696 6060 18748 6069
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 1952 5856 2004 5908
rect 2596 5856 2648 5908
rect 2228 5788 2280 5840
rect 4068 5856 4120 5908
rect 4436 5899 4488 5908
rect 4436 5865 4445 5899
rect 4445 5865 4479 5899
rect 4479 5865 4488 5899
rect 4436 5856 4488 5865
rect 3516 5788 3568 5840
rect 3608 5720 3660 5772
rect 5448 5856 5500 5908
rect 5908 5856 5960 5908
rect 6920 5856 6972 5908
rect 7288 5856 7340 5908
rect 1492 5627 1544 5636
rect 1492 5593 1501 5627
rect 1501 5593 1535 5627
rect 1535 5593 1544 5627
rect 1492 5584 1544 5593
rect 3056 5584 3108 5636
rect 2872 5516 2924 5568
rect 4252 5652 4304 5704
rect 4436 5652 4488 5704
rect 4896 5763 4948 5772
rect 4896 5729 4905 5763
rect 4905 5729 4939 5763
rect 4939 5729 4948 5763
rect 4896 5720 4948 5729
rect 7472 5788 7524 5840
rect 8944 5788 8996 5840
rect 11060 5788 11112 5840
rect 11612 5788 11664 5840
rect 12900 5856 12952 5908
rect 13268 5856 13320 5908
rect 9312 5720 9364 5772
rect 10508 5720 10560 5772
rect 11336 5720 11388 5772
rect 12532 5763 12584 5772
rect 4804 5652 4856 5704
rect 6000 5652 6052 5704
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 8760 5695 8812 5704
rect 7012 5652 7064 5661
rect 6828 5584 6880 5636
rect 8208 5627 8260 5636
rect 8208 5593 8226 5627
rect 8226 5593 8260 5627
rect 8208 5584 8260 5593
rect 8760 5661 8769 5695
rect 8769 5661 8803 5695
rect 8803 5661 8812 5695
rect 8760 5652 8812 5661
rect 9680 5652 9732 5704
rect 12532 5729 12541 5763
rect 12541 5729 12575 5763
rect 12575 5729 12584 5763
rect 12532 5720 12584 5729
rect 14832 5788 14884 5840
rect 15568 5831 15620 5840
rect 15568 5797 15577 5831
rect 15577 5797 15611 5831
rect 15611 5797 15620 5831
rect 15568 5788 15620 5797
rect 17132 5788 17184 5840
rect 14464 5695 14516 5704
rect 14464 5661 14473 5695
rect 14473 5661 14507 5695
rect 14507 5661 14516 5695
rect 14464 5652 14516 5661
rect 3608 5516 3660 5568
rect 3976 5516 4028 5568
rect 4344 5516 4396 5568
rect 5264 5516 5316 5568
rect 5724 5516 5776 5568
rect 7748 5516 7800 5568
rect 8484 5516 8536 5568
rect 8760 5516 8812 5568
rect 9128 5516 9180 5568
rect 9956 5584 10008 5636
rect 10232 5584 10284 5636
rect 10416 5627 10468 5636
rect 10416 5593 10425 5627
rect 10425 5593 10459 5627
rect 10459 5593 10468 5627
rect 10416 5584 10468 5593
rect 12716 5584 12768 5636
rect 12900 5584 12952 5636
rect 13268 5584 13320 5636
rect 15752 5652 15804 5704
rect 17040 5652 17092 5704
rect 11152 5516 11204 5568
rect 11888 5516 11940 5568
rect 13084 5516 13136 5568
rect 13636 5516 13688 5568
rect 16856 5584 16908 5636
rect 17868 5584 17920 5636
rect 18696 5584 18748 5636
rect 14096 5559 14148 5568
rect 14096 5525 14105 5559
rect 14105 5525 14139 5559
rect 14139 5525 14148 5559
rect 14096 5516 14148 5525
rect 14648 5516 14700 5568
rect 17224 5516 17276 5568
rect 19984 5516 20036 5568
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 1584 5355 1636 5364
rect 1584 5321 1593 5355
rect 1593 5321 1627 5355
rect 1627 5321 1636 5355
rect 1584 5312 1636 5321
rect 2688 5312 2740 5364
rect 3332 5312 3384 5364
rect 5540 5312 5592 5364
rect 5632 5312 5684 5364
rect 2136 5244 2188 5296
rect 2044 5176 2096 5228
rect 2596 5176 2648 5228
rect 3332 5176 3384 5228
rect 3792 5244 3844 5296
rect 7012 5312 7064 5364
rect 7196 5312 7248 5364
rect 7932 5312 7984 5364
rect 8116 5312 8168 5364
rect 8576 5355 8628 5364
rect 8576 5321 8585 5355
rect 8585 5321 8619 5355
rect 8619 5321 8628 5355
rect 8576 5312 8628 5321
rect 9772 5312 9824 5364
rect 10416 5355 10468 5364
rect 10416 5321 10425 5355
rect 10425 5321 10459 5355
rect 10459 5321 10468 5355
rect 10416 5312 10468 5321
rect 11152 5312 11204 5364
rect 11244 5312 11296 5364
rect 11888 5312 11940 5364
rect 14096 5355 14148 5364
rect 7288 5244 7340 5296
rect 8300 5244 8352 5296
rect 8668 5244 8720 5296
rect 11060 5244 11112 5296
rect 14096 5321 14105 5355
rect 14105 5321 14139 5355
rect 14139 5321 14148 5355
rect 14096 5312 14148 5321
rect 15200 5355 15252 5364
rect 15200 5321 15209 5355
rect 15209 5321 15243 5355
rect 15243 5321 15252 5355
rect 15200 5312 15252 5321
rect 4436 5219 4488 5228
rect 4436 5185 4445 5219
rect 4445 5185 4479 5219
rect 4479 5185 4488 5219
rect 4436 5176 4488 5185
rect 4804 5219 4856 5228
rect 4804 5185 4813 5219
rect 4813 5185 4847 5219
rect 4847 5185 4856 5219
rect 4804 5176 4856 5185
rect 4896 5176 4948 5228
rect 5356 5176 5408 5228
rect 6460 5176 6512 5228
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 7656 5219 7708 5228
rect 6736 5176 6788 5185
rect 7656 5185 7665 5219
rect 7665 5185 7699 5219
rect 7699 5185 7708 5219
rect 7656 5176 7708 5185
rect 1860 5108 1912 5160
rect 1952 5151 2004 5160
rect 1952 5117 1961 5151
rect 1961 5117 1995 5151
rect 1995 5117 2004 5151
rect 1952 5108 2004 5117
rect 3056 5040 3108 5092
rect 3976 5108 4028 5160
rect 5908 5108 5960 5160
rect 6920 5108 6972 5160
rect 1768 5015 1820 5024
rect 1768 4981 1777 5015
rect 1777 4981 1811 5015
rect 1811 4981 1820 5015
rect 1768 4972 1820 4981
rect 3240 4972 3292 5024
rect 3792 5040 3844 5092
rect 4344 5040 4396 5092
rect 6828 5040 6880 5092
rect 8484 5176 8536 5228
rect 9404 5176 9456 5228
rect 9956 5219 10008 5228
rect 9956 5185 9965 5219
rect 9965 5185 9999 5219
rect 9999 5185 10008 5219
rect 9956 5176 10008 5185
rect 10048 5176 10100 5228
rect 10416 5176 10468 5228
rect 11152 5176 11204 5228
rect 8300 5108 8352 5160
rect 10692 5151 10744 5160
rect 4252 4972 4304 5024
rect 6736 4972 6788 5024
rect 7472 4972 7524 5024
rect 8300 5015 8352 5024
rect 8300 4981 8309 5015
rect 8309 4981 8343 5015
rect 8343 4981 8352 5015
rect 8300 4972 8352 4981
rect 10692 5117 10701 5151
rect 10701 5117 10735 5151
rect 10735 5117 10744 5151
rect 10692 5108 10744 5117
rect 11244 5108 11296 5160
rect 11520 5108 11572 5160
rect 12256 5176 12308 5228
rect 15292 5244 15344 5296
rect 12624 5176 12676 5228
rect 13268 5219 13320 5228
rect 13268 5185 13277 5219
rect 13277 5185 13311 5219
rect 13311 5185 13320 5219
rect 13268 5176 13320 5185
rect 12808 5108 12860 5160
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 13728 5108 13780 5160
rect 14740 5176 14792 5228
rect 15200 5176 15252 5228
rect 17040 5244 17092 5296
rect 17132 5244 17184 5296
rect 17960 5244 18012 5296
rect 9956 4972 10008 5024
rect 10232 4972 10284 5024
rect 10784 4972 10836 5024
rect 10876 4972 10928 5024
rect 11520 4972 11572 5024
rect 12348 4972 12400 5024
rect 12900 5040 12952 5092
rect 15752 5108 15804 5160
rect 17868 5176 17920 5228
rect 19984 5219 20036 5228
rect 17776 5108 17828 5160
rect 19984 5185 19993 5219
rect 19993 5185 20027 5219
rect 20027 5185 20036 5219
rect 19984 5176 20036 5185
rect 14372 5040 14424 5092
rect 14464 5015 14516 5024
rect 14464 4981 14473 5015
rect 14473 4981 14507 5015
rect 14507 4981 14516 5015
rect 14464 4972 14516 4981
rect 14832 5015 14884 5024
rect 14832 4981 14841 5015
rect 14841 4981 14875 5015
rect 14875 4981 14884 5015
rect 14832 4972 14884 4981
rect 16672 4972 16724 5024
rect 18052 5015 18104 5024
rect 18052 4981 18061 5015
rect 18061 4981 18095 5015
rect 18095 4981 18104 5015
rect 18052 4972 18104 4981
rect 20904 4972 20956 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 2044 4768 2096 4820
rect 2320 4768 2372 4820
rect 2964 4768 3016 4820
rect 3884 4768 3936 4820
rect 4160 4768 4212 4820
rect 4436 4768 4488 4820
rect 4988 4768 5040 4820
rect 5264 4768 5316 4820
rect 5816 4768 5868 4820
rect 6828 4768 6880 4820
rect 7656 4768 7708 4820
rect 8208 4768 8260 4820
rect 10692 4768 10744 4820
rect 11428 4811 11480 4820
rect 3056 4700 3108 4752
rect 3148 4700 3200 4752
rect 2504 4632 2556 4684
rect 4712 4700 4764 4752
rect 6552 4700 6604 4752
rect 6736 4700 6788 4752
rect 1584 4564 1636 4616
rect 1676 4564 1728 4616
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 2688 4496 2740 4548
rect 2872 4496 2924 4548
rect 4896 4632 4948 4684
rect 6920 4675 6972 4684
rect 6920 4641 6929 4675
rect 6929 4641 6963 4675
rect 6963 4641 6972 4675
rect 6920 4632 6972 4641
rect 3240 4564 3292 4616
rect 4068 4496 4120 4548
rect 4620 4539 4672 4548
rect 4620 4505 4629 4539
rect 4629 4505 4663 4539
rect 4663 4505 4672 4539
rect 4620 4496 4672 4505
rect 4712 4496 4764 4548
rect 6092 4564 6144 4616
rect 6276 4564 6328 4616
rect 8116 4700 8168 4752
rect 11428 4777 11437 4811
rect 11437 4777 11471 4811
rect 11471 4777 11480 4811
rect 11428 4768 11480 4777
rect 11704 4768 11756 4820
rect 13268 4768 13320 4820
rect 13728 4768 13780 4820
rect 7380 4632 7432 4684
rect 7840 4632 7892 4684
rect 8576 4632 8628 4684
rect 8024 4564 8076 4616
rect 8392 4564 8444 4616
rect 9128 4632 9180 4684
rect 10876 4675 10928 4684
rect 10876 4641 10885 4675
rect 10885 4641 10919 4675
rect 10919 4641 10928 4675
rect 10876 4632 10928 4641
rect 11060 4632 11112 4684
rect 10140 4564 10192 4616
rect 8208 4496 8260 4548
rect 8760 4496 8812 4548
rect 9220 4496 9272 4548
rect 9496 4496 9548 4548
rect 11060 4539 11112 4548
rect 3148 4471 3200 4480
rect 3148 4437 3157 4471
rect 3157 4437 3191 4471
rect 3191 4437 3200 4471
rect 3148 4428 3200 4437
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 3884 4428 3936 4480
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 5448 4428 5500 4480
rect 5724 4428 5776 4480
rect 6552 4428 6604 4480
rect 7748 4428 7800 4480
rect 7840 4428 7892 4480
rect 8300 4428 8352 4480
rect 11060 4505 11069 4539
rect 11069 4505 11103 4539
rect 11103 4505 11112 4539
rect 11060 4496 11112 4505
rect 11428 4496 11480 4548
rect 13912 4700 13964 4752
rect 12716 4675 12768 4684
rect 12716 4641 12725 4675
rect 12725 4641 12759 4675
rect 12759 4641 12768 4675
rect 12716 4632 12768 4641
rect 12808 4632 12860 4684
rect 12532 4564 12584 4616
rect 15660 4675 15712 4684
rect 15660 4641 15669 4675
rect 15669 4641 15703 4675
rect 15703 4641 15712 4675
rect 18052 4768 18104 4820
rect 18144 4700 18196 4752
rect 15660 4632 15712 4641
rect 16672 4632 16724 4684
rect 17960 4675 18012 4684
rect 17960 4641 17969 4675
rect 17969 4641 18003 4675
rect 18003 4641 18012 4675
rect 17960 4632 18012 4641
rect 15476 4564 15528 4616
rect 16948 4564 17000 4616
rect 9680 4471 9732 4480
rect 9680 4437 9689 4471
rect 9689 4437 9723 4471
rect 9723 4437 9732 4471
rect 9680 4428 9732 4437
rect 10048 4428 10100 4480
rect 10324 4428 10376 4480
rect 10692 4428 10744 4480
rect 10876 4428 10928 4480
rect 12992 4539 13044 4548
rect 12992 4505 13001 4539
rect 13001 4505 13035 4539
rect 13035 4505 13044 4539
rect 12992 4496 13044 4505
rect 13728 4496 13780 4548
rect 12348 4428 12400 4480
rect 12440 4471 12492 4480
rect 12440 4437 12449 4471
rect 12449 4437 12483 4471
rect 12483 4437 12492 4471
rect 12440 4428 12492 4437
rect 12624 4428 12676 4480
rect 14188 4428 14240 4480
rect 14556 4471 14608 4480
rect 14556 4437 14565 4471
rect 14565 4437 14599 4471
rect 14599 4437 14608 4471
rect 14924 4471 14976 4480
rect 14556 4428 14608 4437
rect 14924 4437 14933 4471
rect 14933 4437 14967 4471
rect 14967 4437 14976 4471
rect 14924 4428 14976 4437
rect 15568 4428 15620 4480
rect 15844 4471 15896 4480
rect 15844 4437 15853 4471
rect 15853 4437 15887 4471
rect 15887 4437 15896 4471
rect 15844 4428 15896 4437
rect 17776 4539 17828 4548
rect 17776 4505 17785 4539
rect 17785 4505 17819 4539
rect 17819 4505 17828 4539
rect 17776 4496 17828 4505
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 2412 4267 2464 4276
rect 2412 4233 2421 4267
rect 2421 4233 2455 4267
rect 2455 4233 2464 4267
rect 2412 4224 2464 4233
rect 2872 4224 2924 4276
rect 3148 4224 3200 4276
rect 3240 4224 3292 4276
rect 664 4088 716 4140
rect 2044 4131 2096 4140
rect 2044 4097 2053 4131
rect 2053 4097 2087 4131
rect 2087 4097 2096 4131
rect 7104 4224 7156 4276
rect 7472 4224 7524 4276
rect 7748 4224 7800 4276
rect 10876 4267 10928 4276
rect 10876 4233 10885 4267
rect 10885 4233 10919 4267
rect 10919 4233 10928 4267
rect 10876 4224 10928 4233
rect 2044 4088 2096 4097
rect 3148 4088 3200 4140
rect 3240 4020 3292 4072
rect 4068 4088 4120 4140
rect 4436 4156 4488 4208
rect 4896 4156 4948 4208
rect 5264 4156 5316 4208
rect 7012 4156 7064 4208
rect 12716 4224 12768 4276
rect 15476 4224 15528 4276
rect 11060 4156 11112 4208
rect 14188 4156 14240 4208
rect 17960 4156 18012 4208
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 4252 4063 4304 4072
rect 1308 3952 1360 4004
rect 2228 3952 2280 4004
rect 3056 3952 3108 4004
rect 4252 4029 4261 4063
rect 4261 4029 4295 4063
rect 4295 4029 4304 4063
rect 4252 4020 4304 4029
rect 4344 4063 4396 4072
rect 4344 4029 4353 4063
rect 4353 4029 4387 4063
rect 4387 4029 4396 4063
rect 5264 4063 5316 4072
rect 4344 4020 4396 4029
rect 5264 4029 5273 4063
rect 5273 4029 5307 4063
rect 5307 4029 5316 4063
rect 5264 4020 5316 4029
rect 5448 4063 5500 4072
rect 5448 4029 5457 4063
rect 5457 4029 5491 4063
rect 5491 4029 5500 4063
rect 5448 4020 5500 4029
rect 6644 4088 6696 4140
rect 6920 4063 6972 4072
rect 6920 4029 6929 4063
rect 6929 4029 6963 4063
rect 6963 4029 6972 4063
rect 6920 4020 6972 4029
rect 4436 3952 4488 4004
rect 6644 3952 6696 4004
rect 8300 4088 8352 4140
rect 8484 4131 8536 4140
rect 8484 4097 8493 4131
rect 8493 4097 8527 4131
rect 8527 4097 8536 4131
rect 8484 4088 8536 4097
rect 9312 4131 9364 4140
rect 9312 4097 9321 4131
rect 9321 4097 9355 4131
rect 9355 4097 9364 4131
rect 9312 4088 9364 4097
rect 9956 4088 10008 4140
rect 12440 4088 12492 4140
rect 12532 4088 12584 4140
rect 13636 4088 13688 4140
rect 14280 4131 14332 4140
rect 14280 4097 14314 4131
rect 14314 4097 14332 4131
rect 14280 4088 14332 4097
rect 14740 4088 14792 4140
rect 20260 4088 20312 4140
rect 7656 4020 7708 4072
rect 8760 4063 8812 4072
rect 8208 3952 8260 4004
rect 8484 3952 8536 4004
rect 2044 3884 2096 3936
rect 4068 3884 4120 3936
rect 4620 3927 4672 3936
rect 4620 3893 4629 3927
rect 4629 3893 4663 3927
rect 4663 3893 4672 3927
rect 4620 3884 4672 3893
rect 4804 3927 4856 3936
rect 4804 3893 4813 3927
rect 4813 3893 4847 3927
rect 4847 3893 4856 3927
rect 4804 3884 4856 3893
rect 5816 3884 5868 3936
rect 7104 3884 7156 3936
rect 7380 3884 7432 3936
rect 8024 3927 8076 3936
rect 8024 3893 8033 3927
rect 8033 3893 8067 3927
rect 8067 3893 8076 3927
rect 8024 3884 8076 3893
rect 8300 3884 8352 3936
rect 8760 4029 8769 4063
rect 8769 4029 8803 4063
rect 8803 4029 8812 4063
rect 8760 4020 8812 4029
rect 9220 4063 9272 4072
rect 9220 4029 9229 4063
rect 9229 4029 9263 4063
rect 9263 4029 9272 4063
rect 9220 4020 9272 4029
rect 9404 4020 9456 4072
rect 10692 4063 10744 4072
rect 10692 4029 10701 4063
rect 10701 4029 10735 4063
rect 10735 4029 10744 4063
rect 10692 4020 10744 4029
rect 11520 4063 11572 4072
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 9128 3952 9180 4004
rect 13084 4020 13136 4072
rect 13360 4020 13412 4072
rect 15016 4020 15068 4072
rect 16304 4020 16356 4072
rect 16488 4020 16540 4072
rect 10416 3884 10468 3936
rect 10692 3884 10744 3936
rect 11244 3884 11296 3936
rect 12348 3884 12400 3936
rect 13268 3927 13320 3936
rect 13268 3893 13277 3927
rect 13277 3893 13311 3927
rect 13311 3893 13320 3927
rect 13268 3884 13320 3893
rect 13452 3884 13504 3936
rect 13636 3927 13688 3936
rect 13636 3893 13645 3927
rect 13645 3893 13679 3927
rect 13679 3893 13688 3927
rect 13636 3884 13688 3893
rect 13820 3927 13872 3936
rect 13820 3893 13829 3927
rect 13829 3893 13863 3927
rect 13863 3893 13872 3927
rect 13820 3884 13872 3893
rect 15292 3952 15344 4004
rect 15936 3952 15988 4004
rect 15200 3884 15252 3936
rect 15660 3927 15712 3936
rect 15660 3893 15669 3927
rect 15669 3893 15703 3927
rect 15703 3893 15712 3927
rect 15660 3884 15712 3893
rect 16028 3927 16080 3936
rect 16028 3893 16037 3927
rect 16037 3893 16071 3927
rect 16071 3893 16080 3927
rect 16028 3884 16080 3893
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 16672 3927 16724 3936
rect 16672 3893 16681 3927
rect 16681 3893 16715 3927
rect 16715 3893 16724 3927
rect 16672 3884 16724 3893
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 1308 3680 1360 3732
rect 1676 3680 1728 3732
rect 2136 3680 2188 3732
rect 3424 3680 3476 3732
rect 3884 3680 3936 3732
rect 5172 3680 5224 3732
rect 6368 3723 6420 3732
rect 6368 3689 6377 3723
rect 6377 3689 6411 3723
rect 6411 3689 6420 3723
rect 6368 3680 6420 3689
rect 4528 3612 4580 3664
rect 4712 3655 4764 3664
rect 4712 3621 4721 3655
rect 4721 3621 4755 3655
rect 4755 3621 4764 3655
rect 4712 3612 4764 3621
rect 7656 3680 7708 3732
rect 8392 3680 8444 3732
rect 9128 3680 9180 3732
rect 10784 3723 10836 3732
rect 10784 3689 10793 3723
rect 10793 3689 10827 3723
rect 10827 3689 10836 3723
rect 10784 3680 10836 3689
rect 10968 3680 11020 3732
rect 13636 3680 13688 3732
rect 1676 3544 1728 3596
rect 1952 3587 2004 3596
rect 1952 3553 1961 3587
rect 1961 3553 1995 3587
rect 1995 3553 2004 3587
rect 1952 3544 2004 3553
rect 4344 3544 4396 3596
rect 2504 3476 2556 3528
rect 2964 3476 3016 3528
rect 3884 3476 3936 3528
rect 4160 3476 4212 3528
rect 4436 3476 4488 3528
rect 3976 3408 4028 3460
rect 7656 3519 7708 3528
rect 7656 3485 7690 3519
rect 7690 3485 7708 3519
rect 5172 3408 5224 3460
rect 5632 3408 5684 3460
rect 6000 3408 6052 3460
rect 7656 3476 7708 3485
rect 8484 3476 8536 3528
rect 6276 3451 6328 3460
rect 6276 3417 6285 3451
rect 6285 3417 6319 3451
rect 6319 3417 6328 3451
rect 6276 3408 6328 3417
rect 9036 3476 9088 3528
rect 9772 3476 9824 3528
rect 2872 3340 2924 3392
rect 4160 3383 4212 3392
rect 4160 3349 4169 3383
rect 4169 3349 4203 3383
rect 4203 3349 4212 3383
rect 4160 3340 4212 3349
rect 4620 3340 4672 3392
rect 6644 3340 6696 3392
rect 6920 3383 6972 3392
rect 6920 3349 6929 3383
rect 6929 3349 6963 3383
rect 6963 3349 6972 3383
rect 6920 3340 6972 3349
rect 7380 3340 7432 3392
rect 8392 3340 8444 3392
rect 10416 3408 10468 3460
rect 12532 3612 12584 3664
rect 14004 3612 14056 3664
rect 14556 3680 14608 3732
rect 14740 3680 14792 3732
rect 15016 3680 15068 3732
rect 15752 3680 15804 3732
rect 16120 3680 16172 3732
rect 16396 3680 16448 3732
rect 16580 3680 16632 3732
rect 17224 3680 17276 3732
rect 17500 3680 17552 3732
rect 17776 3680 17828 3732
rect 17960 3680 18012 3732
rect 15476 3612 15528 3664
rect 13360 3476 13412 3528
rect 15568 3544 15620 3596
rect 16396 3544 16448 3596
rect 18236 3544 18288 3596
rect 15384 3519 15436 3528
rect 13268 3408 13320 3460
rect 15384 3485 15393 3519
rect 15393 3485 15427 3519
rect 15427 3485 15436 3519
rect 15384 3476 15436 3485
rect 15844 3476 15896 3528
rect 16488 3476 16540 3528
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 22652 3476 22704 3528
rect 15200 3408 15252 3460
rect 16212 3408 16264 3460
rect 19524 3408 19576 3460
rect 10324 3340 10376 3392
rect 10600 3340 10652 3392
rect 10784 3340 10836 3392
rect 13820 3340 13872 3392
rect 14188 3383 14240 3392
rect 14188 3349 14197 3383
rect 14197 3349 14231 3383
rect 14231 3349 14240 3383
rect 14188 3340 14240 3349
rect 15016 3340 15068 3392
rect 15568 3383 15620 3392
rect 15568 3349 15577 3383
rect 15577 3349 15611 3383
rect 15611 3349 15620 3383
rect 15568 3340 15620 3349
rect 15752 3340 15804 3392
rect 16948 3340 17000 3392
rect 19064 3340 19116 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 1676 3179 1728 3188
rect 1676 3145 1685 3179
rect 1685 3145 1719 3179
rect 1719 3145 1728 3179
rect 1676 3136 1728 3145
rect 2044 3136 2096 3188
rect 1952 3068 2004 3120
rect 3240 3136 3292 3188
rect 5172 3136 5224 3188
rect 5356 3179 5408 3188
rect 5356 3145 5365 3179
rect 5365 3145 5399 3179
rect 5399 3145 5408 3179
rect 5356 3136 5408 3145
rect 5908 3179 5960 3188
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 4160 3068 4212 3120
rect 5908 3145 5917 3179
rect 5917 3145 5951 3179
rect 5951 3145 5960 3179
rect 5908 3136 5960 3145
rect 6828 3179 6880 3188
rect 6828 3145 6837 3179
rect 6837 3145 6871 3179
rect 6871 3145 6880 3179
rect 6828 3136 6880 3145
rect 7748 3136 7800 3188
rect 8300 3179 8352 3188
rect 8300 3145 8309 3179
rect 8309 3145 8343 3179
rect 8343 3145 8352 3179
rect 8300 3136 8352 3145
rect 9220 3136 9272 3188
rect 9312 3136 9364 3188
rect 10140 3179 10192 3188
rect 10140 3145 10149 3179
rect 10149 3145 10183 3179
rect 10183 3145 10192 3179
rect 10140 3136 10192 3145
rect 10600 3179 10652 3188
rect 10600 3145 10609 3179
rect 10609 3145 10643 3179
rect 10643 3145 10652 3179
rect 10600 3136 10652 3145
rect 14280 3136 14332 3188
rect 6000 3068 6052 3120
rect 7012 3068 7064 3120
rect 7288 3068 7340 3120
rect 8024 3068 8076 3120
rect 5448 3000 5500 3052
rect 5632 3000 5684 3052
rect 6092 3000 6144 3052
rect 6552 3043 6604 3052
rect 6552 3009 6561 3043
rect 6561 3009 6595 3043
rect 6595 3009 6604 3043
rect 6552 3000 6604 3009
rect 3240 2975 3292 2984
rect 3240 2941 3249 2975
rect 3249 2941 3283 2975
rect 3283 2941 3292 2975
rect 3240 2932 3292 2941
rect 4436 2932 4488 2984
rect 5540 2932 5592 2984
rect 3056 2864 3108 2916
rect 4252 2864 4304 2916
rect 5448 2864 5500 2916
rect 1584 2839 1636 2848
rect 1584 2805 1593 2839
rect 1593 2805 1627 2839
rect 1627 2805 1636 2839
rect 1584 2796 1636 2805
rect 5172 2796 5224 2848
rect 6184 2932 6236 2984
rect 7932 3000 7984 3052
rect 9404 3000 9456 3052
rect 10048 3000 10100 3052
rect 10324 3068 10376 3120
rect 7656 2864 7708 2916
rect 7748 2796 7800 2848
rect 8392 2932 8444 2984
rect 8944 2932 8996 2984
rect 9588 2932 9640 2984
rect 10416 2975 10468 2984
rect 10416 2941 10425 2975
rect 10425 2941 10459 2975
rect 10459 2941 10468 2975
rect 10416 2932 10468 2941
rect 11244 3068 11296 3120
rect 11888 3068 11940 3120
rect 10876 3000 10928 3052
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 11336 2932 11388 2984
rect 12532 3068 12584 3120
rect 15108 3136 15160 3188
rect 12440 3043 12492 3052
rect 12440 3009 12449 3043
rect 12449 3009 12483 3043
rect 12483 3009 12492 3043
rect 12900 3043 12952 3052
rect 12440 3000 12492 3009
rect 12900 3009 12909 3043
rect 12909 3009 12943 3043
rect 12943 3009 12952 3043
rect 12900 3000 12952 3009
rect 13452 3043 13504 3052
rect 13452 3009 13461 3043
rect 13461 3009 13495 3043
rect 13495 3009 13504 3043
rect 13452 3000 13504 3009
rect 14004 3000 14056 3052
rect 14464 3000 14516 3052
rect 15108 3043 15160 3052
rect 15108 3009 15117 3043
rect 15117 3009 15151 3043
rect 15151 3009 15160 3043
rect 15108 3000 15160 3009
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 15752 3068 15804 3120
rect 18052 3136 18104 3188
rect 18604 3136 18656 3188
rect 19984 3136 20036 3188
rect 20260 3179 20312 3188
rect 20260 3145 20269 3179
rect 20269 3145 20303 3179
rect 20303 3145 20312 3179
rect 20260 3136 20312 3145
rect 15844 3000 15896 3052
rect 16120 3000 16172 3052
rect 16396 3000 16448 3052
rect 17040 3000 17092 3052
rect 17224 3043 17276 3052
rect 17224 3009 17233 3043
rect 17233 3009 17267 3043
rect 17267 3009 17276 3043
rect 17224 3000 17276 3009
rect 17500 3043 17552 3052
rect 17500 3009 17509 3043
rect 17509 3009 17543 3043
rect 17543 3009 17552 3043
rect 17500 3000 17552 3009
rect 17960 3000 18012 3052
rect 18236 3000 18288 3052
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 18788 3000 18840 3052
rect 19524 3043 19576 3052
rect 19524 3009 19533 3043
rect 19533 3009 19567 3043
rect 19567 3009 19576 3043
rect 19524 3000 19576 3009
rect 20260 3000 20312 3052
rect 13268 2932 13320 2984
rect 13820 2864 13872 2916
rect 17500 2864 17552 2916
rect 19616 2864 19668 2916
rect 20444 2864 20496 2916
rect 22192 2864 22244 2916
rect 10232 2796 10284 2848
rect 11888 2839 11940 2848
rect 11888 2805 11897 2839
rect 11897 2805 11931 2839
rect 11931 2805 11940 2839
rect 11888 2796 11940 2805
rect 13084 2839 13136 2848
rect 13084 2805 13093 2839
rect 13093 2805 13127 2839
rect 13127 2805 13136 2839
rect 13084 2796 13136 2805
rect 13360 2839 13412 2848
rect 13360 2805 13369 2839
rect 13369 2805 13403 2839
rect 13403 2805 13412 2839
rect 13360 2796 13412 2805
rect 15200 2839 15252 2848
rect 15200 2805 15209 2839
rect 15209 2805 15243 2839
rect 15243 2805 15252 2839
rect 15200 2796 15252 2805
rect 15568 2796 15620 2848
rect 15752 2839 15804 2848
rect 15752 2805 15761 2839
rect 15761 2805 15795 2839
rect 15795 2805 15804 2839
rect 16212 2839 16264 2848
rect 15752 2796 15804 2805
rect 16212 2805 16221 2839
rect 16221 2805 16255 2839
rect 16255 2805 16264 2839
rect 16212 2796 16264 2805
rect 16764 2796 16816 2848
rect 17132 2839 17184 2848
rect 17132 2805 17141 2839
rect 17141 2805 17175 2839
rect 17175 2805 17184 2839
rect 17132 2796 17184 2805
rect 17776 2796 17828 2848
rect 18236 2839 18288 2848
rect 18236 2805 18245 2839
rect 18245 2805 18279 2839
rect 18279 2805 18288 2839
rect 18236 2796 18288 2805
rect 20996 2796 21048 2848
rect 21732 2796 21784 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 3976 2592 4028 2644
rect 5264 2592 5316 2644
rect 5448 2592 5500 2644
rect 6184 2592 6236 2644
rect 6460 2635 6512 2644
rect 6460 2601 6469 2635
rect 6469 2601 6503 2635
rect 6503 2601 6512 2635
rect 6460 2592 6512 2601
rect 6552 2592 6604 2644
rect 6736 2592 6788 2644
rect 7196 2592 7248 2644
rect 7288 2592 7340 2644
rect 7564 2592 7616 2644
rect 7932 2592 7984 2644
rect 9220 2592 9272 2644
rect 9404 2635 9456 2644
rect 9404 2601 9413 2635
rect 9413 2601 9447 2635
rect 9447 2601 9456 2635
rect 9404 2592 9456 2601
rect 9588 2592 9640 2644
rect 12808 2592 12860 2644
rect 15108 2592 15160 2644
rect 2228 2499 2280 2508
rect 2228 2465 2237 2499
rect 2237 2465 2271 2499
rect 2271 2465 2280 2499
rect 2228 2456 2280 2465
rect 4344 2524 4396 2576
rect 7012 2524 7064 2576
rect 1952 2431 2004 2440
rect 1952 2397 1961 2431
rect 1961 2397 1995 2431
rect 1995 2397 2004 2431
rect 1952 2388 2004 2397
rect 3148 2431 3200 2440
rect 3148 2397 3157 2431
rect 3157 2397 3191 2431
rect 3191 2397 3200 2431
rect 3148 2388 3200 2397
rect 4068 2456 4120 2508
rect 5540 2499 5592 2508
rect 5540 2465 5549 2499
rect 5549 2465 5583 2499
rect 5583 2465 5592 2499
rect 5540 2456 5592 2465
rect 4620 2388 4672 2440
rect 8300 2524 8352 2576
rect 10416 2524 10468 2576
rect 8484 2499 8536 2508
rect 8484 2465 8493 2499
rect 8493 2465 8527 2499
rect 8527 2465 8536 2499
rect 8484 2456 8536 2465
rect 8576 2456 8628 2508
rect 9496 2456 9548 2508
rect 10232 2499 10284 2508
rect 10232 2465 10241 2499
rect 10241 2465 10275 2499
rect 10275 2465 10284 2499
rect 10232 2456 10284 2465
rect 10692 2456 10744 2508
rect 13360 2524 13412 2576
rect 12072 2499 12124 2508
rect 12072 2465 12081 2499
rect 12081 2465 12115 2499
rect 12115 2465 12124 2499
rect 12072 2456 12124 2465
rect 12164 2456 12216 2508
rect 3424 2363 3476 2372
rect 3424 2329 3433 2363
rect 3433 2329 3467 2363
rect 3467 2329 3476 2363
rect 3424 2320 3476 2329
rect 5724 2320 5776 2372
rect 4896 2252 4948 2304
rect 6736 2388 6788 2440
rect 7104 2388 7156 2440
rect 7380 2431 7432 2440
rect 7380 2397 7389 2431
rect 7389 2397 7423 2431
rect 7423 2397 7432 2431
rect 7380 2388 7432 2397
rect 7748 2388 7800 2440
rect 8116 2388 8168 2440
rect 10600 2388 10652 2440
rect 11888 2388 11940 2440
rect 13084 2456 13136 2508
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 13728 2524 13780 2576
rect 13820 2388 13872 2440
rect 6092 2363 6144 2372
rect 6092 2329 6101 2363
rect 6101 2329 6135 2363
rect 6135 2329 6144 2363
rect 6092 2320 6144 2329
rect 6184 2320 6236 2372
rect 6552 2363 6604 2372
rect 6552 2329 6561 2363
rect 6561 2329 6595 2363
rect 6595 2329 6604 2363
rect 6552 2320 6604 2329
rect 7656 2320 7708 2372
rect 8668 2320 8720 2372
rect 10416 2320 10468 2372
rect 12440 2320 12492 2372
rect 15200 2388 15252 2440
rect 15568 2431 15620 2440
rect 15568 2397 15577 2431
rect 15577 2397 15611 2431
rect 15611 2397 15620 2431
rect 15568 2388 15620 2397
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 16212 2431 16264 2440
rect 16212 2397 16221 2431
rect 16221 2397 16255 2431
rect 16255 2397 16264 2431
rect 16212 2388 16264 2397
rect 16672 2431 16724 2440
rect 16672 2397 16681 2431
rect 16681 2397 16715 2431
rect 16715 2397 16724 2431
rect 16672 2388 16724 2397
rect 17132 2431 17184 2440
rect 17132 2397 17141 2431
rect 17141 2397 17175 2431
rect 17175 2397 17184 2431
rect 17132 2388 17184 2397
rect 17592 2431 17644 2440
rect 17592 2397 17601 2431
rect 17601 2397 17635 2431
rect 17635 2397 17644 2431
rect 17592 2388 17644 2397
rect 17684 2388 17736 2440
rect 18236 2388 18288 2440
rect 19064 2388 19116 2440
rect 19616 2431 19668 2440
rect 19616 2397 19625 2431
rect 19625 2397 19659 2431
rect 19659 2397 19668 2431
rect 19616 2388 19668 2397
rect 19984 2431 20036 2440
rect 19984 2397 19993 2431
rect 19993 2397 20027 2431
rect 20027 2397 20036 2431
rect 19984 2388 20036 2397
rect 20444 2431 20496 2440
rect 20444 2397 20453 2431
rect 20453 2397 20487 2431
rect 20487 2397 20496 2431
rect 20444 2388 20496 2397
rect 20904 2431 20956 2440
rect 20904 2397 20913 2431
rect 20913 2397 20947 2431
rect 20947 2397 20956 2431
rect 20904 2388 20956 2397
rect 20996 2388 21048 2440
rect 8300 2252 8352 2304
rect 13268 2252 13320 2304
rect 14372 2252 14424 2304
rect 14740 2252 14792 2304
rect 15200 2252 15252 2304
rect 15660 2252 15712 2304
rect 16120 2252 16172 2304
rect 16948 2252 17000 2304
rect 17040 2252 17092 2304
rect 17500 2252 17552 2304
rect 17960 2252 18012 2304
rect 18420 2252 18472 2304
rect 18972 2252 19024 2304
rect 19524 2252 19576 2304
rect 19892 2252 19944 2304
rect 20352 2252 20404 2304
rect 20812 2252 20864 2304
rect 21272 2252 21324 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 3240 2048 3292 2100
rect 6644 2048 6696 2100
rect 6736 2048 6788 2100
rect 14832 2048 14884 2100
rect 1952 1980 2004 2032
rect 7840 1980 7892 2032
rect 7656 1844 7708 1896
rect 8208 1844 8260 1896
rect 8300 1844 8352 1896
rect 12900 1844 12952 1896
rect 5908 1776 5960 1828
rect 6828 1776 6880 1828
rect 15292 1776 15344 1828
rect 1584 1708 1636 1760
rect 14648 1708 14700 1760
rect 6552 1640 6604 1692
rect 6736 1640 6788 1692
rect 14924 1640 14976 1692
rect 3516 1572 3568 1624
rect 14188 1572 14240 1624
rect 4068 1028 4120 1080
rect 6920 1028 6972 1080
<< metal2 >>
rect 202 22200 258 23000
rect 662 22200 718 23000
rect 1122 22200 1178 23000
rect 1582 22200 1638 23000
rect 2042 22200 2098 23000
rect 2318 22672 2374 22681
rect 2318 22607 2374 22616
rect 216 19310 244 22200
rect 676 20505 704 22200
rect 662 20496 718 20505
rect 662 20431 718 20440
rect 1136 19922 1164 22200
rect 1490 21176 1546 21185
rect 1490 21111 1546 21120
rect 1308 20256 1360 20262
rect 1308 20198 1360 20204
rect 1124 19916 1176 19922
rect 1124 19858 1176 19864
rect 204 19304 256 19310
rect 204 19246 256 19252
rect 1214 19272 1270 19281
rect 1214 19207 1270 19216
rect 1228 17066 1256 19207
rect 1216 17060 1268 17066
rect 1216 17002 1268 17008
rect 1320 16522 1348 20198
rect 1400 19440 1452 19446
rect 1400 19382 1452 19388
rect 1308 16516 1360 16522
rect 1308 16458 1360 16464
rect 1412 15434 1440 19382
rect 1504 18970 1532 21111
rect 1492 18964 1544 18970
rect 1492 18906 1544 18912
rect 1596 18850 1624 22200
rect 2056 20618 2084 22200
rect 2056 20590 2176 20618
rect 2148 20466 2176 20590
rect 2044 20460 2096 20466
rect 2044 20402 2096 20408
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 1768 19916 1820 19922
rect 1768 19858 1820 19864
rect 1596 18822 1716 18850
rect 1584 18760 1636 18766
rect 1584 18702 1636 18708
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1504 17921 1532 18022
rect 1490 17912 1546 17921
rect 1490 17847 1546 17856
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17377 1532 17478
rect 1490 17368 1546 17377
rect 1490 17303 1546 17312
rect 1596 17134 1624 18702
rect 1688 17762 1716 18822
rect 1780 18601 1808 19858
rect 1952 19848 2004 19854
rect 1952 19790 2004 19796
rect 1964 19417 1992 19790
rect 1950 19408 2006 19417
rect 2056 19378 2084 20402
rect 1950 19343 2006 19352
rect 2044 19372 2096 19378
rect 2044 19314 2096 19320
rect 1858 18864 1914 18873
rect 1858 18799 1914 18808
rect 1766 18592 1822 18601
rect 1766 18527 1822 18536
rect 1872 17882 1900 18799
rect 2148 18737 2176 20402
rect 2228 19304 2280 19310
rect 2228 19246 2280 19252
rect 2240 18873 2268 19246
rect 2226 18864 2282 18873
rect 2226 18799 2282 18808
rect 2134 18728 2190 18737
rect 2134 18663 2190 18672
rect 2228 18692 2280 18698
rect 2228 18634 2280 18640
rect 2240 18442 2268 18634
rect 2148 18414 2268 18442
rect 2332 18426 2360 22607
rect 2502 22200 2558 23000
rect 2962 22200 3018 23000
rect 3422 22200 3478 23000
rect 3882 22200 3938 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6182 22200 6238 23000
rect 6288 22222 6592 22250
rect 2412 19508 2464 19514
rect 2412 19450 2464 19456
rect 2320 18420 2372 18426
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1860 17876 1912 17882
rect 1860 17818 1912 17824
rect 1688 17734 1808 17762
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1584 17128 1636 17134
rect 1584 17070 1636 17076
rect 1492 16992 1544 16998
rect 1490 16960 1492 16969
rect 1544 16960 1546 16969
rect 1490 16895 1546 16904
rect 1688 16794 1716 17614
rect 1780 17338 1808 17734
rect 1964 17649 1992 18226
rect 2042 17776 2098 17785
rect 2042 17711 2098 17720
rect 1950 17640 2006 17649
rect 1950 17575 2006 17584
rect 2056 17354 2084 17711
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1964 17326 2084 17354
rect 1768 17196 1820 17202
rect 1768 17138 1820 17144
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1492 16448 1544 16454
rect 1490 16416 1492 16425
rect 1544 16416 1546 16425
rect 1490 16351 1546 16360
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1490 16008 1546 16017
rect 1490 15943 1492 15952
rect 1544 15943 1546 15952
rect 1492 15914 1544 15920
rect 1688 15638 1716 16050
rect 1780 15978 1808 17138
rect 1860 16584 1912 16590
rect 1860 16526 1912 16532
rect 1872 16250 1900 16526
rect 1860 16244 1912 16250
rect 1860 16186 1912 16192
rect 1964 16182 1992 17326
rect 2148 17202 2176 18414
rect 2320 18362 2372 18368
rect 2226 18320 2282 18329
rect 2226 18255 2282 18264
rect 2320 18284 2372 18290
rect 2240 17882 2268 18255
rect 2320 18226 2372 18232
rect 2332 18086 2360 18226
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 2228 17876 2280 17882
rect 2228 17818 2280 17824
rect 2228 17672 2280 17678
rect 2228 17614 2280 17620
rect 2044 17196 2096 17202
rect 2044 17138 2096 17144
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 2056 16250 2084 17138
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 1952 16176 2004 16182
rect 1952 16118 2004 16124
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 1768 15972 1820 15978
rect 1768 15914 1820 15920
rect 2148 15706 2176 16050
rect 2240 15978 2268 17614
rect 2318 17232 2374 17241
rect 2318 17167 2374 17176
rect 2332 17066 2360 17167
rect 2320 17060 2372 17066
rect 2320 17002 2372 17008
rect 2424 16590 2452 19450
rect 2516 19446 2544 22200
rect 2778 22128 2834 22137
rect 2976 22114 3004 22200
rect 2976 22086 3096 22114
rect 2778 22063 2834 22072
rect 2688 20392 2740 20398
rect 2688 20334 2740 20340
rect 2594 19816 2650 19825
rect 2594 19751 2650 19760
rect 2504 19440 2556 19446
rect 2504 19382 2556 19388
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2410 16416 2466 16425
rect 2410 16351 2466 16360
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2228 15972 2280 15978
rect 2228 15914 2280 15920
rect 2332 15706 2360 16050
rect 2136 15700 2188 15706
rect 2136 15642 2188 15648
rect 2320 15700 2372 15706
rect 2320 15642 2372 15648
rect 1676 15632 1728 15638
rect 2424 15586 2452 16351
rect 1676 15574 1728 15580
rect 2332 15558 2452 15586
rect 1676 15496 1728 15502
rect 2044 15496 2096 15502
rect 1676 15438 1728 15444
rect 1858 15464 1914 15473
rect 1400 15428 1452 15434
rect 1400 15370 1452 15376
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1504 15065 1532 15302
rect 1688 15162 1716 15438
rect 2044 15438 2096 15444
rect 1858 15399 1914 15408
rect 1872 15366 1900 15399
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1676 15156 1728 15162
rect 1676 15098 1728 15104
rect 1490 15056 1546 15065
rect 1490 14991 1546 15000
rect 1860 15020 1912 15026
rect 1860 14962 1912 14968
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 1768 14952 1820 14958
rect 1768 14894 1820 14900
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1504 14521 1532 14758
rect 1490 14512 1546 14521
rect 1308 14476 1360 14482
rect 1490 14447 1546 14456
rect 1308 14418 1360 14424
rect 1320 12434 1348 14418
rect 1400 14340 1452 14346
rect 1400 14282 1452 14288
rect 1412 13326 1440 14282
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1504 14113 1532 14214
rect 1490 14104 1546 14113
rect 1490 14039 1546 14048
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 1504 13569 1532 13670
rect 1490 13560 1546 13569
rect 1688 13530 1716 13874
rect 1490 13495 1546 13504
rect 1676 13524 1728 13530
rect 1676 13466 1728 13472
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1582 13288 1638 13297
rect 1412 13161 1440 13262
rect 1582 13223 1638 13232
rect 1596 13190 1624 13223
rect 1584 13184 1636 13190
rect 1398 13152 1454 13161
rect 1584 13126 1636 13132
rect 1398 13087 1454 13096
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12617 1440 12786
rect 1584 12640 1636 12646
rect 1398 12608 1454 12617
rect 1584 12582 1636 12588
rect 1398 12543 1454 12552
rect 1228 12406 1348 12434
rect 1122 5536 1178 5545
rect 1122 5471 1178 5480
rect 664 4140 716 4146
rect 664 4082 716 4088
rect 202 2816 258 2825
rect 202 2751 258 2760
rect 216 800 244 2751
rect 676 800 704 4082
rect 1136 800 1164 5471
rect 1228 3369 1256 12406
rect 1412 11354 1440 12543
rect 1492 12232 1544 12238
rect 1490 12200 1492 12209
rect 1544 12200 1546 12209
rect 1490 12135 1546 12144
rect 1400 11348 1452 11354
rect 1400 11290 1452 11296
rect 1398 11112 1454 11121
rect 1398 11047 1454 11056
rect 1412 10674 1440 11047
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1504 10266 1532 12135
rect 1596 11121 1624 12582
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1688 11665 1716 12174
rect 1674 11656 1730 11665
rect 1674 11591 1730 11600
rect 1582 11112 1638 11121
rect 1582 11047 1638 11056
rect 1584 11008 1636 11014
rect 1584 10950 1636 10956
rect 1596 10554 1624 10950
rect 1674 10704 1730 10713
rect 1674 10639 1676 10648
rect 1728 10639 1730 10648
rect 1676 10610 1728 10616
rect 1596 10526 1716 10554
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 1398 9208 1454 9217
rect 1398 9143 1454 9152
rect 1412 8401 1440 9143
rect 1398 8392 1454 8401
rect 1398 8327 1454 8336
rect 1412 7410 1440 8327
rect 1504 8090 1532 9522
rect 1596 9450 1624 9998
rect 1584 9444 1636 9450
rect 1584 9386 1636 9392
rect 1582 8936 1638 8945
rect 1582 8871 1638 8880
rect 1596 8838 1624 8871
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1688 8378 1716 10526
rect 1780 10266 1808 14894
rect 1872 14074 1900 14962
rect 1964 14618 1992 14962
rect 2056 14890 2084 15438
rect 2228 15020 2280 15026
rect 2228 14962 2280 14968
rect 2044 14884 2096 14890
rect 2044 14826 2096 14832
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 2240 14414 2268 14962
rect 2044 14408 2096 14414
rect 2044 14350 2096 14356
rect 2228 14408 2280 14414
rect 2228 14350 2280 14356
rect 2056 14074 2084 14350
rect 1860 14068 1912 14074
rect 1860 14010 1912 14016
rect 2044 14068 2096 14074
rect 2044 14010 2096 14016
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1872 12986 1900 13262
rect 1860 12980 1912 12986
rect 1860 12922 1912 12928
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1952 12096 2004 12102
rect 1952 12038 2004 12044
rect 1872 11801 1900 12038
rect 1964 11830 1992 12038
rect 1952 11824 2004 11830
rect 1858 11792 1914 11801
rect 1952 11766 2004 11772
rect 1858 11727 1914 11736
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 11218 1900 11494
rect 2056 11257 2084 13874
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 2136 13184 2188 13190
rect 2136 13126 2188 13132
rect 2148 12986 2176 13126
rect 2136 12980 2188 12986
rect 2136 12922 2188 12928
rect 2240 12714 2268 13330
rect 2332 13274 2360 15558
rect 2412 15496 2464 15502
rect 2412 15438 2464 15444
rect 2424 15094 2452 15438
rect 2412 15088 2464 15094
rect 2412 15030 2464 15036
rect 2516 14770 2544 18022
rect 2608 17882 2636 19751
rect 2700 19417 2728 20334
rect 2686 19408 2742 19417
rect 2686 19343 2742 19352
rect 2792 18902 2820 22063
rect 2870 21720 2926 21729
rect 2870 21655 2926 21664
rect 2780 18896 2832 18902
rect 2780 18838 2832 18844
rect 2780 18760 2832 18766
rect 2780 18702 2832 18708
rect 2792 18426 2820 18702
rect 2780 18420 2832 18426
rect 2780 18362 2832 18368
rect 2884 18358 2912 21655
rect 3068 20602 3096 22086
rect 3436 20890 3464 22200
rect 3344 20862 3464 20890
rect 3056 20596 3108 20602
rect 3056 20538 3108 20544
rect 3238 20496 3294 20505
rect 3238 20431 3294 20440
rect 3054 20224 3110 20233
rect 3054 20159 3110 20168
rect 2964 19168 3016 19174
rect 2964 19110 3016 19116
rect 2872 18352 2924 18358
rect 2700 18290 2820 18306
rect 2872 18294 2924 18300
rect 2688 18284 2832 18290
rect 2740 18278 2780 18284
rect 2688 18226 2740 18232
rect 2780 18226 2832 18232
rect 2688 18080 2740 18086
rect 2688 18022 2740 18028
rect 2596 17876 2648 17882
rect 2596 17818 2648 17824
rect 2596 17672 2648 17678
rect 2596 17614 2648 17620
rect 2608 15638 2636 17614
rect 2700 16561 2728 18022
rect 2778 17912 2834 17921
rect 2778 17847 2834 17856
rect 2792 17202 2820 17847
rect 2872 17672 2924 17678
rect 2872 17614 2924 17620
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2792 16697 2820 17138
rect 2778 16688 2834 16697
rect 2778 16623 2834 16632
rect 2686 16552 2742 16561
rect 2686 16487 2742 16496
rect 2688 16448 2740 16454
rect 2686 16416 2688 16425
rect 2780 16448 2832 16454
rect 2740 16416 2742 16425
rect 2780 16390 2832 16396
rect 2686 16351 2742 16360
rect 2792 16182 2820 16390
rect 2884 16250 2912 17614
rect 2976 17377 3004 19110
rect 3068 17882 3096 20159
rect 3252 19854 3280 20431
rect 3240 19848 3292 19854
rect 3240 19790 3292 19796
rect 3344 19666 3372 20862
rect 3422 20768 3478 20777
rect 3422 20703 3478 20712
rect 3252 19638 3372 19666
rect 3148 19236 3200 19242
rect 3148 19178 3200 19184
rect 3160 18970 3188 19178
rect 3148 18964 3200 18970
rect 3148 18906 3200 18912
rect 3148 18624 3200 18630
rect 3148 18566 3200 18572
rect 3056 17876 3108 17882
rect 3056 17818 3108 17824
rect 3160 17610 3188 18566
rect 3252 17921 3280 19638
rect 3436 18850 3464 20703
rect 3516 20460 3568 20466
rect 3516 20402 3568 20408
rect 3528 20369 3556 20402
rect 3514 20360 3570 20369
rect 3514 20295 3570 20304
rect 3549 20156 3857 20176
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20080 3857 20100
rect 3514 19952 3570 19961
rect 3514 19887 3570 19896
rect 3528 19854 3556 19887
rect 3516 19848 3568 19854
rect 3516 19790 3568 19796
rect 3700 19712 3752 19718
rect 3700 19654 3752 19660
rect 3712 19417 3740 19654
rect 3698 19408 3754 19417
rect 3698 19343 3754 19352
rect 3549 19068 3857 19088
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 18992 3857 19012
rect 3332 18828 3384 18834
rect 3436 18822 3648 18850
rect 3332 18770 3384 18776
rect 3344 18714 3372 18770
rect 3344 18686 3464 18714
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3344 18193 3372 18566
rect 3436 18290 3464 18686
rect 3424 18284 3476 18290
rect 3424 18226 3476 18232
rect 3330 18184 3386 18193
rect 3620 18170 3648 18822
rect 3792 18420 3844 18426
rect 3896 18408 3924 22200
rect 4066 20496 4122 20505
rect 4066 20431 4122 20440
rect 3976 20256 4028 20262
rect 3974 20224 3976 20233
rect 4028 20224 4030 20233
rect 3974 20159 4030 20168
rect 4080 19825 4108 20431
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 4066 19816 4122 19825
rect 4172 19786 4200 20334
rect 4066 19751 4122 19760
rect 4160 19780 4212 19786
rect 4160 19722 4212 19728
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3844 18380 3924 18408
rect 3792 18362 3844 18368
rect 3330 18119 3386 18128
rect 3436 18142 3648 18170
rect 3238 17912 3294 17921
rect 3436 17882 3464 18142
rect 3549 17980 3857 18000
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17904 3857 17924
rect 3238 17847 3294 17856
rect 3424 17876 3476 17882
rect 3424 17818 3476 17824
rect 3240 17672 3292 17678
rect 3240 17614 3292 17620
rect 3056 17604 3108 17610
rect 3056 17546 3108 17552
rect 3148 17604 3200 17610
rect 3148 17546 3200 17552
rect 2962 17368 3018 17377
rect 2962 17303 3018 17312
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2780 16176 2832 16182
rect 2686 16144 2742 16153
rect 2780 16118 2832 16124
rect 2686 16079 2688 16088
rect 2740 16079 2742 16088
rect 2872 16108 2924 16114
rect 2688 16050 2740 16056
rect 2872 16050 2924 16056
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2596 15496 2648 15502
rect 2596 15438 2648 15444
rect 2608 15162 2636 15438
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2516 14742 2636 14770
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2516 13938 2544 14214
rect 2504 13932 2556 13938
rect 2504 13874 2556 13880
rect 2608 13530 2636 14742
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2596 13524 2648 13530
rect 2596 13466 2648 13472
rect 2332 13246 2636 13274
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2504 13184 2556 13190
rect 2504 13126 2556 13132
rect 2228 12708 2280 12714
rect 2228 12650 2280 12656
rect 2240 11830 2268 12650
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2332 11898 2360 12038
rect 2320 11892 2372 11898
rect 2320 11834 2372 11840
rect 2228 11824 2280 11830
rect 2228 11766 2280 11772
rect 2320 11348 2372 11354
rect 2424 11336 2452 13126
rect 2372 11308 2452 11336
rect 2320 11290 2372 11296
rect 2042 11248 2098 11257
rect 1860 11212 1912 11218
rect 2042 11183 2098 11192
rect 1860 11154 1912 11160
rect 2044 11144 2096 11150
rect 2044 11086 2096 11092
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1872 10169 1900 10610
rect 1952 10532 2004 10538
rect 1952 10474 2004 10480
rect 1858 10160 1914 10169
rect 1964 10146 1992 10474
rect 2056 10470 2084 11086
rect 2516 11014 2544 13126
rect 2608 12918 2636 13246
rect 2596 12912 2648 12918
rect 2596 12854 2648 12860
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 2608 12102 2636 12718
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2596 11212 2648 11218
rect 2596 11154 2648 11160
rect 2504 11008 2556 11014
rect 2504 10950 2556 10956
rect 2320 10668 2372 10674
rect 2320 10610 2372 10616
rect 2134 10568 2190 10577
rect 2134 10503 2136 10512
rect 2188 10503 2190 10512
rect 2136 10474 2188 10480
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2042 10160 2098 10169
rect 1964 10118 2042 10146
rect 1858 10095 1914 10104
rect 2042 10095 2098 10104
rect 2240 9994 2268 10406
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1872 9722 1900 9862
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1768 9648 1820 9654
rect 1768 9590 1820 9596
rect 2042 9616 2098 9625
rect 1596 8350 1716 8378
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1504 7342 1532 8026
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1596 6914 1624 8350
rect 1674 8256 1730 8265
rect 1674 8191 1730 8200
rect 1688 7410 1716 8191
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1674 7304 1730 7313
rect 1780 7290 1808 9590
rect 2042 9551 2098 9560
rect 1952 9036 2004 9042
rect 1952 8978 2004 8984
rect 1964 8634 1992 8978
rect 1952 8628 2004 8634
rect 1952 8570 2004 8576
rect 1860 8356 1912 8362
rect 1860 8298 1912 8304
rect 1730 7262 1808 7290
rect 1674 7239 1730 7248
rect 1504 6886 1624 6914
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1412 6633 1440 6734
rect 1398 6624 1454 6633
rect 1398 6559 1454 6568
rect 1504 6202 1532 6886
rect 1688 6798 1716 7239
rect 1766 6896 1822 6905
rect 1766 6831 1768 6840
rect 1820 6831 1822 6840
rect 1768 6802 1820 6808
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1768 6656 1820 6662
rect 1872 6644 1900 8298
rect 1950 7848 2006 7857
rect 1950 7783 2006 7792
rect 1820 6616 1900 6644
rect 1768 6598 1820 6604
rect 1964 6474 1992 7783
rect 1596 6446 1992 6474
rect 1596 6322 1624 6446
rect 1674 6352 1730 6361
rect 1584 6316 1636 6322
rect 1674 6287 1730 6296
rect 1952 6316 2004 6322
rect 1584 6258 1636 6264
rect 1504 6174 1624 6202
rect 1398 5944 1454 5953
rect 1398 5879 1454 5888
rect 1308 4004 1360 4010
rect 1308 3946 1360 3952
rect 1320 3738 1348 3946
rect 1308 3732 1360 3738
rect 1308 3674 1360 3680
rect 1214 3360 1270 3369
rect 1214 3295 1270 3304
rect 1412 3058 1440 5879
rect 1490 5672 1546 5681
rect 1490 5607 1492 5616
rect 1544 5607 1546 5616
rect 1492 5578 1544 5584
rect 1504 3505 1532 5578
rect 1596 5370 1624 6174
rect 1584 5364 1636 5370
rect 1584 5306 1636 5312
rect 1582 5128 1638 5137
rect 1582 5063 1638 5072
rect 1596 4622 1624 5063
rect 1688 4622 1716 6287
rect 1952 6258 2004 6264
rect 1964 5914 1992 6258
rect 1952 5908 2004 5914
rect 1952 5850 2004 5856
rect 2056 5234 2084 9551
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2148 5302 2176 9318
rect 2240 7886 2268 9318
rect 2332 8566 2360 10610
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2424 10062 2452 10542
rect 2412 10056 2464 10062
rect 2412 9998 2464 10004
rect 2608 9994 2636 11154
rect 2596 9988 2648 9994
rect 2596 9930 2648 9936
rect 2412 9512 2464 9518
rect 2412 9454 2464 9460
rect 2320 8560 2372 8566
rect 2320 8502 2372 8508
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2240 5846 2268 7686
rect 2320 7336 2372 7342
rect 2320 7278 2372 7284
rect 2332 6497 2360 7278
rect 2318 6488 2374 6497
rect 2318 6423 2374 6432
rect 2228 5840 2280 5846
rect 2228 5782 2280 5788
rect 2136 5296 2188 5302
rect 2136 5238 2188 5244
rect 2044 5228 2096 5234
rect 2044 5170 2096 5176
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1952 5160 2004 5166
rect 1952 5102 2004 5108
rect 1768 5024 1820 5030
rect 1768 4966 1820 4972
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1490 3496 1546 3505
rect 1490 3431 1546 3440
rect 1596 3380 1624 4558
rect 1674 3768 1730 3777
rect 1674 3703 1676 3712
rect 1728 3703 1730 3712
rect 1676 3674 1728 3680
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1504 3352 1624 3380
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1412 2009 1440 2994
rect 1398 2000 1454 2009
rect 1398 1935 1454 1944
rect 1504 1193 1532 3352
rect 1688 3194 1716 3538
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1584 2848 1636 2854
rect 1584 2790 1636 2796
rect 1596 1766 1624 2790
rect 1780 2774 1808 4966
rect 1872 3097 1900 5102
rect 1964 3602 1992 5102
rect 2042 4856 2098 4865
rect 2042 4791 2044 4800
rect 2096 4791 2098 4800
rect 2044 4762 2096 4768
rect 2042 4584 2098 4593
rect 2042 4519 2098 4528
rect 2056 4146 2084 4519
rect 2044 4140 2096 4146
rect 2044 4082 2096 4088
rect 2240 4010 2268 5782
rect 2332 4826 2360 6423
rect 2320 4820 2372 4826
rect 2320 4762 2372 4768
rect 2424 4622 2452 9454
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2516 7546 2544 8774
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 2502 7440 2558 7449
rect 2502 7375 2558 7384
rect 2516 7274 2544 7375
rect 2608 7342 2636 9930
rect 2700 9450 2728 13806
rect 2884 13462 2912 16050
rect 2872 13456 2924 13462
rect 2872 13398 2924 13404
rect 2780 13388 2832 13394
rect 2780 13330 2832 13336
rect 2792 11218 2820 13330
rect 2976 13326 3004 16934
rect 3068 16674 3096 17546
rect 3252 16794 3280 17614
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 3240 16788 3292 16794
rect 3240 16730 3292 16736
rect 3068 16646 3280 16674
rect 3056 16584 3108 16590
rect 3056 16526 3108 16532
rect 3068 15434 3096 16526
rect 3146 16008 3202 16017
rect 3146 15943 3202 15952
rect 3160 15910 3188 15943
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 3056 15428 3108 15434
rect 3056 15370 3108 15376
rect 3068 14090 3096 15370
rect 3160 15162 3188 15438
rect 3148 15156 3200 15162
rect 3148 15098 3200 15104
rect 3252 14906 3280 16646
rect 3344 16046 3372 17274
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 3436 16726 3464 17138
rect 3549 16892 3857 16912
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16816 3857 16836
rect 3424 16720 3476 16726
rect 3424 16662 3476 16668
rect 3884 16720 3936 16726
rect 3884 16662 3936 16668
rect 3896 16114 3924 16662
rect 3988 16590 4016 19654
rect 4160 19440 4212 19446
rect 4212 19417 4292 19428
rect 4212 19408 4306 19417
rect 4212 19400 4250 19408
rect 4160 19382 4212 19388
rect 4250 19343 4306 19352
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4068 17876 4120 17882
rect 4068 17818 4120 17824
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3976 16448 4028 16454
rect 3976 16390 4028 16396
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3884 16108 3936 16114
rect 3884 16050 3936 16056
rect 3332 16040 3384 16046
rect 3332 15982 3384 15988
rect 3332 15904 3384 15910
rect 3332 15846 3384 15852
rect 3344 15570 3372 15846
rect 3436 15706 3464 16050
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3549 15804 3857 15824
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15728 3857 15748
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3514 15600 3570 15609
rect 3332 15564 3384 15570
rect 3514 15535 3516 15544
rect 3332 15506 3384 15512
rect 3568 15535 3570 15544
rect 3516 15506 3568 15512
rect 3896 15502 3924 15914
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3988 15366 4016 16390
rect 4080 15434 4108 17818
rect 4172 17202 4200 18566
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4264 18193 4292 18362
rect 4250 18184 4306 18193
rect 4250 18119 4306 18128
rect 4356 17218 4384 22200
rect 4620 20596 4672 20602
rect 4620 20538 4672 20544
rect 4632 20398 4660 20538
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 4816 20346 4844 22200
rect 4896 20596 4948 20602
rect 4896 20538 4948 20544
rect 4908 20466 4936 20538
rect 5172 20528 5224 20534
rect 5170 20496 5172 20505
rect 5224 20496 5226 20505
rect 4896 20460 4948 20466
rect 5170 20431 5226 20440
rect 4896 20402 4948 20408
rect 5172 20392 5224 20398
rect 4528 19780 4580 19786
rect 4528 19722 4580 19728
rect 4540 19514 4568 19722
rect 4436 19508 4488 19514
rect 4436 19450 4488 19456
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4448 19378 4476 19450
rect 4436 19372 4488 19378
rect 4436 19314 4488 19320
rect 4436 18624 4488 18630
rect 4436 18566 4488 18572
rect 4448 18426 4476 18566
rect 4436 18420 4488 18426
rect 4436 18362 4488 18368
rect 4434 18320 4490 18329
rect 4540 18290 4568 19450
rect 4632 19145 4660 20334
rect 4816 20318 4936 20346
rect 5172 20334 5224 20340
rect 4804 20256 4856 20262
rect 4804 20198 4856 20204
rect 4816 19553 4844 20198
rect 4802 19544 4858 19553
rect 4802 19479 4858 19488
rect 4618 19136 4674 19145
rect 4618 19071 4674 19080
rect 4908 18748 4936 20318
rect 4988 18760 5040 18766
rect 4908 18720 4988 18748
rect 4988 18702 5040 18708
rect 4712 18692 4764 18698
rect 4712 18634 4764 18640
rect 4434 18255 4490 18264
rect 4528 18284 4580 18290
rect 4160 17196 4212 17202
rect 4160 17138 4212 17144
rect 4264 17190 4384 17218
rect 4160 17060 4212 17066
rect 4160 17002 4212 17008
rect 4172 16794 4200 17002
rect 4160 16788 4212 16794
rect 4160 16730 4212 16736
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 4172 15570 4200 16050
rect 4264 15706 4292 17190
rect 4344 17128 4396 17134
rect 4344 17070 4396 17076
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4356 15638 4384 17070
rect 4448 16572 4476 18255
rect 4528 18226 4580 18232
rect 4540 17678 4568 18226
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4632 17921 4660 18022
rect 4618 17912 4674 17921
rect 4618 17847 4674 17856
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 4540 16726 4568 17614
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4528 16720 4580 16726
rect 4528 16662 4580 16668
rect 4448 16544 4568 16572
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4448 15706 4476 16390
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4344 15632 4396 15638
rect 4250 15600 4306 15609
rect 4160 15564 4212 15570
rect 4344 15574 4396 15580
rect 4250 15535 4306 15544
rect 4160 15506 4212 15512
rect 4068 15428 4120 15434
rect 4068 15370 4120 15376
rect 4264 15366 4292 15535
rect 4540 15484 4568 16544
rect 4356 15456 4568 15484
rect 3976 15360 4028 15366
rect 3976 15302 4028 15308
rect 4252 15360 4304 15366
rect 4252 15302 4304 15308
rect 3424 15088 3476 15094
rect 3424 15030 3476 15036
rect 3160 14878 3280 14906
rect 3332 14952 3384 14958
rect 3332 14894 3384 14900
rect 3160 14385 3188 14878
rect 3240 14816 3292 14822
rect 3240 14758 3292 14764
rect 3146 14376 3202 14385
rect 3146 14311 3202 14320
rect 3252 14278 3280 14758
rect 3344 14618 3372 14894
rect 3332 14612 3384 14618
rect 3332 14554 3384 14560
rect 3332 14340 3384 14346
rect 3332 14282 3384 14288
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 3068 14062 3280 14090
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 2964 12436 3016 12442
rect 2964 12378 3016 12384
rect 2976 12102 3004 12378
rect 2964 12096 3016 12102
rect 2964 12038 3016 12044
rect 3160 11898 3188 12786
rect 3252 12434 3280 14062
rect 3344 13938 3372 14282
rect 3436 14074 3464 15030
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3700 14952 3752 14958
rect 3514 14920 3570 14929
rect 3752 14900 3924 14906
rect 3700 14894 3924 14900
rect 3712 14878 3924 14894
rect 3514 14855 3516 14864
rect 3568 14855 3570 14864
rect 3516 14826 3568 14832
rect 3549 14716 3857 14736
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14640 3857 14660
rect 3896 14618 3924 14878
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3882 14376 3938 14385
rect 3882 14311 3938 14320
rect 3896 14278 3924 14311
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3620 14074 3648 14214
rect 3988 14074 4016 14962
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4080 14482 4108 14894
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4172 13938 4200 14010
rect 3332 13932 3384 13938
rect 3332 13874 3384 13880
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 3516 13864 3568 13870
rect 3436 13824 3516 13852
rect 3436 13530 3464 13824
rect 3516 13806 3568 13812
rect 3549 13628 3857 13648
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13552 3857 13572
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3436 13394 3464 13466
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 4264 12730 4292 15302
rect 3988 12702 4292 12730
rect 3549 12540 3857 12560
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12464 3857 12484
rect 3332 12436 3384 12442
rect 3252 12406 3332 12434
rect 3332 12378 3384 12384
rect 3332 12232 3384 12238
rect 3332 12174 3384 12180
rect 3148 11892 3200 11898
rect 3148 11834 3200 11840
rect 3344 11694 3372 12174
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3056 11620 3108 11626
rect 3056 11562 3108 11568
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2976 9994 3004 11494
rect 3068 11218 3096 11562
rect 3549 11452 3857 11472
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11376 3857 11396
rect 3424 11280 3476 11286
rect 3424 11222 3476 11228
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 3332 11076 3384 11082
rect 3332 11018 3384 11024
rect 3240 10668 3292 10674
rect 3240 10610 3292 10616
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2778 9752 2834 9761
rect 2778 9687 2834 9696
rect 3056 9716 3108 9722
rect 2688 9444 2740 9450
rect 2688 9386 2740 9392
rect 2792 9178 2820 9687
rect 3056 9658 3108 9664
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2780 9172 2832 9178
rect 2780 9114 2832 9120
rect 2884 9110 2912 9522
rect 2872 9104 2924 9110
rect 2872 9046 2924 9052
rect 3068 9042 3096 9658
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 3056 9036 3108 9042
rect 3056 8978 3108 8984
rect 2872 8968 2924 8974
rect 2872 8910 2924 8916
rect 2964 8968 3016 8974
rect 2964 8910 3016 8916
rect 2884 8090 2912 8910
rect 2976 8809 3004 8910
rect 2962 8800 3018 8809
rect 2962 8735 3018 8744
rect 3068 8566 3096 8978
rect 3056 8560 3108 8566
rect 3056 8502 3108 8508
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2872 8084 2924 8090
rect 2872 8026 2924 8032
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2686 7712 2742 7721
rect 2686 7647 2742 7656
rect 2596 7336 2648 7342
rect 2596 7278 2648 7284
rect 2504 7268 2556 7274
rect 2504 7210 2556 7216
rect 2504 6860 2556 6866
rect 2504 6802 2556 6808
rect 2516 4690 2544 6802
rect 2700 6610 2728 7647
rect 2608 6582 2728 6610
rect 2608 6458 2636 6582
rect 2792 6474 2820 7822
rect 2596 6452 2648 6458
rect 2596 6394 2648 6400
rect 2700 6446 2820 6474
rect 2700 6390 2728 6446
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 2596 5908 2648 5914
rect 2700 5896 2728 6326
rect 2792 6118 2820 6326
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2884 5930 2912 7890
rect 2976 7342 3004 8434
rect 3056 7540 3108 7546
rect 3160 7528 3188 9522
rect 3252 8974 3280 10610
rect 3344 10470 3372 11018
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3436 9500 3464 11222
rect 3988 11218 4016 12702
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 4080 12102 4108 12582
rect 4356 12434 4384 15456
rect 4632 14498 4660 17138
rect 4448 14470 4660 14498
rect 4448 13530 4476 14470
rect 4528 14408 4580 14414
rect 4528 14350 4580 14356
rect 4436 13524 4488 13530
rect 4436 13466 4488 13472
rect 4264 12406 4384 12434
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4080 11626 4108 12038
rect 4068 11620 4120 11626
rect 4068 11562 4120 11568
rect 3608 11212 3660 11218
rect 3608 11154 3660 11160
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3620 11014 3648 11154
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 3792 11008 3844 11014
rect 3988 10985 4016 11154
rect 3792 10950 3844 10956
rect 3974 10976 4030 10985
rect 3804 10674 3832 10950
rect 3974 10911 4030 10920
rect 3792 10668 3844 10674
rect 4080 10656 4108 11562
rect 3792 10610 3844 10616
rect 3988 10628 4108 10656
rect 3988 10538 4016 10628
rect 3976 10532 4028 10538
rect 3976 10474 4028 10480
rect 4068 10532 4120 10538
rect 4068 10474 4120 10480
rect 3884 10464 3936 10470
rect 3884 10406 3936 10412
rect 3549 10364 3857 10384
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10288 3857 10308
rect 3896 10266 3924 10406
rect 3884 10260 3936 10266
rect 3884 10202 3936 10208
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3620 10033 3648 10066
rect 3606 10024 3662 10033
rect 3344 9472 3464 9500
rect 3528 9982 3606 10010
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 7886 3280 8774
rect 3344 7886 3372 9472
rect 3528 9364 3556 9982
rect 3606 9959 3662 9968
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3804 9466 3832 9862
rect 3896 9586 3924 10202
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3804 9438 3924 9466
rect 3436 9336 3556 9364
rect 3436 8974 3464 9336
rect 3549 9276 3857 9296
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9200 3857 9220
rect 3896 8974 3924 9438
rect 3988 9178 4016 10202
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3884 8968 3936 8974
rect 3884 8910 3936 8916
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3436 7954 3464 8434
rect 3549 8188 3857 8208
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8112 3857 8132
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3514 7848 3570 7857
rect 3344 7750 3372 7822
rect 3514 7783 3570 7792
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3528 7546 3556 7783
rect 3108 7500 3188 7528
rect 3240 7540 3292 7546
rect 3056 7482 3108 7488
rect 3240 7482 3292 7488
rect 3516 7540 3568 7546
rect 3516 7482 3568 7488
rect 2964 7336 3016 7342
rect 3016 7296 3096 7324
rect 2964 7278 3016 7284
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2648 5868 2728 5896
rect 2792 5902 2912 5930
rect 2596 5850 2648 5856
rect 2792 5409 2820 5902
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2778 5400 2834 5409
rect 2688 5364 2740 5370
rect 2778 5335 2834 5344
rect 2688 5306 2740 5312
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2504 4684 2556 4690
rect 2504 4626 2556 4632
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2410 4312 2466 4321
rect 2410 4247 2412 4256
rect 2464 4247 2466 4256
rect 2412 4218 2464 4224
rect 2228 4004 2280 4010
rect 2228 3946 2280 3952
rect 2044 3936 2096 3942
rect 2240 3913 2268 3946
rect 2044 3878 2096 3884
rect 2226 3904 2282 3913
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 1964 3126 1992 3538
rect 2056 3194 2084 3878
rect 2226 3839 2282 3848
rect 2136 3732 2188 3738
rect 2136 3674 2188 3680
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 1952 3120 2004 3126
rect 1858 3088 1914 3097
rect 1952 3062 2004 3068
rect 1858 3023 1914 3032
rect 2148 2774 2176 3674
rect 2516 3534 2544 4626
rect 2504 3528 2556 3534
rect 2226 3496 2282 3505
rect 2504 3470 2556 3476
rect 2226 3431 2282 3440
rect 2240 2825 2268 3431
rect 1688 2746 1808 2774
rect 2056 2746 2176 2774
rect 2226 2816 2282 2825
rect 2608 2774 2636 5170
rect 2700 4729 2728 5306
rect 2778 5264 2834 5273
rect 2778 5199 2834 5208
rect 2686 4720 2742 4729
rect 2686 4655 2742 4664
rect 2700 4554 2728 4655
rect 2688 4548 2740 4554
rect 2688 4490 2740 4496
rect 2792 4457 2820 5199
rect 2884 4672 2912 5510
rect 2976 4826 3004 6598
rect 3068 6186 3096 7296
rect 3252 6746 3280 7482
rect 3896 7478 3924 8774
rect 3988 8401 4016 8842
rect 3974 8392 4030 8401
rect 3974 8327 4030 8336
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3344 7002 3372 7278
rect 3332 6996 3384 7002
rect 3436 6984 3464 7278
rect 3549 7100 3857 7120
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7024 3857 7044
rect 3436 6956 3556 6984
rect 3332 6938 3384 6944
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3160 6718 3280 6746
rect 3160 6458 3188 6718
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3056 6180 3108 6186
rect 3056 6122 3108 6128
rect 3054 5808 3110 5817
rect 3054 5743 3110 5752
rect 3068 5642 3096 5743
rect 3056 5636 3108 5642
rect 3056 5578 3108 5584
rect 3252 5114 3280 6598
rect 3344 5370 3372 6598
rect 3436 6254 3464 6802
rect 3424 6248 3476 6254
rect 3424 6190 3476 6196
rect 3528 6100 3556 6956
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3712 6186 3740 6734
rect 3792 6656 3844 6662
rect 3792 6598 3844 6604
rect 3804 6458 3832 6598
rect 3792 6452 3844 6458
rect 3792 6394 3844 6400
rect 3700 6180 3752 6186
rect 3700 6122 3752 6128
rect 3436 6072 3556 6100
rect 3332 5364 3384 5370
rect 3332 5306 3384 5312
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3056 5092 3108 5098
rect 3056 5034 3108 5040
rect 3160 5086 3280 5114
rect 2964 4820 3016 4826
rect 2964 4762 3016 4768
rect 3068 4758 3096 5034
rect 3160 4758 3188 5086
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 3148 4752 3200 4758
rect 3148 4694 3200 4700
rect 2884 4644 3004 4672
rect 2872 4548 2924 4554
rect 2872 4490 2924 4496
rect 2778 4448 2834 4457
rect 2778 4383 2834 4392
rect 2884 4282 2912 4490
rect 2872 4276 2924 4282
rect 2872 4218 2924 4224
rect 2870 4040 2926 4049
rect 2976 4026 3004 4644
rect 2926 3998 3004 4026
rect 3068 4010 3096 4694
rect 3252 4622 3280 4966
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3160 4282 3188 4422
rect 3252 4282 3280 4422
rect 3148 4276 3200 4282
rect 3148 4218 3200 4224
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3146 4176 3202 4185
rect 3146 4111 3148 4120
rect 3200 4111 3202 4120
rect 3148 4082 3200 4088
rect 3240 4072 3292 4078
rect 3240 4014 3292 4020
rect 3056 4004 3108 4010
rect 2870 3975 2926 3984
rect 3056 3946 3108 3952
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2872 3392 2924 3398
rect 2872 3334 2924 3340
rect 2226 2751 2282 2760
rect 1584 1760 1636 1766
rect 1584 1702 1636 1708
rect 1688 1578 1716 2746
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 1964 2038 1992 2382
rect 1952 2032 2004 2038
rect 1952 1974 2004 1980
rect 1596 1550 1716 1578
rect 1490 1184 1546 1193
rect 1490 1119 1546 1128
rect 1596 800 1624 1550
rect 2056 800 2084 2746
rect 2240 2514 2268 2751
rect 2516 2746 2636 2774
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2516 800 2544 2746
rect 2884 2553 2912 3334
rect 2870 2544 2926 2553
rect 2870 2479 2926 2488
rect 2976 1465 3004 3470
rect 3068 2922 3096 3946
rect 3252 3194 3280 4014
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3240 2984 3292 2990
rect 3238 2952 3240 2961
rect 3292 2952 3294 2961
rect 3056 2916 3108 2922
rect 3238 2887 3294 2896
rect 3056 2858 3108 2864
rect 3344 2774 3372 5170
rect 3436 4593 3464 6072
rect 3549 6012 3857 6032
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5936 3857 5956
rect 3516 5840 3568 5846
rect 3516 5782 3568 5788
rect 3528 5409 3556 5782
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3620 5574 3648 5714
rect 3608 5568 3660 5574
rect 3608 5510 3660 5516
rect 3514 5400 3570 5409
rect 3514 5335 3570 5344
rect 3620 5273 3648 5510
rect 3792 5296 3844 5302
rect 3606 5264 3662 5273
rect 3792 5238 3844 5244
rect 3606 5199 3662 5208
rect 3804 5098 3832 5238
rect 3792 5092 3844 5098
rect 3792 5034 3844 5040
rect 3549 4924 3857 4944
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4848 3857 4868
rect 3896 4826 3924 7278
rect 3988 6934 4016 7346
rect 3976 6928 4028 6934
rect 3976 6870 4028 6876
rect 3974 6624 4030 6633
rect 3974 6559 4030 6568
rect 3988 5574 4016 6559
rect 4080 5914 4108 10474
rect 4172 9654 4200 12106
rect 4264 11558 4292 12406
rect 4252 11552 4304 11558
rect 4252 11494 4304 11500
rect 4448 11286 4476 13466
rect 4436 11280 4488 11286
rect 4436 11222 4488 11228
rect 4540 11098 4568 14350
rect 4620 14340 4672 14346
rect 4620 14282 4672 14288
rect 4448 11070 4568 11098
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4160 9648 4212 9654
rect 4160 9590 4212 9596
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4172 8634 4200 8774
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 4172 8401 4200 8434
rect 4158 8392 4214 8401
rect 4158 8327 4214 8336
rect 4264 8090 4292 8774
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4252 7744 4304 7750
rect 4250 7712 4252 7721
rect 4304 7712 4306 7721
rect 4250 7647 4306 7656
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4264 7206 4292 7346
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4160 6996 4212 7002
rect 4160 6938 4212 6944
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3976 5160 4028 5166
rect 3976 5102 4028 5108
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3422 4584 3478 4593
rect 3422 4519 3478 4528
rect 3436 3738 3464 4519
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3549 3836 3857 3856
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3760 3857 3780
rect 3896 3738 3924 4422
rect 3424 3732 3476 3738
rect 3424 3674 3476 3680
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3422 3088 3478 3097
rect 3422 3023 3478 3032
rect 3252 2746 3372 2774
rect 3054 2544 3110 2553
rect 3054 2479 3110 2488
rect 3068 1601 3096 2479
rect 3148 2440 3200 2446
rect 3146 2408 3148 2417
rect 3200 2408 3202 2417
rect 3146 2343 3202 2352
rect 3252 2258 3280 2746
rect 3436 2530 3464 3023
rect 3549 2748 3857 2768
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2672 3857 2692
rect 3436 2502 3556 2530
rect 3422 2408 3478 2417
rect 3160 2230 3280 2258
rect 3344 2352 3422 2360
rect 3344 2332 3424 2352
rect 3160 1873 3188 2230
rect 3240 2100 3292 2106
rect 3240 2042 3292 2048
rect 3146 1864 3202 1873
rect 3146 1799 3202 1808
rect 3252 1737 3280 2042
rect 3238 1728 3294 1737
rect 3238 1663 3294 1672
rect 3054 1592 3110 1601
rect 3054 1527 3110 1536
rect 2962 1456 3018 1465
rect 2962 1391 3018 1400
rect 2976 800 3004 1391
rect 202 0 258 800
rect 662 0 718 800
rect 1122 0 1178 800
rect 1582 0 1638 800
rect 2042 0 2098 800
rect 2502 0 2558 800
rect 2962 0 3018 800
rect 3344 649 3372 2332
rect 3476 2343 3478 2352
rect 3424 2314 3476 2320
rect 3422 1864 3478 1873
rect 3422 1799 3478 1808
rect 3436 800 3464 1799
rect 3528 1630 3556 2502
rect 3516 1624 3568 1630
rect 3516 1566 3568 1572
rect 3896 800 3924 3470
rect 3988 3466 4016 5102
rect 4080 4554 4108 5850
rect 4172 4826 4200 6938
rect 4356 6866 4384 10746
rect 4448 9654 4476 11070
rect 4632 10538 4660 14282
rect 4724 12696 4752 18634
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4816 17814 4844 18226
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4908 18086 4936 18158
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4804 17808 4856 17814
rect 4856 17768 4936 17796
rect 4804 17750 4856 17756
rect 4802 17096 4858 17105
rect 4802 17031 4804 17040
rect 4856 17031 4858 17040
rect 4804 17002 4856 17008
rect 4804 16652 4856 16658
rect 4804 16594 4856 16600
rect 4816 16250 4844 16594
rect 4804 16244 4856 16250
rect 4804 16186 4856 16192
rect 4908 14600 4936 17768
rect 5000 15638 5028 18702
rect 5080 18624 5132 18630
rect 5080 18566 5132 18572
rect 5092 18222 5120 18566
rect 5080 18216 5132 18222
rect 5080 18158 5132 18164
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 5092 17134 5120 17478
rect 5080 17128 5132 17134
rect 5080 17070 5132 17076
rect 5080 16584 5132 16590
rect 5080 16526 5132 16532
rect 5092 15706 5120 16526
rect 5080 15700 5132 15706
rect 5080 15642 5132 15648
rect 4988 15632 5040 15638
rect 4988 15574 5040 15580
rect 5184 15473 5212 20334
rect 5276 19281 5304 22200
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5460 19961 5488 20402
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5632 20392 5684 20398
rect 5632 20334 5684 20340
rect 5552 20058 5580 20334
rect 5540 20052 5592 20058
rect 5540 19994 5592 20000
rect 5446 19952 5502 19961
rect 5446 19887 5502 19896
rect 5540 19780 5592 19786
rect 5540 19722 5592 19728
rect 5356 19712 5408 19718
rect 5356 19654 5408 19660
rect 5262 19272 5318 19281
rect 5262 19207 5318 19216
rect 5264 17672 5316 17678
rect 5264 17614 5316 17620
rect 5276 16250 5304 17614
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5170 15464 5226 15473
rect 5170 15399 5226 15408
rect 4908 14572 5120 14600
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4908 13530 4936 14214
rect 5000 14074 5028 14418
rect 4988 14068 5040 14074
rect 4988 14010 5040 14016
rect 4896 13524 4948 13530
rect 4896 13466 4948 13472
rect 4896 12844 4948 12850
rect 4896 12786 4948 12792
rect 4804 12708 4856 12714
rect 4724 12668 4804 12696
rect 4804 12650 4856 12656
rect 4712 12096 4764 12102
rect 4712 12038 4764 12044
rect 4724 11898 4752 12038
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4724 11558 4752 11834
rect 4816 11665 4844 12650
rect 4802 11656 4858 11665
rect 4802 11591 4858 11600
rect 4712 11552 4764 11558
rect 4710 11520 4712 11529
rect 4804 11552 4856 11558
rect 4764 11520 4766 11529
rect 4804 11494 4856 11500
rect 4710 11455 4766 11464
rect 4712 11076 4764 11082
rect 4712 11018 4764 11024
rect 4620 10532 4672 10538
rect 4620 10474 4672 10480
rect 4724 10418 4752 11018
rect 4540 10390 4752 10418
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 4448 8498 4476 9590
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4448 7002 4476 7142
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4250 6760 4306 6769
rect 4250 6695 4306 6704
rect 4264 6225 4292 6695
rect 4540 6662 4568 10390
rect 4816 9586 4844 11494
rect 4908 11218 4936 12786
rect 5092 12646 5120 14572
rect 5368 14278 5396 19654
rect 5552 19496 5580 19722
rect 5644 19514 5672 20334
rect 5736 20097 5764 22200
rect 6196 22114 6224 22200
rect 6288 22114 6316 22222
rect 6196 22086 6316 22114
rect 6148 20700 6456 20720
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20624 6456 20644
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 5908 20324 5960 20330
rect 5908 20266 5960 20272
rect 5816 20256 5868 20262
rect 5816 20198 5868 20204
rect 5722 20088 5778 20097
rect 5722 20023 5778 20032
rect 5460 19468 5580 19496
rect 5632 19508 5684 19514
rect 5460 19174 5488 19468
rect 5632 19450 5684 19456
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5552 19174 5580 19314
rect 5448 19168 5500 19174
rect 5448 19110 5500 19116
rect 5540 19168 5592 19174
rect 5540 19110 5592 19116
rect 5632 18216 5684 18222
rect 5632 18158 5684 18164
rect 5540 17740 5592 17746
rect 5540 17682 5592 17688
rect 5552 17626 5580 17682
rect 5460 17598 5580 17626
rect 5460 16998 5488 17598
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5448 16992 5500 16998
rect 5448 16934 5500 16940
rect 5552 16590 5580 17478
rect 5540 16584 5592 16590
rect 5540 16526 5592 16532
rect 5644 16182 5672 18158
rect 5722 17368 5778 17377
rect 5722 17303 5778 17312
rect 5632 16176 5684 16182
rect 5632 16118 5684 16124
rect 5448 16108 5500 16114
rect 5448 16050 5500 16056
rect 5460 15065 5488 16050
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5552 15570 5580 15642
rect 5540 15564 5592 15570
rect 5540 15506 5592 15512
rect 5446 15056 5502 15065
rect 5446 14991 5502 15000
rect 5460 14890 5488 14991
rect 5448 14884 5500 14890
rect 5448 14826 5500 14832
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5448 14340 5500 14346
rect 5448 14282 5500 14288
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5080 12640 5132 12646
rect 5080 12582 5132 12588
rect 4986 11792 5042 11801
rect 4986 11727 5042 11736
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4908 10742 4936 11154
rect 5000 10996 5028 11727
rect 5092 11354 5120 12582
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5080 11348 5132 11354
rect 5080 11290 5132 11296
rect 5080 11008 5132 11014
rect 5000 10968 5080 10996
rect 5080 10950 5132 10956
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 4988 10668 5040 10674
rect 4988 10610 5040 10616
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 5000 9382 5028 10610
rect 5080 9988 5132 9994
rect 5080 9930 5132 9936
rect 5092 9654 5120 9930
rect 5080 9648 5132 9654
rect 5080 9590 5132 9596
rect 4988 9376 5040 9382
rect 4894 9344 4950 9353
rect 4988 9318 5040 9324
rect 4894 9279 4950 9288
rect 4712 8900 4764 8906
rect 4632 8860 4712 8888
rect 4632 8498 4660 8860
rect 4712 8842 4764 8848
rect 4908 8616 4936 9279
rect 5184 8650 5212 11834
rect 5276 10742 5304 14214
rect 5356 13932 5408 13938
rect 5460 13920 5488 14282
rect 5408 13892 5488 13920
rect 5540 13932 5592 13938
rect 5356 13874 5408 13880
rect 5540 13874 5592 13880
rect 5552 13394 5580 13874
rect 5644 13852 5672 14350
rect 5736 13954 5764 17303
rect 5828 15994 5856 20198
rect 5920 19378 5948 20266
rect 6380 19922 6408 20402
rect 6564 20369 6592 22222
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7562 22200 7618 23000
rect 8022 22200 8078 23000
rect 8482 22200 8538 23000
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9862 22200 9918 23000
rect 10322 22200 10378 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12162 22200 12218 23000
rect 12622 22200 12678 23000
rect 13082 22200 13138 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14462 22200 14518 23000
rect 14922 22200 14978 23000
rect 15382 22200 15438 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 17222 22200 17278 23000
rect 17682 22200 17738 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 19062 22200 19118 23000
rect 19522 22200 19578 23000
rect 19982 22200 20038 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21362 22200 21418 23000
rect 21822 22200 21878 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 6656 20602 6684 22200
rect 7116 20618 7144 22200
rect 6644 20596 6696 20602
rect 6644 20538 6696 20544
rect 7024 20590 7144 20618
rect 7576 20602 7604 22200
rect 7564 20596 7616 20602
rect 6550 20360 6606 20369
rect 6550 20295 6606 20304
rect 6368 19916 6420 19922
rect 6368 19858 6420 19864
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 5908 19372 5960 19378
rect 5908 19314 5960 19320
rect 6012 18426 6040 19790
rect 6148 19612 6456 19632
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19536 6456 19556
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6182 19272 6238 19281
rect 6182 19207 6184 19216
rect 6236 19207 6238 19216
rect 6184 19178 6236 19184
rect 6472 18766 6500 19314
rect 6552 19304 6604 19310
rect 6552 19246 6604 19252
rect 6564 18834 6592 19246
rect 6656 18850 6684 20538
rect 6826 20496 6882 20505
rect 6826 20431 6882 20440
rect 6734 20088 6790 20097
rect 6734 20023 6790 20032
rect 6748 18970 6776 20023
rect 6840 19854 6868 20431
rect 6828 19848 6880 19854
rect 6828 19790 6880 19796
rect 6828 19712 6880 19718
rect 6880 19660 6960 19666
rect 6828 19654 6960 19660
rect 6840 19638 6960 19654
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6552 18828 6604 18834
rect 6656 18822 6776 18850
rect 6552 18770 6604 18776
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6644 18760 6696 18766
rect 6644 18702 6696 18708
rect 6552 18692 6604 18698
rect 6552 18634 6604 18640
rect 6148 18524 6456 18544
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18448 6456 18468
rect 6000 18420 6052 18426
rect 6000 18362 6052 18368
rect 6564 18290 6592 18634
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6564 17921 6592 18226
rect 6550 17912 6606 17921
rect 6550 17847 6606 17856
rect 6656 17746 6684 18702
rect 6644 17740 6696 17746
rect 6644 17682 6696 17688
rect 6748 17626 6776 18822
rect 6840 18426 6868 19110
rect 6932 19009 6960 19638
rect 6918 19000 6974 19009
rect 6918 18935 6974 18944
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 6828 18284 6880 18290
rect 6828 18226 6880 18232
rect 6564 17598 6776 17626
rect 6148 17436 6456 17456
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17360 6456 17380
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 6092 17128 6144 17134
rect 6092 17070 6144 17076
rect 6104 16794 6132 17070
rect 6196 16998 6224 17138
rect 6184 16992 6236 16998
rect 6184 16934 6236 16940
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6104 16590 6132 16730
rect 6092 16584 6144 16590
rect 6288 16561 6316 17138
rect 6092 16526 6144 16532
rect 6274 16552 6330 16561
rect 6274 16487 6330 16496
rect 6148 16348 6456 16368
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16272 6456 16292
rect 6564 16182 6592 17598
rect 6644 17536 6696 17542
rect 6644 17478 6696 17484
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6656 17270 6684 17478
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6748 16266 6776 17478
rect 6840 17202 6868 18226
rect 6932 18222 6960 18935
rect 7024 18698 7052 20590
rect 7564 20538 7616 20544
rect 7104 20460 7156 20466
rect 7104 20402 7156 20408
rect 7116 19922 7144 20402
rect 7576 20398 7604 20538
rect 7564 20392 7616 20398
rect 8036 20380 8064 22200
rect 8300 20392 8352 20398
rect 8036 20352 8300 20380
rect 7564 20334 7616 20340
rect 8352 20352 8432 20380
rect 8300 20334 8352 20340
rect 7840 20256 7892 20262
rect 7840 20198 7892 20204
rect 7104 19916 7156 19922
rect 7104 19858 7156 19864
rect 7116 19514 7144 19858
rect 7380 19712 7432 19718
rect 7380 19654 7432 19660
rect 7104 19508 7156 19514
rect 7104 19450 7156 19456
rect 7012 18692 7064 18698
rect 7012 18634 7064 18640
rect 7102 18592 7158 18601
rect 7102 18527 7158 18536
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6826 16688 6882 16697
rect 6826 16623 6882 16632
rect 6840 16522 6868 16623
rect 6828 16516 6880 16522
rect 6828 16458 6880 16464
rect 6656 16238 6776 16266
rect 6552 16176 6604 16182
rect 6552 16118 6604 16124
rect 6552 16040 6604 16046
rect 5828 15966 5948 15994
rect 6552 15982 6604 15988
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 5828 14414 5856 15846
rect 5816 14408 5868 14414
rect 5816 14350 5868 14356
rect 5736 13926 5856 13954
rect 5724 13864 5776 13870
rect 5644 13824 5724 13852
rect 5724 13806 5776 13812
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 12481 5488 13262
rect 5446 12472 5502 12481
rect 5552 12442 5580 13330
rect 5632 13252 5684 13258
rect 5632 13194 5684 13200
rect 5446 12407 5502 12416
rect 5540 12436 5592 12442
rect 5460 12322 5488 12407
rect 5540 12378 5592 12384
rect 5644 12345 5672 13194
rect 5736 13190 5764 13806
rect 5828 13190 5856 13926
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5736 12918 5764 13126
rect 5828 12986 5856 13126
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 5630 12336 5686 12345
rect 5460 12306 5580 12322
rect 5460 12300 5592 12306
rect 5460 12294 5540 12300
rect 5630 12271 5686 12280
rect 5540 12242 5592 12248
rect 5736 12238 5764 12854
rect 5920 12434 5948 15966
rect 6000 15360 6052 15366
rect 6000 15302 6052 15308
rect 6012 15162 6040 15302
rect 6148 15260 6456 15280
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15184 6456 15204
rect 6564 15162 6592 15982
rect 6000 15156 6052 15162
rect 6000 15098 6052 15104
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6656 14618 6684 16238
rect 6736 16108 6788 16114
rect 6736 16050 6788 16056
rect 6932 16096 6960 18158
rect 7012 18148 7064 18154
rect 7012 18090 7064 18096
rect 7024 17542 7052 18090
rect 7116 18057 7144 18527
rect 7196 18080 7248 18086
rect 7102 18048 7158 18057
rect 7196 18022 7248 18028
rect 7102 17983 7158 17992
rect 7208 17678 7236 18022
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7012 17536 7064 17542
rect 7012 17478 7064 17484
rect 7024 16590 7052 17478
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7116 16998 7144 17274
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 7012 16108 7064 16114
rect 6932 16068 7012 16096
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6148 14172 6456 14192
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14096 6456 14116
rect 6552 13796 6604 13802
rect 6552 13738 6604 13744
rect 6148 13084 6456 13104
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13008 6456 13028
rect 6564 12714 6592 13738
rect 6644 13320 6696 13326
rect 6644 13262 6696 13268
rect 6552 12708 6604 12714
rect 6552 12650 6604 12656
rect 5920 12406 6040 12434
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5644 11830 5672 12106
rect 5632 11824 5684 11830
rect 5632 11766 5684 11772
rect 5448 11756 5500 11762
rect 5448 11698 5500 11704
rect 5540 11756 5592 11762
rect 5540 11698 5592 11704
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5368 10810 5396 11630
rect 5460 11354 5488 11698
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5552 11082 5580 11698
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5816 11620 5868 11626
rect 5816 11562 5868 11568
rect 5632 11552 5684 11558
rect 5632 11494 5684 11500
rect 5540 11076 5592 11082
rect 5540 11018 5592 11024
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5552 10198 5580 10542
rect 5540 10192 5592 10198
rect 5540 10134 5592 10140
rect 5264 10056 5316 10062
rect 5448 10056 5500 10062
rect 5264 9998 5316 10004
rect 5368 10016 5448 10044
rect 5276 9722 5304 9998
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5264 9376 5316 9382
rect 5262 9344 5264 9353
rect 5316 9344 5318 9353
rect 5262 9279 5318 9288
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 4816 8588 4936 8616
rect 4988 8628 5040 8634
rect 4620 8492 4672 8498
rect 4620 8434 4672 8440
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4344 6452 4396 6458
rect 4344 6394 4396 6400
rect 4250 6216 4306 6225
rect 4250 6151 4306 6160
rect 4264 5710 4292 6151
rect 4252 5704 4304 5710
rect 4252 5646 4304 5652
rect 4356 5574 4384 6394
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4448 5914 4476 6122
rect 4540 6089 4568 6258
rect 4526 6080 4582 6089
rect 4526 6015 4582 6024
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4436 5704 4488 5710
rect 4436 5646 4488 5652
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4448 5352 4476 5646
rect 4356 5324 4476 5352
rect 4356 5098 4384 5324
rect 4434 5264 4490 5273
rect 4434 5199 4436 5208
rect 4488 5199 4490 5208
rect 4436 5170 4488 5176
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4160 4820 4212 4826
rect 4160 4762 4212 4768
rect 4158 4584 4214 4593
rect 4068 4548 4120 4554
rect 4158 4519 4214 4528
rect 4068 4490 4120 4496
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 4080 4049 4108 4082
rect 4066 4040 4122 4049
rect 4066 3975 4122 3984
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3976 3460 4028 3466
rect 3976 3402 4028 3408
rect 3974 2680 4030 2689
rect 3974 2615 3976 2624
rect 4028 2615 4030 2624
rect 3976 2586 4028 2592
rect 4080 2514 4108 3878
rect 4172 3534 4200 4519
rect 4264 4486 4292 4966
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4356 4078 4384 5034
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4448 4214 4476 4762
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4252 4072 4304 4078
rect 4252 4014 4304 4020
rect 4344 4072 4396 4078
rect 4344 4014 4396 4020
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4160 3392 4212 3398
rect 4160 3334 4212 3340
rect 4172 3126 4200 3334
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4264 2922 4292 4014
rect 4436 4004 4488 4010
rect 4436 3946 4488 3952
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 4356 2582 4384 3538
rect 4448 3534 4476 3946
rect 4540 3670 4568 6015
rect 4632 5137 4660 8434
rect 4712 8424 4764 8430
rect 4816 8412 4844 8588
rect 4988 8570 5040 8576
rect 5092 8622 5212 8650
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4764 8384 4844 8412
rect 4712 8366 4764 8372
rect 4712 7744 4764 7750
rect 4712 7686 4764 7692
rect 4618 5128 4674 5137
rect 4618 5063 4674 5072
rect 4618 4992 4674 5001
rect 4618 4927 4674 4936
rect 4632 4554 4660 4927
rect 4724 4758 4752 7686
rect 4802 7304 4858 7313
rect 4802 7239 4858 7248
rect 4816 6458 4844 7239
rect 4908 6866 4936 8434
rect 5000 7546 5028 8570
rect 5092 7970 5120 8622
rect 5170 8392 5226 8401
rect 5170 8327 5226 8336
rect 5184 8090 5212 8327
rect 5172 8084 5224 8090
rect 5172 8026 5224 8032
rect 5092 7942 5212 7970
rect 5080 7812 5132 7818
rect 5080 7754 5132 7760
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 5000 6769 5028 6870
rect 4986 6760 5042 6769
rect 4986 6695 5042 6704
rect 4894 6488 4950 6497
rect 4804 6452 4856 6458
rect 4894 6423 4950 6432
rect 4804 6394 4856 6400
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4816 5710 4844 6190
rect 4908 5817 4936 6423
rect 5000 5953 5028 6695
rect 4986 5944 5042 5953
rect 4986 5879 5042 5888
rect 4894 5808 4950 5817
rect 4894 5743 4896 5752
rect 4948 5743 4950 5752
rect 4896 5714 4948 5720
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4816 5409 4844 5646
rect 4802 5400 4858 5409
rect 4802 5335 4858 5344
rect 4816 5234 4844 5335
rect 4804 5228 4856 5234
rect 4804 5170 4856 5176
rect 4896 5228 4948 5234
rect 5000 5216 5028 5879
rect 4948 5188 5028 5216
rect 4896 5170 4948 5176
rect 4712 4752 4764 4758
rect 4712 4694 4764 4700
rect 4908 4690 4936 5170
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4896 4684 4948 4690
rect 4896 4626 4948 4632
rect 4620 4548 4672 4554
rect 4620 4490 4672 4496
rect 4712 4548 4764 4554
rect 4712 4490 4764 4496
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4632 3398 4660 3878
rect 4724 3670 4752 4490
rect 4896 4208 4948 4214
rect 4896 4150 4948 4156
rect 4804 3936 4856 3942
rect 4804 3878 4856 3884
rect 4712 3664 4764 3670
rect 4712 3606 4764 3612
rect 4620 3392 4672 3398
rect 4816 3369 4844 3878
rect 4908 3505 4936 4150
rect 4894 3496 4950 3505
rect 4894 3431 4950 3440
rect 4620 3334 4672 3340
rect 4802 3360 4858 3369
rect 4802 3295 4858 3304
rect 5000 3210 5028 4762
rect 4632 3182 5028 3210
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 4344 2576 4396 2582
rect 4344 2518 4396 2524
rect 4068 2508 4120 2514
rect 4068 2450 4120 2456
rect 4448 1442 4476 2926
rect 4632 2446 4660 3182
rect 5092 2774 5120 7754
rect 5184 7002 5212 7942
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5172 6112 5224 6118
rect 5276 6089 5304 9114
rect 5368 7410 5396 10016
rect 5644 10033 5672 11494
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5736 10962 5764 11154
rect 5828 11082 5856 11562
rect 5920 11150 5948 11630
rect 6012 11370 6040 12406
rect 6564 12170 6592 12650
rect 6656 12646 6684 13262
rect 6748 12986 6776 16050
rect 6828 15428 6880 15434
rect 6828 15370 6880 15376
rect 6840 14346 6868 15370
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6644 12640 6696 12646
rect 6644 12582 6696 12588
rect 6644 12436 6696 12442
rect 6644 12378 6696 12384
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6148 11996 6456 12016
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11920 6456 11940
rect 6012 11354 6132 11370
rect 6012 11348 6144 11354
rect 6012 11342 6092 11348
rect 6092 11290 6144 11296
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 6656 11014 6684 12378
rect 6840 12170 6868 12650
rect 6828 12164 6880 12170
rect 6828 12106 6880 12112
rect 6840 11218 6868 12106
rect 6932 11778 6960 16068
rect 7012 16050 7064 16056
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 7104 15428 7156 15434
rect 7104 15370 7156 15376
rect 7024 13326 7052 15370
rect 7116 14822 7144 15370
rect 7104 14816 7156 14822
rect 7104 14758 7156 14764
rect 7196 14544 7248 14550
rect 7196 14486 7248 14492
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 7012 12776 7064 12782
rect 7012 12718 7064 12724
rect 7024 12442 7052 12718
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7116 11898 7144 13670
rect 7208 12782 7236 14486
rect 7288 13932 7340 13938
rect 7288 13874 7340 13880
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7300 12102 7328 13874
rect 7392 12442 7420 19654
rect 7562 18864 7618 18873
rect 7562 18799 7618 18808
rect 7576 18329 7604 18799
rect 7852 18698 7880 20198
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8128 19446 8156 19654
rect 8116 19440 8168 19446
rect 8116 19382 8168 19388
rect 7840 18692 7892 18698
rect 7840 18634 7892 18640
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 7562 18320 7618 18329
rect 8128 18290 8156 18566
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 7562 18255 7618 18264
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 7472 17740 7524 17746
rect 7472 17682 7524 17688
rect 7564 17740 7616 17746
rect 7564 17682 7616 17688
rect 7484 16794 7512 17682
rect 7576 17542 7604 17682
rect 7564 17536 7616 17542
rect 7564 17478 7616 17484
rect 8312 17320 8340 18362
rect 8220 17292 8340 17320
rect 7472 16788 7524 16794
rect 7472 16730 7524 16736
rect 8220 16538 8248 17292
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8312 16590 8340 17138
rect 8404 16726 8432 20352
rect 8496 19394 8524 22200
rect 8668 20324 8720 20330
rect 8956 20312 8984 22200
rect 9416 20618 9444 22200
rect 9312 20596 9364 20602
rect 9416 20590 9628 20618
rect 9312 20538 9364 20544
rect 9324 20398 9352 20538
rect 9404 20460 9456 20466
rect 9456 20420 9536 20448
rect 9404 20402 9456 20408
rect 9312 20392 9364 20398
rect 9312 20334 9364 20340
rect 8956 20284 9168 20312
rect 8668 20266 8720 20272
rect 8680 19938 8708 20266
rect 8747 20156 9055 20176
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20080 9055 20100
rect 8680 19910 8800 19938
rect 8668 19848 8720 19854
rect 8668 19790 8720 19796
rect 8680 19514 8708 19790
rect 8668 19508 8720 19514
rect 8668 19450 8720 19456
rect 8496 19366 8616 19394
rect 8484 19304 8536 19310
rect 8484 19246 8536 19252
rect 8496 18766 8524 19246
rect 8588 18766 8616 19366
rect 8772 19334 8800 19910
rect 8680 19306 8800 19334
rect 8484 18760 8536 18766
rect 8484 18702 8536 18708
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8484 17604 8536 17610
rect 8484 17546 8536 17552
rect 8392 16720 8444 16726
rect 8392 16662 8444 16668
rect 8496 16658 8524 17546
rect 8588 16794 8616 18702
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8484 16652 8536 16658
rect 8484 16594 8536 16600
rect 8128 16510 8248 16538
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8128 16153 8156 16510
rect 8208 16448 8260 16454
rect 8208 16390 8260 16396
rect 8220 16250 8248 16390
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8300 16176 8352 16182
rect 8114 16144 8170 16153
rect 8300 16118 8352 16124
rect 8114 16079 8170 16088
rect 8208 16108 8260 16114
rect 8208 16050 8260 16056
rect 7840 16040 7892 16046
rect 7654 16008 7710 16017
rect 7840 15982 7892 15988
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 7654 15943 7710 15952
rect 7472 15904 7524 15910
rect 7472 15846 7524 15852
rect 7484 15366 7512 15846
rect 7472 15360 7524 15366
rect 7472 15302 7524 15308
rect 7472 15020 7524 15026
rect 7524 14980 7604 15008
rect 7472 14962 7524 14968
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7484 14618 7512 14758
rect 7576 14618 7604 14980
rect 7472 14612 7524 14618
rect 7472 14554 7524 14560
rect 7564 14612 7616 14618
rect 7564 14554 7616 14560
rect 7472 14272 7524 14278
rect 7472 14214 7524 14220
rect 7564 14272 7616 14278
rect 7564 14214 7616 14220
rect 7484 13920 7512 14214
rect 7576 14074 7604 14214
rect 7668 14074 7696 15943
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7760 15026 7788 15438
rect 7852 15162 7880 15982
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7748 15020 7800 15026
rect 7748 14962 7800 14968
rect 7748 14612 7800 14618
rect 7748 14554 7800 14560
rect 7564 14068 7616 14074
rect 7564 14010 7616 14016
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7484 13892 7696 13920
rect 7472 13796 7524 13802
rect 7472 13738 7524 13744
rect 7564 13796 7616 13802
rect 7564 13738 7616 13744
rect 7484 12850 7512 13738
rect 7576 13433 7604 13738
rect 7562 13424 7618 13433
rect 7562 13359 7618 13368
rect 7576 13258 7604 13359
rect 7564 13252 7616 13258
rect 7564 13194 7616 13200
rect 7472 12844 7524 12850
rect 7472 12786 7524 12792
rect 7380 12436 7432 12442
rect 7380 12378 7432 12384
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 6932 11762 7052 11778
rect 6932 11756 7064 11762
rect 6932 11750 7012 11756
rect 7012 11698 7064 11704
rect 7300 11694 7328 12038
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7392 11558 7420 12378
rect 7576 11898 7604 13194
rect 7668 12442 7696 13892
rect 7760 12986 7788 14554
rect 7944 14550 7972 15982
rect 8220 15502 8248 16050
rect 8312 15570 8340 16118
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8300 15564 8352 15570
rect 8300 15506 8352 15512
rect 8208 15496 8260 15502
rect 8208 15438 8260 15444
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 8036 14618 8064 14894
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 7932 14544 7984 14550
rect 7932 14486 7984 14492
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 8036 14362 8064 14418
rect 8404 14396 8432 15982
rect 8484 15972 8536 15978
rect 8484 15914 8536 15920
rect 8496 15706 8524 15914
rect 8484 15700 8536 15706
rect 8484 15642 8536 15648
rect 8588 15366 8616 16050
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8576 15020 8628 15026
rect 8576 14962 8628 14968
rect 8588 14550 8616 14962
rect 8576 14544 8628 14550
rect 8576 14486 8628 14492
rect 8404 14368 8524 14396
rect 7944 14334 8064 14362
rect 7944 13734 7972 14334
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8208 14272 8260 14278
rect 8208 14214 8260 14220
rect 8392 14272 8444 14278
rect 8392 14214 8444 14220
rect 8128 14074 8156 14214
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 7932 13728 7984 13734
rect 7932 13670 7984 13676
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7852 12986 7880 13126
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7840 12980 7892 12986
rect 7840 12922 7892 12928
rect 7944 12918 7972 13670
rect 8036 13462 8064 13874
rect 8220 13530 8248 14214
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8208 13524 8260 13530
rect 8208 13466 8260 13472
rect 8024 13456 8076 13462
rect 8312 13410 8340 13874
rect 8024 13398 8076 13404
rect 8220 13394 8340 13410
rect 8208 13388 8340 13394
rect 8260 13382 8340 13388
rect 8208 13330 8260 13336
rect 7932 12912 7984 12918
rect 7932 12854 7984 12860
rect 8208 12844 8260 12850
rect 8208 12786 8260 12792
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 7564 11892 7616 11898
rect 7564 11834 7616 11840
rect 7564 11620 7616 11626
rect 7564 11562 7616 11568
rect 7380 11552 7432 11558
rect 7380 11494 7432 11500
rect 6920 11348 6972 11354
rect 6920 11290 6972 11296
rect 6828 11212 6880 11218
rect 6828 11154 6880 11160
rect 6736 11144 6788 11150
rect 6736 11086 6788 11092
rect 6826 11112 6882 11121
rect 6000 11008 6052 11014
rect 5736 10934 5856 10962
rect 6000 10950 6052 10956
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5736 10130 5764 10610
rect 5828 10130 5856 10934
rect 6012 10792 6040 10950
rect 6148 10908 6456 10928
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10832 6456 10852
rect 6012 10764 6408 10792
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5920 10266 5948 10406
rect 5908 10260 5960 10266
rect 5908 10202 5960 10208
rect 5724 10124 5776 10130
rect 5724 10066 5776 10072
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5448 9998 5500 10004
rect 5630 10024 5686 10033
rect 5630 9959 5686 9968
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5460 7546 5488 9522
rect 5552 7818 5580 9862
rect 5644 8634 5672 9862
rect 5736 9042 5764 10066
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5724 9036 5776 9042
rect 5724 8978 5776 8984
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5736 8566 5764 8978
rect 5828 8634 5856 9522
rect 5920 9518 5948 9930
rect 6012 9625 6040 10406
rect 6380 9908 6408 10764
rect 6564 10266 6592 10950
rect 6748 10742 6776 11086
rect 6826 11047 6882 11056
rect 6840 10742 6868 11047
rect 6736 10736 6788 10742
rect 6736 10678 6788 10684
rect 6828 10736 6880 10742
rect 6828 10678 6880 10684
rect 6644 10668 6696 10674
rect 6644 10610 6696 10616
rect 6656 10470 6684 10610
rect 6644 10464 6696 10470
rect 6644 10406 6696 10412
rect 6552 10260 6604 10266
rect 6552 10202 6604 10208
rect 6656 10146 6684 10406
rect 6564 10130 6684 10146
rect 6552 10124 6684 10130
rect 6604 10118 6684 10124
rect 6552 10066 6604 10072
rect 6644 9920 6696 9926
rect 6380 9880 6592 9908
rect 6148 9820 6456 9840
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9744 6456 9764
rect 6564 9674 6592 9880
rect 6644 9862 6696 9868
rect 6104 9646 6592 9674
rect 5998 9616 6054 9625
rect 5998 9551 6054 9560
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 6000 9512 6052 9518
rect 6000 9454 6052 9460
rect 5920 9178 5948 9454
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5736 8090 5764 8502
rect 5920 8362 5948 8842
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5356 7404 5408 7410
rect 5356 7346 5408 7352
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5368 6633 5396 6870
rect 5460 6866 5488 7278
rect 5538 7168 5594 7177
rect 5538 7103 5594 7112
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5354 6624 5410 6633
rect 5354 6559 5410 6568
rect 5460 6390 5488 6802
rect 5552 6662 5580 7103
rect 5644 6798 5672 7890
rect 5724 7336 5776 7342
rect 5724 7278 5776 7284
rect 5736 7002 5764 7278
rect 5724 6996 5776 7002
rect 5724 6938 5776 6944
rect 5632 6792 5684 6798
rect 5632 6734 5684 6740
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 5172 6054 5224 6060
rect 5262 6080 5318 6089
rect 5184 5137 5212 6054
rect 5262 6015 5318 6024
rect 5262 5944 5318 5953
rect 5460 5914 5488 6326
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5262 5879 5318 5888
rect 5448 5908 5500 5914
rect 5276 5574 5304 5879
rect 5448 5850 5500 5856
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5170 5128 5226 5137
rect 5170 5063 5226 5072
rect 5276 4826 5304 5510
rect 5552 5370 5580 6054
rect 5644 5370 5672 6734
rect 5828 6390 5856 8026
rect 5920 7324 5948 8298
rect 6012 7546 6040 9454
rect 6104 9081 6132 9646
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6090 9072 6146 9081
rect 6090 9007 6146 9016
rect 6148 8732 6456 8752
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8656 6456 8676
rect 6564 8022 6592 9318
rect 6656 8974 6684 9862
rect 6748 9654 6776 10678
rect 6932 10588 6960 11290
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 6840 10560 6960 10588
rect 6736 9648 6788 9654
rect 6736 9590 6788 9596
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6748 8838 6776 9318
rect 6736 8832 6788 8838
rect 6736 8774 6788 8780
rect 6644 8560 6696 8566
rect 6644 8502 6696 8508
rect 6552 8016 6604 8022
rect 6552 7958 6604 7964
rect 6552 7744 6604 7750
rect 6550 7712 6552 7721
rect 6604 7712 6606 7721
rect 6148 7644 6456 7664
rect 6550 7647 6606 7656
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7568 6456 7588
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6000 7336 6052 7342
rect 5920 7296 6000 7324
rect 6000 7278 6052 7284
rect 6104 7002 6132 7346
rect 6552 7336 6604 7342
rect 6552 7278 6604 7284
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 6000 6792 6052 6798
rect 6000 6734 6052 6740
rect 5816 6384 5868 6390
rect 5816 6326 5868 6332
rect 5724 5568 5776 5574
rect 5828 5545 5856 6326
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5724 5510 5776 5516
rect 5814 5536 5870 5545
rect 5540 5364 5592 5370
rect 5540 5306 5592 5312
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 5736 5250 5764 5510
rect 5814 5471 5870 5480
rect 5356 5228 5408 5234
rect 5356 5170 5408 5176
rect 5552 5222 5764 5250
rect 5264 4820 5316 4826
rect 5264 4762 5316 4768
rect 5262 4312 5318 4321
rect 5262 4247 5318 4256
rect 5276 4214 5304 4247
rect 5264 4208 5316 4214
rect 5264 4150 5316 4156
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5184 3738 5212 4082
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 5184 3194 5212 3402
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5184 2854 5212 3130
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 5000 2746 5120 2774
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4896 2304 4948 2310
rect 4896 2246 4948 2252
rect 4356 1414 4476 1442
rect 4068 1080 4120 1086
rect 4068 1022 4120 1028
rect 3330 640 3386 649
rect 3330 575 3386 584
rect 3422 0 3478 800
rect 3882 0 3938 800
rect 4080 241 4108 1022
rect 4356 800 4384 1414
rect 4908 800 4936 2246
rect 4066 232 4122 241
rect 4066 167 4122 176
rect 4342 0 4398 800
rect 4894 0 4950 800
rect 5000 762 5028 2746
rect 5276 2650 5304 4014
rect 5368 3194 5396 5170
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5460 4078 5488 4422
rect 5448 4072 5500 4078
rect 5448 4014 5500 4020
rect 5356 3188 5408 3194
rect 5356 3130 5408 3136
rect 5460 3058 5488 4014
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5552 2990 5580 5222
rect 5920 5166 5948 5850
rect 6012 5710 6040 6734
rect 6564 6730 6592 7278
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6148 6556 6456 6576
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6480 6456 6500
rect 6564 6458 6592 6666
rect 6656 6662 6684 8502
rect 6840 7750 6868 10560
rect 7484 10198 7512 10746
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 6920 10124 6972 10130
rect 6920 10066 6972 10072
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 6932 9518 6960 10066
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 7024 9353 7052 9998
rect 7116 9722 7144 10066
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7010 9344 7066 9353
rect 7010 9279 7066 9288
rect 7472 8832 7524 8838
rect 7472 8774 7524 8780
rect 7484 8498 7512 8774
rect 7576 8634 7604 11562
rect 8128 11354 8156 12038
rect 8220 11778 8248 12786
rect 8404 12374 8432 14214
rect 8496 12850 8524 14368
rect 8680 14278 8708 19306
rect 8747 19068 9055 19088
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 18992 9055 19012
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8956 18290 8984 18566
rect 9140 18290 9168 20284
rect 9312 20256 9364 20262
rect 9312 20198 9364 20204
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9220 19780 9272 19786
rect 9220 19722 9272 19728
rect 8944 18284 8996 18290
rect 8944 18226 8996 18232
rect 9128 18284 9180 18290
rect 9128 18226 9180 18232
rect 8747 17980 9055 18000
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17904 9055 17924
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 9048 17202 9076 17682
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 8747 16892 9055 16912
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16816 9055 16836
rect 9140 16794 9168 18226
rect 9232 18154 9260 19722
rect 9324 19446 9352 20198
rect 9312 19440 9364 19446
rect 9312 19382 9364 19388
rect 9416 18834 9444 20198
rect 9508 19718 9536 20420
rect 9600 20312 9628 20590
rect 9680 20324 9732 20330
rect 9600 20284 9680 20312
rect 9680 20266 9732 20272
rect 9586 19952 9642 19961
rect 9586 19887 9642 19896
rect 9496 19712 9548 19718
rect 9496 19654 9548 19660
rect 9508 18834 9536 19654
rect 9600 19496 9628 19887
rect 9876 19786 9904 22200
rect 10232 20800 10284 20806
rect 10232 20742 10284 20748
rect 10244 20602 10272 20742
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10140 20460 10192 20466
rect 10140 20402 10192 20408
rect 10048 20392 10100 20398
rect 10048 20334 10100 20340
rect 10060 20262 10088 20334
rect 10048 20256 10100 20262
rect 10048 20198 10100 20204
rect 10152 20058 10180 20402
rect 10140 20052 10192 20058
rect 10140 19994 10192 20000
rect 9864 19780 9916 19786
rect 9864 19722 9916 19728
rect 10140 19712 10192 19718
rect 10140 19654 10192 19660
rect 9864 19508 9916 19514
rect 9600 19468 9720 19496
rect 9586 19408 9642 19417
rect 9586 19343 9642 19352
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9496 18828 9548 18834
rect 9496 18770 9548 18776
rect 9404 18692 9456 18698
rect 9404 18634 9456 18640
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9324 18426 9352 18566
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9220 18148 9272 18154
rect 9220 18090 9272 18096
rect 9416 17626 9444 18634
rect 9494 18592 9550 18601
rect 9494 18527 9550 18536
rect 9508 18057 9536 18527
rect 9600 18426 9628 19343
rect 9692 18426 9720 19468
rect 9864 19450 9916 19456
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9494 18048 9550 18057
rect 9494 17983 9550 17992
rect 9680 17740 9732 17746
rect 9680 17682 9732 17688
rect 9232 17598 9444 17626
rect 9128 16788 9180 16794
rect 9128 16730 9180 16736
rect 8758 16688 8814 16697
rect 8758 16623 8760 16632
rect 8812 16623 8814 16632
rect 8760 16594 8812 16600
rect 9126 16008 9182 16017
rect 9126 15943 9182 15952
rect 8747 15804 9055 15824
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15728 9055 15748
rect 9034 15464 9090 15473
rect 9034 15399 9090 15408
rect 8758 15056 8814 15065
rect 9048 15026 9076 15399
rect 9140 15162 9168 15943
rect 9128 15156 9180 15162
rect 9128 15098 9180 15104
rect 8758 14991 8814 15000
rect 9036 15020 9088 15026
rect 8772 14958 8800 14991
rect 9036 14962 9088 14968
rect 8760 14952 8812 14958
rect 8760 14894 8812 14900
rect 8747 14716 9055 14736
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14640 9055 14660
rect 9140 14618 9168 15098
rect 9128 14612 9180 14618
rect 9128 14554 9180 14560
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8747 13628 9055 13648
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13552 9055 13572
rect 9140 13530 9168 14554
rect 9128 13524 9180 13530
rect 9128 13466 9180 13472
rect 8576 13456 8628 13462
rect 8576 13398 8628 13404
rect 8484 12844 8536 12850
rect 8484 12786 8536 12792
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8392 12164 8444 12170
rect 8392 12106 8444 12112
rect 8220 11750 8340 11778
rect 8208 11688 8260 11694
rect 8208 11630 8260 11636
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7852 10810 7880 11018
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7852 10606 7880 10746
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7852 9178 7880 9862
rect 8128 9738 8156 10950
rect 8220 10538 8248 11630
rect 8208 10532 8260 10538
rect 8208 10474 8260 10480
rect 8128 9710 8248 9738
rect 8220 9586 8248 9710
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 8036 8634 8064 9522
rect 8312 9194 8340 11750
rect 8404 10810 8432 12106
rect 8496 11354 8524 12242
rect 8588 11898 8616 13398
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 9036 13388 9088 13394
rect 9036 13330 9088 13336
rect 8680 12918 8708 13330
rect 8668 12912 8720 12918
rect 8668 12854 8720 12860
rect 8668 12640 8720 12646
rect 9048 12628 9076 13330
rect 9140 13190 9168 13466
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 9232 12714 9260 17598
rect 9404 17536 9456 17542
rect 9404 17478 9456 17484
rect 9310 17232 9366 17241
rect 9310 17167 9366 17176
rect 9324 15162 9352 17167
rect 9416 16182 9444 17478
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9508 16250 9536 16390
rect 9496 16244 9548 16250
rect 9496 16186 9548 16192
rect 9404 16176 9456 16182
rect 9404 16118 9456 16124
rect 9312 15156 9364 15162
rect 9312 15098 9364 15104
rect 9588 15156 9640 15162
rect 9588 15098 9640 15104
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 9312 14000 9364 14006
rect 9364 13960 9444 13988
rect 9312 13942 9364 13948
rect 9312 13864 9364 13870
rect 9312 13806 9364 13812
rect 9324 12850 9352 13806
rect 9416 13394 9444 13960
rect 9508 13938 9536 14962
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9508 13462 9536 13874
rect 9496 13456 9548 13462
rect 9496 13398 9548 13404
rect 9404 13388 9456 13394
rect 9404 13330 9456 13336
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9312 12844 9364 12850
rect 9312 12786 9364 12792
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9048 12600 9168 12628
rect 8668 12582 8720 12588
rect 8680 12238 8708 12582
rect 8747 12540 9055 12560
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12464 9055 12484
rect 8760 12368 8812 12374
rect 8760 12310 8812 12316
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8680 11762 8708 12174
rect 8668 11756 8720 11762
rect 8668 11698 8720 11704
rect 8772 11642 8800 12310
rect 9048 11898 9076 12310
rect 9140 11898 9168 12600
rect 9036 11892 9088 11898
rect 9036 11834 9088 11840
rect 9128 11892 9180 11898
rect 9128 11834 9180 11840
rect 9048 11694 9076 11834
rect 8588 11614 8800 11642
rect 9036 11688 9088 11694
rect 9036 11630 9088 11636
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8392 10804 8444 10810
rect 8392 10746 8444 10752
rect 8496 10062 8524 11290
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8220 9166 8340 9194
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 8024 8628 8076 8634
rect 8024 8570 8076 8576
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7116 8090 7144 8434
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7564 7880 7616 7886
rect 7564 7822 7616 7828
rect 7012 7812 7064 7818
rect 7012 7754 7064 7760
rect 6828 7744 6880 7750
rect 6828 7686 6880 7692
rect 6734 7576 6790 7585
rect 6734 7511 6790 7520
rect 6748 7313 6776 7511
rect 6920 7472 6972 7478
rect 6920 7414 6972 7420
rect 6734 7304 6790 7313
rect 6734 7239 6790 7248
rect 6826 7168 6882 7177
rect 6826 7103 6882 7112
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6734 6624 6790 6633
rect 6734 6559 6790 6568
rect 6552 6452 6604 6458
rect 6552 6394 6604 6400
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6000 5704 6052 5710
rect 6000 5646 6052 5652
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5816 4820 5868 4826
rect 5816 4762 5868 4768
rect 5724 4480 5776 4486
rect 5724 4422 5776 4428
rect 5630 3768 5686 3777
rect 5630 3703 5686 3712
rect 5644 3466 5672 3703
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5630 3224 5686 3233
rect 5630 3159 5686 3168
rect 5644 3058 5672 3159
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5540 2984 5592 2990
rect 5540 2926 5592 2932
rect 5448 2916 5500 2922
rect 5448 2858 5500 2864
rect 5460 2650 5488 2858
rect 5538 2680 5594 2689
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5448 2644 5500 2650
rect 5538 2615 5594 2624
rect 5448 2586 5500 2592
rect 5552 2514 5580 2615
rect 5540 2508 5592 2514
rect 5540 2450 5592 2456
rect 5736 2378 5764 4422
rect 5828 4185 5856 4762
rect 6012 4604 6040 5646
rect 6148 5468 6456 5488
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5392 6456 5412
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6472 5137 6500 5170
rect 6458 5128 6514 5137
rect 6458 5063 6514 5072
rect 6274 4856 6330 4865
rect 6274 4791 6330 4800
rect 6288 4622 6316 4791
rect 6564 4758 6592 6054
rect 6552 4752 6604 4758
rect 6552 4694 6604 4700
rect 6092 4616 6144 4622
rect 6012 4576 6092 4604
rect 5814 4176 5870 4185
rect 5814 4111 5870 4120
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5906 3904 5962 3913
rect 5724 2372 5776 2378
rect 5724 2314 5776 2320
rect 5828 1737 5856 3878
rect 5906 3839 5962 3848
rect 5920 3194 5948 3839
rect 6012 3466 6040 4576
rect 6092 4558 6144 4564
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6552 4480 6604 4486
rect 6550 4448 6552 4457
rect 6604 4448 6606 4457
rect 6148 4380 6456 4400
rect 6550 4383 6606 4392
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4304 6456 4324
rect 6550 4176 6606 4185
rect 6656 4146 6684 6054
rect 6748 5953 6776 6559
rect 6734 5944 6790 5953
rect 6734 5879 6790 5888
rect 6840 5642 6868 7103
rect 6932 6186 6960 7414
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6828 5636 6880 5642
rect 6828 5578 6880 5584
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6748 5030 6776 5170
rect 6932 5166 6960 5850
rect 7024 5710 7052 7754
rect 7288 7336 7340 7342
rect 7288 7278 7340 7284
rect 7104 7200 7156 7206
rect 7104 7142 7156 7148
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 7116 6458 7144 7142
rect 7208 7002 7236 7142
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7300 6798 7328 7278
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7194 6488 7250 6497
rect 7104 6452 7156 6458
rect 7194 6423 7250 6432
rect 7104 6394 7156 6400
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6840 4826 6868 5034
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6736 4752 6788 4758
rect 6736 4694 6788 4700
rect 6550 4111 6606 4120
rect 6644 4140 6696 4146
rect 6366 3904 6422 3913
rect 6366 3839 6422 3848
rect 6380 3738 6408 3839
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6564 3482 6592 4111
rect 6644 4082 6696 4088
rect 6644 4004 6696 4010
rect 6644 3946 6696 3952
rect 6288 3466 6592 3482
rect 6000 3460 6052 3466
rect 6000 3402 6052 3408
rect 6276 3460 6592 3466
rect 6328 3454 6592 3460
rect 6276 3402 6328 3408
rect 6148 3292 6456 3312
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 5998 3224 6054 3233
rect 5908 3188 5960 3194
rect 6148 3216 6456 3236
rect 6564 3210 6592 3454
rect 6656 3398 6684 3946
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6748 3346 6776 4694
rect 6920 4684 6972 4690
rect 6920 4626 6972 4632
rect 6932 4078 6960 4626
rect 7024 4214 7052 5306
rect 7116 4282 7144 6054
rect 7208 5370 7236 6423
rect 7300 5914 7328 6734
rect 7392 6254 7420 6938
rect 7472 6860 7524 6866
rect 7472 6802 7524 6808
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7288 5908 7340 5914
rect 7288 5850 7340 5856
rect 7484 5846 7512 6802
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7196 5364 7248 5370
rect 7196 5306 7248 5312
rect 7288 5296 7340 5302
rect 7288 5238 7340 5244
rect 7300 5137 7328 5238
rect 7286 5128 7342 5137
rect 7286 5063 7342 5072
rect 7194 4584 7250 4593
rect 7194 4519 7250 4528
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 7012 4208 7064 4214
rect 7012 4150 7064 4156
rect 6920 4072 6972 4078
rect 7208 4026 7236 4519
rect 6920 4014 6972 4020
rect 6932 3777 6960 4014
rect 7024 3998 7236 4026
rect 6918 3768 6974 3777
rect 6918 3703 6974 3712
rect 6920 3392 6972 3398
rect 6748 3340 6920 3346
rect 6748 3334 6972 3340
rect 6748 3318 6960 3334
rect 6826 3224 6882 3233
rect 6564 3182 6684 3210
rect 5998 3159 6054 3168
rect 5908 3130 5960 3136
rect 5920 3097 5948 3130
rect 6012 3126 6040 3159
rect 6000 3120 6052 3126
rect 5906 3088 5962 3097
rect 6000 3062 6052 3068
rect 5906 3023 5962 3032
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 6552 3052 6604 3058
rect 6552 2994 6604 3000
rect 6104 2961 6132 2994
rect 6184 2984 6236 2990
rect 6090 2952 6146 2961
rect 6184 2926 6236 2932
rect 6090 2887 6146 2896
rect 6196 2774 6224 2926
rect 6104 2746 6224 2774
rect 6104 2378 6132 2746
rect 6458 2680 6514 2689
rect 6184 2644 6236 2650
rect 6564 2650 6592 2994
rect 6458 2615 6460 2624
rect 6184 2586 6236 2592
rect 6512 2615 6514 2624
rect 6552 2644 6604 2650
rect 6460 2586 6512 2592
rect 6552 2586 6604 2592
rect 6196 2378 6224 2586
rect 6092 2372 6144 2378
rect 6012 2332 6092 2360
rect 5908 1828 5960 1834
rect 5908 1770 5960 1776
rect 5814 1728 5870 1737
rect 5814 1663 5870 1672
rect 5920 1578 5948 1770
rect 5828 1550 5948 1578
rect 5276 870 5396 898
rect 5276 762 5304 870
rect 5368 800 5396 870
rect 5828 800 5856 1550
rect 5000 734 5304 762
rect 5354 0 5410 800
rect 5814 0 5870 800
rect 6012 762 6040 2332
rect 6092 2314 6144 2320
rect 6184 2372 6236 2378
rect 6184 2314 6236 2320
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 6148 2204 6456 2224
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2128 6456 2148
rect 6564 1698 6592 2314
rect 6656 2106 6684 3182
rect 6826 3159 6828 3168
rect 6880 3159 6882 3168
rect 6828 3130 6880 3136
rect 7024 3126 7052 3998
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 7024 2774 7052 3062
rect 6932 2746 7052 2774
rect 7116 2774 7144 3878
rect 7300 3126 7328 5063
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7392 3942 7420 4626
rect 7484 4282 7512 4966
rect 7472 4276 7524 4282
rect 7472 4218 7524 4224
rect 7470 4040 7526 4049
rect 7470 3975 7526 3984
rect 7380 3936 7432 3942
rect 7380 3878 7432 3884
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7288 3120 7340 3126
rect 7288 3062 7340 3068
rect 7116 2746 7236 2774
rect 6736 2644 6788 2650
rect 6736 2586 6788 2592
rect 6748 2530 6776 2586
rect 6748 2502 6868 2530
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 6748 2106 6776 2382
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6736 2100 6788 2106
rect 6736 2042 6788 2048
rect 6840 1834 6868 2502
rect 6828 1828 6880 1834
rect 6828 1770 6880 1776
rect 6552 1692 6604 1698
rect 6552 1634 6604 1640
rect 6736 1692 6788 1698
rect 6736 1634 6788 1640
rect 6196 870 6316 898
rect 6196 762 6224 870
rect 6288 800 6316 870
rect 6748 800 6776 1634
rect 6932 1086 6960 2746
rect 7208 2650 7236 2746
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7012 2576 7064 2582
rect 7300 2530 7328 2586
rect 7064 2524 7328 2530
rect 7012 2518 7328 2524
rect 7024 2502 7328 2518
rect 7392 2446 7420 3334
rect 7104 2440 7156 2446
rect 7104 2382 7156 2388
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7116 2258 7144 2382
rect 7484 2258 7512 3975
rect 7576 2650 7604 7822
rect 7748 6860 7800 6866
rect 7748 6802 7800 6808
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7668 6458 7696 6598
rect 7656 6452 7708 6458
rect 7656 6394 7708 6400
rect 7760 6322 7788 6802
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7760 5574 7788 6258
rect 7748 5568 7800 5574
rect 7748 5510 7800 5516
rect 7656 5228 7708 5234
rect 7656 5170 7708 5176
rect 7668 4826 7696 5170
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7852 4690 7880 8570
rect 7932 7880 7984 7886
rect 7932 7822 7984 7828
rect 7944 7002 7972 7822
rect 8220 7546 8248 9166
rect 8300 9104 8352 9110
rect 8300 9046 8352 9052
rect 8312 8634 8340 9046
rect 8300 8628 8352 8634
rect 8300 8570 8352 8576
rect 8208 7540 8260 7546
rect 8208 7482 8260 7488
rect 8404 7392 8432 9930
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8496 8838 8524 9590
rect 8588 9178 8616 11614
rect 8668 11552 8720 11558
rect 8668 11494 8720 11500
rect 8680 10810 8708 11494
rect 8747 11452 9055 11472
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11376 9055 11396
rect 9140 10810 9168 11834
rect 9218 11792 9274 11801
rect 9218 11727 9274 11736
rect 8668 10804 8720 10810
rect 8668 10746 8720 10752
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 8747 10364 9055 10384
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10288 9055 10308
rect 9126 10160 9182 10169
rect 9126 10095 9182 10104
rect 9140 9722 9168 10095
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 8747 9276 9055 9296
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9200 9055 9220
rect 8576 9172 8628 9178
rect 8576 9114 8628 9120
rect 8588 8974 8616 9114
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 9140 8906 9168 9318
rect 8760 8900 8812 8906
rect 8760 8842 8812 8848
rect 9128 8900 9180 8906
rect 9128 8842 9180 8848
rect 8484 8832 8536 8838
rect 8482 8800 8484 8809
rect 8536 8800 8538 8809
rect 8482 8735 8538 8744
rect 8772 8430 8800 8842
rect 9232 8673 9260 11727
rect 9312 10464 9364 10470
rect 9312 10406 9364 10412
rect 9218 8664 9274 8673
rect 9324 8634 9352 10406
rect 9416 9761 9444 13126
rect 9496 12844 9548 12850
rect 9496 12786 9548 12792
rect 9508 12442 9536 12786
rect 9496 12436 9548 12442
rect 9600 12434 9628 15098
rect 9692 14822 9720 17682
rect 9784 17066 9812 18226
rect 9772 17060 9824 17066
rect 9772 17002 9824 17008
rect 9784 16046 9812 17002
rect 9772 16040 9824 16046
rect 9772 15982 9824 15988
rect 9680 14816 9732 14822
rect 9680 14758 9732 14764
rect 9876 14618 9904 19450
rect 10048 19440 10100 19446
rect 10048 19382 10100 19388
rect 9954 19000 10010 19009
rect 9954 18935 10010 18944
rect 9968 18630 9996 18935
rect 9956 18624 10008 18630
rect 9956 18566 10008 18572
rect 9968 18465 9996 18566
rect 9954 18456 10010 18465
rect 9954 18391 10010 18400
rect 10060 17814 10088 19382
rect 10048 17808 10100 17814
rect 10048 17750 10100 17756
rect 10046 17640 10102 17649
rect 10046 17575 10102 17584
rect 10060 17542 10088 17575
rect 10048 17536 10100 17542
rect 10048 17478 10100 17484
rect 10152 17082 10180 19654
rect 10336 19446 10364 22200
rect 10416 20392 10468 20398
rect 10600 20392 10652 20398
rect 10416 20334 10468 20340
rect 10520 20352 10600 20380
rect 10428 19990 10456 20334
rect 10416 19984 10468 19990
rect 10416 19926 10468 19932
rect 10520 19514 10548 20352
rect 10600 20334 10652 20340
rect 10796 20210 10824 22200
rect 11256 20806 11284 22200
rect 11244 20800 11296 20806
rect 11244 20742 11296 20748
rect 11256 20534 11284 20742
rect 11346 20700 11654 20720
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20624 11654 20644
rect 11244 20528 11296 20534
rect 11244 20470 11296 20476
rect 11152 20392 11204 20398
rect 11152 20334 11204 20340
rect 10876 20324 10928 20330
rect 10876 20266 10928 20272
rect 11060 20324 11112 20330
rect 11060 20266 11112 20272
rect 10612 20182 10824 20210
rect 10508 19508 10560 19514
rect 10508 19450 10560 19456
rect 10324 19440 10376 19446
rect 10376 19400 10456 19428
rect 10324 19382 10376 19388
rect 10428 19310 10456 19400
rect 10508 19372 10560 19378
rect 10508 19314 10560 19320
rect 10324 19304 10376 19310
rect 10324 19246 10376 19252
rect 10416 19304 10468 19310
rect 10416 19246 10468 19252
rect 10336 18970 10364 19246
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 10244 18873 10272 18906
rect 10230 18864 10286 18873
rect 10230 18799 10286 18808
rect 10232 17672 10284 17678
rect 10232 17614 10284 17620
rect 10060 17054 10180 17082
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9968 15978 9996 16390
rect 10060 16250 10088 17054
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10152 16658 10180 16934
rect 10140 16652 10192 16658
rect 10140 16594 10192 16600
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 10152 16250 10180 16458
rect 10048 16244 10100 16250
rect 10048 16186 10100 16192
rect 10140 16244 10192 16250
rect 10140 16186 10192 16192
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 10152 15026 10180 15982
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 9864 14612 9916 14618
rect 9864 14554 9916 14560
rect 9876 14521 9904 14554
rect 10048 14544 10100 14550
rect 9862 14512 9918 14521
rect 10048 14486 10100 14492
rect 9862 14447 9918 14456
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9692 13977 9720 14282
rect 9678 13968 9734 13977
rect 9678 13903 9734 13912
rect 9692 13546 9720 13903
rect 9784 13734 9812 14350
rect 9864 14272 9916 14278
rect 9864 14214 9916 14220
rect 9876 14006 9904 14214
rect 9864 14000 9916 14006
rect 9864 13942 9916 13948
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9876 13546 9904 13806
rect 9692 13530 9904 13546
rect 9680 13524 9904 13530
rect 9732 13518 9904 13524
rect 9680 13466 9732 13472
rect 9864 13184 9916 13190
rect 9864 13126 9916 13132
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9876 12442 9904 13126
rect 9864 12436 9916 12442
rect 9600 12406 9720 12434
rect 9496 12378 9548 12384
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9508 11898 9536 12106
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9494 11248 9550 11257
rect 9494 11183 9550 11192
rect 9508 9874 9536 11183
rect 9692 11150 9720 12406
rect 9864 12378 9916 12384
rect 9968 11354 9996 13126
rect 10060 12102 10088 14486
rect 10152 14482 10180 14962
rect 10244 14929 10272 17614
rect 10336 17270 10364 18906
rect 10520 18902 10548 19314
rect 10508 18896 10560 18902
rect 10508 18838 10560 18844
rect 10612 18222 10640 20182
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10704 19258 10732 19994
rect 10704 19230 10824 19258
rect 10888 19242 10916 20266
rect 11072 19922 11100 20266
rect 11164 20058 11192 20334
rect 11716 20058 11744 22200
rect 12176 20448 12204 22200
rect 12440 20460 12492 20466
rect 12176 20420 12440 20448
rect 12440 20402 12492 20408
rect 12440 20324 12492 20330
rect 12440 20266 12492 20272
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11704 20052 11756 20058
rect 11704 19994 11756 20000
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 10968 19780 11020 19786
rect 10968 19722 11020 19728
rect 10692 19168 10744 19174
rect 10692 19110 10744 19116
rect 10704 18290 10732 19110
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10600 18216 10652 18222
rect 10600 18158 10652 18164
rect 10416 18080 10468 18086
rect 10416 18022 10468 18028
rect 10508 18080 10560 18086
rect 10508 18022 10560 18028
rect 10324 17264 10376 17270
rect 10324 17206 10376 17212
rect 10428 17202 10456 18022
rect 10520 17785 10548 18022
rect 10796 17882 10824 19230
rect 10876 19236 10928 19242
rect 10876 19178 10928 19184
rect 10980 18086 11008 19722
rect 11346 19612 11654 19632
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19536 11654 19556
rect 11060 19304 11112 19310
rect 11060 19246 11112 19252
rect 11072 18222 11100 19246
rect 11704 19168 11756 19174
rect 11704 19110 11756 19116
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11164 18426 11192 18566
rect 11152 18420 11204 18426
rect 11152 18362 11204 18368
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10784 17876 10836 17882
rect 10784 17818 10836 17824
rect 10506 17776 10562 17785
rect 10796 17746 10824 17818
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 10506 17711 10562 17720
rect 10784 17740 10836 17746
rect 10784 17682 10836 17688
rect 10784 17536 10836 17542
rect 10784 17478 10836 17484
rect 10796 17338 10824 17478
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10324 16176 10376 16182
rect 10324 16118 10376 16124
rect 10230 14920 10286 14929
rect 10230 14855 10286 14864
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 10232 13932 10284 13938
rect 10232 13874 10284 13880
rect 10048 12096 10100 12102
rect 10048 12038 10100 12044
rect 9956 11348 10008 11354
rect 9956 11290 10008 11296
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9600 10266 9628 11018
rect 9692 10674 9720 11086
rect 10060 11082 10088 12038
rect 10244 11830 10272 13874
rect 10232 11824 10284 11830
rect 10232 11766 10284 11772
rect 10336 11098 10364 16118
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 10428 13326 10456 15370
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10612 14006 10640 14758
rect 10796 14618 10824 16390
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10704 14074 10732 14214
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10600 14000 10652 14006
rect 10600 13942 10652 13948
rect 10508 13388 10560 13394
rect 10508 13330 10560 13336
rect 10416 13320 10468 13326
rect 10416 13262 10468 13268
rect 10428 11898 10456 13262
rect 10520 12442 10548 13330
rect 10600 12640 10652 12646
rect 10600 12582 10652 12588
rect 10508 12436 10560 12442
rect 10508 12378 10560 12384
rect 10612 12306 10640 12582
rect 10784 12368 10836 12374
rect 10782 12336 10784 12345
rect 10836 12336 10838 12345
rect 10600 12300 10652 12306
rect 10782 12271 10838 12280
rect 10600 12242 10652 12248
rect 10612 12170 10640 12242
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10416 11892 10468 11898
rect 10416 11834 10468 11840
rect 10048 11076 10100 11082
rect 10048 11018 10100 11024
rect 10244 11070 10364 11098
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9956 10600 10008 10606
rect 9956 10542 10008 10548
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9680 9920 9732 9926
rect 9508 9846 9628 9874
rect 9680 9862 9732 9868
rect 9402 9752 9458 9761
rect 9402 9687 9458 9696
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 9402 8664 9458 8673
rect 9218 8599 9274 8608
rect 9312 8628 9364 8634
rect 9402 8599 9458 8608
rect 9312 8570 9364 8576
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8747 8188 9055 8208
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8112 9055 8132
rect 9140 8090 9168 8434
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 8668 8016 8720 8022
rect 8668 7958 8720 7964
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8036 7364 8432 7392
rect 7932 6996 7984 7002
rect 7932 6938 7984 6944
rect 7932 6724 7984 6730
rect 7932 6666 7984 6672
rect 7944 6497 7972 6666
rect 7930 6488 7986 6497
rect 7930 6423 7986 6432
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 7944 5370 7972 6054
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7840 4684 7892 4690
rect 7840 4626 7892 4632
rect 8036 4622 8064 7364
rect 8298 7304 8354 7313
rect 8298 7239 8354 7248
rect 8206 7032 8262 7041
rect 8206 6967 8262 6976
rect 8220 6730 8248 6967
rect 8208 6724 8260 6730
rect 8208 6666 8260 6672
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8128 5370 8156 6598
rect 8220 6322 8248 6666
rect 8312 6361 8340 7239
rect 8390 7168 8446 7177
rect 8390 7103 8446 7112
rect 8404 6798 8432 7103
rect 8496 6934 8524 7482
rect 8588 7478 8616 7686
rect 8576 7472 8628 7478
rect 8576 7414 8628 7420
rect 8484 6928 8536 6934
rect 8536 6888 8616 6916
rect 8484 6870 8536 6876
rect 8392 6792 8444 6798
rect 8392 6734 8444 6740
rect 8588 6458 8616 6888
rect 8680 6848 8708 7958
rect 9128 7948 9180 7954
rect 9128 7890 9180 7896
rect 9140 7750 9168 7890
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 7177 9168 7686
rect 9232 7478 9260 8502
rect 9310 8120 9366 8129
rect 9310 8055 9366 8064
rect 9220 7472 9272 7478
rect 9324 7449 9352 8055
rect 9416 7954 9444 8599
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9508 7546 9536 9658
rect 9600 7834 9628 9846
rect 9692 9654 9720 9862
rect 9968 9654 9996 10542
rect 10244 9926 10272 11070
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10336 10606 10364 10950
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9968 7954 9996 9590
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10048 9444 10100 9450
rect 10048 9386 10100 9392
rect 9956 7948 10008 7954
rect 9956 7890 10008 7896
rect 9600 7806 9720 7834
rect 9588 7744 9640 7750
rect 9588 7686 9640 7692
rect 9496 7540 9548 7546
rect 9496 7482 9548 7488
rect 9220 7414 9272 7420
rect 9310 7440 9366 7449
rect 9310 7375 9366 7384
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9220 7200 9272 7206
rect 9126 7168 9182 7177
rect 8747 7100 9055 7120
rect 9220 7142 9272 7148
rect 9126 7103 9182 7112
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7024 9055 7044
rect 9126 7032 9182 7041
rect 9126 6967 9128 6976
rect 9180 6967 9182 6976
rect 9128 6938 9180 6944
rect 8944 6928 8996 6934
rect 8944 6870 8996 6876
rect 8760 6860 8812 6866
rect 8680 6820 8760 6848
rect 8760 6802 8812 6808
rect 8668 6724 8720 6730
rect 8668 6666 8720 6672
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8298 6352 8354 6361
rect 8208 6316 8260 6322
rect 8680 6338 8708 6666
rect 8850 6488 8906 6497
rect 8760 6452 8812 6458
rect 8850 6423 8906 6432
rect 8760 6394 8812 6400
rect 8298 6287 8354 6296
rect 8404 6310 8708 6338
rect 8208 6258 8260 6264
rect 8300 6248 8352 6254
rect 8404 6236 8432 6310
rect 8352 6208 8432 6236
rect 8576 6248 8628 6254
rect 8300 6190 8352 6196
rect 8576 6190 8628 6196
rect 8484 6180 8536 6186
rect 8484 6122 8536 6128
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8220 4826 8248 5578
rect 8312 5302 8340 6054
rect 8496 5574 8524 6122
rect 8484 5568 8536 5574
rect 8484 5510 8536 5516
rect 8588 5370 8616 6190
rect 8772 6100 8800 6394
rect 8864 6186 8892 6423
rect 8956 6361 8984 6870
rect 8942 6352 8998 6361
rect 8942 6287 8998 6296
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 8852 6180 8904 6186
rect 8852 6122 8904 6128
rect 8680 6072 8800 6100
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8300 5296 8352 5302
rect 8300 5238 8352 5244
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8300 5160 8352 5166
rect 8298 5128 8300 5137
rect 8352 5128 8354 5137
rect 8298 5063 8354 5072
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8208 4820 8260 4826
rect 8208 4762 8260 4768
rect 8116 4752 8168 4758
rect 8116 4694 8168 4700
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7748 4480 7800 4486
rect 7748 4422 7800 4428
rect 7840 4480 7892 4486
rect 7840 4422 7892 4428
rect 7760 4282 7788 4422
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7668 3738 7696 4014
rect 7656 3732 7708 3738
rect 7656 3674 7708 3680
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 2922 7696 3470
rect 7760 3194 7788 4218
rect 7852 3505 7880 4422
rect 8024 3936 8076 3942
rect 8024 3878 8076 3884
rect 7838 3496 7894 3505
rect 7838 3431 7894 3440
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 7656 2916 7708 2922
rect 7656 2858 7708 2864
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 7760 2446 7788 2790
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 7116 2230 7512 2258
rect 6920 1080 6972 1086
rect 6920 1022 6972 1028
rect 7208 800 7236 2230
rect 7668 1902 7696 2314
rect 7852 2038 7880 3431
rect 8036 3126 8064 3878
rect 8128 3754 8156 4694
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 8220 4010 8248 4490
rect 8312 4486 8340 4966
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8312 4146 8340 4422
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8128 3726 8248 3754
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7944 2650 7972 2994
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 7840 2032 7892 2038
rect 7840 1974 7892 1980
rect 7656 1896 7708 1902
rect 7656 1838 7708 1844
rect 7668 800 7696 1838
rect 8128 800 8156 2382
rect 8220 1902 8248 3726
rect 8312 3194 8340 3878
rect 8404 3738 8432 4558
rect 8496 4434 8524 5170
rect 8588 4690 8616 5306
rect 8680 5302 8708 6072
rect 8747 6012 9055 6032
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5936 9055 5956
rect 8944 5840 8996 5846
rect 8944 5782 8996 5788
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8772 5574 8800 5646
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 8956 5012 8984 5782
rect 9140 5574 9168 6258
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 8680 4984 8984 5012
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8496 4406 8616 4434
rect 8482 4312 8538 4321
rect 8482 4247 8538 4256
rect 8496 4146 8524 4247
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8484 4004 8536 4010
rect 8484 3946 8536 3952
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8496 3534 8524 3946
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8392 3392 8444 3398
rect 8392 3334 8444 3340
rect 8482 3360 8538 3369
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8404 2990 8432 3334
rect 8482 3295 8538 3304
rect 8392 2984 8444 2990
rect 8392 2926 8444 2932
rect 8404 2774 8432 2926
rect 8312 2746 8432 2774
rect 8312 2582 8340 2746
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8496 2514 8524 3295
rect 8588 2514 8616 4406
rect 8484 2508 8536 2514
rect 8484 2450 8536 2456
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8680 2378 8708 4984
rect 8747 4924 9055 4944
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4848 9055 4868
rect 9140 4690 9168 5510
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9232 4554 9260 7142
rect 9508 6730 9536 7278
rect 9600 6798 9628 7686
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9496 6724 9548 6730
rect 9496 6666 9548 6672
rect 9312 6656 9364 6662
rect 9692 6610 9720 7806
rect 9770 7712 9826 7721
rect 9770 7647 9826 7656
rect 9312 6598 9364 6604
rect 9324 6497 9352 6598
rect 9508 6582 9720 6610
rect 9310 6488 9366 6497
rect 9310 6423 9366 6432
rect 9508 6372 9536 6582
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9324 6344 9536 6372
rect 9324 5778 9352 6344
rect 9404 6248 9456 6254
rect 9404 6190 9456 6196
rect 9312 5772 9364 5778
rect 9312 5714 9364 5720
rect 9416 5234 9444 6190
rect 9404 5228 9456 5234
rect 9404 5170 9456 5176
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 9220 4548 9272 4554
rect 9496 4548 9548 4554
rect 9220 4490 9272 4496
rect 9416 4508 9496 4536
rect 8772 4078 8800 4490
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 9220 4072 9272 4078
rect 9220 4014 9272 4020
rect 9128 4004 9180 4010
rect 9128 3946 9180 3952
rect 8747 3836 9055 3856
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3760 9055 3780
rect 9140 3738 9168 3946
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9140 3618 9168 3674
rect 8956 3590 9168 3618
rect 8956 2990 8984 3590
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 9048 2938 9076 3470
rect 9232 3194 9260 4014
rect 9324 3194 9352 4082
rect 9416 4078 9444 4508
rect 9496 4490 9548 4496
rect 9600 4434 9628 6394
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9692 5710 9720 6258
rect 9680 5704 9732 5710
rect 9680 5646 9732 5652
rect 9784 5370 9812 7647
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9876 7410 9904 7482
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9968 7274 9996 7890
rect 10060 7546 10088 9386
rect 10140 9376 10192 9382
rect 10140 9318 10192 9324
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10152 8634 10180 9318
rect 10244 8906 10272 9318
rect 10232 8900 10284 8906
rect 10232 8842 10284 8848
rect 10336 8634 10364 9454
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10428 7886 10456 11834
rect 10612 11694 10640 12106
rect 10600 11688 10652 11694
rect 10600 11630 10652 11636
rect 10612 11218 10640 11630
rect 10600 11212 10652 11218
rect 10600 11154 10652 11160
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10508 10192 10560 10198
rect 10508 10134 10560 10140
rect 10520 9722 10548 10134
rect 10612 10130 10640 10950
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10600 10124 10652 10130
rect 10600 10066 10652 10072
rect 10704 9926 10732 10542
rect 10692 9920 10744 9926
rect 10692 9862 10744 9868
rect 10508 9716 10560 9722
rect 10508 9658 10560 9664
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10520 9178 10548 9522
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10612 8974 10640 9046
rect 10600 8968 10652 8974
rect 10600 8910 10652 8916
rect 10600 8832 10652 8838
rect 10600 8774 10652 8780
rect 10612 8430 10640 8774
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10600 8288 10652 8294
rect 10600 8230 10652 8236
rect 10416 7880 10468 7886
rect 10416 7822 10468 7828
rect 10232 7744 10284 7750
rect 10232 7686 10284 7692
rect 10244 7546 10272 7686
rect 10048 7540 10100 7546
rect 10048 7482 10100 7488
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9954 7168 10010 7177
rect 9954 7103 10010 7112
rect 9864 6860 9916 6866
rect 9864 6802 9916 6808
rect 9876 6322 9904 6802
rect 9968 6662 9996 7103
rect 10048 6996 10100 7002
rect 10048 6938 10100 6944
rect 9956 6656 10008 6662
rect 9956 6598 10008 6604
rect 9864 6316 9916 6322
rect 9864 6258 9916 6264
rect 10060 6225 10088 6938
rect 10152 6866 10180 7278
rect 10324 6928 10376 6934
rect 10324 6870 10376 6876
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10232 6860 10284 6866
rect 10232 6802 10284 6808
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10046 6216 10102 6225
rect 10046 6151 10102 6160
rect 9864 6112 9916 6118
rect 9864 6054 9916 6060
rect 9772 5364 9824 5370
rect 9772 5306 9824 5312
rect 9770 5264 9826 5273
rect 9770 5199 9826 5208
rect 9680 4480 9732 4486
rect 9508 4406 9628 4434
rect 9678 4448 9680 4457
rect 9732 4448 9734 4457
rect 9404 4072 9456 4078
rect 9404 4014 9456 4020
rect 9220 3188 9272 3194
rect 9220 3130 9272 3136
rect 9312 3188 9364 3194
rect 9312 3130 9364 3136
rect 9416 3058 9444 4014
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 9048 2910 9168 2938
rect 8747 2748 9055 2768
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2672 9055 2692
rect 8668 2372 8720 2378
rect 8588 2332 8668 2360
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 8312 1902 8340 2246
rect 8208 1896 8260 1902
rect 8208 1838 8260 1844
rect 8300 1896 8352 1902
rect 8300 1838 8352 1844
rect 8588 800 8616 2332
rect 8668 2314 8720 2320
rect 9140 1442 9168 2910
rect 9218 2816 9274 2825
rect 9218 2751 9274 2760
rect 9232 2650 9260 2751
rect 9402 2680 9458 2689
rect 9220 2644 9272 2650
rect 9402 2615 9404 2624
rect 9220 2586 9272 2592
rect 9456 2615 9458 2624
rect 9404 2586 9456 2592
rect 9508 2514 9536 4406
rect 9678 4383 9734 4392
rect 9784 3534 9812 5199
rect 9876 5137 9904 6054
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 9968 5273 9996 5578
rect 9954 5264 10010 5273
rect 9954 5199 9956 5208
rect 10008 5199 10010 5208
rect 10048 5228 10100 5234
rect 9956 5170 10008 5176
rect 10048 5170 10100 5176
rect 9968 5139 9996 5170
rect 9862 5128 9918 5137
rect 9862 5063 9918 5072
rect 9956 5024 10008 5030
rect 9956 4966 10008 4972
rect 9968 4146 9996 4966
rect 10060 4486 10088 5170
rect 10152 4622 10180 6598
rect 10244 6118 10272 6802
rect 10232 6112 10284 6118
rect 10232 6054 10284 6060
rect 10244 5642 10272 6054
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10232 5024 10284 5030
rect 10232 4966 10284 4972
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10048 4480 10100 4486
rect 10048 4422 10100 4428
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 10138 3768 10194 3777
rect 10138 3703 10194 3712
rect 9772 3528 9824 3534
rect 9772 3470 9824 3476
rect 10152 3194 10180 3703
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9600 2650 9628 2926
rect 10060 2825 10088 2994
rect 10244 2854 10272 4966
rect 10336 4486 10364 6870
rect 10428 5642 10456 7822
rect 10506 6760 10562 6769
rect 10506 6695 10562 6704
rect 10520 6089 10548 6695
rect 10506 6080 10562 6089
rect 10506 6015 10562 6024
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10414 5400 10470 5409
rect 10414 5335 10416 5344
rect 10468 5335 10470 5344
rect 10416 5306 10468 5312
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10428 5001 10456 5170
rect 10414 4992 10470 5001
rect 10414 4927 10470 4936
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10428 3942 10456 4927
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10416 3460 10468 3466
rect 10416 3402 10468 3408
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10336 3126 10364 3334
rect 10324 3120 10376 3126
rect 10324 3062 10376 3068
rect 10428 2990 10456 3402
rect 10416 2984 10468 2990
rect 10416 2926 10468 2932
rect 10232 2848 10284 2854
rect 10046 2816 10102 2825
rect 10232 2790 10284 2796
rect 10046 2751 10102 2760
rect 10230 2680 10286 2689
rect 9588 2644 9640 2650
rect 10230 2615 10286 2624
rect 9588 2586 9640 2592
rect 10244 2514 10272 2615
rect 10428 2582 10456 2926
rect 10416 2576 10468 2582
rect 10416 2518 10468 2524
rect 9496 2508 9548 2514
rect 9496 2450 9548 2456
rect 10232 2508 10284 2514
rect 10232 2450 10284 2456
rect 9508 1714 9536 2450
rect 10416 2372 10468 2378
rect 10520 2360 10548 5714
rect 10612 3398 10640 8230
rect 10888 7546 10916 17750
rect 11256 17678 11284 18906
rect 11610 18864 11666 18873
rect 11610 18799 11612 18808
rect 11664 18799 11666 18808
rect 11612 18770 11664 18776
rect 11346 18524 11654 18544
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18448 11654 18468
rect 11612 18352 11664 18358
rect 11612 18294 11664 18300
rect 11624 18193 11652 18294
rect 11716 18290 11744 19110
rect 11794 18864 11850 18873
rect 11794 18799 11850 18808
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 11610 18184 11666 18193
rect 11610 18119 11666 18128
rect 11808 18057 11836 18799
rect 11794 18048 11850 18057
rect 11794 17983 11850 17992
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11704 17604 11756 17610
rect 11704 17546 11756 17552
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11164 16794 11192 17478
rect 11346 17436 11654 17456
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17360 11654 17380
rect 11716 17066 11744 17546
rect 11796 17264 11848 17270
rect 11796 17206 11848 17212
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 11152 16788 11204 16794
rect 11152 16730 11204 16736
rect 11716 16658 11744 17002
rect 11244 16652 11296 16658
rect 11244 16594 11296 16600
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11072 15162 11100 16526
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 11164 16250 11192 16390
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11152 16040 11204 16046
rect 11152 15982 11204 15988
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 10980 14278 11008 14486
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 11072 13870 11100 15098
rect 11164 14482 11192 15982
rect 11256 14618 11284 16594
rect 11808 16454 11836 17206
rect 11900 16794 11928 20198
rect 12348 19848 12400 19854
rect 12348 19790 12400 19796
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 11980 19304 12032 19310
rect 11980 19246 12032 19252
rect 11992 18902 12020 19246
rect 11980 18896 12032 18902
rect 11980 18838 12032 18844
rect 11992 18766 12020 18838
rect 11980 18760 12032 18766
rect 11980 18702 12032 18708
rect 12084 17524 12112 19314
rect 12256 19304 12308 19310
rect 12256 19246 12308 19252
rect 12164 19236 12216 19242
rect 12164 19178 12216 19184
rect 12176 18766 12204 19178
rect 12164 18760 12216 18766
rect 12164 18702 12216 18708
rect 12268 18630 12296 19246
rect 12360 18970 12388 19790
rect 12452 19446 12480 20266
rect 12636 19938 12664 22200
rect 13096 20602 13124 22200
rect 13556 20602 13584 22200
rect 14016 20602 14044 22200
rect 14476 20602 14504 22200
rect 14936 20618 14964 22200
rect 14936 20602 15240 20618
rect 15396 20602 15424 22200
rect 15856 20602 15884 22200
rect 16316 20602 16344 22200
rect 16776 20890 16804 22200
rect 16776 20862 16988 20890
rect 16544 20700 16852 20720
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20624 16852 20644
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13544 20596 13596 20602
rect 13544 20538 13596 20544
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 14464 20596 14516 20602
rect 14936 20596 15252 20602
rect 14936 20590 15200 20596
rect 14464 20538 14516 20544
rect 15200 20538 15252 20544
rect 15384 20596 15436 20602
rect 15384 20538 15436 20544
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 16304 20596 16356 20602
rect 16304 20538 16356 20544
rect 12636 19910 12848 19938
rect 12532 19848 12584 19854
rect 12532 19790 12584 19796
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12452 19174 12480 19382
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12348 18964 12400 18970
rect 12348 18906 12400 18912
rect 12256 18624 12308 18630
rect 12256 18566 12308 18572
rect 12164 18420 12216 18426
rect 12268 18408 12296 18566
rect 12216 18380 12296 18408
rect 12164 18362 12216 18368
rect 12360 18358 12388 18906
rect 12348 18352 12400 18358
rect 12348 18294 12400 18300
rect 12254 17912 12310 17921
rect 12254 17847 12310 17856
rect 11992 17496 12112 17524
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11796 16448 11848 16454
rect 11796 16390 11848 16396
rect 11346 16348 11654 16368
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16272 11654 16292
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11704 15496 11756 15502
rect 11704 15438 11756 15444
rect 11346 15260 11654 15280
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15184 11654 15204
rect 11244 14612 11296 14618
rect 11244 14554 11296 14560
rect 11152 14476 11204 14482
rect 11152 14418 11204 14424
rect 11346 14172 11654 14192
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14096 11654 14116
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11164 12986 11192 13874
rect 11716 13530 11744 15438
rect 11796 15156 11848 15162
rect 11796 15098 11848 15104
rect 11808 15026 11836 15098
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11808 13870 11836 14214
rect 11900 14074 11928 16050
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11796 13864 11848 13870
rect 11796 13806 11848 13812
rect 11704 13524 11756 13530
rect 11704 13466 11756 13472
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11152 12980 11204 12986
rect 11152 12922 11204 12928
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 11072 12238 11100 12718
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11256 12102 11284 13126
rect 11346 13084 11654 13104
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13008 11654 13028
rect 11716 12986 11744 13126
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11348 12238 11376 12854
rect 11704 12640 11756 12646
rect 11704 12582 11756 12588
rect 11336 12232 11388 12238
rect 11336 12174 11388 12180
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11346 11996 11654 12016
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11920 11654 11940
rect 11242 11656 11298 11665
rect 11242 11591 11298 11600
rect 10966 11248 11022 11257
rect 10966 11183 11022 11192
rect 11152 11212 11204 11218
rect 10980 11014 11008 11183
rect 11152 11154 11204 11160
rect 10968 11008 11020 11014
rect 10968 10950 11020 10956
rect 11060 9988 11112 9994
rect 11060 9930 11112 9936
rect 11072 9654 11100 9930
rect 11164 9926 11192 11154
rect 11152 9920 11204 9926
rect 11152 9862 11204 9868
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 11072 9042 11100 9590
rect 11164 9042 11192 9862
rect 11060 9036 11112 9042
rect 11060 8978 11112 8984
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10980 8634 11008 8774
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11060 8628 11112 8634
rect 11060 8570 11112 8576
rect 11072 8498 11100 8570
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11058 7848 11114 7857
rect 11058 7783 11114 7792
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10876 7540 10928 7546
rect 10876 7482 10928 7488
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10704 6322 10732 7210
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10796 6662 10824 7142
rect 10888 7002 10916 7142
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 10980 6882 11008 7686
rect 10888 6854 11008 6882
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10692 6316 10744 6322
rect 10692 6258 10744 6264
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10704 5166 10732 6258
rect 10692 5160 10744 5166
rect 10692 5102 10744 5108
rect 10704 4826 10732 5102
rect 10796 5030 10824 6258
rect 10888 5030 10916 6854
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10784 5024 10836 5030
rect 10784 4966 10836 4972
rect 10876 5024 10928 5030
rect 10876 4966 10928 4972
rect 10692 4820 10744 4826
rect 10692 4762 10744 4768
rect 10888 4690 10916 4966
rect 10876 4684 10928 4690
rect 10796 4644 10876 4672
rect 10692 4480 10744 4486
rect 10690 4448 10692 4457
rect 10744 4448 10746 4457
rect 10690 4383 10746 4392
rect 10796 4298 10824 4644
rect 10876 4626 10928 4632
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10704 4270 10824 4298
rect 10888 4282 10916 4422
rect 10876 4276 10928 4282
rect 10704 4078 10732 4270
rect 10876 4218 10928 4224
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10782 4040 10838 4049
rect 10782 3975 10838 3984
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10612 2446 10640 3130
rect 10704 2514 10732 3878
rect 10796 3738 10824 3975
rect 10980 3890 11008 6734
rect 11072 6186 11100 7783
rect 11256 7290 11284 11591
rect 11520 11552 11572 11558
rect 11520 11494 11572 11500
rect 11532 11393 11560 11494
rect 11518 11384 11574 11393
rect 11518 11319 11574 11328
rect 11346 10908 11654 10928
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10832 11654 10852
rect 11612 10668 11664 10674
rect 11612 10610 11664 10616
rect 11624 10470 11652 10610
rect 11612 10464 11664 10470
rect 11612 10406 11664 10412
rect 11716 10033 11744 12582
rect 11808 11762 11836 13806
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11900 12345 11928 13670
rect 11886 12336 11942 12345
rect 11886 12271 11942 12280
rect 11796 11756 11848 11762
rect 11796 11698 11848 11704
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11808 11150 11836 11698
rect 11900 11558 11928 11698
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11992 11200 12020 17496
rect 12268 15366 12296 17847
rect 12360 15978 12388 18294
rect 12544 17338 12572 19790
rect 12624 19780 12676 19786
rect 12624 19722 12676 19728
rect 12636 18970 12664 19722
rect 12820 19378 12848 19910
rect 12912 19514 12940 20538
rect 13268 20460 13320 20466
rect 13268 20402 13320 20408
rect 13544 20460 13596 20466
rect 13544 20402 13596 20408
rect 13636 20460 13688 20466
rect 13636 20402 13688 20408
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 14280 20460 14332 20466
rect 14280 20402 14332 20408
rect 14832 20460 14884 20466
rect 14832 20402 14884 20408
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 12900 19508 12952 19514
rect 12900 19450 12952 19456
rect 13082 19408 13138 19417
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12808 19372 12860 19378
rect 13082 19343 13084 19352
rect 12808 19314 12860 19320
rect 13136 19343 13138 19352
rect 13084 19314 13136 19320
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12624 18692 12676 18698
rect 12624 18634 12676 18640
rect 12636 18290 12664 18634
rect 12624 18284 12676 18290
rect 12624 18226 12676 18232
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12532 17332 12584 17338
rect 12452 17292 12532 17320
rect 12348 15972 12400 15978
rect 12348 15914 12400 15920
rect 12360 15570 12388 15914
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 12256 15360 12308 15366
rect 12256 15302 12308 15308
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 12162 14240 12218 14249
rect 12084 13938 12112 14214
rect 12162 14175 12218 14184
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 12084 12442 12112 12786
rect 12072 12436 12124 12442
rect 12072 12378 12124 12384
rect 12176 11830 12204 14175
rect 12164 11824 12216 11830
rect 12164 11766 12216 11772
rect 12268 11694 12296 15302
rect 12360 15094 12388 15506
rect 12348 15088 12400 15094
rect 12348 15030 12400 15036
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 12360 14074 12388 14350
rect 12348 14068 12400 14074
rect 12348 14010 12400 14016
rect 12360 13734 12388 14010
rect 12348 13728 12400 13734
rect 12348 13670 12400 13676
rect 12452 12434 12480 17292
rect 12532 17274 12584 17280
rect 12530 16688 12586 16697
rect 12530 16623 12586 16632
rect 12544 14362 12572 16623
rect 12636 16522 12664 17478
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12636 14482 12664 14962
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12544 14334 12664 14362
rect 12636 14278 12664 14334
rect 12624 14272 12676 14278
rect 12624 14214 12676 14220
rect 12636 13977 12664 14214
rect 12622 13968 12678 13977
rect 12622 13903 12678 13912
rect 12728 12442 12756 19314
rect 12820 18902 12848 19314
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 12808 18896 12860 18902
rect 12808 18838 12860 18844
rect 12912 18766 12940 19110
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12900 18760 12952 18766
rect 12900 18702 12952 18708
rect 12820 14006 12848 18702
rect 13004 17882 13032 19110
rect 13280 18902 13308 20402
rect 13452 20324 13504 20330
rect 13452 20266 13504 20272
rect 13360 19848 13412 19854
rect 13360 19790 13412 19796
rect 13372 18970 13400 19790
rect 13464 19514 13492 20266
rect 13556 20058 13584 20402
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13544 19780 13596 19786
rect 13544 19722 13596 19728
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13450 19136 13506 19145
rect 13450 19071 13506 19080
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13268 18896 13320 18902
rect 13268 18838 13320 18844
rect 13268 18352 13320 18358
rect 13266 18320 13268 18329
rect 13320 18320 13322 18329
rect 13084 18284 13136 18290
rect 13464 18290 13492 19071
rect 13266 18255 13322 18264
rect 13452 18284 13504 18290
rect 13084 18226 13136 18232
rect 13452 18226 13504 18232
rect 13096 17882 13124 18226
rect 12992 17876 13044 17882
rect 12992 17818 13044 17824
rect 13084 17876 13136 17882
rect 13084 17818 13136 17824
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13372 17338 13400 17614
rect 13360 17332 13412 17338
rect 13360 17274 13412 17280
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13188 16794 13216 17138
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 13556 16574 13584 19722
rect 13648 19514 13676 20402
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13636 19508 13688 19514
rect 13636 19450 13688 19456
rect 13740 19242 13768 19790
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13634 19000 13690 19009
rect 13634 18935 13636 18944
rect 13688 18935 13690 18944
rect 13636 18906 13688 18912
rect 13832 17882 13860 20402
rect 13945 20156 14253 20176
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20080 14253 20100
rect 14292 20058 14320 20402
rect 14646 20360 14702 20369
rect 14372 20324 14424 20330
rect 14646 20295 14702 20304
rect 14372 20266 14424 20272
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14384 19990 14412 20266
rect 14372 19984 14424 19990
rect 14372 19926 14424 19932
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14372 19848 14424 19854
rect 14372 19790 14424 19796
rect 14292 19174 14320 19790
rect 14384 19514 14412 19790
rect 14462 19680 14518 19689
rect 14462 19615 14518 19624
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 13945 19068 14253 19088
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 18992 14253 19012
rect 13912 18896 13964 18902
rect 13910 18864 13912 18873
rect 13964 18864 13966 18873
rect 13910 18799 13966 18808
rect 13945 17980 14253 18000
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17904 14253 17924
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13945 16892 14253 16912
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16816 14253 16836
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13372 16546 13584 16574
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 13096 16250 13124 16390
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 13004 15570 13032 16050
rect 12992 15564 13044 15570
rect 12992 15506 13044 15512
rect 12900 15156 12952 15162
rect 13004 15144 13032 15506
rect 13176 15360 13228 15366
rect 13176 15302 13228 15308
rect 13188 15162 13216 15302
rect 12952 15116 13032 15144
rect 13176 15156 13228 15162
rect 12900 15098 12952 15104
rect 13176 15098 13228 15104
rect 13268 14544 13320 14550
rect 13268 14486 13320 14492
rect 13280 14278 13308 14486
rect 13268 14272 13320 14278
rect 13268 14214 13320 14220
rect 12808 14000 12860 14006
rect 12808 13942 12860 13948
rect 12808 13796 12860 13802
rect 12808 13738 12860 13744
rect 12820 13190 12848 13738
rect 13372 13410 13400 16546
rect 13544 16448 13596 16454
rect 13544 16390 13596 16396
rect 13556 15706 13584 16390
rect 13832 16250 13860 16594
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13945 15804 14253 15824
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15728 14253 15748
rect 13544 15700 13596 15706
rect 13544 15642 13596 15648
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 13832 15162 13860 15370
rect 13820 15156 13872 15162
rect 13820 15098 13872 15104
rect 13728 15020 13780 15026
rect 13728 14962 13780 14968
rect 13452 14952 13504 14958
rect 13452 14894 13504 14900
rect 13280 13382 13400 13410
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12912 12986 12940 13262
rect 13176 13184 13228 13190
rect 13176 13126 13228 13132
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 12716 12436 12768 12442
rect 12452 12406 12664 12434
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12360 11393 12388 11698
rect 12346 11384 12402 11393
rect 12346 11319 12402 11328
rect 12530 11384 12586 11393
rect 12636 11370 12664 12406
rect 12716 12378 12768 12384
rect 12912 12306 12940 12922
rect 13188 12782 13216 13126
rect 13176 12776 13228 12782
rect 13176 12718 13228 12724
rect 13280 12434 13308 13382
rect 13358 13288 13414 13297
rect 13358 13223 13414 13232
rect 13372 12986 13400 13223
rect 13464 12986 13492 14894
rect 13740 14618 13768 14962
rect 13820 14884 13872 14890
rect 13820 14826 13872 14832
rect 13728 14612 13780 14618
rect 13728 14554 13780 14560
rect 13832 14482 13860 14826
rect 13945 14716 14253 14736
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14640 14253 14660
rect 13820 14476 13872 14482
rect 13820 14418 13872 14424
rect 13636 14272 13688 14278
rect 13636 14214 13688 14220
rect 13360 12980 13412 12986
rect 13360 12922 13412 12928
rect 13452 12980 13504 12986
rect 13452 12922 13504 12928
rect 13372 12646 13400 12922
rect 13452 12776 13504 12782
rect 13452 12718 13504 12724
rect 13360 12640 13412 12646
rect 13360 12582 13412 12588
rect 13188 12406 13308 12434
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 12636 11342 12940 11370
rect 12530 11319 12586 11328
rect 11992 11172 12112 11200
rect 11796 11144 11848 11150
rect 11796 11086 11848 11092
rect 11808 10810 11836 11086
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11796 10804 11848 10810
rect 11796 10746 11848 10752
rect 11796 10600 11848 10606
rect 11796 10542 11848 10548
rect 11702 10024 11758 10033
rect 11702 9959 11758 9968
rect 11704 9920 11756 9926
rect 11704 9862 11756 9868
rect 11346 9820 11654 9840
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9744 11654 9764
rect 11716 9518 11744 9862
rect 11704 9512 11756 9518
rect 11704 9454 11756 9460
rect 11704 9036 11756 9042
rect 11704 8978 11756 8984
rect 11346 8732 11654 8752
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8656 11654 8676
rect 11716 8430 11744 8978
rect 11808 8974 11836 10542
rect 11888 9580 11940 9586
rect 11888 9522 11940 9528
rect 11900 9178 11928 9522
rect 11888 9172 11940 9178
rect 11888 9114 11940 9120
rect 11796 8968 11848 8974
rect 11796 8910 11848 8916
rect 11704 8424 11756 8430
rect 11796 8424 11848 8430
rect 11704 8366 11756 8372
rect 11794 8392 11796 8401
rect 11848 8392 11850 8401
rect 11794 8327 11850 8336
rect 11346 7644 11654 7664
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7568 11654 7588
rect 11164 7262 11284 7290
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 11060 5840 11112 5846
rect 11060 5782 11112 5788
rect 11072 5545 11100 5782
rect 11164 5574 11192 7262
rect 11886 7032 11942 7041
rect 11886 6967 11942 6976
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11152 5568 11204 5574
rect 11058 5536 11114 5545
rect 11152 5510 11204 5516
rect 11058 5471 11114 5480
rect 11256 5370 11284 6598
rect 11346 6556 11654 6576
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6480 11654 6500
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11348 5778 11376 6054
rect 11624 5846 11652 6054
rect 11612 5840 11664 5846
rect 11612 5782 11664 5788
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11346 5468 11654 5488
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5392 11654 5412
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11244 5364 11296 5370
rect 11244 5306 11296 5312
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 11072 4690 11100 5238
rect 11164 5234 11192 5306
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11520 5160 11572 5166
rect 11520 5102 11572 5108
rect 11060 4684 11112 4690
rect 11112 4644 11192 4672
rect 11060 4626 11112 4632
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 11072 4214 11100 4490
rect 11060 4208 11112 4214
rect 11060 4150 11112 4156
rect 10888 3862 11008 3890
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10888 3505 10916 3862
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10874 3496 10930 3505
rect 10874 3431 10930 3440
rect 10784 3392 10836 3398
rect 10784 3334 10836 3340
rect 10692 2508 10744 2514
rect 10692 2450 10744 2456
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10468 2332 10548 2360
rect 10416 2314 10468 2320
rect 10520 1714 10548 2332
rect 9508 1686 9628 1714
rect 9048 1414 9168 1442
rect 9048 800 9076 1414
rect 9600 800 9628 1686
rect 10428 1686 10548 1714
rect 10060 870 10180 898
rect 10060 800 10088 870
rect 6012 734 6224 762
rect 6274 0 6330 800
rect 6734 0 6790 800
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8574 0 8630 800
rect 9034 0 9090 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10152 762 10180 870
rect 10428 762 10456 1686
rect 10520 870 10640 898
rect 10520 800 10548 870
rect 10152 734 10456 762
rect 10506 0 10562 800
rect 10612 762 10640 870
rect 10796 762 10824 3334
rect 10888 3058 10916 3431
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10980 800 11008 3674
rect 11060 3052 11112 3058
rect 11164 3040 11192 4644
rect 11256 3942 11284 5102
rect 11532 5030 11560 5102
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11716 4826 11744 6598
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11704 4820 11756 4826
rect 11704 4762 11756 4768
rect 11440 4554 11468 4762
rect 11428 4548 11480 4554
rect 11428 4490 11480 4496
rect 11346 4380 11654 4400
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4304 11654 4324
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 11532 3777 11560 4014
rect 11518 3768 11574 3777
rect 11518 3703 11574 3712
rect 11346 3292 11654 3312
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3216 11654 3236
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 11112 3012 11192 3040
rect 11060 2994 11112 3000
rect 11256 2088 11284 3062
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11348 2825 11376 2926
rect 11334 2816 11390 2825
rect 11808 2774 11836 6598
rect 11900 6458 11928 6967
rect 11992 6914 12020 11018
rect 12084 10470 12112 11172
rect 12256 11008 12308 11014
rect 12256 10950 12308 10956
rect 12268 10810 12296 10950
rect 12256 10804 12308 10810
rect 12256 10746 12308 10752
rect 12440 10600 12492 10606
rect 12440 10542 12492 10548
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 12072 9512 12124 9518
rect 12072 9454 12124 9460
rect 12084 8634 12112 9454
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12176 8566 12204 9998
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12176 7818 12204 8502
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12176 7478 12204 7754
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 12268 7324 12296 10406
rect 12452 10266 12480 10542
rect 12440 10260 12492 10266
rect 12440 10202 12492 10208
rect 12544 7857 12572 11319
rect 12808 11212 12860 11218
rect 12808 11154 12860 11160
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12636 9450 12664 10610
rect 12820 10062 12848 11154
rect 12808 10056 12860 10062
rect 12808 9998 12860 10004
rect 12624 9444 12676 9450
rect 12624 9386 12676 9392
rect 12808 8900 12860 8906
rect 12808 8842 12860 8848
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12728 8362 12756 8570
rect 12716 8356 12768 8362
rect 12716 8298 12768 8304
rect 12820 7886 12848 8842
rect 12912 8090 12940 11342
rect 13188 11257 13216 12406
rect 13268 12096 13320 12102
rect 13268 12038 13320 12044
rect 13280 11558 13308 12038
rect 13360 11688 13412 11694
rect 13360 11630 13412 11636
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13174 11248 13230 11257
rect 13174 11183 13230 11192
rect 13372 10577 13400 11630
rect 13358 10568 13414 10577
rect 13358 10503 13414 10512
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 12992 8900 13044 8906
rect 12992 8842 13044 8848
rect 13004 8537 13032 8842
rect 12990 8528 13046 8537
rect 12990 8463 13046 8472
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12990 7984 13046 7993
rect 12990 7919 13046 7928
rect 12808 7880 12860 7886
rect 12530 7848 12586 7857
rect 12808 7822 12860 7828
rect 12530 7783 12586 7792
rect 12544 7546 12572 7783
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12176 7296 12296 7324
rect 11992 6886 12112 6914
rect 11978 6760 12034 6769
rect 11978 6695 12034 6704
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11992 6390 12020 6695
rect 11980 6384 12032 6390
rect 11980 6326 12032 6332
rect 11888 6112 11940 6118
rect 11888 6054 11940 6060
rect 11900 5817 11928 6054
rect 11886 5808 11942 5817
rect 11886 5743 11942 5752
rect 11888 5568 11940 5574
rect 11888 5510 11940 5516
rect 11900 5370 11928 5510
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 11886 4856 11942 4865
rect 11886 4791 11942 4800
rect 11900 4185 11928 4791
rect 11886 4176 11942 4185
rect 11886 4111 11942 4120
rect 11886 3224 11942 3233
rect 11886 3159 11942 3168
rect 11900 3126 11928 3159
rect 11888 3120 11940 3126
rect 11888 3062 11940 3068
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 11334 2751 11390 2760
rect 11716 2746 11836 2774
rect 11346 2204 11654 2224
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2128 11654 2148
rect 11256 2060 11468 2088
rect 11440 800 11468 2060
rect 11716 1873 11744 2746
rect 11900 2446 11928 2790
rect 12084 2514 12112 6886
rect 12176 2514 12204 7296
rect 12346 7168 12402 7177
rect 12346 7103 12402 7112
rect 12360 6798 12388 7103
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12348 6112 12400 6118
rect 12348 6054 12400 6060
rect 12254 5264 12310 5273
rect 12254 5199 12256 5208
rect 12308 5199 12310 5208
rect 12256 5170 12308 5176
rect 12360 5114 12388 6054
rect 12268 5086 12388 5114
rect 12268 3097 12296 5086
rect 12348 5024 12400 5030
rect 12348 4966 12400 4972
rect 12360 4486 12388 4966
rect 12452 4486 12480 7482
rect 12636 7410 12664 7686
rect 12624 7404 12676 7410
rect 12624 7346 12676 7352
rect 12806 6896 12862 6905
rect 12806 6831 12808 6840
rect 12860 6831 12862 6840
rect 12900 6860 12952 6866
rect 12808 6802 12860 6808
rect 12900 6802 12952 6808
rect 12912 6390 12940 6802
rect 13004 6458 13032 7919
rect 13084 7744 13136 7750
rect 13084 7686 13136 7692
rect 13096 7342 13124 7686
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 12992 6452 13044 6458
rect 12992 6394 13044 6400
rect 12900 6384 12952 6390
rect 12820 6332 12900 6338
rect 12820 6326 12952 6332
rect 12532 6316 12584 6322
rect 12532 6258 12584 6264
rect 12820 6310 12940 6326
rect 12544 5778 12572 6258
rect 12820 5794 12848 6310
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12912 5914 12940 6190
rect 13096 5930 13124 7278
rect 13280 6882 13308 9658
rect 13372 7546 13400 10503
rect 13464 8974 13492 12718
rect 13544 12164 13596 12170
rect 13544 12106 13596 12112
rect 13556 11898 13584 12106
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13544 11620 13596 11626
rect 13544 11562 13596 11568
rect 13556 11082 13584 11562
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13544 10260 13596 10266
rect 13544 10202 13596 10208
rect 13556 9586 13584 10202
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13452 8968 13504 8974
rect 13450 8936 13452 8945
rect 13504 8936 13506 8945
rect 13648 8906 13676 14214
rect 13832 14074 13860 14418
rect 14292 14414 14320 19110
rect 14384 17134 14412 19450
rect 14476 18426 14504 19615
rect 14660 18970 14688 20295
rect 14844 20058 14872 20402
rect 15120 20058 15148 20402
rect 15948 20058 15976 20402
rect 14832 20052 14884 20058
rect 14832 19994 14884 20000
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 16684 19990 16712 20402
rect 16960 20330 16988 20862
rect 17236 20602 17264 22200
rect 17696 20618 17724 22200
rect 17696 20602 18000 20618
rect 18156 20602 18184 22200
rect 18616 20602 18644 22200
rect 17224 20596 17276 20602
rect 17696 20596 18012 20602
rect 17696 20590 17960 20596
rect 17224 20538 17276 20544
rect 17960 20538 18012 20544
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 18604 20596 18656 20602
rect 19076 20584 19104 22200
rect 19536 20602 19564 22200
rect 19996 20602 20024 22200
rect 20456 20602 20484 22200
rect 20916 20602 20944 22200
rect 21376 21026 21404 22200
rect 21376 20998 21496 21026
rect 19340 20596 19392 20602
rect 19076 20556 19340 20584
rect 18604 20538 18656 20544
rect 19340 20538 19392 20544
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 20444 20596 20496 20602
rect 20444 20538 20496 20544
rect 20904 20596 20956 20602
rect 20904 20538 20956 20544
rect 17040 20460 17092 20466
rect 17040 20402 17092 20408
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17684 20460 17736 20466
rect 17684 20402 17736 20408
rect 17960 20460 18012 20466
rect 17960 20402 18012 20408
rect 18328 20460 18380 20466
rect 18328 20402 18380 20408
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 19708 20460 19760 20466
rect 19708 20402 19760 20408
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 21180 20460 21232 20466
rect 21180 20402 21232 20408
rect 16948 20324 17000 20330
rect 16948 20266 17000 20272
rect 17052 20058 17080 20402
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 16672 19984 16724 19990
rect 15212 19910 15424 19938
rect 16672 19926 16724 19932
rect 14740 19848 14792 19854
rect 14740 19790 14792 19796
rect 14752 19514 14780 19790
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14740 19372 14792 19378
rect 14740 19314 14792 19320
rect 15016 19372 15068 19378
rect 15016 19314 15068 19320
rect 14648 18964 14700 18970
rect 14648 18906 14700 18912
rect 14464 18420 14516 18426
rect 14464 18362 14516 18368
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14280 14408 14332 14414
rect 14280 14350 14332 14356
rect 13820 14068 13872 14074
rect 13820 14010 13872 14016
rect 13728 13932 13780 13938
rect 13728 13874 13780 13880
rect 13740 13190 13768 13874
rect 13945 13628 14253 13648
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13552 14253 13572
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13945 12540 14253 12560
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12464 14253 12484
rect 14384 11830 14412 17070
rect 14464 16720 14516 16726
rect 14464 16662 14516 16668
rect 14476 16574 14504 16662
rect 14752 16574 14780 19314
rect 14830 18728 14886 18737
rect 14830 18663 14832 18672
rect 14884 18663 14886 18672
rect 14832 18634 14884 18640
rect 14832 18080 14884 18086
rect 14832 18022 14884 18028
rect 14476 16546 14596 16574
rect 14464 12776 14516 12782
rect 14464 12718 14516 12724
rect 14476 11898 14504 12718
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 13820 11824 13872 11830
rect 13820 11766 13872 11772
rect 14372 11824 14424 11830
rect 14372 11766 14424 11772
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13450 8871 13506 8880
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13740 8634 13768 11494
rect 13832 11150 13860 11766
rect 13945 11452 14253 11472
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11376 14253 11396
rect 14568 11234 14596 16546
rect 14660 16546 14780 16574
rect 14660 12986 14688 16546
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14752 15502 14780 16390
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14752 13870 14780 14214
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14752 13394 14780 13806
rect 14740 13388 14792 13394
rect 14740 13330 14792 13336
rect 14648 12980 14700 12986
rect 14648 12922 14700 12928
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14384 11206 14596 11234
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 14188 10668 14240 10674
rect 14188 10610 14240 10616
rect 14200 10554 14228 10610
rect 14200 10526 14320 10554
rect 13945 10364 14253 10384
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10288 14253 10308
rect 14292 9722 14320 10526
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14384 9654 14412 11206
rect 14464 11144 14516 11150
rect 14660 11098 14688 12378
rect 14752 12170 14780 13330
rect 14844 12730 14872 18022
rect 14924 14272 14976 14278
rect 14924 14214 14976 14220
rect 14936 14074 14964 14214
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14844 12702 14964 12730
rect 14832 12640 14884 12646
rect 14832 12582 14884 12588
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14464 11086 14516 11092
rect 14476 10674 14504 11086
rect 14568 11070 14688 11098
rect 14568 10810 14596 11070
rect 14648 11008 14700 11014
rect 14648 10950 14700 10956
rect 14660 10810 14688 10950
rect 14556 10804 14608 10810
rect 14556 10746 14608 10752
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14464 10668 14516 10674
rect 14464 10610 14516 10616
rect 14372 9648 14424 9654
rect 14372 9590 14424 9596
rect 14372 9512 14424 9518
rect 14372 9454 14424 9460
rect 13945 9276 14253 9296
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9200 14253 9220
rect 13820 9036 13872 9042
rect 13820 8978 13872 8984
rect 13728 8628 13780 8634
rect 13728 8570 13780 8576
rect 13832 8498 13860 8978
rect 14384 8974 14412 9454
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14280 8832 14332 8838
rect 14280 8774 14332 8780
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13832 7954 13860 8298
rect 13945 8188 14253 8208
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8112 14253 8132
rect 14292 7954 14320 8774
rect 14476 8634 14504 10610
rect 14752 10606 14780 12106
rect 14740 10600 14792 10606
rect 14740 10542 14792 10548
rect 14752 10130 14780 10542
rect 14740 10124 14792 10130
rect 14740 10066 14792 10072
rect 14648 10056 14700 10062
rect 14648 9998 14700 10004
rect 14556 8832 14608 8838
rect 14556 8774 14608 8780
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 14280 7948 14332 7954
rect 14280 7890 14332 7896
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13360 7540 13412 7546
rect 13360 7482 13412 7488
rect 13452 7404 13504 7410
rect 13452 7346 13504 7352
rect 13464 7002 13492 7346
rect 13452 6996 13504 7002
rect 13452 6938 13504 6944
rect 13280 6854 13492 6882
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13372 6322 13400 6734
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13268 6180 13320 6186
rect 13268 6122 13320 6128
rect 13176 6112 13228 6118
rect 13176 6054 13228 6060
rect 12900 5908 12952 5914
rect 12900 5850 12952 5856
rect 13004 5902 13124 5930
rect 12532 5772 12584 5778
rect 12820 5766 12940 5794
rect 12532 5714 12584 5720
rect 12912 5642 12940 5766
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12532 4616 12584 4622
rect 12530 4584 12532 4593
rect 12584 4584 12586 4593
rect 12530 4519 12586 4528
rect 12636 4486 12664 5170
rect 12728 4690 12756 5578
rect 12806 5264 12862 5273
rect 12806 5199 12862 5208
rect 12820 5166 12848 5199
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12900 5092 12952 5098
rect 12900 5034 12952 5040
rect 12806 4856 12862 4865
rect 12806 4791 12862 4800
rect 12820 4690 12848 4791
rect 12716 4684 12768 4690
rect 12716 4626 12768 4632
rect 12808 4684 12860 4690
rect 12808 4626 12860 4632
rect 12348 4480 12400 4486
rect 12440 4480 12492 4486
rect 12348 4422 12400 4428
rect 12438 4448 12440 4457
rect 12624 4480 12676 4486
rect 12492 4448 12494 4457
rect 12624 4422 12676 4428
rect 12438 4383 12494 4392
rect 12452 4146 12480 4383
rect 12728 4282 12756 4626
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12348 3936 12400 3942
rect 12348 3878 12400 3884
rect 12254 3088 12310 3097
rect 12254 3023 12310 3032
rect 12360 3040 12388 3878
rect 12544 3670 12572 4082
rect 12532 3664 12584 3670
rect 12532 3606 12584 3612
rect 12544 3126 12572 3606
rect 12532 3120 12584 3126
rect 12532 3062 12584 3068
rect 12912 3058 12940 5034
rect 13004 5012 13032 5902
rect 13188 5681 13216 6054
rect 13280 5914 13308 6122
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13174 5672 13230 5681
rect 13174 5607 13230 5616
rect 13268 5636 13320 5642
rect 13268 5578 13320 5584
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 13096 5166 13124 5510
rect 13280 5386 13308 5578
rect 13188 5358 13308 5386
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13004 4984 13124 5012
rect 12990 4856 13046 4865
rect 12990 4791 13046 4800
rect 13004 4554 13032 4791
rect 12992 4548 13044 4554
rect 12992 4490 13044 4496
rect 13096 4078 13124 4984
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 12440 3052 12492 3058
rect 12360 3012 12440 3040
rect 12440 2994 12492 3000
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 13188 2938 13216 5358
rect 13268 5228 13320 5234
rect 13268 5170 13320 5176
rect 13280 4826 13308 5170
rect 13268 4820 13320 4826
rect 13268 4762 13320 4768
rect 13372 4078 13400 6258
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13268 3936 13320 3942
rect 13268 3878 13320 3884
rect 13280 3466 13308 3878
rect 13372 3534 13400 4014
rect 13464 3942 13492 6854
rect 13648 6798 13676 7822
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13740 7546 13768 7754
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13832 7342 13860 7890
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 14384 7324 14412 8230
rect 14476 7954 14504 8570
rect 14464 7948 14516 7954
rect 14464 7890 14516 7896
rect 14568 7818 14596 8774
rect 14556 7812 14608 7818
rect 14556 7754 14608 7760
rect 14464 7336 14516 7342
rect 14384 7296 14464 7324
rect 13945 7100 14253 7120
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7024 14253 7044
rect 14384 6934 14412 7296
rect 14464 7278 14516 7284
rect 14372 6928 14424 6934
rect 14372 6870 14424 6876
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13924 6458 13952 6598
rect 13912 6452 13964 6458
rect 13912 6394 13964 6400
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13648 5574 13676 6258
rect 14660 6254 14688 9998
rect 14740 9648 14792 9654
rect 14740 9590 14792 9596
rect 14752 6746 14780 9590
rect 14844 8974 14872 12582
rect 14936 12322 14964 12702
rect 15028 12442 15056 19314
rect 15108 14952 15160 14958
rect 15108 14894 15160 14900
rect 15120 14006 15148 14894
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15016 12436 15068 12442
rect 15016 12378 15068 12384
rect 14936 12294 15056 12322
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14936 11898 14964 12174
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 15028 11801 15056 12294
rect 15014 11792 15070 11801
rect 15014 11727 15070 11736
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14924 8900 14976 8906
rect 14924 8842 14976 8848
rect 14936 8090 14964 8842
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 15028 7274 15056 8774
rect 15016 7268 15068 7274
rect 15016 7210 15068 7216
rect 14752 6718 14964 6746
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14648 6248 14700 6254
rect 14648 6190 14700 6196
rect 13945 6012 14253 6032
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5936 14253 5956
rect 14462 5944 14518 5953
rect 14462 5879 14518 5888
rect 14476 5710 14504 5879
rect 14464 5704 14516 5710
rect 14464 5646 14516 5652
rect 14660 5574 14688 6190
rect 14752 6118 14780 6598
rect 14740 6112 14792 6118
rect 14740 6054 14792 6060
rect 14832 6112 14884 6118
rect 14832 6054 14884 6060
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 14096 5568 14148 5574
rect 14096 5510 14148 5516
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14108 5370 14136 5510
rect 14096 5364 14148 5370
rect 14096 5306 14148 5312
rect 13728 5160 13780 5166
rect 13728 5102 13780 5108
rect 13740 4826 13768 5102
rect 14372 5092 14424 5098
rect 14372 5034 14424 5040
rect 13945 4924 14253 4944
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4848 14253 4868
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13912 4752 13964 4758
rect 13910 4720 13912 4729
rect 13964 4720 13966 4729
rect 13910 4655 13966 4664
rect 13728 4548 13780 4554
rect 13728 4490 13780 4496
rect 13636 4140 13688 4146
rect 13636 4082 13688 4088
rect 13648 3942 13676 4082
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13636 3936 13688 3942
rect 13636 3878 13688 3884
rect 13648 3738 13676 3878
rect 13636 3732 13688 3738
rect 13636 3674 13688 3680
rect 13360 3528 13412 3534
rect 13360 3470 13412 3476
rect 13268 3460 13320 3466
rect 13268 3402 13320 3408
rect 13452 3052 13504 3058
rect 13452 2994 13504 3000
rect 12912 2910 13216 2938
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 12808 2644 12860 2650
rect 12808 2586 12860 2592
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 11702 1864 11758 1873
rect 11702 1799 11758 1808
rect 11900 800 11928 2382
rect 12440 2372 12492 2378
rect 12360 2332 12440 2360
rect 12360 800 12388 2332
rect 12440 2314 12492 2320
rect 12820 800 12848 2586
rect 12912 1902 12940 2910
rect 13084 2848 13136 2854
rect 13084 2790 13136 2796
rect 13096 2514 13124 2790
rect 13084 2508 13136 2514
rect 13084 2450 13136 2456
rect 13280 2446 13308 2926
rect 13360 2848 13412 2854
rect 13360 2790 13412 2796
rect 13372 2582 13400 2790
rect 13360 2576 13412 2582
rect 13360 2518 13412 2524
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 12900 1896 12952 1902
rect 12900 1838 12952 1844
rect 13280 800 13308 2246
rect 13464 1737 13492 2994
rect 13740 2961 13768 4490
rect 14188 4480 14240 4486
rect 14188 4422 14240 4428
rect 14200 4214 14228 4422
rect 14188 4208 14240 4214
rect 14188 4150 14240 4156
rect 14280 4140 14332 4146
rect 14280 4082 14332 4088
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13832 3398 13860 3878
rect 13945 3836 14253 3856
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3760 14253 3780
rect 14004 3664 14056 3670
rect 14004 3606 14056 3612
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 14016 3058 14044 3606
rect 14188 3392 14240 3398
rect 14186 3360 14188 3369
rect 14240 3360 14242 3369
rect 14186 3295 14242 3304
rect 14292 3194 14320 4082
rect 14280 3188 14332 3194
rect 14280 3130 14332 3136
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 13726 2952 13782 2961
rect 13726 2887 13782 2896
rect 13820 2916 13872 2922
rect 13820 2858 13872 2864
rect 13728 2576 13780 2582
rect 13728 2518 13780 2524
rect 13450 1728 13506 1737
rect 13450 1663 13506 1672
rect 13740 800 13768 2518
rect 13832 2446 13860 2858
rect 14384 2774 14412 5034
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14476 3058 14504 4966
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14568 3738 14596 4422
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14464 3052 14516 3058
rect 14464 2994 14516 3000
rect 13945 2748 14253 2768
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2672 14253 2692
rect 14292 2746 14412 2774
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 14292 2360 14320 2746
rect 14200 2332 14320 2360
rect 14200 1630 14228 2332
rect 14372 2304 14424 2310
rect 14292 2264 14372 2292
rect 14188 1624 14240 1630
rect 14188 1566 14240 1572
rect 14292 800 14320 2264
rect 14372 2246 14424 2252
rect 14660 1766 14688 5510
rect 14752 5234 14780 6054
rect 14844 5846 14872 6054
rect 14832 5840 14884 5846
rect 14832 5782 14884 5788
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14936 5114 14964 6718
rect 14752 5086 14964 5114
rect 14752 4146 14780 5086
rect 14832 5024 14884 5030
rect 14832 4966 14884 4972
rect 14740 4140 14792 4146
rect 14740 4082 14792 4088
rect 14752 3738 14780 4082
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14740 2304 14792 2310
rect 14740 2246 14792 2252
rect 14648 1760 14700 1766
rect 14648 1702 14700 1708
rect 14752 800 14780 2246
rect 14844 2106 14872 4966
rect 14924 4480 14976 4486
rect 14924 4422 14976 4428
rect 14832 2100 14884 2106
rect 14832 2042 14884 2048
rect 14936 1698 14964 4422
rect 15016 4072 15068 4078
rect 15014 4040 15016 4049
rect 15068 4040 15070 4049
rect 15014 3975 15070 3984
rect 15016 3732 15068 3738
rect 15016 3674 15068 3680
rect 15028 3398 15056 3674
rect 15016 3392 15068 3398
rect 15016 3334 15068 3340
rect 15120 3194 15148 13466
rect 15212 13190 15240 19910
rect 15396 19854 15424 19910
rect 15292 19848 15344 19854
rect 15292 19790 15344 19796
rect 15384 19848 15436 19854
rect 15384 19790 15436 19796
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 16578 19816 16634 19825
rect 15304 19174 15332 19790
rect 15948 19514 15976 19790
rect 16578 19751 16580 19760
rect 16632 19751 16634 19760
rect 16948 19780 17000 19786
rect 16580 19722 16632 19728
rect 16948 19722 17000 19728
rect 16304 19712 16356 19718
rect 16304 19654 16356 19660
rect 16316 19514 16344 19654
rect 16544 19612 16852 19632
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19536 16852 19556
rect 16960 19514 16988 19722
rect 17144 19514 17172 20402
rect 17696 20058 17724 20402
rect 17972 20058 18000 20402
rect 18340 20058 18368 20402
rect 18420 20324 18472 20330
rect 18420 20266 18472 20272
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17960 20052 18012 20058
rect 17960 19994 18012 20000
rect 18328 20052 18380 20058
rect 18328 19994 18380 20000
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17500 19848 17552 19854
rect 17500 19790 17552 19796
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 16304 19508 16356 19514
rect 16304 19450 16356 19456
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 17040 19440 17092 19446
rect 17040 19382 17092 19388
rect 15474 19272 15530 19281
rect 15474 19207 15476 19216
rect 15528 19207 15530 19216
rect 15476 19178 15528 19184
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15660 19168 15712 19174
rect 15660 19110 15712 19116
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15304 15026 15332 19110
rect 15672 18737 15700 19110
rect 15658 18728 15714 18737
rect 15658 18663 15714 18672
rect 15764 15910 15792 19110
rect 16544 18524 16852 18544
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18448 16852 18468
rect 16544 17436 16852 17456
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17360 16852 17380
rect 16544 16348 16852 16368
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16272 16852 16292
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15580 14822 15608 14962
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15580 13818 15608 14758
rect 15672 14414 15700 15302
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15580 13790 15700 13818
rect 15568 13728 15620 13734
rect 15568 13670 15620 13676
rect 15476 13456 15528 13462
rect 15476 13398 15528 13404
rect 15200 13184 15252 13190
rect 15200 13126 15252 13132
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15212 12714 15240 13126
rect 15200 12708 15252 12714
rect 15200 12650 15252 12656
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15200 8016 15252 8022
rect 15304 7993 15332 9862
rect 15396 9625 15424 13126
rect 15488 12986 15516 13398
rect 15580 12986 15608 13670
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15568 12980 15620 12986
rect 15568 12922 15620 12928
rect 15568 12776 15620 12782
rect 15568 12718 15620 12724
rect 15580 12102 15608 12718
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15580 11762 15608 12038
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15476 10736 15528 10742
rect 15476 10678 15528 10684
rect 15382 9616 15438 9625
rect 15382 9551 15438 9560
rect 15384 8832 15436 8838
rect 15384 8774 15436 8780
rect 15200 7958 15252 7964
rect 15290 7984 15346 7993
rect 15212 7546 15240 7958
rect 15290 7919 15346 7928
rect 15200 7540 15252 7546
rect 15200 7482 15252 7488
rect 15198 7304 15254 7313
rect 15198 7239 15254 7248
rect 15212 5370 15240 7239
rect 15304 6390 15332 7919
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15292 5296 15344 5302
rect 15292 5238 15344 5244
rect 15200 5228 15252 5234
rect 15200 5170 15252 5176
rect 15212 3942 15240 5170
rect 15304 4185 15332 5238
rect 15290 4176 15346 4185
rect 15290 4111 15346 4120
rect 15292 4004 15344 4010
rect 15292 3946 15344 3952
rect 15200 3936 15252 3942
rect 15200 3878 15252 3884
rect 15200 3460 15252 3466
rect 15200 3402 15252 3408
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15108 3052 15160 3058
rect 15212 3040 15240 3402
rect 15160 3012 15240 3040
rect 15108 2994 15160 3000
rect 15120 2650 15148 2994
rect 15200 2848 15252 2854
rect 15200 2790 15252 2796
rect 15108 2644 15160 2650
rect 15108 2586 15160 2592
rect 15212 2446 15240 2790
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 14924 1692 14976 1698
rect 14924 1634 14976 1640
rect 15212 800 15240 2246
rect 15304 1834 15332 3946
rect 15396 3534 15424 8774
rect 15488 8514 15516 10678
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15580 8634 15608 8978
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15488 8486 15608 8514
rect 15474 6760 15530 6769
rect 15474 6695 15476 6704
rect 15528 6695 15530 6704
rect 15476 6666 15528 6672
rect 15580 6390 15608 8486
rect 15672 7002 15700 13790
rect 15764 13326 15792 15846
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16224 14482 16252 15438
rect 16544 15260 16852 15280
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15184 16852 15204
rect 16212 14476 16264 14482
rect 16212 14418 16264 14424
rect 16948 14408 17000 14414
rect 16316 14346 16528 14362
rect 16948 14350 17000 14356
rect 16316 14340 16540 14346
rect 16316 14334 16488 14340
rect 16316 13938 16344 14334
rect 16488 14282 16540 14288
rect 16396 14272 16448 14278
rect 16396 14214 16448 14220
rect 16408 14074 16436 14214
rect 16544 14172 16852 14192
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14096 16852 14116
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16304 13796 16356 13802
rect 16304 13738 16356 13744
rect 16316 13530 16344 13738
rect 16304 13524 16356 13530
rect 16304 13466 16356 13472
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 15752 13320 15804 13326
rect 15752 13262 15804 13268
rect 16408 12918 16436 13466
rect 16960 13326 16988 14350
rect 17052 13530 17080 19382
rect 17224 19372 17276 19378
rect 17224 19314 17276 19320
rect 17236 19174 17264 19314
rect 17420 19310 17448 19790
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 17224 19168 17276 19174
rect 17224 19110 17276 19116
rect 17408 19168 17460 19174
rect 17512 19122 17540 19790
rect 17788 19174 17816 19790
rect 18432 19718 18460 20266
rect 18800 20058 18828 20402
rect 19143 20156 19451 20176
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20080 19451 20100
rect 19720 20058 19748 20402
rect 20548 20058 20576 20402
rect 20904 20256 20956 20262
rect 20904 20198 20956 20204
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 19708 20052 19760 20058
rect 19708 19994 19760 20000
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20916 19854 20944 20198
rect 21192 20058 21220 20402
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21180 20052 21232 20058
rect 21180 19994 21232 20000
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 18420 19712 18472 19718
rect 18420 19654 18472 19660
rect 18604 19712 18656 19718
rect 18604 19654 18656 19660
rect 18512 19372 18564 19378
rect 18512 19314 18564 19320
rect 18524 19174 18552 19314
rect 17460 19116 17540 19122
rect 17408 19110 17540 19116
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16544 13084 16852 13104
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13008 16852 13028
rect 16396 12912 16448 12918
rect 16396 12854 16448 12860
rect 15752 12844 15804 12850
rect 15752 12786 15804 12792
rect 15764 11898 15792 12786
rect 16960 12170 16988 13262
rect 16948 12164 17000 12170
rect 16948 12106 17000 12112
rect 16396 12096 16448 12102
rect 16396 12038 16448 12044
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 16120 11756 16172 11762
rect 16120 11698 16172 11704
rect 16132 10810 16160 11698
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16224 10266 16252 11630
rect 16408 11082 16436 12038
rect 16544 11996 16852 12016
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11920 16852 11940
rect 16960 11830 16988 12106
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 17236 11354 17264 19110
rect 17420 19094 17540 19110
rect 17420 16182 17448 19094
rect 17788 18086 17816 19110
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 17776 18080 17828 18086
rect 17776 18022 17828 18028
rect 17408 16176 17460 16182
rect 17408 16118 17460 16124
rect 17224 11348 17276 11354
rect 17224 11290 17276 11296
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16544 10908 16852 10928
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10832 16852 10852
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 16544 9820 16852 9840
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9744 16852 9764
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16408 7886 16436 8774
rect 16544 8732 16852 8752
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8656 16852 8676
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16948 7744 17000 7750
rect 16948 7686 17000 7692
rect 16544 7644 16852 7664
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7568 16852 7588
rect 15936 7540 15988 7546
rect 15936 7482 15988 7488
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15672 6662 15700 6734
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15568 6384 15620 6390
rect 15568 6326 15620 6332
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 15488 4622 15516 6258
rect 15580 5846 15608 6326
rect 15660 6112 15712 6118
rect 15660 6054 15712 6060
rect 15672 5953 15700 6054
rect 15658 5944 15714 5953
rect 15658 5879 15714 5888
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15764 5710 15792 6802
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15752 5160 15804 5166
rect 15658 5128 15714 5137
rect 15752 5102 15804 5108
rect 15658 5063 15714 5072
rect 15672 4690 15700 5063
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15476 4616 15528 4622
rect 15476 4558 15528 4564
rect 15488 4282 15516 4558
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 15474 4176 15530 4185
rect 15474 4111 15530 4120
rect 15488 3670 15516 4111
rect 15476 3664 15528 3670
rect 15476 3606 15528 3612
rect 15384 3528 15436 3534
rect 15384 3470 15436 3476
rect 15384 3052 15436 3058
rect 15488 3040 15516 3606
rect 15580 3602 15608 4422
rect 15660 3936 15712 3942
rect 15660 3878 15712 3884
rect 15568 3596 15620 3602
rect 15568 3538 15620 3544
rect 15672 3505 15700 3878
rect 15764 3738 15792 5102
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15856 4321 15884 4422
rect 15842 4312 15898 4321
rect 15842 4247 15898 4256
rect 15948 4128 15976 7482
rect 16304 7472 16356 7478
rect 16304 7414 16356 7420
rect 16210 6760 16266 6769
rect 16210 6695 16212 6704
rect 16264 6695 16266 6704
rect 16212 6666 16264 6672
rect 16210 4448 16266 4457
rect 16210 4383 16266 4392
rect 15856 4100 15976 4128
rect 15752 3732 15804 3738
rect 15752 3674 15804 3680
rect 15856 3618 15884 4100
rect 15936 4004 15988 4010
rect 15936 3946 15988 3952
rect 15764 3590 15884 3618
rect 15658 3496 15714 3505
rect 15658 3431 15714 3440
rect 15764 3398 15792 3590
rect 15844 3528 15896 3534
rect 15844 3470 15896 3476
rect 15568 3392 15620 3398
rect 15568 3334 15620 3340
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15580 3097 15608 3334
rect 15764 3126 15792 3334
rect 15752 3120 15804 3126
rect 15436 3012 15516 3040
rect 15566 3088 15622 3097
rect 15752 3062 15804 3068
rect 15856 3058 15884 3470
rect 15566 3023 15622 3032
rect 15844 3052 15896 3058
rect 15384 2994 15436 3000
rect 15844 2994 15896 3000
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15752 2848 15804 2854
rect 15752 2790 15804 2796
rect 15580 2446 15608 2790
rect 15764 2446 15792 2790
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 15660 2304 15712 2310
rect 15660 2246 15712 2252
rect 15292 1828 15344 1834
rect 15292 1770 15344 1776
rect 15672 800 15700 2246
rect 15948 2009 15976 3946
rect 16028 3936 16080 3942
rect 16028 3878 16080 3884
rect 15934 2000 15990 2009
rect 15934 1935 15990 1944
rect 16040 1465 16068 3878
rect 16120 3732 16172 3738
rect 16120 3674 16172 3680
rect 16132 3058 16160 3674
rect 16224 3466 16252 4383
rect 16316 4078 16344 7414
rect 16396 7200 16448 7206
rect 16396 7142 16448 7148
rect 16408 6458 16436 7142
rect 16544 6556 16852 6576
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6480 16852 6500
rect 16396 6452 16448 6458
rect 16396 6394 16448 6400
rect 16960 6202 16988 7686
rect 16868 6174 16988 6202
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 16868 5642 16896 6174
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16856 5636 16908 5642
rect 16856 5578 16908 5584
rect 16544 5468 16852 5488
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5392 16852 5412
rect 16672 5024 16724 5030
rect 16394 4992 16450 5001
rect 16672 4966 16724 4972
rect 16394 4927 16450 4936
rect 16304 4072 16356 4078
rect 16304 4014 16356 4020
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16212 3460 16264 3466
rect 16212 3402 16264 3408
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 16212 2848 16264 2854
rect 16212 2790 16264 2796
rect 16224 2446 16252 2790
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16026 1456 16082 1465
rect 16026 1391 16082 1400
rect 16132 800 16160 2246
rect 16316 1601 16344 3878
rect 16408 3738 16436 4927
rect 16684 4690 16712 4966
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16960 4622 16988 6054
rect 17236 5930 17264 6190
rect 17144 5902 17264 5930
rect 17144 5846 17172 5902
rect 17132 5840 17184 5846
rect 17132 5782 17184 5788
rect 17222 5808 17278 5817
rect 17040 5704 17092 5710
rect 17040 5646 17092 5652
rect 17052 5302 17080 5646
rect 17144 5302 17172 5782
rect 17222 5743 17278 5752
rect 17236 5574 17264 5743
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 17132 5296 17184 5302
rect 17132 5238 17184 5244
rect 17788 5166 17816 9046
rect 17868 5636 17920 5642
rect 17868 5578 17920 5584
rect 17880 5234 17908 5578
rect 17972 5302 18000 18634
rect 18524 11558 18552 19110
rect 18616 16017 18644 19654
rect 18602 16008 18658 16017
rect 18602 15943 18658 15952
rect 19076 14618 19104 19790
rect 19628 19514 19656 19790
rect 19616 19508 19668 19514
rect 19616 19450 19668 19456
rect 19143 19068 19451 19088
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 18992 19451 19012
rect 19143 17980 19451 18000
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17904 19451 17924
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 21100 17105 21128 17478
rect 21086 17096 21142 17105
rect 21086 17031 21142 17040
rect 19143 16892 19451 16912
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16816 19451 16836
rect 19143 15804 19451 15824
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15728 19451 15748
rect 19143 14716 19451 14736
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14640 19451 14660
rect 19064 14612 19116 14618
rect 19064 14554 19116 14560
rect 21376 13938 21404 20198
rect 21468 20058 21496 20998
rect 21456 20052 21508 20058
rect 21456 19994 21508 20000
rect 21836 19990 21864 22200
rect 21824 19984 21876 19990
rect 21824 19926 21876 19932
rect 22296 19310 22324 22200
rect 22756 20466 22784 22200
rect 22744 20460 22796 20466
rect 22744 20402 22796 20408
rect 22284 19304 22336 19310
rect 22284 19246 22336 19252
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21468 17241 21496 17478
rect 21454 17232 21510 17241
rect 21454 17167 21510 17176
rect 21364 13932 21416 13938
rect 21364 13874 21416 13880
rect 19143 13628 19451 13648
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13552 19451 13572
rect 21364 13252 21416 13258
rect 21364 13194 21416 13200
rect 19143 12540 19451 12560
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12464 19451 12484
rect 18512 11552 18564 11558
rect 18512 11494 18564 11500
rect 19143 11452 19451 11472
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11376 19451 11396
rect 19143 10364 19451 10384
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10288 19451 10308
rect 19143 9276 19451 9296
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9200 19451 9220
rect 19143 8188 19451 8208
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8112 19451 8132
rect 19143 7100 19451 7120
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7024 19451 7044
rect 21376 6458 21404 13194
rect 21364 6452 21416 6458
rect 21364 6394 21416 6400
rect 18052 6316 18104 6322
rect 18052 6258 18104 6264
rect 21548 6316 21600 6322
rect 21548 6258 21600 6264
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 17868 5228 17920 5234
rect 17868 5170 17920 5176
rect 17776 5160 17828 5166
rect 17776 5102 17828 5108
rect 16948 4616 17000 4622
rect 16948 4558 17000 4564
rect 17788 4554 17816 5102
rect 17972 4690 18000 5238
rect 18064 5030 18092 6258
rect 18786 6216 18842 6225
rect 18236 6180 18288 6186
rect 18786 6151 18842 6160
rect 18236 6122 18288 6128
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 18064 4826 18092 4966
rect 18052 4820 18104 4826
rect 18052 4762 18104 4768
rect 18144 4752 18196 4758
rect 18144 4694 18196 4700
rect 17960 4684 18012 4690
rect 18012 4644 18092 4672
rect 17960 4626 18012 4632
rect 17776 4548 17828 4554
rect 17776 4490 17828 4496
rect 16544 4380 16852 4400
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4304 16852 4324
rect 16488 4072 16540 4078
rect 16488 4014 16540 4020
rect 16500 3890 16528 4014
rect 16672 3936 16724 3942
rect 16500 3862 16620 3890
rect 16672 3878 16724 3884
rect 16592 3738 16620 3862
rect 16396 3732 16448 3738
rect 16580 3732 16632 3738
rect 16448 3692 16528 3720
rect 16396 3674 16448 3680
rect 16396 3596 16448 3602
rect 16396 3538 16448 3544
rect 16408 3058 16436 3538
rect 16500 3534 16528 3692
rect 16580 3674 16632 3680
rect 16684 3641 16712 3878
rect 17788 3738 17816 4490
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 17972 3738 18000 4150
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 17500 3732 17552 3738
rect 17500 3674 17552 3680
rect 17776 3732 17828 3738
rect 17776 3674 17828 3680
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 16670 3632 16726 3641
rect 16670 3567 16726 3576
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16544 3292 16852 3312
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3216 16852 3236
rect 16396 3052 16448 3058
rect 16396 2994 16448 3000
rect 16764 2848 16816 2854
rect 16684 2808 16764 2836
rect 16684 2446 16712 2808
rect 16764 2790 16816 2796
rect 16672 2440 16724 2446
rect 16960 2417 16988 3334
rect 17038 3088 17094 3097
rect 17236 3058 17264 3674
rect 17512 3058 17540 3674
rect 18064 3194 18092 4644
rect 18156 3534 18184 4694
rect 18248 3602 18276 6122
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18708 5642 18736 6054
rect 18696 5636 18748 5642
rect 18696 5578 18748 5584
rect 18602 5264 18658 5273
rect 18602 5199 18658 5208
rect 18236 3596 18288 3602
rect 18236 3538 18288 3544
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18052 3188 18104 3194
rect 18052 3130 18104 3136
rect 17038 3023 17040 3032
rect 17092 3023 17094 3032
rect 17224 3052 17276 3058
rect 17040 2994 17092 3000
rect 17224 2994 17276 3000
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17960 3052 18012 3058
rect 18064 3040 18092 3130
rect 18248 3058 18276 3538
rect 18616 3194 18644 5199
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18616 3058 18644 3130
rect 18800 3058 18828 6151
rect 19143 6012 19451 6032
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5936 19451 5956
rect 21560 5817 21588 6258
rect 21546 5808 21602 5817
rect 21546 5743 21602 5752
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19996 5234 20024 5510
rect 19984 5228 20036 5234
rect 19984 5170 20036 5176
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 19143 4924 19451 4944
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4848 19451 4868
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 19143 3836 19451 3856
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3760 19451 3780
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19064 3392 19116 3398
rect 19064 3334 19116 3340
rect 18012 3012 18092 3040
rect 18236 3052 18288 3058
rect 17960 2994 18012 3000
rect 18236 2994 18288 3000
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 18788 3052 18840 3058
rect 18788 2994 18840 3000
rect 17500 2916 17552 2922
rect 17500 2858 17552 2864
rect 17132 2848 17184 2854
rect 17132 2790 17184 2796
rect 17144 2446 17172 2790
rect 17512 2774 17540 2858
rect 17776 2848 17828 2854
rect 17696 2808 17776 2836
rect 17512 2746 17632 2774
rect 17604 2446 17632 2746
rect 17696 2446 17724 2808
rect 17776 2790 17828 2796
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 18248 2446 18276 2790
rect 19076 2446 19104 3334
rect 19536 3058 19564 3402
rect 20272 3194 20300 4082
rect 19984 3188 20036 3194
rect 19984 3130 20036 3136
rect 20260 3188 20312 3194
rect 20260 3130 20312 3136
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19616 2916 19668 2922
rect 19616 2858 19668 2864
rect 19143 2748 19451 2768
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2672 19451 2692
rect 19628 2446 19656 2858
rect 19996 2446 20024 3130
rect 20272 3058 20300 3130
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 20444 2916 20496 2922
rect 20444 2858 20496 2864
rect 20456 2446 20484 2858
rect 20916 2446 20944 4966
rect 22652 3528 22704 3534
rect 22652 3470 22704 3476
rect 22192 2916 22244 2922
rect 22192 2858 22244 2864
rect 20996 2848 21048 2854
rect 20996 2790 21048 2796
rect 21732 2848 21784 2854
rect 21732 2790 21784 2796
rect 21008 2446 21036 2790
rect 17132 2440 17184 2446
rect 16672 2382 16724 2388
rect 16946 2408 17002 2417
rect 17132 2382 17184 2388
rect 17592 2440 17644 2446
rect 17592 2382 17644 2388
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 18236 2440 18288 2446
rect 18236 2382 18288 2388
rect 19064 2440 19116 2446
rect 19064 2382 19116 2388
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 20444 2440 20496 2446
rect 20444 2382 20496 2388
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 20996 2440 21048 2446
rect 20996 2382 21048 2388
rect 16946 2343 17002 2352
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 17500 2304 17552 2310
rect 17500 2246 17552 2252
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 18420 2304 18472 2310
rect 18420 2246 18472 2252
rect 18972 2304 19024 2310
rect 19524 2304 19576 2310
rect 18972 2246 19024 2252
rect 19444 2264 19524 2292
rect 16544 2204 16852 2224
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2128 16852 2148
rect 16302 1592 16358 1601
rect 16302 1527 16358 1536
rect 16592 870 16712 898
rect 16592 800 16620 870
rect 10612 734 10824 762
rect 10966 0 11022 800
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13266 0 13322 800
rect 13726 0 13782 800
rect 14278 0 14334 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16578 0 16634 800
rect 16684 762 16712 870
rect 16960 762 16988 2246
rect 17052 800 17080 2246
rect 17512 800 17540 2246
rect 17972 800 18000 2246
rect 18432 800 18460 2246
rect 18984 800 19012 2246
rect 19444 800 19472 2264
rect 19524 2246 19576 2252
rect 19892 2304 19944 2310
rect 19892 2246 19944 2252
rect 20352 2304 20404 2310
rect 20352 2246 20404 2252
rect 20812 2304 20864 2310
rect 20812 2246 20864 2252
rect 21272 2304 21324 2310
rect 21272 2246 21324 2252
rect 19904 800 19932 2246
rect 20364 800 20392 2246
rect 20824 800 20852 2246
rect 21284 800 21312 2246
rect 21744 800 21772 2790
rect 22204 800 22232 2858
rect 22664 800 22692 3470
rect 16684 734 16988 762
rect 17038 0 17094 800
rect 17498 0 17554 800
rect 17958 0 18014 800
rect 18418 0 18474 800
rect 18970 0 19026 800
rect 19430 0 19486 800
rect 19890 0 19946 800
rect 20350 0 20406 800
rect 20810 0 20866 800
rect 21270 0 21326 800
rect 21730 0 21786 800
rect 22190 0 22246 800
rect 22650 0 22706 800
<< via2 >>
rect 2318 22616 2374 22672
rect 662 20440 718 20496
rect 1490 21120 1546 21176
rect 1214 19216 1270 19272
rect 1490 17856 1546 17912
rect 1490 17312 1546 17368
rect 1950 19352 2006 19408
rect 1858 18808 1914 18864
rect 1766 18536 1822 18592
rect 2226 18808 2282 18864
rect 2134 18672 2190 18728
rect 1490 16940 1492 16960
rect 1492 16940 1544 16960
rect 1544 16940 1546 16960
rect 1490 16904 1546 16940
rect 2042 17720 2098 17776
rect 1950 17584 2006 17640
rect 1490 16396 1492 16416
rect 1492 16396 1544 16416
rect 1544 16396 1546 16416
rect 1490 16360 1546 16396
rect 1490 15972 1546 16008
rect 1490 15952 1492 15972
rect 1492 15952 1544 15972
rect 1544 15952 1546 15972
rect 2226 18264 2282 18320
rect 2318 17176 2374 17232
rect 2778 22072 2834 22128
rect 2594 19760 2650 19816
rect 2410 16360 2466 16416
rect 1858 15408 1914 15464
rect 1490 15000 1546 15056
rect 1490 14456 1546 14512
rect 1490 14048 1546 14104
rect 1490 13504 1546 13560
rect 1582 13232 1638 13288
rect 1398 13096 1454 13152
rect 1398 12552 1454 12608
rect 1122 5480 1178 5536
rect 202 2760 258 2816
rect 1490 12180 1492 12200
rect 1492 12180 1544 12200
rect 1544 12180 1546 12200
rect 1490 12144 1546 12180
rect 1398 11056 1454 11112
rect 1674 11600 1730 11656
rect 1582 11056 1638 11112
rect 1674 10668 1730 10704
rect 1674 10648 1676 10668
rect 1676 10648 1728 10668
rect 1728 10648 1730 10668
rect 1398 9152 1454 9208
rect 1398 8336 1454 8392
rect 1582 8880 1638 8936
rect 1858 11736 1914 11792
rect 2686 19352 2742 19408
rect 2870 21664 2926 21720
rect 3238 20440 3294 20496
rect 3054 20168 3110 20224
rect 2778 17856 2834 17912
rect 2778 16632 2834 16688
rect 2686 16496 2742 16552
rect 2686 16396 2688 16416
rect 2688 16396 2740 16416
rect 2740 16396 2742 16416
rect 2686 16360 2742 16396
rect 3422 20712 3478 20768
rect 3514 20304 3570 20360
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3514 19896 3570 19952
rect 3698 19352 3754 19408
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3330 18128 3386 18184
rect 4066 20440 4122 20496
rect 3974 20204 3976 20224
rect 3976 20204 4028 20224
rect 4028 20204 4030 20224
rect 3974 20168 4030 20204
rect 4066 19760 4122 19816
rect 3238 17856 3294 17912
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 2962 17312 3018 17368
rect 2686 16108 2742 16144
rect 2686 16088 2688 16108
rect 2688 16088 2740 16108
rect 2740 16088 2742 16108
rect 2042 11192 2098 11248
rect 1858 10104 1914 10160
rect 2134 10532 2190 10568
rect 2134 10512 2136 10532
rect 2136 10512 2188 10532
rect 2188 10512 2190 10532
rect 2042 10104 2098 10160
rect 1674 8200 1730 8256
rect 1674 7248 1730 7304
rect 2042 9560 2098 9616
rect 1398 6568 1454 6624
rect 1766 6860 1822 6896
rect 1766 6840 1768 6860
rect 1768 6840 1820 6860
rect 1820 6840 1822 6860
rect 1950 7792 2006 7848
rect 1674 6296 1730 6352
rect 1398 5888 1454 5944
rect 1214 3304 1270 3360
rect 1490 5636 1546 5672
rect 1490 5616 1492 5636
rect 1492 5616 1544 5636
rect 1544 5616 1546 5636
rect 1582 5072 1638 5128
rect 2318 6432 2374 6488
rect 1490 3440 1546 3496
rect 1674 3732 1730 3768
rect 1674 3712 1676 3732
rect 1676 3712 1728 3732
rect 1728 3712 1730 3732
rect 1398 1944 1454 2000
rect 2042 4820 2098 4856
rect 2042 4800 2044 4820
rect 2044 4800 2096 4820
rect 2096 4800 2098 4820
rect 2042 4528 2098 4584
rect 2502 7384 2558 7440
rect 3146 15952 3202 16008
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 4250 19352 4306 19408
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3514 15564 3570 15600
rect 3514 15544 3516 15564
rect 3516 15544 3568 15564
rect 3568 15544 3570 15564
rect 4250 18128 4306 18184
rect 5170 20476 5172 20496
rect 5172 20476 5224 20496
rect 5224 20476 5226 20496
rect 5170 20440 5226 20476
rect 4434 18264 4490 18320
rect 4802 19488 4858 19544
rect 4618 19080 4674 19136
rect 4618 17856 4674 17912
rect 4250 15544 4306 15600
rect 3146 14320 3202 14376
rect 3514 14884 3570 14920
rect 3514 14864 3516 14884
rect 3516 14864 3568 14884
rect 3568 14864 3570 14884
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3882 14320 3938 14376
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 2778 9696 2834 9752
rect 2962 8744 3018 8800
rect 2686 7656 2742 7712
rect 3974 10920 4030 10976
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3606 9968 3662 10024
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3514 7792 3570 7848
rect 2778 5344 2834 5400
rect 2410 4276 2466 4312
rect 2410 4256 2412 4276
rect 2412 4256 2464 4276
rect 2464 4256 2466 4276
rect 2226 3848 2282 3904
rect 1858 3032 1914 3088
rect 2226 3440 2282 3496
rect 2226 2760 2282 2816
rect 2778 5208 2834 5264
rect 2686 4664 2742 4720
rect 3974 8336 4030 8392
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3054 5752 3110 5808
rect 2778 4392 2834 4448
rect 2870 3984 2926 4040
rect 3146 4140 3202 4176
rect 3146 4120 3148 4140
rect 3148 4120 3200 4140
rect 3200 4120 3202 4140
rect 1490 1128 1546 1184
rect 2870 2488 2926 2544
rect 3238 2932 3240 2952
rect 3240 2932 3292 2952
rect 3292 2932 3294 2952
rect 3238 2896 3294 2932
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3514 5344 3570 5400
rect 3606 5208 3662 5264
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3974 6568 4030 6624
rect 4158 8336 4214 8392
rect 4250 7692 4252 7712
rect 4252 7692 4304 7712
rect 4304 7692 4306 7712
rect 4250 7656 4306 7692
rect 3422 4528 3478 4584
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3422 3032 3478 3088
rect 3054 2488 3110 2544
rect 3146 2388 3148 2408
rect 3148 2388 3200 2408
rect 3200 2388 3202 2408
rect 3146 2352 3202 2388
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 3422 2372 3478 2408
rect 3422 2352 3424 2372
rect 3424 2352 3476 2372
rect 3476 2352 3478 2372
rect 3146 1808 3202 1864
rect 3238 1672 3294 1728
rect 3054 1536 3110 1592
rect 2962 1400 3018 1456
rect 3422 1808 3478 1864
rect 4802 17060 4858 17096
rect 4802 17040 4804 17060
rect 4804 17040 4856 17060
rect 4856 17040 4858 17060
rect 5446 19896 5502 19952
rect 5262 19216 5318 19272
rect 5170 15408 5226 15464
rect 4802 11600 4858 11656
rect 4710 11500 4712 11520
rect 4712 11500 4764 11520
rect 4764 11500 4766 11520
rect 4710 11464 4766 11500
rect 4250 6704 4306 6760
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 5722 20032 5778 20088
rect 5722 17312 5778 17368
rect 5446 15000 5502 15056
rect 4986 11736 5042 11792
rect 4894 9288 4950 9344
rect 6550 20304 6606 20360
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 6182 19236 6238 19272
rect 6182 19216 6184 19236
rect 6184 19216 6236 19236
rect 6236 19216 6238 19236
rect 6826 20440 6882 20496
rect 6734 20032 6790 20088
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6550 17856 6606 17912
rect 6918 18944 6974 19000
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6274 16496 6330 16552
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 7102 18536 7158 18592
rect 6826 16632 6882 16688
rect 5446 12416 5502 12472
rect 5630 12280 5686 12336
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 7102 17992 7158 18048
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 5262 9324 5264 9344
rect 5264 9324 5316 9344
rect 5316 9324 5318 9344
rect 5262 9288 5318 9324
rect 4250 6160 4306 6216
rect 4526 6024 4582 6080
rect 4434 5228 4490 5264
rect 4434 5208 4436 5228
rect 4436 5208 4488 5228
rect 4488 5208 4490 5228
rect 4158 4528 4214 4584
rect 4066 3984 4122 4040
rect 3974 2644 4030 2680
rect 3974 2624 3976 2644
rect 3976 2624 4028 2644
rect 4028 2624 4030 2644
rect 4618 5072 4674 5128
rect 4618 4936 4674 4992
rect 4802 7248 4858 7304
rect 5170 8336 5226 8392
rect 4986 6704 5042 6760
rect 4894 6432 4950 6488
rect 4986 5888 5042 5944
rect 4894 5772 4950 5808
rect 4894 5752 4896 5772
rect 4896 5752 4948 5772
rect 4948 5752 4950 5772
rect 4802 5344 4858 5400
rect 4894 3440 4950 3496
rect 4802 3304 4858 3360
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 7562 18808 7618 18864
rect 7562 18264 7618 18320
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8114 16088 8170 16144
rect 7654 15952 7710 16008
rect 7562 13368 7618 13424
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 5630 9968 5686 10024
rect 6826 11056 6882 11112
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 5998 9560 6054 9616
rect 5538 7112 5594 7168
rect 5354 6568 5410 6624
rect 5262 6024 5318 6080
rect 5262 5888 5318 5944
rect 5170 5072 5226 5128
rect 6090 9016 6146 9072
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6550 7692 6552 7712
rect 6552 7692 6604 7712
rect 6604 7692 6606 7712
rect 6550 7656 6606 7692
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 5814 5480 5870 5536
rect 5262 4256 5318 4312
rect 3330 584 3386 640
rect 4066 176 4122 232
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 7010 9288 7066 9344
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 9586 19896 9642 19952
rect 9586 19352 9642 19408
rect 9494 18536 9550 18592
rect 9494 17992 9550 18048
rect 8758 16652 8814 16688
rect 8758 16632 8760 16652
rect 8760 16632 8812 16652
rect 8812 16632 8814 16652
rect 9126 15952 9182 16008
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 9034 15408 9090 15464
rect 8758 15000 8814 15056
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 9310 17176 9366 17232
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 6734 7520 6790 7576
rect 6734 7248 6790 7304
rect 6826 7112 6882 7168
rect 6734 6568 6790 6624
rect 5630 3712 5686 3768
rect 5630 3168 5686 3224
rect 5538 2624 5594 2680
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6458 5072 6514 5128
rect 6274 4800 6330 4856
rect 5814 4120 5870 4176
rect 5906 3848 5962 3904
rect 6550 4428 6552 4448
rect 6552 4428 6604 4448
rect 6604 4428 6606 4448
rect 6550 4392 6606 4428
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6550 4120 6606 4176
rect 6734 5888 6790 5944
rect 7194 6432 7250 6488
rect 6366 3848 6422 3904
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 5998 3168 6054 3224
rect 7286 5072 7342 5128
rect 7194 4528 7250 4584
rect 6918 3712 6974 3768
rect 5906 3032 5962 3088
rect 6090 2896 6146 2952
rect 6458 2644 6514 2680
rect 6458 2624 6460 2644
rect 6460 2624 6512 2644
rect 6512 2624 6514 2644
rect 5814 1672 5870 1728
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 6826 3188 6882 3224
rect 6826 3168 6828 3188
rect 6828 3168 6880 3188
rect 6880 3168 6882 3188
rect 7470 3984 7526 4040
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 9218 11736 9274 11792
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 9126 10104 9182 10160
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8482 8780 8484 8800
rect 8484 8780 8536 8800
rect 8536 8780 8538 8800
rect 8482 8744 8538 8780
rect 9218 8608 9274 8664
rect 9954 18944 10010 19000
rect 9954 18400 10010 18456
rect 10046 17584 10102 17640
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 10230 18808 10286 18864
rect 9862 14456 9918 14512
rect 9678 13912 9734 13968
rect 9494 11192 9550 11248
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 10506 17720 10562 17776
rect 10230 14864 10286 14920
rect 10782 12316 10784 12336
rect 10784 12316 10836 12336
rect 10836 12316 10838 12336
rect 10782 12280 10838 12316
rect 9402 9696 9458 9752
rect 9402 8608 9458 8664
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 7930 6432 7986 6488
rect 8298 7248 8354 7304
rect 8206 6976 8262 7032
rect 8390 7112 8446 7168
rect 9310 8064 9366 8120
rect 9310 7384 9366 7440
rect 9126 7112 9182 7168
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 9126 6996 9182 7032
rect 9126 6976 9128 6996
rect 9128 6976 9180 6996
rect 9180 6976 9182 6996
rect 8298 6296 8354 6352
rect 8850 6432 8906 6488
rect 8942 6296 8998 6352
rect 8298 5108 8300 5128
rect 8300 5108 8352 5128
rect 8352 5108 8354 5128
rect 8298 5072 8354 5108
rect 7838 3440 7894 3496
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8482 4256 8538 4312
rect 8482 3304 8538 3360
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 9770 7656 9826 7712
rect 9310 6432 9366 6488
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 9954 7112 10010 7168
rect 10046 6160 10102 6216
rect 9770 5208 9826 5264
rect 9678 4428 9680 4448
rect 9680 4428 9732 4448
rect 9732 4428 9734 4448
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9218 2760 9274 2816
rect 9402 2644 9458 2680
rect 9402 2624 9404 2644
rect 9404 2624 9456 2644
rect 9456 2624 9458 2644
rect 9678 4392 9734 4428
rect 9954 5228 10010 5264
rect 9954 5208 9956 5228
rect 9956 5208 10008 5228
rect 10008 5208 10010 5228
rect 9862 5072 9918 5128
rect 10138 3712 10194 3768
rect 10506 6704 10562 6760
rect 10506 6024 10562 6080
rect 10414 5364 10470 5400
rect 10414 5344 10416 5364
rect 10416 5344 10468 5364
rect 10468 5344 10470 5364
rect 10414 4936 10470 4992
rect 10046 2760 10102 2816
rect 10230 2624 10286 2680
rect 11610 18828 11666 18864
rect 11610 18808 11612 18828
rect 11612 18808 11664 18828
rect 11664 18808 11666 18828
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11794 18808 11850 18864
rect 11610 18128 11666 18184
rect 11794 17992 11850 18048
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 12254 17856 12310 17912
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11242 11600 11298 11656
rect 10966 11192 11022 11248
rect 11058 7792 11114 7848
rect 10690 4428 10692 4448
rect 10692 4428 10744 4448
rect 10744 4428 10746 4448
rect 10690 4392 10746 4428
rect 10782 3984 10838 4040
rect 11518 11328 11574 11384
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11886 12280 11942 12336
rect 13082 19372 13138 19408
rect 13082 19352 13084 19372
rect 13084 19352 13136 19372
rect 13136 19352 13138 19372
rect 12162 14184 12218 14240
rect 12530 16632 12586 16688
rect 12622 13912 12678 13968
rect 13450 19080 13506 19136
rect 13266 18300 13268 18320
rect 13268 18300 13320 18320
rect 13320 18300 13322 18320
rect 13266 18264 13322 18300
rect 13634 18964 13690 19000
rect 13634 18944 13636 18964
rect 13636 18944 13688 18964
rect 13688 18944 13690 18964
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 14646 20304 14702 20360
rect 14462 19624 14518 19680
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13910 18844 13912 18864
rect 13912 18844 13964 18864
rect 13964 18844 13966 18864
rect 13910 18808 13966 18844
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 12346 11328 12402 11384
rect 12530 11328 12586 11384
rect 13358 13232 13414 13288
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 11702 9968 11758 10024
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11794 8372 11796 8392
rect 11796 8372 11848 8392
rect 11848 8372 11850 8392
rect 11794 8336 11850 8372
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11886 6976 11942 7032
rect 11058 5480 11114 5536
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 10874 3440 10930 3496
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11518 3712 11574 3768
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11334 2760 11390 2816
rect 13174 11192 13230 11248
rect 13358 10512 13414 10568
rect 12990 8472 13046 8528
rect 12990 7928 13046 7984
rect 12530 7792 12586 7848
rect 11978 6704 12034 6760
rect 11886 5752 11942 5808
rect 11886 4800 11942 4856
rect 11886 4120 11942 4176
rect 11886 3168 11942 3224
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12346 7112 12402 7168
rect 12254 5228 12310 5264
rect 12254 5208 12256 5228
rect 12256 5208 12308 5228
rect 12308 5208 12310 5228
rect 12806 6860 12862 6896
rect 12806 6840 12808 6860
rect 12808 6840 12860 6860
rect 12860 6840 12862 6860
rect 13450 8916 13452 8936
rect 13452 8916 13504 8936
rect 13504 8916 13506 8936
rect 13450 8880 13506 8916
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 14830 18692 14886 18728
rect 14830 18672 14832 18692
rect 14832 18672 14884 18692
rect 14884 18672 14886 18692
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 12530 4564 12532 4584
rect 12532 4564 12584 4584
rect 12584 4564 12586 4584
rect 12530 4528 12586 4564
rect 12806 5208 12862 5264
rect 12806 4800 12862 4856
rect 12438 4428 12440 4448
rect 12440 4428 12492 4448
rect 12492 4428 12494 4448
rect 12438 4392 12494 4428
rect 12254 3032 12310 3088
rect 13174 5616 13230 5672
rect 12990 4800 13046 4856
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 15014 11736 15070 11792
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 14462 5888 14518 5944
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13910 4700 13912 4720
rect 13912 4700 13964 4720
rect 13964 4700 13966 4720
rect 13910 4664 13966 4700
rect 11702 1808 11758 1864
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 14186 3340 14188 3360
rect 14188 3340 14240 3360
rect 14240 3340 14242 3360
rect 14186 3304 14242 3340
rect 13726 2896 13782 2952
rect 13450 1672 13506 1728
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 15014 4020 15016 4040
rect 15016 4020 15068 4040
rect 15068 4020 15070 4040
rect 15014 3984 15070 4020
rect 16578 19780 16634 19816
rect 16578 19760 16580 19780
rect 16580 19760 16632 19780
rect 16632 19760 16634 19780
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 15474 19236 15530 19272
rect 15474 19216 15476 19236
rect 15476 19216 15528 19236
rect 15528 19216 15530 19236
rect 15658 18672 15714 18728
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 15382 9560 15438 9616
rect 15290 7928 15346 7984
rect 15198 7248 15254 7304
rect 15290 4120 15346 4176
rect 15474 6724 15530 6760
rect 15474 6704 15476 6724
rect 15476 6704 15528 6724
rect 15528 6704 15530 6724
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 15658 5888 15714 5944
rect 15658 5072 15714 5128
rect 15474 4120 15530 4176
rect 15842 4256 15898 4312
rect 16210 6724 16266 6760
rect 16210 6704 16212 6724
rect 16212 6704 16264 6724
rect 16264 6704 16266 6724
rect 16210 4392 16266 4448
rect 15658 3440 15714 3496
rect 15566 3032 15622 3088
rect 15934 1944 15990 2000
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16394 4936 16450 4992
rect 16026 1400 16082 1456
rect 17222 5752 17278 5808
rect 18602 15952 18658 16008
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 21086 17040 21142 17096
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 21454 17176 21510 17232
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 18786 6160 18842 6216
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16670 3576 16726 3632
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 17038 3052 17094 3088
rect 18602 5208 18658 5264
rect 17038 3032 17040 3052
rect 17040 3032 17092 3052
rect 17092 3032 17094 3052
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 21546 5752 21602 5808
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 16946 2352 17002 2408
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 16302 1536 16358 1592
<< metal3 >>
rect 0 22674 800 22704
rect 2313 22674 2379 22677
rect 0 22672 2379 22674
rect 0 22616 2318 22672
rect 2374 22616 2379 22672
rect 0 22614 2379 22616
rect 0 22584 800 22614
rect 2313 22611 2379 22614
rect 0 22130 800 22160
rect 2773 22130 2839 22133
rect 0 22128 2839 22130
rect 0 22072 2778 22128
rect 2834 22072 2839 22128
rect 0 22070 2839 22072
rect 0 22040 800 22070
rect 2773 22067 2839 22070
rect 0 21722 800 21752
rect 2865 21722 2931 21725
rect 0 21720 2931 21722
rect 0 21664 2870 21720
rect 2926 21664 2931 21720
rect 0 21662 2931 21664
rect 0 21632 800 21662
rect 2865 21659 2931 21662
rect 0 21178 800 21208
rect 1485 21178 1551 21181
rect 0 21176 1551 21178
rect 0 21120 1490 21176
rect 1546 21120 1551 21176
rect 0 21118 1551 21120
rect 0 21088 800 21118
rect 1485 21115 1551 21118
rect 0 20770 800 20800
rect 3417 20770 3483 20773
rect 0 20768 3483 20770
rect 0 20712 3422 20768
rect 3478 20712 3483 20768
rect 0 20710 3483 20712
rect 0 20680 800 20710
rect 3417 20707 3483 20710
rect 6142 20704 6462 20705
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 20639 6462 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 16538 20704 16858 20705
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 20639 16858 20640
rect 657 20498 723 20501
rect 3233 20498 3299 20501
rect 4061 20498 4127 20501
rect 657 20496 4127 20498
rect 657 20440 662 20496
rect 718 20440 3238 20496
rect 3294 20440 4066 20496
rect 4122 20440 4127 20496
rect 657 20438 4127 20440
rect 657 20435 723 20438
rect 3233 20435 3299 20438
rect 4061 20435 4127 20438
rect 5165 20498 5231 20501
rect 6821 20498 6887 20501
rect 5165 20496 6887 20498
rect 5165 20440 5170 20496
rect 5226 20440 6826 20496
rect 6882 20440 6887 20496
rect 5165 20438 6887 20440
rect 5165 20435 5231 20438
rect 6821 20435 6887 20438
rect 3509 20362 3575 20365
rect 6545 20362 6611 20365
rect 14641 20362 14707 20365
rect 3509 20360 14707 20362
rect 3509 20304 3514 20360
rect 3570 20304 6550 20360
rect 6606 20304 14646 20360
rect 14702 20304 14707 20360
rect 3509 20302 14707 20304
rect 3509 20299 3575 20302
rect 6545 20299 6611 20302
rect 14641 20299 14707 20302
rect 0 20226 800 20256
rect 3049 20226 3115 20229
rect 0 20224 3115 20226
rect 0 20168 3054 20224
rect 3110 20168 3115 20224
rect 0 20166 3115 20168
rect 0 20136 800 20166
rect 3049 20163 3115 20166
rect 3969 20226 4035 20229
rect 7414 20226 7420 20228
rect 3969 20224 7420 20226
rect 3969 20168 3974 20224
rect 4030 20168 7420 20224
rect 3969 20166 7420 20168
rect 3969 20163 4035 20166
rect 7414 20164 7420 20166
rect 7484 20164 7490 20228
rect 3543 20160 3863 20161
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 20095 3863 20096
rect 8741 20160 9061 20161
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 20095 9061 20096
rect 13939 20160 14259 20161
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 20095 14259 20096
rect 19137 20160 19457 20161
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 20095 19457 20096
rect 5717 20090 5783 20093
rect 6729 20090 6795 20093
rect 3926 20088 6795 20090
rect 3926 20032 5722 20088
rect 5778 20032 6734 20088
rect 6790 20032 6795 20088
rect 3926 20030 6795 20032
rect 3509 19954 3575 19957
rect 3926 19954 3986 20030
rect 5717 20027 5783 20030
rect 6729 20027 6795 20030
rect 3509 19952 3986 19954
rect 3509 19896 3514 19952
rect 3570 19896 3986 19952
rect 3509 19894 3986 19896
rect 5441 19954 5507 19957
rect 9581 19954 9647 19957
rect 5441 19952 9647 19954
rect 5441 19896 5446 19952
rect 5502 19896 9586 19952
rect 9642 19896 9647 19952
rect 5441 19894 9647 19896
rect 3509 19891 3575 19894
rect 5441 19891 5507 19894
rect 9581 19891 9647 19894
rect 0 19818 800 19848
rect 2589 19818 2655 19821
rect 0 19816 2655 19818
rect 0 19760 2594 19816
rect 2650 19760 2655 19816
rect 0 19758 2655 19760
rect 0 19728 800 19758
rect 2589 19755 2655 19758
rect 4061 19818 4127 19821
rect 4061 19816 12450 19818
rect 4061 19760 4066 19816
rect 4122 19760 12450 19816
rect 4061 19758 12450 19760
rect 4061 19755 4127 19758
rect 12390 19682 12450 19758
rect 12934 19756 12940 19820
rect 13004 19818 13010 19820
rect 16573 19818 16639 19821
rect 13004 19816 16639 19818
rect 13004 19760 16578 19816
rect 16634 19760 16639 19816
rect 13004 19758 16639 19760
rect 13004 19756 13010 19758
rect 16573 19755 16639 19758
rect 14457 19682 14523 19685
rect 12390 19680 14523 19682
rect 12390 19624 14462 19680
rect 14518 19624 14523 19680
rect 12390 19622 14523 19624
rect 14457 19619 14523 19622
rect 6142 19616 6462 19617
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 19551 6462 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 16538 19616 16858 19617
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 19551 16858 19552
rect 1894 19484 1900 19548
rect 1964 19546 1970 19548
rect 4797 19546 4863 19549
rect 1964 19544 4863 19546
rect 1964 19488 4802 19544
rect 4858 19488 4863 19544
rect 1964 19486 4863 19488
rect 1964 19484 1970 19486
rect 4797 19483 4863 19486
rect 1710 19348 1716 19412
rect 1780 19410 1786 19412
rect 1945 19410 2011 19413
rect 2681 19412 2747 19413
rect 2630 19410 2636 19412
rect 1780 19408 2011 19410
rect 1780 19352 1950 19408
rect 2006 19352 2011 19408
rect 1780 19350 2011 19352
rect 2590 19350 2636 19410
rect 2700 19408 2747 19412
rect 2742 19352 2747 19408
rect 1780 19348 1786 19350
rect 1945 19347 2011 19350
rect 2630 19348 2636 19350
rect 2700 19348 2747 19352
rect 2681 19347 2747 19348
rect 3693 19410 3759 19413
rect 4102 19410 4108 19412
rect 3693 19408 4108 19410
rect 3693 19352 3698 19408
rect 3754 19352 4108 19408
rect 3693 19350 4108 19352
rect 3693 19347 3759 19350
rect 4102 19348 4108 19350
rect 4172 19348 4178 19412
rect 4245 19410 4311 19413
rect 9581 19410 9647 19413
rect 4245 19408 9647 19410
rect 4245 19352 4250 19408
rect 4306 19352 9586 19408
rect 9642 19352 9647 19408
rect 4245 19350 9647 19352
rect 4245 19347 4311 19350
rect 9581 19347 9647 19350
rect 12750 19348 12756 19412
rect 12820 19410 12826 19412
rect 13077 19410 13143 19413
rect 12820 19408 13143 19410
rect 12820 19352 13082 19408
rect 13138 19352 13143 19408
rect 12820 19350 13143 19352
rect 12820 19348 12826 19350
rect 13077 19347 13143 19350
rect 0 19274 800 19304
rect 1209 19274 1275 19277
rect 0 19272 1275 19274
rect 0 19216 1214 19272
rect 1270 19216 1275 19272
rect 0 19214 1275 19216
rect 0 19184 800 19214
rect 1209 19211 1275 19214
rect 5257 19274 5323 19277
rect 6177 19274 6243 19277
rect 15469 19274 15535 19277
rect 5257 19272 6243 19274
rect 5257 19216 5262 19272
rect 5318 19216 6182 19272
rect 6238 19216 6243 19272
rect 5257 19214 6243 19216
rect 5257 19211 5323 19214
rect 6177 19211 6243 19214
rect 6318 19272 15535 19274
rect 6318 19216 15474 19272
rect 15530 19216 15535 19272
rect 6318 19214 15535 19216
rect 4613 19138 4679 19141
rect 6318 19138 6378 19214
rect 15469 19211 15535 19214
rect 13445 19138 13511 19141
rect 4613 19136 6378 19138
rect 4613 19080 4618 19136
rect 4674 19080 6378 19136
rect 4613 19078 6378 19080
rect 9262 19136 13511 19138
rect 9262 19080 13450 19136
rect 13506 19080 13511 19136
rect 9262 19078 13511 19080
rect 4613 19075 4679 19078
rect 3543 19072 3863 19073
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 19007 3863 19008
rect 8741 19072 9061 19073
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 19007 9061 19008
rect 6913 19002 6979 19005
rect 6913 19000 7850 19002
rect 6913 18944 6918 19000
rect 6974 18944 7850 19000
rect 6913 18942 7850 18944
rect 6913 18939 6979 18942
rect 0 18866 800 18896
rect 1853 18866 1919 18869
rect 0 18864 1919 18866
rect 0 18808 1858 18864
rect 1914 18808 1919 18864
rect 0 18806 1919 18808
rect 0 18776 800 18806
rect 1853 18803 1919 18806
rect 2221 18866 2287 18869
rect 7557 18866 7623 18869
rect 2221 18864 7623 18866
rect 2221 18808 2226 18864
rect 2282 18808 7562 18864
rect 7618 18808 7623 18864
rect 2221 18806 7623 18808
rect 7790 18866 7850 18942
rect 9262 18866 9322 19078
rect 13445 19075 13511 19078
rect 13939 19072 14259 19073
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 19007 14259 19008
rect 19137 19072 19457 19073
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 19007 19457 19008
rect 9949 19002 10015 19005
rect 13629 19002 13695 19005
rect 9949 19000 13695 19002
rect 9949 18944 9954 19000
rect 10010 18944 13634 19000
rect 13690 18944 13695 19000
rect 9949 18942 13695 18944
rect 9949 18939 10015 18942
rect 13629 18939 13695 18942
rect 7790 18806 9322 18866
rect 10225 18866 10291 18869
rect 11605 18866 11671 18869
rect 10225 18864 11671 18866
rect 10225 18808 10230 18864
rect 10286 18808 11610 18864
rect 11666 18808 11671 18864
rect 10225 18806 11671 18808
rect 2221 18803 2287 18806
rect 7557 18803 7623 18806
rect 10225 18803 10291 18806
rect 11605 18803 11671 18806
rect 11789 18866 11855 18869
rect 13905 18866 13971 18869
rect 11789 18864 13971 18866
rect 11789 18808 11794 18864
rect 11850 18808 13910 18864
rect 13966 18808 13971 18864
rect 11789 18806 13971 18808
rect 11789 18803 11855 18806
rect 13905 18803 13971 18806
rect 2129 18730 2195 18733
rect 2262 18730 2268 18732
rect 2129 18728 2268 18730
rect 2129 18672 2134 18728
rect 2190 18672 2268 18728
rect 2129 18670 2268 18672
rect 2129 18667 2195 18670
rect 2262 18668 2268 18670
rect 2332 18668 2338 18732
rect 14825 18730 14891 18733
rect 2454 18728 14891 18730
rect 2454 18672 14830 18728
rect 14886 18672 14891 18728
rect 2454 18670 14891 18672
rect 1761 18594 1827 18597
rect 2454 18594 2514 18670
rect 14825 18667 14891 18670
rect 15142 18668 15148 18732
rect 15212 18730 15218 18732
rect 15653 18730 15719 18733
rect 15212 18728 15719 18730
rect 15212 18672 15658 18728
rect 15714 18672 15719 18728
rect 15212 18670 15719 18672
rect 15212 18668 15218 18670
rect 15653 18667 15719 18670
rect 1761 18592 2514 18594
rect 1761 18536 1766 18592
rect 1822 18536 2514 18592
rect 1761 18534 2514 18536
rect 7097 18594 7163 18597
rect 9489 18594 9555 18597
rect 7097 18592 9555 18594
rect 7097 18536 7102 18592
rect 7158 18536 9494 18592
rect 9550 18536 9555 18592
rect 7097 18534 9555 18536
rect 1761 18531 1827 18534
rect 7097 18531 7163 18534
rect 9489 18531 9555 18534
rect 6142 18528 6462 18529
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 18463 6462 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 16538 18528 16858 18529
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 18463 16858 18464
rect 9949 18458 10015 18461
rect 7422 18456 10015 18458
rect 7422 18400 9954 18456
rect 10010 18400 10015 18456
rect 7422 18398 10015 18400
rect 0 18322 800 18352
rect 2221 18322 2287 18325
rect 0 18320 2287 18322
rect 0 18264 2226 18320
rect 2282 18264 2287 18320
rect 0 18262 2287 18264
rect 0 18232 800 18262
rect 2221 18259 2287 18262
rect 4429 18322 4495 18325
rect 7422 18322 7482 18398
rect 9949 18395 10015 18398
rect 4429 18320 7482 18322
rect 4429 18264 4434 18320
rect 4490 18264 7482 18320
rect 4429 18262 7482 18264
rect 7557 18322 7623 18325
rect 13261 18322 13327 18325
rect 7557 18320 13327 18322
rect 7557 18264 7562 18320
rect 7618 18264 13266 18320
rect 13322 18264 13327 18320
rect 7557 18262 13327 18264
rect 4429 18259 4495 18262
rect 7557 18259 7623 18262
rect 13261 18259 13327 18262
rect 3325 18188 3391 18189
rect 3325 18186 3372 18188
rect 3244 18184 3372 18186
rect 3436 18186 3442 18188
rect 4245 18186 4311 18189
rect 11605 18186 11671 18189
rect 3244 18128 3330 18184
rect 3244 18126 3372 18128
rect 3325 18124 3372 18126
rect 3436 18126 3986 18186
rect 3436 18124 3442 18126
rect 3325 18123 3391 18124
rect 3926 18050 3986 18126
rect 4245 18184 11671 18186
rect 4245 18128 4250 18184
rect 4306 18128 11610 18184
rect 11666 18128 11671 18184
rect 4245 18126 11671 18128
rect 4245 18123 4311 18126
rect 11605 18123 11671 18126
rect 7097 18050 7163 18053
rect 3926 18048 7163 18050
rect 3926 17992 7102 18048
rect 7158 17992 7163 18048
rect 3926 17990 7163 17992
rect 7097 17987 7163 17990
rect 9489 18050 9555 18053
rect 11789 18050 11855 18053
rect 9489 18048 11855 18050
rect 9489 17992 9494 18048
rect 9550 17992 11794 18048
rect 11850 17992 11855 18048
rect 9489 17990 11855 17992
rect 9489 17987 9555 17990
rect 11789 17987 11855 17990
rect 3543 17984 3863 17985
rect 0 17914 800 17944
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 17919 3863 17920
rect 8741 17984 9061 17985
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 17919 9061 17920
rect 13939 17984 14259 17985
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 17919 14259 17920
rect 19137 17984 19457 17985
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 17919 19457 17920
rect 1485 17914 1551 17917
rect 0 17912 1551 17914
rect 0 17856 1490 17912
rect 1546 17856 1551 17912
rect 0 17854 1551 17856
rect 0 17824 800 17854
rect 1485 17851 1551 17854
rect 2773 17914 2839 17917
rect 3233 17914 3299 17917
rect 2773 17912 3299 17914
rect 2773 17856 2778 17912
rect 2834 17856 3238 17912
rect 3294 17856 3299 17912
rect 2773 17854 3299 17856
rect 2773 17851 2839 17854
rect 3233 17851 3299 17854
rect 4613 17914 4679 17917
rect 6545 17914 6611 17917
rect 4613 17912 6611 17914
rect 4613 17856 4618 17912
rect 4674 17856 6550 17912
rect 6606 17856 6611 17912
rect 4613 17854 6611 17856
rect 4613 17851 4679 17854
rect 6545 17851 6611 17854
rect 12249 17914 12315 17917
rect 12750 17914 12756 17916
rect 12249 17912 12756 17914
rect 12249 17856 12254 17912
rect 12310 17856 12756 17912
rect 12249 17854 12756 17856
rect 12249 17851 12315 17854
rect 12750 17852 12756 17854
rect 12820 17852 12826 17916
rect 2037 17778 2103 17781
rect 10501 17778 10567 17781
rect 2037 17776 10567 17778
rect 2037 17720 2042 17776
rect 2098 17720 10506 17776
rect 10562 17720 10567 17776
rect 2037 17718 10567 17720
rect 2037 17715 2103 17718
rect 10501 17715 10567 17718
rect 1945 17642 2011 17645
rect 10041 17642 10107 17645
rect 1945 17640 10107 17642
rect 1945 17584 1950 17640
rect 2006 17584 10046 17640
rect 10102 17584 10107 17640
rect 1945 17582 10107 17584
rect 1945 17579 2011 17582
rect 10041 17579 10107 17582
rect 6142 17440 6462 17441
rect 0 17370 800 17400
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 17375 6462 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 16538 17440 16858 17441
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 17375 16858 17376
rect 1485 17370 1551 17373
rect 0 17368 1551 17370
rect 0 17312 1490 17368
rect 1546 17312 1551 17368
rect 0 17310 1551 17312
rect 0 17280 800 17310
rect 1485 17307 1551 17310
rect 2957 17370 3023 17373
rect 5717 17370 5783 17373
rect 2957 17368 5783 17370
rect 2957 17312 2962 17368
rect 3018 17312 5722 17368
rect 5778 17312 5783 17368
rect 2957 17310 5783 17312
rect 2957 17307 3023 17310
rect 5717 17307 5783 17310
rect 2313 17234 2379 17237
rect 9305 17234 9371 17237
rect 2313 17232 9371 17234
rect 2313 17176 2318 17232
rect 2374 17176 9310 17232
rect 9366 17176 9371 17232
rect 2313 17174 9371 17176
rect 2313 17171 2379 17174
rect 9305 17171 9371 17174
rect 21449 17234 21515 17237
rect 22200 17234 23000 17264
rect 21449 17232 23000 17234
rect 21449 17176 21454 17232
rect 21510 17176 23000 17232
rect 21449 17174 23000 17176
rect 21449 17171 21515 17174
rect 22200 17144 23000 17174
rect 4797 17098 4863 17101
rect 21081 17098 21147 17101
rect 4797 17096 21147 17098
rect 4797 17040 4802 17096
rect 4858 17040 21086 17096
rect 21142 17040 21147 17096
rect 4797 17038 21147 17040
rect 4797 17035 4863 17038
rect 21081 17035 21147 17038
rect 0 16962 800 16992
rect 1485 16962 1551 16965
rect 0 16960 1551 16962
rect 0 16904 1490 16960
rect 1546 16904 1551 16960
rect 0 16902 1551 16904
rect 0 16872 800 16902
rect 1485 16899 1551 16902
rect 3543 16896 3863 16897
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 16831 3863 16832
rect 8741 16896 9061 16897
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 16831 9061 16832
rect 13939 16896 14259 16897
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 16831 14259 16832
rect 19137 16896 19457 16897
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 16831 19457 16832
rect 2773 16690 2839 16693
rect 6821 16690 6887 16693
rect 2773 16688 6887 16690
rect 2773 16632 2778 16688
rect 2834 16632 6826 16688
rect 6882 16632 6887 16688
rect 2773 16630 6887 16632
rect 2773 16627 2839 16630
rect 6821 16627 6887 16630
rect 8753 16690 8819 16693
rect 12525 16690 12591 16693
rect 8753 16688 12591 16690
rect 8753 16632 8758 16688
rect 8814 16632 12530 16688
rect 12586 16632 12591 16688
rect 8753 16630 12591 16632
rect 8753 16627 8819 16630
rect 12525 16627 12591 16630
rect 2681 16554 2747 16557
rect 6269 16554 6335 16557
rect 2454 16552 2747 16554
rect 2454 16496 2686 16552
rect 2742 16496 2747 16552
rect 2454 16494 2747 16496
rect 0 16418 800 16448
rect 2454 16421 2514 16494
rect 2681 16491 2747 16494
rect 4662 16552 6335 16554
rect 4662 16496 6274 16552
rect 6330 16496 6335 16552
rect 4662 16494 6335 16496
rect 1485 16418 1551 16421
rect 0 16416 1551 16418
rect 0 16360 1490 16416
rect 1546 16360 1551 16416
rect 0 16358 1551 16360
rect 0 16328 800 16358
rect 1485 16355 1551 16358
rect 2405 16416 2514 16421
rect 2405 16360 2410 16416
rect 2466 16360 2514 16416
rect 2405 16358 2514 16360
rect 2681 16418 2747 16421
rect 4662 16418 4722 16494
rect 6269 16491 6335 16494
rect 2681 16416 4722 16418
rect 2681 16360 2686 16416
rect 2742 16360 4722 16416
rect 2681 16358 4722 16360
rect 2405 16355 2471 16358
rect 2681 16355 2747 16358
rect 6142 16352 6462 16353
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 16287 6462 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 16538 16352 16858 16353
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 16287 16858 16288
rect 2681 16146 2747 16149
rect 8109 16146 8175 16149
rect 2681 16144 8175 16146
rect 2681 16088 2686 16144
rect 2742 16088 8114 16144
rect 8170 16088 8175 16144
rect 2681 16086 8175 16088
rect 2681 16083 2747 16086
rect 8109 16083 8175 16086
rect 0 16010 800 16040
rect 1485 16010 1551 16013
rect 0 16008 1551 16010
rect 0 15952 1490 16008
rect 1546 15952 1551 16008
rect 0 15950 1551 15952
rect 0 15920 800 15950
rect 1485 15947 1551 15950
rect 3141 16010 3207 16013
rect 7649 16010 7715 16013
rect 3141 16008 7715 16010
rect 3141 15952 3146 16008
rect 3202 15952 7654 16008
rect 7710 15952 7715 16008
rect 3141 15950 7715 15952
rect 3141 15947 3207 15950
rect 7649 15947 7715 15950
rect 9121 16010 9187 16013
rect 18597 16010 18663 16013
rect 9121 16008 18663 16010
rect 9121 15952 9126 16008
rect 9182 15952 18602 16008
rect 18658 15952 18663 16008
rect 9121 15950 18663 15952
rect 9121 15947 9187 15950
rect 18597 15947 18663 15950
rect 3543 15808 3863 15809
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 15743 3863 15744
rect 8741 15808 9061 15809
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 15743 9061 15744
rect 13939 15808 14259 15809
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 15743 14259 15744
rect 19137 15808 19457 15809
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 15743 19457 15744
rect 3366 15540 3372 15604
rect 3436 15602 3442 15604
rect 3509 15602 3575 15605
rect 4245 15602 4311 15605
rect 3436 15600 4311 15602
rect 3436 15544 3514 15600
rect 3570 15544 4250 15600
rect 4306 15544 4311 15600
rect 3436 15542 4311 15544
rect 3436 15540 3442 15542
rect 3509 15539 3575 15542
rect 4245 15539 4311 15542
rect 0 15466 800 15496
rect 1853 15466 1919 15469
rect 0 15464 1919 15466
rect 0 15408 1858 15464
rect 1914 15408 1919 15464
rect 0 15406 1919 15408
rect 0 15376 800 15406
rect 1853 15403 1919 15406
rect 5165 15466 5231 15469
rect 9029 15466 9095 15469
rect 5165 15464 9095 15466
rect 5165 15408 5170 15464
rect 5226 15408 9034 15464
rect 9090 15408 9095 15464
rect 5165 15406 9095 15408
rect 5165 15403 5231 15406
rect 9029 15403 9095 15406
rect 6142 15264 6462 15265
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 15199 6462 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 16538 15264 16858 15265
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 15199 16858 15200
rect 0 15058 800 15088
rect 1485 15058 1551 15061
rect 0 15056 1551 15058
rect 0 15000 1490 15056
rect 1546 15000 1551 15056
rect 0 14998 1551 15000
rect 0 14968 800 14998
rect 1485 14995 1551 14998
rect 5441 15058 5507 15061
rect 8753 15058 8819 15061
rect 5441 15056 8819 15058
rect 5441 15000 5446 15056
rect 5502 15000 8758 15056
rect 8814 15000 8819 15056
rect 5441 14998 8819 15000
rect 5441 14995 5507 14998
rect 8753 14995 8819 14998
rect 3509 14922 3575 14925
rect 10225 14922 10291 14925
rect 3509 14920 10291 14922
rect 3509 14864 3514 14920
rect 3570 14864 10230 14920
rect 10286 14864 10291 14920
rect 3509 14862 10291 14864
rect 3509 14859 3575 14862
rect 10225 14859 10291 14862
rect 3543 14720 3863 14721
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 14655 3863 14656
rect 8741 14720 9061 14721
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 14655 9061 14656
rect 13939 14720 14259 14721
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 14655 14259 14656
rect 19137 14720 19457 14721
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 14655 19457 14656
rect 0 14514 800 14544
rect 1485 14514 1551 14517
rect 0 14512 1551 14514
rect 0 14456 1490 14512
rect 1546 14456 1551 14512
rect 0 14454 1551 14456
rect 0 14424 800 14454
rect 1485 14451 1551 14454
rect 9857 14514 9923 14517
rect 10542 14514 10548 14516
rect 9857 14512 10548 14514
rect 9857 14456 9862 14512
rect 9918 14456 10548 14512
rect 9857 14454 10548 14456
rect 9857 14451 9923 14454
rect 10542 14452 10548 14454
rect 10612 14452 10618 14516
rect 3141 14378 3207 14381
rect 3877 14378 3943 14381
rect 3141 14376 3943 14378
rect 3141 14320 3146 14376
rect 3202 14320 3882 14376
rect 3938 14320 3943 14376
rect 3141 14318 3943 14320
rect 3141 14315 3207 14318
rect 3877 14315 3943 14318
rect 12157 14242 12223 14245
rect 12934 14242 12940 14244
rect 12157 14240 12940 14242
rect 12157 14184 12162 14240
rect 12218 14184 12940 14240
rect 12157 14182 12940 14184
rect 12157 14179 12223 14182
rect 12934 14180 12940 14182
rect 13004 14180 13010 14244
rect 6142 14176 6462 14177
rect 0 14106 800 14136
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 14111 6462 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 16538 14176 16858 14177
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 14111 16858 14112
rect 1485 14106 1551 14109
rect 0 14104 1551 14106
rect 0 14048 1490 14104
rect 1546 14048 1551 14104
rect 0 14046 1551 14048
rect 0 14016 800 14046
rect 1485 14043 1551 14046
rect 2630 13908 2636 13972
rect 2700 13970 2706 13972
rect 9673 13970 9739 13973
rect 2700 13968 9739 13970
rect 2700 13912 9678 13968
rect 9734 13912 9739 13968
rect 2700 13910 9739 13912
rect 2700 13908 2706 13910
rect 9673 13907 9739 13910
rect 10910 13908 10916 13972
rect 10980 13970 10986 13972
rect 12617 13970 12683 13973
rect 10980 13968 12683 13970
rect 10980 13912 12622 13968
rect 12678 13912 12683 13968
rect 10980 13910 12683 13912
rect 10980 13908 10986 13910
rect 12617 13907 12683 13910
rect 3543 13632 3863 13633
rect 0 13562 800 13592
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 13567 3863 13568
rect 8741 13632 9061 13633
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 13567 9061 13568
rect 13939 13632 14259 13633
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 13567 14259 13568
rect 19137 13632 19457 13633
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 13567 19457 13568
rect 1485 13562 1551 13565
rect 0 13560 1551 13562
rect 0 13504 1490 13560
rect 1546 13504 1551 13560
rect 0 13502 1551 13504
rect 0 13472 800 13502
rect 1485 13499 1551 13502
rect 1710 13364 1716 13428
rect 1780 13426 1786 13428
rect 7557 13426 7623 13429
rect 1780 13424 7623 13426
rect 1780 13368 7562 13424
rect 7618 13368 7623 13424
rect 1780 13366 7623 13368
rect 1780 13364 1786 13366
rect 7557 13363 7623 13366
rect 1577 13290 1643 13293
rect 13353 13290 13419 13293
rect 1577 13288 13419 13290
rect 1577 13232 1582 13288
rect 1638 13232 13358 13288
rect 13414 13232 13419 13288
rect 1577 13230 13419 13232
rect 1577 13227 1643 13230
rect 13353 13227 13419 13230
rect 0 13154 800 13184
rect 1393 13154 1459 13157
rect 0 13152 1459 13154
rect 0 13096 1398 13152
rect 1454 13096 1459 13152
rect 0 13094 1459 13096
rect 0 13064 800 13094
rect 1393 13091 1459 13094
rect 6142 13088 6462 13089
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 13023 6462 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 16538 13088 16858 13089
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 13023 16858 13024
rect 0 12610 800 12640
rect 1393 12610 1459 12613
rect 0 12608 1459 12610
rect 0 12552 1398 12608
rect 1454 12552 1459 12608
rect 0 12550 1459 12552
rect 0 12520 800 12550
rect 1393 12547 1459 12550
rect 3543 12544 3863 12545
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 12479 3863 12480
rect 8741 12544 9061 12545
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 12479 9061 12480
rect 13939 12544 14259 12545
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 12479 14259 12480
rect 19137 12544 19457 12545
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 12479 19457 12480
rect 4470 12412 4476 12476
rect 4540 12474 4546 12476
rect 5441 12474 5507 12477
rect 4540 12472 5507 12474
rect 4540 12416 5446 12472
rect 5502 12416 5507 12472
rect 4540 12414 5507 12416
rect 4540 12412 4546 12414
rect 5441 12411 5507 12414
rect 5625 12338 5691 12341
rect 10777 12338 10843 12341
rect 11881 12338 11947 12341
rect 5625 12336 9276 12338
rect 5625 12280 5630 12336
rect 5686 12280 9276 12336
rect 5625 12278 9276 12280
rect 5625 12275 5691 12278
rect 0 12202 800 12232
rect 1485 12202 1551 12205
rect 0 12200 1551 12202
rect 0 12144 1490 12200
rect 1546 12144 1551 12200
rect 0 12142 1551 12144
rect 0 12112 800 12142
rect 1485 12139 1551 12142
rect 6142 12000 6462 12001
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 11935 6462 11936
rect 9216 11797 9276 12278
rect 10777 12336 11947 12338
rect 10777 12280 10782 12336
rect 10838 12280 11886 12336
rect 11942 12280 11947 12336
rect 10777 12278 11947 12280
rect 10777 12275 10843 12278
rect 11881 12275 11947 12278
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 16538 12000 16858 12001
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 11935 16858 11936
rect 1853 11794 1919 11797
rect 4981 11794 5047 11797
rect 9213 11794 9279 11797
rect 15009 11794 15075 11797
rect 1853 11792 5047 11794
rect 1853 11736 1858 11792
rect 1914 11736 4986 11792
rect 5042 11736 5047 11792
rect 1853 11734 5047 11736
rect 9086 11792 15075 11794
rect 9086 11736 9218 11792
rect 9274 11736 15014 11792
rect 15070 11736 15075 11792
rect 9086 11734 15075 11736
rect 1853 11731 1919 11734
rect 4981 11731 5047 11734
rect 9213 11731 9279 11734
rect 15009 11731 15075 11734
rect 0 11658 800 11688
rect 1669 11658 1735 11661
rect 0 11656 1735 11658
rect 0 11600 1674 11656
rect 1730 11600 1735 11656
rect 0 11598 1735 11600
rect 0 11568 800 11598
rect 1669 11595 1735 11598
rect 4797 11658 4863 11661
rect 11237 11658 11303 11661
rect 4797 11656 11303 11658
rect 4797 11600 4802 11656
rect 4858 11600 11242 11656
rect 11298 11600 11303 11656
rect 4797 11598 11303 11600
rect 4797 11595 4863 11598
rect 11237 11595 11303 11598
rect 4705 11522 4771 11525
rect 5574 11522 5580 11524
rect 4705 11520 5580 11522
rect 4705 11464 4710 11520
rect 4766 11464 5580 11520
rect 4705 11462 5580 11464
rect 4705 11459 4771 11462
rect 5574 11460 5580 11462
rect 5644 11460 5650 11524
rect 3543 11456 3863 11457
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 11391 3863 11392
rect 8741 11456 9061 11457
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 11391 9061 11392
rect 13939 11456 14259 11457
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 11391 14259 11392
rect 19137 11456 19457 11457
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 11391 19457 11392
rect 9438 11324 9444 11388
rect 9508 11386 9514 11388
rect 11513 11386 11579 11389
rect 9508 11384 11579 11386
rect 9508 11328 11518 11384
rect 11574 11328 11579 11384
rect 9508 11326 11579 11328
rect 9508 11324 9514 11326
rect 11513 11323 11579 11326
rect 12341 11386 12407 11389
rect 12525 11386 12591 11389
rect 12341 11384 12591 11386
rect 12341 11328 12346 11384
rect 12402 11328 12530 11384
rect 12586 11328 12591 11384
rect 12341 11326 12591 11328
rect 12341 11323 12407 11326
rect 12525 11323 12591 11326
rect 2037 11250 2103 11253
rect 9489 11250 9555 11253
rect 2037 11248 9555 11250
rect 2037 11192 2042 11248
rect 2098 11192 9494 11248
rect 9550 11192 9555 11248
rect 2037 11190 9555 11192
rect 2037 11187 2103 11190
rect 9489 11187 9555 11190
rect 10961 11250 11027 11253
rect 13169 11250 13235 11253
rect 10961 11248 13235 11250
rect 10961 11192 10966 11248
rect 11022 11192 13174 11248
rect 13230 11192 13235 11248
rect 10961 11190 13235 11192
rect 10961 11187 11027 11190
rect 13169 11187 13235 11190
rect 0 11114 800 11144
rect 1393 11114 1459 11117
rect 0 11112 1459 11114
rect 0 11056 1398 11112
rect 1454 11056 1459 11112
rect 0 11054 1459 11056
rect 0 11024 800 11054
rect 1393 11051 1459 11054
rect 1577 11114 1643 11117
rect 6821 11114 6887 11117
rect 1577 11112 6887 11114
rect 1577 11056 1582 11112
rect 1638 11056 6826 11112
rect 6882 11056 6887 11112
rect 1577 11054 6887 11056
rect 1577 11051 1643 11054
rect 6821 11051 6887 11054
rect 3969 10978 4035 10981
rect 5206 10978 5212 10980
rect 3969 10976 5212 10978
rect 3969 10920 3974 10976
rect 4030 10920 5212 10976
rect 3969 10918 5212 10920
rect 3969 10915 4035 10918
rect 5206 10916 5212 10918
rect 5276 10916 5282 10980
rect 6142 10912 6462 10913
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 10847 6462 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 16538 10912 16858 10913
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 10847 16858 10848
rect 0 10706 800 10736
rect 1669 10706 1735 10709
rect 0 10704 1735 10706
rect 0 10648 1674 10704
rect 1730 10648 1735 10704
rect 0 10646 1735 10648
rect 0 10616 800 10646
rect 1669 10643 1735 10646
rect 2129 10570 2195 10573
rect 13353 10570 13419 10573
rect 2129 10568 13419 10570
rect 2129 10512 2134 10568
rect 2190 10512 13358 10568
rect 13414 10512 13419 10568
rect 2129 10510 13419 10512
rect 2129 10507 2195 10510
rect 13353 10507 13419 10510
rect 3543 10368 3863 10369
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 10303 3863 10304
rect 8741 10368 9061 10369
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 10303 9061 10304
rect 13939 10368 14259 10369
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 10303 14259 10304
rect 19137 10368 19457 10369
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 10303 19457 10304
rect 0 10162 800 10192
rect 1853 10162 1919 10165
rect 0 10160 1919 10162
rect 0 10104 1858 10160
rect 1914 10104 1919 10160
rect 0 10102 1919 10104
rect 0 10072 800 10102
rect 1853 10099 1919 10102
rect 2037 10162 2103 10165
rect 9121 10162 9187 10165
rect 2037 10160 9187 10162
rect 2037 10104 2042 10160
rect 2098 10104 9126 10160
rect 9182 10104 9187 10160
rect 2037 10102 9187 10104
rect 2037 10099 2103 10102
rect 9121 10099 9187 10102
rect 3601 10026 3667 10029
rect 5625 10026 5691 10029
rect 5758 10026 5764 10028
rect 3601 10024 5764 10026
rect 3601 9968 3606 10024
rect 3662 9968 5630 10024
rect 5686 9968 5764 10024
rect 3601 9966 5764 9968
rect 3601 9963 3667 9966
rect 5625 9963 5691 9966
rect 5758 9964 5764 9966
rect 5828 9964 5834 10028
rect 6678 9964 6684 10028
rect 6748 10026 6754 10028
rect 11697 10026 11763 10029
rect 6748 10024 11763 10026
rect 6748 9968 11702 10024
rect 11758 9968 11763 10024
rect 6748 9966 11763 9968
rect 6748 9964 6754 9966
rect 11697 9963 11763 9966
rect 6142 9824 6462 9825
rect 0 9754 800 9784
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 9759 6462 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 16538 9824 16858 9825
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 9759 16858 9760
rect 2773 9754 2839 9757
rect 0 9752 2839 9754
rect 0 9696 2778 9752
rect 2834 9696 2839 9752
rect 0 9694 2839 9696
rect 0 9664 800 9694
rect 2773 9691 2839 9694
rect 9397 9754 9463 9757
rect 10358 9754 10364 9756
rect 9397 9752 10364 9754
rect 9397 9696 9402 9752
rect 9458 9696 10364 9752
rect 9397 9694 10364 9696
rect 9397 9691 9463 9694
rect 10358 9692 10364 9694
rect 10428 9692 10434 9756
rect 2037 9618 2103 9621
rect 5993 9618 6059 9621
rect 2037 9616 6059 9618
rect 2037 9560 2042 9616
rect 2098 9560 5998 9616
rect 6054 9560 6059 9616
rect 2037 9558 6059 9560
rect 2037 9555 2103 9558
rect 5993 9555 6059 9558
rect 12014 9556 12020 9620
rect 12084 9618 12090 9620
rect 15377 9618 15443 9621
rect 12084 9616 15443 9618
rect 12084 9560 15382 9616
rect 15438 9560 15443 9616
rect 12084 9558 15443 9560
rect 12084 9556 12090 9558
rect 15377 9555 15443 9558
rect 4889 9346 4955 9349
rect 5257 9346 5323 9349
rect 5942 9346 5948 9348
rect 4889 9344 5948 9346
rect 4889 9288 4894 9344
rect 4950 9288 5262 9344
rect 5318 9288 5948 9344
rect 4889 9286 5948 9288
rect 4889 9283 4955 9286
rect 5257 9283 5323 9286
rect 5942 9284 5948 9286
rect 6012 9346 6018 9348
rect 7005 9346 7071 9349
rect 6012 9344 7071 9346
rect 6012 9288 7010 9344
rect 7066 9288 7071 9344
rect 6012 9286 7071 9288
rect 6012 9284 6018 9286
rect 7005 9283 7071 9286
rect 3543 9280 3863 9281
rect 0 9210 800 9240
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 9215 3863 9216
rect 8741 9280 9061 9281
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 9215 9061 9216
rect 13939 9280 14259 9281
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 9215 14259 9216
rect 19137 9280 19457 9281
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 9215 19457 9216
rect 1393 9210 1459 9213
rect 0 9208 1459 9210
rect 0 9152 1398 9208
rect 1454 9152 1459 9208
rect 0 9150 1459 9152
rect 0 9120 800 9150
rect 1393 9147 1459 9150
rect 5390 9012 5396 9076
rect 5460 9074 5466 9076
rect 6085 9074 6151 9077
rect 5460 9072 6151 9074
rect 5460 9016 6090 9072
rect 6146 9016 6151 9072
rect 5460 9014 6151 9016
rect 5460 9012 5466 9014
rect 6085 9011 6151 9014
rect 1577 8938 1643 8941
rect 13445 8938 13511 8941
rect 1577 8936 13511 8938
rect 1577 8880 1582 8936
rect 1638 8880 13450 8936
rect 13506 8880 13511 8936
rect 1577 8878 13511 8880
rect 1577 8875 1643 8878
rect 13445 8875 13511 8878
rect 0 8802 800 8832
rect 1342 8802 1348 8804
rect 0 8742 1348 8802
rect 0 8712 800 8742
rect 1342 8740 1348 8742
rect 1412 8740 1418 8804
rect 2630 8740 2636 8804
rect 2700 8802 2706 8804
rect 2957 8802 3023 8805
rect 8477 8804 8543 8805
rect 8477 8802 8524 8804
rect 2700 8800 3023 8802
rect 2700 8744 2962 8800
rect 3018 8744 3023 8800
rect 2700 8742 3023 8744
rect 8432 8800 8524 8802
rect 8432 8744 8482 8800
rect 8432 8742 8524 8744
rect 2700 8740 2706 8742
rect 2957 8739 3023 8742
rect 8477 8740 8524 8742
rect 8588 8740 8594 8804
rect 8477 8739 8543 8740
rect 6142 8736 6462 8737
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 8671 6462 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 16538 8736 16858 8737
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 8671 16858 8672
rect 9213 8666 9279 8669
rect 9397 8666 9463 8669
rect 9213 8664 9463 8666
rect 9213 8608 9218 8664
rect 9274 8608 9402 8664
rect 9458 8608 9463 8664
rect 9213 8606 9463 8608
rect 9213 8603 9279 8606
rect 9397 8603 9463 8606
rect 2078 8468 2084 8532
rect 2148 8530 2154 8532
rect 12985 8530 13051 8533
rect 2148 8528 13051 8530
rect 2148 8472 12990 8528
rect 13046 8472 13051 8528
rect 2148 8470 13051 8472
rect 2148 8468 2154 8470
rect 12985 8467 13051 8470
rect 1393 8394 1459 8397
rect 3969 8394 4035 8397
rect 4153 8394 4219 8397
rect 1393 8392 4035 8394
rect 1393 8336 1398 8392
rect 1454 8336 3974 8392
rect 4030 8336 4035 8392
rect 1393 8334 4035 8336
rect 1393 8331 1459 8334
rect 3969 8331 4035 8334
rect 4110 8392 4219 8394
rect 4110 8336 4158 8392
rect 4214 8336 4219 8392
rect 4110 8331 4219 8336
rect 5165 8394 5231 8397
rect 8334 8394 8340 8396
rect 5165 8392 8340 8394
rect 5165 8336 5170 8392
rect 5226 8336 8340 8392
rect 5165 8334 8340 8336
rect 5165 8331 5231 8334
rect 8334 8332 8340 8334
rect 8404 8394 8410 8396
rect 11789 8394 11855 8397
rect 8404 8392 11855 8394
rect 8404 8336 11794 8392
rect 11850 8336 11855 8392
rect 8404 8334 11855 8336
rect 8404 8332 8410 8334
rect 11789 8331 11855 8334
rect 0 8258 800 8288
rect 1669 8258 1735 8261
rect 4110 8260 4170 8331
rect 0 8256 1735 8258
rect 0 8200 1674 8256
rect 1730 8200 1735 8256
rect 0 8198 1735 8200
rect 0 8168 800 8198
rect 1669 8195 1735 8198
rect 4102 8196 4108 8260
rect 4172 8196 4178 8260
rect 3543 8192 3863 8193
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 8127 3863 8128
rect 8741 8192 9061 8193
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 8127 9061 8128
rect 13939 8192 14259 8193
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 8127 14259 8128
rect 19137 8192 19457 8193
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 8127 19457 8128
rect 9305 8122 9371 8125
rect 9305 8120 13738 8122
rect 9305 8064 9310 8120
rect 9366 8064 13738 8120
rect 9305 8062 13738 8064
rect 9305 8059 9371 8062
rect 12985 7986 13051 7989
rect 2730 7984 13051 7986
rect 2730 7928 12990 7984
rect 13046 7928 13051 7984
rect 2730 7926 13051 7928
rect 13678 7986 13738 8062
rect 15285 7986 15351 7989
rect 13678 7984 15351 7986
rect 13678 7928 15290 7984
rect 15346 7928 15351 7984
rect 13678 7926 15351 7928
rect 0 7850 800 7880
rect 1945 7850 2011 7853
rect 2730 7850 2790 7926
rect 12985 7923 13051 7926
rect 15285 7923 15351 7926
rect 0 7848 2790 7850
rect 0 7792 1950 7848
rect 2006 7792 2790 7848
rect 0 7790 2790 7792
rect 3509 7850 3575 7853
rect 11053 7850 11119 7853
rect 12525 7850 12591 7853
rect 3509 7848 11119 7850
rect 3509 7792 3514 7848
rect 3570 7792 11058 7848
rect 11114 7792 11119 7848
rect 3509 7790 11119 7792
rect 0 7760 800 7790
rect 1945 7787 2011 7790
rect 3509 7787 3575 7790
rect 11053 7787 11119 7790
rect 12390 7848 12591 7850
rect 12390 7792 12530 7848
rect 12586 7792 12591 7848
rect 12390 7790 12591 7792
rect 2681 7714 2747 7717
rect 4245 7716 4311 7717
rect 4245 7714 4292 7716
rect 2681 7712 4292 7714
rect 2681 7656 2686 7712
rect 2742 7656 4250 7712
rect 2681 7654 4292 7656
rect 2681 7651 2747 7654
rect 4245 7652 4292 7654
rect 4356 7652 4362 7716
rect 6545 7714 6611 7717
rect 9765 7714 9831 7717
rect 6545 7712 9831 7714
rect 6545 7656 6550 7712
rect 6606 7656 9770 7712
rect 9826 7656 9831 7712
rect 6545 7654 9831 7656
rect 4245 7651 4311 7652
rect 6545 7651 6611 7654
rect 9765 7651 9831 7654
rect 6142 7648 6462 7649
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 7583 6462 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 6729 7578 6795 7581
rect 6729 7576 9506 7578
rect 6729 7520 6734 7576
rect 6790 7520 9506 7576
rect 6729 7518 9506 7520
rect 6729 7515 6795 7518
rect 2497 7442 2563 7445
rect 9305 7442 9371 7445
rect 2497 7440 9371 7442
rect 2497 7384 2502 7440
rect 2558 7384 9310 7440
rect 9366 7384 9371 7440
rect 2497 7382 9371 7384
rect 9446 7442 9506 7518
rect 12390 7442 12450 7790
rect 12525 7787 12591 7790
rect 16538 7648 16858 7649
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 7583 16858 7584
rect 9446 7382 12450 7442
rect 2497 7379 2563 7382
rect 9305 7379 9371 7382
rect 0 7306 800 7336
rect 1669 7306 1735 7309
rect 0 7304 1735 7306
rect 0 7248 1674 7304
rect 1730 7248 1735 7304
rect 0 7246 1735 7248
rect 0 7216 800 7246
rect 1669 7243 1735 7246
rect 4797 7306 4863 7309
rect 6729 7306 6795 7309
rect 4797 7304 6795 7306
rect 4797 7248 4802 7304
rect 4858 7248 6734 7304
rect 6790 7248 6795 7304
rect 4797 7246 6795 7248
rect 4797 7243 4863 7246
rect 6729 7243 6795 7246
rect 8293 7306 8359 7309
rect 15193 7306 15259 7309
rect 8293 7304 15259 7306
rect 8293 7248 8298 7304
rect 8354 7248 15198 7304
rect 15254 7248 15259 7304
rect 8293 7246 15259 7248
rect 8293 7243 8359 7246
rect 15193 7243 15259 7246
rect 5390 7108 5396 7172
rect 5460 7170 5466 7172
rect 5533 7170 5599 7173
rect 5460 7168 5599 7170
rect 5460 7112 5538 7168
rect 5594 7112 5599 7168
rect 5460 7110 5599 7112
rect 5460 7108 5466 7110
rect 5533 7107 5599 7110
rect 6821 7170 6887 7173
rect 8385 7170 8451 7173
rect 6821 7168 8451 7170
rect 6821 7112 6826 7168
rect 6882 7112 8390 7168
rect 8446 7112 8451 7168
rect 6821 7110 8451 7112
rect 6821 7107 6887 7110
rect 8385 7107 8451 7110
rect 9121 7170 9187 7173
rect 9254 7170 9260 7172
rect 9121 7168 9260 7170
rect 9121 7112 9126 7168
rect 9182 7112 9260 7168
rect 9121 7110 9260 7112
rect 9121 7107 9187 7110
rect 9254 7108 9260 7110
rect 9324 7108 9330 7172
rect 9949 7170 10015 7173
rect 12341 7170 12407 7173
rect 9949 7168 12407 7170
rect 9949 7112 9954 7168
rect 10010 7112 12346 7168
rect 12402 7112 12407 7168
rect 9949 7110 12407 7112
rect 9949 7107 10015 7110
rect 12341 7107 12407 7110
rect 3543 7104 3863 7105
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 7039 3863 7040
rect 8741 7104 9061 7105
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 7039 9061 7040
rect 13939 7104 14259 7105
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 7039 14259 7040
rect 19137 7104 19457 7105
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 7039 19457 7040
rect 4286 6972 4292 7036
rect 4356 7034 4362 7036
rect 8201 7034 8267 7037
rect 4356 7032 8267 7034
rect 4356 6976 8206 7032
rect 8262 6976 8267 7032
rect 4356 6974 8267 6976
rect 4356 6972 4362 6974
rect 8201 6971 8267 6974
rect 9121 7034 9187 7037
rect 11881 7034 11947 7037
rect 9121 7032 11947 7034
rect 9121 6976 9126 7032
rect 9182 6976 11886 7032
rect 11942 6976 11947 7032
rect 9121 6974 11947 6976
rect 9121 6971 9187 6974
rect 11881 6971 11947 6974
rect 0 6898 800 6928
rect 1761 6898 1827 6901
rect 12801 6898 12867 6901
rect 0 6838 1456 6898
rect 0 6808 800 6838
rect 1396 6762 1456 6838
rect 1761 6896 12867 6898
rect 1761 6840 1766 6896
rect 1822 6840 12806 6896
rect 12862 6840 12867 6896
rect 1761 6838 12867 6840
rect 1761 6835 1827 6838
rect 12801 6835 12867 6838
rect 4245 6762 4311 6765
rect 1396 6760 4311 6762
rect 1396 6704 4250 6760
rect 4306 6704 4311 6760
rect 1396 6702 4311 6704
rect 4245 6699 4311 6702
rect 4981 6762 5047 6765
rect 10501 6762 10567 6765
rect 11973 6762 12039 6765
rect 4981 6760 10567 6762
rect 4981 6704 4986 6760
rect 5042 6704 10506 6760
rect 10562 6704 10567 6760
rect 4981 6702 10567 6704
rect 4981 6699 5047 6702
rect 10501 6699 10567 6702
rect 10734 6760 12039 6762
rect 10734 6704 11978 6760
rect 12034 6704 12039 6760
rect 10734 6702 12039 6704
rect 1393 6628 1459 6629
rect 1342 6564 1348 6628
rect 1412 6626 1459 6628
rect 3969 6626 4035 6629
rect 5349 6626 5415 6629
rect 1412 6624 1504 6626
rect 1454 6568 1504 6624
rect 1412 6566 1504 6568
rect 3969 6624 5415 6626
rect 3969 6568 3974 6624
rect 4030 6568 5354 6624
rect 5410 6568 5415 6624
rect 3969 6566 5415 6568
rect 1412 6564 1459 6566
rect 1393 6563 1459 6564
rect 3969 6563 4035 6566
rect 5349 6563 5415 6566
rect 6729 6626 6795 6629
rect 10734 6626 10794 6702
rect 11973 6699 12039 6702
rect 15469 6762 15535 6765
rect 16205 6762 16271 6765
rect 15469 6760 16271 6762
rect 15469 6704 15474 6760
rect 15530 6704 16210 6760
rect 16266 6704 16271 6760
rect 15469 6702 16271 6704
rect 15469 6699 15535 6702
rect 16205 6699 16271 6702
rect 6729 6624 10794 6626
rect 6729 6568 6734 6624
rect 6790 6568 10794 6624
rect 6729 6566 10794 6568
rect 6729 6563 6795 6566
rect 6142 6560 6462 6561
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 6495 6462 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 16538 6560 16858 6561
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 6495 16858 6496
rect 2313 6490 2379 6493
rect 4889 6490 4955 6493
rect 2313 6488 4955 6490
rect 2313 6432 2318 6488
rect 2374 6432 4894 6488
rect 4950 6432 4955 6488
rect 2313 6430 4955 6432
rect 2313 6427 2379 6430
rect 4889 6427 4955 6430
rect 7189 6490 7255 6493
rect 7925 6490 7991 6493
rect 7189 6488 7991 6490
rect 7189 6432 7194 6488
rect 7250 6432 7930 6488
rect 7986 6432 7991 6488
rect 7189 6430 7991 6432
rect 7189 6427 7255 6430
rect 7925 6427 7991 6430
rect 8845 6490 8911 6493
rect 9305 6490 9371 6493
rect 8845 6488 9371 6490
rect 8845 6432 8850 6488
rect 8906 6432 9310 6488
rect 9366 6432 9371 6488
rect 8845 6430 9371 6432
rect 8845 6427 8911 6430
rect 9305 6427 9371 6430
rect 0 6354 800 6384
rect 1669 6354 1735 6357
rect 8293 6354 8359 6357
rect 0 6352 8359 6354
rect 0 6296 1674 6352
rect 1730 6296 8298 6352
rect 8354 6296 8359 6352
rect 0 6294 8359 6296
rect 0 6264 800 6294
rect 1669 6291 1735 6294
rect 8293 6291 8359 6294
rect 8937 6354 9003 6357
rect 8937 6352 10978 6354
rect 8937 6296 8942 6352
rect 8998 6296 10978 6352
rect 8937 6294 10978 6296
rect 8937 6291 9003 6294
rect 4245 6218 4311 6221
rect 10041 6218 10107 6221
rect 4245 6216 10107 6218
rect 4245 6160 4250 6216
rect 4306 6160 10046 6216
rect 10102 6160 10107 6216
rect 4245 6158 10107 6160
rect 10918 6218 10978 6294
rect 18781 6218 18847 6221
rect 10918 6216 18847 6218
rect 10918 6160 18786 6216
rect 18842 6160 18847 6216
rect 10918 6158 18847 6160
rect 4245 6155 4311 6158
rect 10041 6155 10107 6158
rect 18781 6155 18847 6158
rect 4521 6082 4587 6085
rect 5257 6082 5323 6085
rect 4521 6080 5323 6082
rect 4521 6024 4526 6080
rect 4582 6024 5262 6080
rect 5318 6024 5323 6080
rect 4521 6022 5323 6024
rect 4521 6019 4587 6022
rect 5257 6019 5323 6022
rect 10501 6082 10567 6085
rect 10501 6080 12450 6082
rect 10501 6024 10506 6080
rect 10562 6024 12450 6080
rect 10501 6022 12450 6024
rect 10501 6019 10567 6022
rect 3543 6016 3863 6017
rect 0 5946 800 5976
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 5951 3863 5952
rect 8741 6016 9061 6017
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 5951 9061 5952
rect 1393 5946 1459 5949
rect 4981 5946 5047 5949
rect 5257 5948 5323 5949
rect 0 5944 1459 5946
rect 0 5888 1398 5944
rect 1454 5888 1459 5944
rect 0 5886 1459 5888
rect 0 5856 800 5886
rect 1393 5883 1459 5886
rect 3926 5944 5047 5946
rect 3926 5888 4986 5944
rect 5042 5888 5047 5944
rect 3926 5886 5047 5888
rect 3049 5810 3115 5813
rect 3926 5810 3986 5886
rect 4981 5883 5047 5886
rect 5206 5884 5212 5948
rect 5276 5946 5323 5948
rect 6729 5946 6795 5949
rect 5276 5944 6795 5946
rect 5318 5888 6734 5944
rect 6790 5888 6795 5944
rect 5276 5886 6795 5888
rect 5276 5884 5323 5886
rect 5257 5883 5323 5884
rect 6729 5883 6795 5886
rect 3049 5808 3986 5810
rect 3049 5752 3054 5808
rect 3110 5752 3986 5808
rect 3049 5750 3986 5752
rect 4889 5810 4955 5813
rect 11881 5810 11947 5813
rect 4889 5808 11947 5810
rect 4889 5752 4894 5808
rect 4950 5752 11886 5808
rect 11942 5752 11947 5808
rect 4889 5750 11947 5752
rect 12390 5810 12450 6022
rect 13939 6016 14259 6017
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 5951 14259 5952
rect 19137 6016 19457 6017
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 5951 19457 5952
rect 14457 5946 14523 5949
rect 15653 5946 15719 5949
rect 14457 5944 15719 5946
rect 14457 5888 14462 5944
rect 14518 5888 15658 5944
rect 15714 5888 15719 5944
rect 14457 5886 15719 5888
rect 14457 5883 14523 5886
rect 15653 5883 15719 5886
rect 17217 5810 17283 5813
rect 12390 5808 17283 5810
rect 12390 5752 17222 5808
rect 17278 5752 17283 5808
rect 12390 5750 17283 5752
rect 3049 5747 3115 5750
rect 4889 5747 4955 5750
rect 11881 5747 11947 5750
rect 17217 5747 17283 5750
rect 21541 5810 21607 5813
rect 22200 5810 23000 5840
rect 21541 5808 23000 5810
rect 21541 5752 21546 5808
rect 21602 5752 23000 5808
rect 21541 5750 23000 5752
rect 21541 5747 21607 5750
rect 22200 5720 23000 5750
rect 1485 5674 1551 5677
rect 13169 5674 13235 5677
rect 1485 5672 13235 5674
rect 1485 5616 1490 5672
rect 1546 5616 13174 5672
rect 13230 5616 13235 5672
rect 1485 5614 13235 5616
rect 1485 5611 1551 5614
rect 13169 5611 13235 5614
rect 1117 5538 1183 5541
rect 5809 5538 5875 5541
rect 11053 5538 11119 5541
rect 1117 5536 5875 5538
rect 1117 5480 1122 5536
rect 1178 5480 5814 5536
rect 5870 5480 5875 5536
rect 1117 5478 5875 5480
rect 1117 5475 1183 5478
rect 5809 5475 5875 5478
rect 8158 5536 11119 5538
rect 8158 5480 11058 5536
rect 11114 5480 11119 5536
rect 8158 5478 11119 5480
rect 6142 5472 6462 5473
rect 0 5402 800 5432
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 5407 6462 5408
rect 2773 5402 2839 5405
rect 0 5400 2839 5402
rect 0 5344 2778 5400
rect 2834 5344 2839 5400
rect 0 5342 2839 5344
rect 0 5312 800 5342
rect 2773 5339 2839 5342
rect 3366 5340 3372 5404
rect 3436 5402 3442 5404
rect 3509 5402 3575 5405
rect 4797 5402 4863 5405
rect 3436 5400 4863 5402
rect 3436 5344 3514 5400
rect 3570 5344 4802 5400
rect 4858 5344 4863 5400
rect 3436 5342 4863 5344
rect 3436 5340 3442 5342
rect 3509 5339 3575 5342
rect 4797 5339 4863 5342
rect 2773 5266 2839 5269
rect 3601 5266 3667 5269
rect 4429 5268 4495 5269
rect 4429 5266 4476 5268
rect 2773 5264 3667 5266
rect 2773 5208 2778 5264
rect 2834 5208 3606 5264
rect 3662 5208 3667 5264
rect 2773 5206 3667 5208
rect 4384 5264 4476 5266
rect 4540 5266 4546 5268
rect 8158 5266 8218 5478
rect 11053 5475 11119 5478
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 16538 5472 16858 5473
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 5407 16858 5408
rect 10409 5402 10475 5405
rect 10542 5402 10548 5404
rect 10409 5400 10548 5402
rect 10409 5344 10414 5400
rect 10470 5344 10548 5400
rect 10409 5342 10548 5344
rect 10409 5339 10475 5342
rect 10542 5340 10548 5342
rect 10612 5340 10618 5404
rect 4384 5208 4434 5264
rect 4384 5206 4476 5208
rect 2773 5203 2839 5206
rect 3601 5203 3667 5206
rect 4429 5204 4476 5206
rect 4540 5206 8218 5266
rect 9765 5266 9831 5269
rect 9949 5266 10015 5269
rect 9765 5264 10015 5266
rect 9765 5208 9770 5264
rect 9826 5208 9954 5264
rect 10010 5208 10015 5264
rect 9765 5206 10015 5208
rect 4540 5204 4546 5206
rect 4429 5203 4495 5204
rect 9765 5203 9831 5206
rect 9949 5203 10015 5206
rect 10726 5204 10732 5268
rect 10796 5266 10802 5268
rect 12249 5266 12315 5269
rect 10796 5264 12315 5266
rect 10796 5208 12254 5264
rect 12310 5208 12315 5264
rect 10796 5206 12315 5208
rect 10796 5204 10802 5206
rect 12249 5203 12315 5206
rect 12801 5266 12867 5269
rect 18597 5266 18663 5269
rect 12801 5264 18663 5266
rect 12801 5208 12806 5264
rect 12862 5208 18602 5264
rect 18658 5208 18663 5264
rect 12801 5206 18663 5208
rect 12801 5203 12867 5206
rect 18597 5203 18663 5206
rect 1577 5130 1643 5133
rect 1710 5130 1716 5132
rect 1577 5128 1716 5130
rect 1577 5072 1582 5128
rect 1638 5072 1716 5128
rect 1577 5070 1716 5072
rect 1577 5067 1643 5070
rect 1710 5068 1716 5070
rect 1780 5068 1786 5132
rect 4613 5130 4679 5133
rect 2730 5128 4679 5130
rect 2730 5072 4618 5128
rect 4674 5072 4679 5128
rect 2730 5070 4679 5072
rect 0 4994 800 5024
rect 2730 4994 2790 5070
rect 4613 5067 4679 5070
rect 5165 5130 5231 5133
rect 6453 5130 6519 5133
rect 7281 5130 7347 5133
rect 5165 5128 7347 5130
rect 5165 5072 5170 5128
rect 5226 5072 6458 5128
rect 6514 5072 7286 5128
rect 7342 5072 7347 5128
rect 5165 5070 7347 5072
rect 5165 5067 5231 5070
rect 6453 5067 6519 5070
rect 7281 5067 7347 5070
rect 7414 5068 7420 5132
rect 7484 5130 7490 5132
rect 8293 5130 8359 5133
rect 7484 5128 8359 5130
rect 7484 5072 8298 5128
rect 8354 5072 8359 5128
rect 7484 5070 8359 5072
rect 7484 5068 7490 5070
rect 8293 5067 8359 5070
rect 9857 5130 9923 5133
rect 9857 5128 15072 5130
rect 9857 5072 9862 5128
rect 9918 5072 15072 5128
rect 9857 5070 15072 5072
rect 9857 5067 9923 5070
rect 0 4934 2790 4994
rect 4613 4994 4679 4997
rect 6678 4994 6684 4996
rect 4613 4992 6684 4994
rect 4613 4936 4618 4992
rect 4674 4936 6684 4992
rect 4613 4934 6684 4936
rect 0 4904 800 4934
rect 4613 4931 4679 4934
rect 6678 4932 6684 4934
rect 6748 4932 6754 4996
rect 10409 4994 10475 4997
rect 15012 4994 15072 5070
rect 15142 5068 15148 5132
rect 15212 5130 15218 5132
rect 15653 5130 15719 5133
rect 15212 5128 15719 5130
rect 15212 5072 15658 5128
rect 15714 5072 15719 5128
rect 15212 5070 15719 5072
rect 15212 5068 15218 5070
rect 15653 5067 15719 5070
rect 16389 4994 16455 4997
rect 10409 4992 13002 4994
rect 10409 4936 10414 4992
rect 10470 4936 13002 4992
rect 10409 4934 13002 4936
rect 15012 4992 16455 4994
rect 15012 4936 16394 4992
rect 16450 4936 16455 4992
rect 15012 4934 16455 4936
rect 10409 4931 10475 4934
rect 3543 4928 3863 4929
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 4863 3863 4864
rect 8741 4928 9061 4929
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 4863 9061 4864
rect 12942 4861 13002 4934
rect 16389 4931 16455 4934
rect 13939 4928 14259 4929
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 4863 14259 4864
rect 19137 4928 19457 4929
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 4863 19457 4864
rect 2037 4860 2103 4861
rect 2037 4858 2084 4860
rect 1992 4856 2084 4858
rect 1992 4800 2042 4856
rect 1992 4798 2084 4800
rect 2037 4796 2084 4798
rect 2148 4796 2154 4860
rect 4102 4796 4108 4860
rect 4172 4858 4178 4860
rect 6269 4858 6335 4861
rect 4172 4856 6335 4858
rect 4172 4800 6274 4856
rect 6330 4800 6335 4856
rect 4172 4798 6335 4800
rect 4172 4796 4178 4798
rect 2037 4795 2103 4796
rect 6269 4795 6335 4798
rect 11881 4858 11947 4861
rect 12801 4858 12867 4861
rect 11881 4856 12867 4858
rect 11881 4800 11886 4856
rect 11942 4800 12806 4856
rect 12862 4800 12867 4856
rect 11881 4798 12867 4800
rect 12942 4856 13051 4861
rect 12942 4800 12990 4856
rect 13046 4800 13051 4856
rect 12942 4798 13051 4800
rect 11881 4795 11947 4798
rect 12801 4795 12867 4798
rect 12985 4795 13051 4798
rect 2681 4722 2747 4725
rect 13905 4722 13971 4725
rect 2681 4720 13971 4722
rect 2681 4664 2686 4720
rect 2742 4664 13910 4720
rect 13966 4664 13971 4720
rect 2681 4662 13971 4664
rect 2681 4659 2747 4662
rect 13905 4659 13971 4662
rect 2037 4586 2103 4589
rect 3417 4586 3483 4589
rect 2037 4584 3483 4586
rect 2037 4528 2042 4584
rect 2098 4528 3422 4584
rect 3478 4528 3483 4584
rect 2037 4526 3483 4528
rect 2037 4523 2103 4526
rect 3417 4523 3483 4526
rect 4153 4586 4219 4589
rect 7189 4586 7255 4589
rect 12525 4586 12591 4589
rect 4153 4584 7114 4586
rect 4153 4528 4158 4584
rect 4214 4528 7114 4584
rect 4153 4526 7114 4528
rect 4153 4523 4219 4526
rect 0 4450 800 4480
rect 2773 4450 2839 4453
rect 0 4448 2839 4450
rect 0 4392 2778 4448
rect 2834 4392 2839 4448
rect 0 4390 2839 4392
rect 0 4360 800 4390
rect 2773 4387 2839 4390
rect 6545 4450 6611 4453
rect 6678 4450 6684 4452
rect 6545 4448 6684 4450
rect 6545 4392 6550 4448
rect 6606 4392 6684 4448
rect 6545 4390 6684 4392
rect 6545 4387 6611 4390
rect 6678 4388 6684 4390
rect 6748 4388 6754 4452
rect 7054 4450 7114 4526
rect 7189 4584 12591 4586
rect 7189 4528 7194 4584
rect 7250 4528 12530 4584
rect 12586 4528 12591 4584
rect 7189 4526 12591 4528
rect 7189 4523 7255 4526
rect 12525 4523 12591 4526
rect 9673 4450 9739 4453
rect 10685 4452 10751 4453
rect 10685 4450 10732 4452
rect 7054 4448 9739 4450
rect 7054 4392 9678 4448
rect 9734 4392 9739 4448
rect 7054 4390 9739 4392
rect 10640 4448 10732 4450
rect 10640 4392 10690 4448
rect 10640 4390 10732 4392
rect 9673 4387 9739 4390
rect 10685 4388 10732 4390
rect 10796 4388 10802 4452
rect 12433 4450 12499 4453
rect 16205 4450 16271 4453
rect 12433 4448 16271 4450
rect 12433 4392 12438 4448
rect 12494 4392 16210 4448
rect 16266 4392 16271 4448
rect 12433 4390 16271 4392
rect 10685 4387 10751 4388
rect 12433 4387 12499 4390
rect 16205 4387 16271 4390
rect 6142 4384 6462 4385
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 4319 6462 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 16538 4384 16858 4385
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 4319 16858 4320
rect 2405 4316 2471 4317
rect 2405 4314 2452 4316
rect 2360 4312 2452 4314
rect 2360 4256 2410 4312
rect 2360 4254 2452 4256
rect 2405 4252 2452 4254
rect 2516 4252 2522 4316
rect 5257 4314 5323 4317
rect 3006 4312 5323 4314
rect 3006 4256 5262 4312
rect 5318 4256 5323 4312
rect 3006 4254 5323 4256
rect 2405 4251 2471 4252
rect 0 4042 800 4072
rect 2865 4042 2931 4045
rect 0 4040 2931 4042
rect 0 3984 2870 4040
rect 2926 3984 2931 4040
rect 0 3982 2931 3984
rect 0 3952 800 3982
rect 2865 3979 2931 3982
rect 2221 3906 2287 3909
rect 3006 3906 3066 4254
rect 5257 4251 5323 4254
rect 8334 4252 8340 4316
rect 8404 4314 8410 4316
rect 8477 4314 8543 4317
rect 8404 4312 8543 4314
rect 8404 4256 8482 4312
rect 8538 4256 8543 4312
rect 8404 4254 8543 4256
rect 8404 4252 8410 4254
rect 8477 4251 8543 4254
rect 15142 4252 15148 4316
rect 15212 4314 15218 4316
rect 15837 4314 15903 4317
rect 15212 4312 15903 4314
rect 15212 4256 15842 4312
rect 15898 4256 15903 4312
rect 15212 4254 15903 4256
rect 15212 4252 15218 4254
rect 15837 4251 15903 4254
rect 3141 4178 3207 4181
rect 5809 4178 5875 4181
rect 3141 4176 5875 4178
rect 3141 4120 3146 4176
rect 3202 4120 5814 4176
rect 5870 4120 5875 4176
rect 3141 4118 5875 4120
rect 3141 4115 3207 4118
rect 5809 4115 5875 4118
rect 6545 4178 6611 4181
rect 11881 4178 11947 4181
rect 6545 4176 11947 4178
rect 6545 4120 6550 4176
rect 6606 4120 11886 4176
rect 11942 4120 11947 4176
rect 6545 4118 11947 4120
rect 6545 4115 6611 4118
rect 11881 4115 11947 4118
rect 15285 4178 15351 4181
rect 15469 4178 15535 4181
rect 15285 4176 15535 4178
rect 15285 4120 15290 4176
rect 15346 4120 15474 4176
rect 15530 4120 15535 4176
rect 15285 4118 15535 4120
rect 15285 4115 15351 4118
rect 15469 4115 15535 4118
rect 4061 4042 4127 4045
rect 7230 4042 7236 4044
rect 4061 4040 7236 4042
rect 4061 3984 4066 4040
rect 4122 3984 7236 4040
rect 4061 3982 7236 3984
rect 4061 3979 4127 3982
rect 7230 3980 7236 3982
rect 7300 3980 7306 4044
rect 7465 4042 7531 4045
rect 10777 4042 10843 4045
rect 10910 4042 10916 4044
rect 7465 4040 9276 4042
rect 7465 3984 7470 4040
rect 7526 3984 9276 4040
rect 7465 3982 9276 3984
rect 7465 3979 7531 3982
rect 2221 3904 3066 3906
rect 2221 3848 2226 3904
rect 2282 3848 3066 3904
rect 2221 3846 3066 3848
rect 2221 3843 2287 3846
rect 5758 3844 5764 3908
rect 5828 3906 5834 3908
rect 5901 3906 5967 3909
rect 6361 3906 6427 3909
rect 5828 3904 6427 3906
rect 5828 3848 5906 3904
rect 5962 3848 6366 3904
rect 6422 3848 6427 3904
rect 5828 3846 6427 3848
rect 9216 3906 9276 3982
rect 10777 4040 10916 4042
rect 10777 3984 10782 4040
rect 10838 3984 10916 4040
rect 10777 3982 10916 3984
rect 10777 3979 10843 3982
rect 10910 3980 10916 3982
rect 10980 3980 10986 4044
rect 15009 4042 15075 4045
rect 12390 4040 15075 4042
rect 12390 3984 15014 4040
rect 15070 3984 15075 4040
rect 12390 3982 15075 3984
rect 12390 3906 12450 3982
rect 15009 3979 15075 3982
rect 9216 3846 12450 3906
rect 5828 3844 5834 3846
rect 5901 3843 5967 3846
rect 6361 3843 6427 3846
rect 3543 3840 3863 3841
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 3775 3863 3776
rect 8741 3840 9061 3841
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 3775 9061 3776
rect 13939 3840 14259 3841
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 3775 14259 3776
rect 19137 3840 19457 3841
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 3775 19457 3776
rect 1669 3770 1735 3773
rect 2630 3770 2636 3772
rect 1669 3768 2636 3770
rect 1669 3712 1674 3768
rect 1730 3712 2636 3768
rect 1669 3710 2636 3712
rect 1669 3707 1735 3710
rect 2630 3708 2636 3710
rect 2700 3708 2706 3772
rect 5625 3770 5691 3773
rect 6913 3770 6979 3773
rect 5625 3768 6979 3770
rect 5625 3712 5630 3768
rect 5686 3712 6918 3768
rect 6974 3712 6979 3768
rect 5625 3710 6979 3712
rect 5625 3707 5691 3710
rect 6913 3707 6979 3710
rect 10133 3770 10199 3773
rect 11513 3770 11579 3773
rect 10133 3768 11579 3770
rect 10133 3712 10138 3768
rect 10194 3712 11518 3768
rect 11574 3712 11579 3768
rect 10133 3710 11579 3712
rect 10133 3707 10199 3710
rect 11513 3707 11579 3710
rect 16665 3634 16731 3637
rect 2730 3632 16731 3634
rect 2730 3576 16670 3632
rect 16726 3576 16731 3632
rect 2730 3574 16731 3576
rect 0 3498 800 3528
rect 1485 3498 1551 3501
rect 0 3496 1551 3498
rect 0 3440 1490 3496
rect 1546 3440 1551 3496
rect 0 3438 1551 3440
rect 0 3408 800 3438
rect 1485 3435 1551 3438
rect 2221 3498 2287 3501
rect 2730 3498 2790 3574
rect 16665 3571 16731 3574
rect 2221 3496 2790 3498
rect 2221 3440 2226 3496
rect 2282 3440 2790 3496
rect 2221 3438 2790 3440
rect 4889 3498 4955 3501
rect 7833 3498 7899 3501
rect 10869 3498 10935 3501
rect 15653 3498 15719 3501
rect 4889 3496 6746 3498
rect 4889 3440 4894 3496
rect 4950 3440 6746 3496
rect 4889 3438 6746 3440
rect 2221 3435 2287 3438
rect 4889 3435 4955 3438
rect 1209 3362 1275 3365
rect 4797 3362 4863 3365
rect 1209 3360 4863 3362
rect 1209 3304 1214 3360
rect 1270 3304 4802 3360
rect 4858 3304 4863 3360
rect 1209 3302 4863 3304
rect 1209 3299 1275 3302
rect 4797 3299 4863 3302
rect 6142 3296 6462 3297
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 3231 6462 3232
rect 2630 3164 2636 3228
rect 2700 3226 2706 3228
rect 5625 3226 5691 3229
rect 5993 3228 6059 3229
rect 5942 3226 5948 3228
rect 2700 3224 5691 3226
rect 2700 3168 5630 3224
rect 5686 3168 5691 3224
rect 2700 3166 5691 3168
rect 5902 3166 5948 3226
rect 6012 3224 6059 3228
rect 6054 3168 6059 3224
rect 2700 3164 2706 3166
rect 5625 3163 5691 3166
rect 5942 3164 5948 3166
rect 6012 3164 6059 3168
rect 6686 3226 6746 3438
rect 7833 3496 10935 3498
rect 7833 3440 7838 3496
rect 7894 3440 10874 3496
rect 10930 3440 10935 3496
rect 7833 3438 10935 3440
rect 7833 3435 7899 3438
rect 10869 3435 10935 3438
rect 11102 3496 15719 3498
rect 11102 3440 15658 3496
rect 15714 3440 15719 3496
rect 11102 3438 15719 3440
rect 8477 3364 8543 3365
rect 8477 3360 8524 3364
rect 8588 3362 8594 3364
rect 8477 3304 8482 3360
rect 8477 3300 8524 3304
rect 8588 3302 8634 3362
rect 8588 3300 8594 3302
rect 8477 3299 8543 3300
rect 6821 3226 6887 3229
rect 11102 3226 11162 3438
rect 15653 3435 15719 3438
rect 14181 3362 14247 3365
rect 14406 3362 14412 3364
rect 14181 3360 14412 3362
rect 14181 3304 14186 3360
rect 14242 3304 14412 3360
rect 14181 3302 14412 3304
rect 14181 3299 14247 3302
rect 14406 3300 14412 3302
rect 14476 3300 14482 3364
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 16538 3296 16858 3297
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 3231 16858 3232
rect 6686 3224 11162 3226
rect 6686 3168 6826 3224
rect 6882 3168 11162 3224
rect 6686 3166 11162 3168
rect 11881 3226 11947 3229
rect 12014 3226 12020 3228
rect 11881 3224 12020 3226
rect 11881 3168 11886 3224
rect 11942 3168 12020 3224
rect 11881 3166 12020 3168
rect 5993 3163 6059 3164
rect 6821 3163 6887 3166
rect 11881 3163 11947 3166
rect 12014 3164 12020 3166
rect 12084 3164 12090 3228
rect 0 3090 800 3120
rect 1853 3090 1919 3093
rect 3417 3090 3483 3093
rect 0 3088 3483 3090
rect 0 3032 1858 3088
rect 1914 3032 3422 3088
rect 3478 3032 3483 3088
rect 0 3030 3483 3032
rect 0 3000 800 3030
rect 1853 3027 1919 3030
rect 3417 3027 3483 3030
rect 5901 3090 5967 3093
rect 12249 3090 12315 3093
rect 5901 3088 12315 3090
rect 5901 3032 5906 3088
rect 5962 3032 12254 3088
rect 12310 3032 12315 3088
rect 5901 3030 12315 3032
rect 5901 3027 5967 3030
rect 12249 3027 12315 3030
rect 15561 3090 15627 3093
rect 17033 3090 17099 3093
rect 15561 3088 17099 3090
rect 15561 3032 15566 3088
rect 15622 3032 17038 3088
rect 17094 3032 17099 3088
rect 15561 3030 17099 3032
rect 15561 3027 15627 3030
rect 17033 3027 17099 3030
rect 3233 2954 3299 2957
rect 3366 2954 3372 2956
rect 3233 2952 3372 2954
rect 3233 2896 3238 2952
rect 3294 2896 3372 2952
rect 3233 2894 3372 2896
rect 3233 2891 3299 2894
rect 3366 2892 3372 2894
rect 3436 2892 3442 2956
rect 6085 2954 6151 2957
rect 13721 2954 13787 2957
rect 6085 2952 13787 2954
rect 6085 2896 6090 2952
rect 6146 2896 13726 2952
rect 13782 2896 13787 2952
rect 6085 2894 13787 2896
rect 6085 2891 6151 2894
rect 13721 2891 13787 2894
rect 197 2818 263 2821
rect 2221 2818 2287 2821
rect 197 2816 2287 2818
rect 197 2760 202 2816
rect 258 2760 2226 2816
rect 2282 2760 2287 2816
rect 197 2758 2287 2760
rect 197 2755 263 2758
rect 2221 2755 2287 2758
rect 9213 2820 9279 2821
rect 9213 2816 9260 2820
rect 9324 2818 9330 2820
rect 10041 2818 10107 2821
rect 11329 2818 11395 2821
rect 9213 2760 9218 2816
rect 9213 2756 9260 2760
rect 9324 2758 9370 2818
rect 10041 2816 11395 2818
rect 10041 2760 10046 2816
rect 10102 2760 11334 2816
rect 11390 2760 11395 2816
rect 10041 2758 11395 2760
rect 9324 2756 9330 2758
rect 9213 2755 9279 2756
rect 10041 2755 10107 2758
rect 11329 2755 11395 2758
rect 3543 2752 3863 2753
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2687 3863 2688
rect 8741 2752 9061 2753
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2687 9061 2688
rect 13939 2752 14259 2753
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2687 14259 2688
rect 19137 2752 19457 2753
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2687 19457 2688
rect 3969 2682 4035 2685
rect 5533 2684 5599 2685
rect 4102 2682 4108 2684
rect 3969 2680 4108 2682
rect 3969 2624 3974 2680
rect 4030 2624 4108 2680
rect 3969 2622 4108 2624
rect 3969 2619 4035 2622
rect 4102 2620 4108 2622
rect 4172 2620 4178 2684
rect 5533 2680 5580 2684
rect 5644 2682 5650 2684
rect 6453 2682 6519 2685
rect 9397 2684 9463 2685
rect 6678 2682 6684 2684
rect 5533 2624 5538 2680
rect 5533 2620 5580 2624
rect 5644 2622 5690 2682
rect 6453 2680 6684 2682
rect 6453 2624 6458 2680
rect 6514 2624 6684 2680
rect 6453 2622 6684 2624
rect 5644 2620 5650 2622
rect 5533 2619 5599 2620
rect 6453 2619 6519 2622
rect 6678 2620 6684 2622
rect 6748 2620 6754 2684
rect 9397 2680 9444 2684
rect 9508 2682 9514 2684
rect 10225 2682 10291 2685
rect 10358 2682 10364 2684
rect 9397 2624 9402 2680
rect 9397 2620 9444 2624
rect 9508 2622 9554 2682
rect 10225 2680 10364 2682
rect 10225 2624 10230 2680
rect 10286 2624 10364 2680
rect 10225 2622 10364 2624
rect 9508 2620 9514 2622
rect 9397 2619 9463 2620
rect 10225 2619 10291 2622
rect 10358 2620 10364 2622
rect 10428 2620 10434 2684
rect 0 2546 800 2576
rect 2865 2546 2931 2549
rect 3049 2546 3115 2549
rect 15142 2546 15148 2548
rect 0 2544 3115 2546
rect 0 2488 2870 2544
rect 2926 2488 3054 2544
rect 3110 2488 3115 2544
rect 0 2486 3115 2488
rect 0 2456 800 2486
rect 2865 2483 2931 2486
rect 3049 2483 3115 2486
rect 3190 2486 15148 2546
rect 3190 2413 3250 2486
rect 15142 2484 15148 2486
rect 15212 2484 15218 2548
rect 3141 2410 3250 2413
rect 3060 2408 3250 2410
rect 3060 2352 3146 2408
rect 3202 2352 3250 2408
rect 3060 2350 3250 2352
rect 3141 2347 3250 2350
rect 3417 2410 3483 2413
rect 16941 2410 17007 2413
rect 3417 2408 17007 2410
rect 3417 2352 3422 2408
rect 3478 2352 16946 2408
rect 17002 2352 17007 2408
rect 3417 2350 17007 2352
rect 3417 2347 3483 2350
rect 16941 2347 17007 2350
rect 0 2138 800 2168
rect 3190 2138 3250 2347
rect 6142 2208 6462 2209
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2143 6462 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 16538 2208 16858 2209
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2143 16858 2144
rect 0 2078 3250 2138
rect 0 2048 800 2078
rect 1393 2002 1459 2005
rect 15929 2002 15995 2005
rect 1393 2000 15995 2002
rect 1393 1944 1398 2000
rect 1454 1944 15934 2000
rect 15990 1944 15995 2000
rect 1393 1942 15995 1944
rect 1393 1939 1459 1942
rect 15929 1939 15995 1942
rect 3141 1866 3207 1869
rect 3417 1866 3483 1869
rect 11697 1866 11763 1869
rect 3141 1864 11763 1866
rect 3141 1808 3146 1864
rect 3202 1808 3422 1864
rect 3478 1808 11702 1864
rect 11758 1808 11763 1864
rect 3141 1806 11763 1808
rect 3141 1803 3207 1806
rect 3417 1803 3483 1806
rect 11697 1803 11763 1806
rect 3233 1730 3299 1733
rect 2638 1728 3299 1730
rect 2638 1672 3238 1728
rect 3294 1672 3299 1728
rect 2638 1670 3299 1672
rect 0 1594 800 1624
rect 2638 1594 2698 1670
rect 3233 1667 3299 1670
rect 5809 1730 5875 1733
rect 13445 1730 13511 1733
rect 5809 1728 13511 1730
rect 5809 1672 5814 1728
rect 5870 1672 13450 1728
rect 13506 1672 13511 1728
rect 5809 1670 13511 1672
rect 5809 1667 5875 1670
rect 13445 1667 13511 1670
rect 0 1534 2698 1594
rect 3049 1594 3115 1597
rect 16297 1594 16363 1597
rect 3049 1592 16363 1594
rect 3049 1536 3054 1592
rect 3110 1536 16302 1592
rect 16358 1536 16363 1592
rect 3049 1534 16363 1536
rect 0 1504 800 1534
rect 3049 1531 3115 1534
rect 16297 1531 16363 1534
rect 2957 1458 3023 1461
rect 16021 1458 16087 1461
rect 2957 1456 16087 1458
rect 2957 1400 2962 1456
rect 3018 1400 16026 1456
rect 16082 1400 16087 1456
rect 2957 1398 16087 1400
rect 2957 1395 3023 1398
rect 16021 1395 16087 1398
rect 0 1186 800 1216
rect 1485 1186 1551 1189
rect 0 1184 1551 1186
rect 0 1128 1490 1184
rect 1546 1128 1551 1184
rect 0 1126 1551 1128
rect 0 1096 800 1126
rect 1485 1123 1551 1126
rect 0 642 800 672
rect 3325 642 3391 645
rect 0 640 3391 642
rect 0 584 3330 640
rect 3386 584 3391 640
rect 0 582 3391 584
rect 0 552 800 582
rect 3325 579 3391 582
rect 0 234 800 264
rect 4061 234 4127 237
rect 0 232 4127 234
rect 0 176 4066 232
rect 4122 176 4127 232
rect 0 174 4127 176
rect 0 144 800 174
rect 4061 171 4127 174
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 7420 20164 7484 20228
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 12940 19756 13004 19820
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 1900 19484 1964 19548
rect 1716 19348 1780 19412
rect 2636 19408 2700 19412
rect 2636 19352 2686 19408
rect 2686 19352 2700 19408
rect 2636 19348 2700 19352
rect 4108 19348 4172 19412
rect 12756 19348 12820 19412
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 2268 18668 2332 18732
rect 15148 18668 15212 18732
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 3372 18184 3436 18188
rect 3372 18128 3386 18184
rect 3386 18128 3436 18184
rect 3372 18124 3436 18128
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 12756 17852 12820 17916
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 3372 15540 3436 15604
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 10548 14452 10612 14516
rect 12940 14180 13004 14244
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 2636 13908 2700 13972
rect 10916 13908 10980 13972
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 1716 13364 1780 13428
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 4476 12412 4540 12476
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 5580 11460 5644 11524
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 9444 11324 9508 11388
rect 5212 10916 5276 10980
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 5764 9964 5828 10028
rect 6684 9964 6748 10028
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 10364 9692 10428 9756
rect 12020 9556 12084 9620
rect 5948 9284 6012 9348
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 5396 9012 5460 9076
rect 1348 8740 1412 8804
rect 2636 8740 2700 8804
rect 8524 8800 8588 8804
rect 8524 8744 8538 8800
rect 8538 8744 8588 8800
rect 8524 8740 8588 8744
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 2084 8468 2148 8532
rect 8340 8332 8404 8396
rect 4108 8196 4172 8260
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 4292 7712 4356 7716
rect 4292 7656 4306 7712
rect 4306 7656 4356 7712
rect 4292 7652 4356 7656
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 5396 7108 5460 7172
rect 9260 7108 9324 7172
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 4292 6972 4356 7036
rect 1348 6624 1412 6628
rect 1348 6568 1398 6624
rect 1398 6568 1412 6624
rect 1348 6564 1412 6568
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 5212 5944 5276 5948
rect 5212 5888 5262 5944
rect 5262 5888 5276 5944
rect 5212 5884 5276 5888
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 3372 5340 3436 5404
rect 4476 5264 4540 5268
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 10548 5340 10612 5404
rect 4476 5208 4490 5264
rect 4490 5208 4540 5264
rect 4476 5204 4540 5208
rect 10732 5204 10796 5268
rect 1716 5068 1780 5132
rect 7420 5068 7484 5132
rect 6684 4932 6748 4996
rect 15148 5068 15212 5132
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 2084 4856 2148 4860
rect 2084 4800 2098 4856
rect 2098 4800 2148 4856
rect 2084 4796 2148 4800
rect 4108 4796 4172 4860
rect 6684 4388 6748 4452
rect 10732 4448 10796 4452
rect 10732 4392 10746 4448
rect 10746 4392 10796 4448
rect 10732 4388 10796 4392
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 2452 4312 2516 4316
rect 2452 4256 2466 4312
rect 2466 4256 2516 4312
rect 2452 4252 2516 4256
rect 8340 4252 8404 4316
rect 15148 4252 15212 4316
rect 7236 3980 7300 4044
rect 5764 3844 5828 3908
rect 10916 3980 10980 4044
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 2636 3708 2700 3772
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 2636 3164 2700 3228
rect 5948 3224 6012 3228
rect 5948 3168 5998 3224
rect 5998 3168 6012 3224
rect 5948 3164 6012 3168
rect 8524 3360 8588 3364
rect 8524 3304 8538 3360
rect 8538 3304 8588 3360
rect 8524 3300 8588 3304
rect 14412 3300 14476 3364
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 12020 3164 12084 3228
rect 3372 2892 3436 2956
rect 9260 2816 9324 2820
rect 9260 2760 9274 2816
rect 9274 2760 9324 2816
rect 9260 2756 9324 2760
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 4108 2620 4172 2684
rect 5580 2680 5644 2684
rect 5580 2624 5594 2680
rect 5594 2624 5644 2680
rect 5580 2620 5644 2624
rect 6684 2620 6748 2684
rect 9444 2680 9508 2684
rect 9444 2624 9458 2680
rect 9458 2624 9508 2680
rect 9444 2620 9508 2624
rect 10364 2620 10428 2684
rect 15148 2484 15212 2548
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 1899 19548 1965 19549
rect 1899 19484 1900 19548
rect 1964 19484 1965 19548
rect 1899 19483 1965 19484
rect 1715 19412 1781 19413
rect 1715 19348 1716 19412
rect 1780 19348 1781 19412
rect 1715 19347 1781 19348
rect 1718 13429 1778 19347
rect 1902 16590 1962 19483
rect 2635 19412 2701 19413
rect 2635 19348 2636 19412
rect 2700 19348 2701 19412
rect 2635 19347 2701 19348
rect 1902 16530 2514 16590
rect 1715 13428 1781 13429
rect 1715 13364 1716 13428
rect 1780 13364 1781 13428
rect 1715 13363 1781 13364
rect 1347 8804 1413 8805
rect 1347 8740 1348 8804
rect 1412 8740 1413 8804
rect 1347 8739 1413 8740
rect 1350 6629 1410 8739
rect 2083 8532 2149 8533
rect 2083 8468 2084 8532
rect 2148 8468 2149 8532
rect 2083 8467 2149 8468
rect 1347 6628 1413 6629
rect 1347 6564 1348 6628
rect 1412 6564 1413 6628
rect 1347 6563 1413 6564
rect 2086 4861 2146 8467
rect 2083 4860 2149 4861
rect 2083 4796 2084 4860
rect 2148 4796 2149 4860
rect 2083 4795 2149 4796
rect 2454 4317 2514 16530
rect 2638 13973 2698 19347
rect 3543 19072 3863 20096
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 7419 20228 7485 20229
rect 7419 20164 7420 20228
rect 7484 20164 7485 20228
rect 7419 20163 7485 20164
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 4107 19412 4173 19413
rect 4107 19348 4108 19412
rect 4172 19348 4173 19412
rect 4107 19347 4173 19348
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3371 18188 3437 18189
rect 3371 18124 3372 18188
rect 3436 18124 3437 18188
rect 3371 18123 3437 18124
rect 3374 15605 3434 18123
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3371 15604 3437 15605
rect 3371 15540 3372 15604
rect 3436 15540 3437 15604
rect 3371 15539 3437 15540
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 2635 13972 2701 13973
rect 2635 13908 2636 13972
rect 2700 13908 2701 13972
rect 2635 13907 2701 13908
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 4110 12450 4170 19347
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 4475 12476 4541 12477
rect 4110 12390 4354 12450
rect 4475 12412 4476 12476
rect 4540 12412 4541 12476
rect 4475 12411 4541 12412
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 2635 8804 2701 8805
rect 2635 8740 2636 8804
rect 2700 8740 2701 8804
rect 2635 8739 2701 8740
rect 2451 4316 2517 4317
rect 2451 4252 2452 4316
rect 2516 4252 2517 4316
rect 2451 4251 2517 4252
rect 2454 3770 2514 4251
rect 2638 3773 2698 8739
rect 3543 8192 3863 9216
rect 4107 8260 4173 8261
rect 4107 8196 4108 8260
rect 4172 8196 4173 8260
rect 4107 8195 4173 8196
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3371 5404 3437 5405
rect 3371 5340 3372 5404
rect 3436 5340 3437 5404
rect 3371 5339 3437 5340
rect 2050 3710 2514 3770
rect 2635 3772 2701 3773
rect 2635 3708 2636 3772
rect 2700 3708 2701 3772
rect 2635 3707 2701 3708
rect 2638 3229 2698 3707
rect 2635 3228 2701 3229
rect 2635 3164 2636 3228
rect 2700 3164 2701 3228
rect 2635 3163 2701 3164
rect 3374 2957 3434 5339
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 4110 4861 4170 8195
rect 4294 7717 4354 12390
rect 4291 7716 4357 7717
rect 4291 7652 4292 7716
rect 4356 7652 4357 7716
rect 4291 7651 4357 7652
rect 4294 7037 4354 7651
rect 4291 7036 4357 7037
rect 4291 6972 4292 7036
rect 4356 6972 4357 7036
rect 4291 6971 4357 6972
rect 4478 5269 4538 12411
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 5579 11524 5645 11525
rect 5579 11460 5580 11524
rect 5644 11460 5645 11524
rect 5579 11459 5645 11460
rect 5211 10980 5277 10981
rect 5211 10916 5212 10980
rect 5276 10916 5277 10980
rect 5211 10915 5277 10916
rect 5214 5949 5274 10915
rect 5395 9076 5461 9077
rect 5395 9012 5396 9076
rect 5460 9012 5461 9076
rect 5395 9011 5461 9012
rect 5398 7173 5458 9011
rect 5395 7172 5461 7173
rect 5395 7108 5396 7172
rect 5460 7108 5461 7172
rect 5395 7107 5461 7108
rect 5211 5948 5277 5949
rect 5211 5884 5212 5948
rect 5276 5884 5277 5948
rect 5211 5883 5277 5884
rect 4475 5268 4541 5269
rect 4475 5204 4476 5268
rect 4540 5204 4541 5268
rect 4475 5203 4541 5204
rect 4107 4860 4173 4861
rect 4107 4796 4108 4860
rect 4172 4796 4173 4860
rect 4107 4795 4173 4796
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3371 2956 3437 2957
rect 3371 2892 3372 2956
rect 3436 2892 3437 2956
rect 3371 2891 3437 2892
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 4110 2685 4170 4795
rect 5582 2685 5642 11459
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 5763 10028 5829 10029
rect 5763 9964 5764 10028
rect 5828 9964 5829 10028
rect 5763 9963 5829 9964
rect 5766 3909 5826 9963
rect 6142 9824 6462 10848
rect 6683 10028 6749 10029
rect 6683 9964 6684 10028
rect 6748 9964 6749 10028
rect 6683 9963 6749 9964
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 5947 9348 6013 9349
rect 5947 9284 5948 9348
rect 6012 9284 6013 9348
rect 5947 9283 6013 9284
rect 5763 3908 5829 3909
rect 5763 3844 5764 3908
rect 5828 3844 5829 3908
rect 5763 3843 5829 3844
rect 5950 3229 6010 9283
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6686 4997 6746 9963
rect 7422 5133 7482 20163
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 12939 19820 13005 19821
rect 12939 19756 12940 19820
rect 13004 19756 13005 19820
rect 12939 19755 13005 19756
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 12755 19412 12821 19413
rect 12755 19348 12756 19412
rect 12820 19348 12821 19412
rect 12755 19347 12821 19348
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 12758 17917 12818 19347
rect 12755 17916 12821 17917
rect 12755 17852 12756 17916
rect 12820 17852 12821 17916
rect 12755 17851 12821 17852
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 10547 14516 10613 14517
rect 10547 14452 10548 14516
rect 10612 14452 10613 14516
rect 10547 14451 10613 14452
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 9443 11388 9509 11389
rect 9443 11324 9444 11388
rect 9508 11324 9509 11388
rect 9443 11323 9509 11324
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8523 8804 8589 8805
rect 8523 8740 8524 8804
rect 8588 8740 8589 8804
rect 8523 8739 8589 8740
rect 8339 8396 8405 8397
rect 8339 8332 8340 8396
rect 8404 8332 8405 8396
rect 8339 8331 8405 8332
rect 7419 5132 7485 5133
rect 7419 5130 7420 5132
rect 7238 5070 7420 5130
rect 6683 4996 6749 4997
rect 6683 4932 6684 4996
rect 6748 4932 6749 4996
rect 6683 4931 6749 4932
rect 6686 4453 6746 4931
rect 6683 4452 6749 4453
rect 6683 4388 6684 4452
rect 6748 4388 6749 4452
rect 6683 4387 6749 4388
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 5947 3228 6013 3229
rect 5947 3164 5948 3228
rect 6012 3164 6013 3228
rect 5947 3163 6013 3164
rect 4107 2684 4173 2685
rect 4107 2620 4108 2684
rect 4172 2620 4173 2684
rect 4107 2619 4173 2620
rect 5579 2684 5645 2685
rect 5579 2620 5580 2684
rect 5644 2620 5645 2684
rect 5579 2619 5645 2620
rect 6142 2208 6462 3232
rect 6686 2685 6746 4387
rect 7238 4045 7298 5070
rect 7419 5068 7420 5070
rect 7484 5068 7485 5132
rect 7419 5067 7485 5068
rect 8342 4317 8402 8331
rect 8339 4316 8405 4317
rect 8339 4252 8340 4316
rect 8404 4252 8405 4316
rect 8339 4251 8405 4252
rect 7235 4044 7301 4045
rect 7235 3980 7236 4044
rect 7300 3980 7301 4044
rect 7235 3979 7301 3980
rect 8526 3365 8586 8739
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 9259 7172 9325 7173
rect 9259 7108 9260 7172
rect 9324 7108 9325 7172
rect 9259 7107 9325 7108
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8523 3364 8589 3365
rect 8523 3300 8524 3364
rect 8588 3300 8589 3364
rect 8523 3299 8589 3300
rect 8741 2752 9061 3776
rect 9262 2821 9322 7107
rect 9259 2820 9325 2821
rect 9259 2756 9260 2820
rect 9324 2756 9325 2820
rect 9259 2755 9325 2756
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 6683 2684 6749 2685
rect 6683 2620 6684 2684
rect 6748 2620 6749 2684
rect 6683 2619 6749 2620
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 2128 9061 2688
rect 9446 2685 9506 11323
rect 10363 9756 10429 9757
rect 10363 9692 10364 9756
rect 10428 9692 10429 9756
rect 10363 9691 10429 9692
rect 10366 2685 10426 9691
rect 10550 5405 10610 14451
rect 11340 14176 11660 15200
rect 12942 14245 13002 19755
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 12939 14244 13005 14245
rect 12939 14180 12940 14244
rect 13004 14180 13005 14244
rect 12939 14179 13005 14180
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 10915 13972 10981 13973
rect 10915 13908 10916 13972
rect 10980 13908 10981 13972
rect 10915 13907 10981 13908
rect 10547 5404 10613 5405
rect 10547 5340 10548 5404
rect 10612 5340 10613 5404
rect 10547 5339 10613 5340
rect 10731 5268 10797 5269
rect 10731 5204 10732 5268
rect 10796 5204 10797 5268
rect 10731 5203 10797 5204
rect 10734 4453 10794 5203
rect 10731 4452 10797 4453
rect 10731 4388 10732 4452
rect 10796 4388 10797 4452
rect 10731 4387 10797 4388
rect 10918 4045 10978 13907
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 12019 9620 12085 9621
rect 12019 9556 12020 9620
rect 12084 9556 12085 9620
rect 12019 9555 12085 9556
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 10915 4044 10981 4045
rect 10915 3980 10916 4044
rect 10980 3980 10981 4044
rect 10915 3979 10981 3980
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 9443 2684 9509 2685
rect 9443 2620 9444 2684
rect 9508 2620 9509 2684
rect 9443 2619 9509 2620
rect 10363 2684 10429 2685
rect 10363 2620 10364 2684
rect 10428 2620 10429 2684
rect 10363 2619 10429 2620
rect 11340 2208 11660 3232
rect 12022 3229 12082 9555
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 15147 4316 15213 4317
rect 15147 4252 15148 4316
rect 15212 4252 15213 4316
rect 15147 4251 15213 4252
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 12019 3228 12085 3229
rect 12019 3164 12020 3228
rect 12084 3164 12085 3228
rect 12019 3163 12085 3164
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 2752 14259 3776
rect 14414 3365 14474 3622
rect 14411 3364 14477 3365
rect 14411 3300 14412 3364
rect 14476 3300 14477 3364
rect 14411 3299 14477 3300
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 15150 2549 15210 4251
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 15147 2548 15213 2549
rect 15147 2484 15148 2548
rect 15212 2484 15213 2548
rect 15147 2483 15213 2484
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
<< via4 >>
rect 2182 18732 2418 18818
rect 2182 18668 2268 18732
rect 2268 18668 2332 18732
rect 2332 18668 2418 18732
rect 2182 18582 2418 18668
rect 1630 5132 1866 5218
rect 1630 5068 1716 5132
rect 1716 5068 1780 5132
rect 1780 5068 1866 5132
rect 1630 4982 1866 5068
rect 1814 3622 2050 3858
rect 15062 18732 15298 18818
rect 15062 18668 15148 18732
rect 15148 18668 15212 18732
rect 15212 18668 15298 18732
rect 15062 18582 15298 18668
rect 15062 5132 15298 5218
rect 15062 5068 15148 5132
rect 15148 5068 15212 5132
rect 15212 5068 15298 5132
rect 15062 4982 15298 5068
rect 14326 3622 14562 3858
<< metal5 >>
rect 2140 18818 15340 18860
rect 2140 18582 2182 18818
rect 2418 18582 15062 18818
rect 15298 18582 15340 18818
rect 2140 18540 15340 18582
rect 1588 5218 15340 5260
rect 1588 4982 1630 5218
rect 1866 4982 15062 5218
rect 15298 4982 15340 5218
rect 1588 4940 15340 4982
rect 1772 3858 14604 3900
rect 1772 3622 1814 3858
rect 2050 3622 14326 3858
rect 14562 3622 14604 3858
rect 1772 3580 14604 3622
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform -1 0 16192 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1649977179
transform -1 0 16376 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1649977179
transform 1 0 16560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform 1 0 17020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1649977179
transform 1 0 17296 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A
timestamp 1649977179
transform 1 0 17848 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1649977179
transform -1 0 19044 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1649977179
transform -1 0 19504 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1649977179
transform -1 0 19964 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1649977179
transform -1 0 20424 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__A
timestamp 1649977179
transform 1 0 16376 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1649977179
transform -1 0 18492 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1649977179
transform 1 0 14168 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1649977179
transform -1 0 15640 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__A
timestamp 1649977179
transform 1 0 15272 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1649977179
transform -1 0 16376 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform -1 0 17388 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A
timestamp 1649977179
transform 1 0 17388 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1649977179
transform -1 0 18768 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A
timestamp 1649977179
transform -1 0 13984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1649977179
transform -1 0 20056 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1649977179
transform 1 0 15824 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1649977179
transform 1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1649977179
transform -1 0 14168 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 16836 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform 1 0 7360 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 9292 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 1932 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 8648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 6256 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 16192 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 11960 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 21344 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 21344 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 12420 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 12972 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 4048 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 4232 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 4140 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 3956 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 1564 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 1564 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 1932 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 3680 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 6808 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 16560 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 15272 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 11040 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 5060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 13156 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 11408 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 12420 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 4784 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 11408 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 13984 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 13800 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 12052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 13892 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 15824 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 8832 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 14904 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 5704 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 15640 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 12788 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 15088 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 16008 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 13616 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 11684 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 13800 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 9384 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 14260 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 13432 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 8372 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 8096 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 10948 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 13616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 13248 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 3956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 9384 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 14628 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 14812 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 9568 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 4416 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 16468 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 9568 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform -1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1649977179
transform -1 0 16928 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1649977179
transform -1 0 15824 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1649977179
transform -1 0 13984 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1649977179
transform -1 0 16008 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1649977179
transform -1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1649977179
transform -1 0 15088 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1649977179
transform -1 0 13340 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1649977179
transform -1 0 14168 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1649977179
transform -1 0 13984 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1649977179
transform -1 0 14996 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1649977179
transform -1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1649977179
transform -1 0 15824 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1649977179
transform -1 0 3588 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1649977179
transform -1 0 15640 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1649977179
transform -1 0 10212 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1649977179
transform -1 0 20884 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8372 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15088 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 14904 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 15640 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13800 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12880 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17940 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17756 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11684 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4416 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 4508 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 2208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 1840 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 5060 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 4140 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 4324 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14536 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 15824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12788 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12052 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 15640 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15272 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 15272 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 12604 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 7176 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 4416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8464 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 4416 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 5520 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 5428 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3404 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9016 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9200 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 8556 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9016 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9844 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10212 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7636 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 12236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13616 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13248 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 13984 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 14996 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4600 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 14444 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13432 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1649977179
transform -1 0 3680 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 9384 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 10304 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 10396 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_4__A0
timestamp 1649977179
transform -1 0 15640 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A0
timestamp 1649977179
transform -1 0 13984 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_5__A1
timestamp 1649977179
transform 1 0 12696 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15640 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15824 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 15824 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 14260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 15364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 11316 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13616 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9016 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.sky130_fd_sc_hd__buf_4_0__A
timestamp 1649977179
transform 1 0 18492 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1649977179
transform -1 0 21252 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 17756 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3220 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_158
timestamp 1649977179
transform 1 0 15640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_163
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_178
timestamp 1649977179
transform 1 0 17480 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_183
timestamp 1649977179
transform 1 0 17940 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_188
timestamp 1649977179
transform 1 0 18400 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_214
timestamp 1649977179
transform 1 0 20792 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_22
timestamp 1649977179
transform 1 0 3128 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_213 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_154
timestamp 1649977179
transform 1 0 15272 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_172
timestamp 1649977179
transform 1 0 16928 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_175
timestamp 1649977179
transform 1 0 17204 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_178 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_184
timestamp 1649977179
transform 1 0 18032 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_188 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_217
timestamp 1649977179
transform 1 0 21068 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_49
timestamp 1649977179
transform 1 0 5612 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_66
timestamp 1649977179
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_171
timestamp 1649977179
transform 1 0 16836 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_183
timestamp 1649977179
transform 1 0 17940 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_195
timestamp 1649977179
transform 1 0 19044 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_207
timestamp 1649977179
transform 1 0 20148 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_219
timestamp 1649977179
transform 1 0 21252 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_79
timestamp 1649977179
transform 1 0 8372 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_124
timestamp 1649977179
transform 1 0 12512 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_162
timestamp 1649977179
transform 1 0 16008 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_166
timestamp 1649977179
transform 1 0 16376 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_179
timestamp 1649977179
transform 1 0 17572 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_185
timestamp 1649977179
transform 1 0 18124 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 1649977179
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_66
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_100
timestamp 1649977179
transform 1 0 10304 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_127
timestamp 1649977179
transform 1 0 12788 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_154
timestamp 1649977179
transform 1 0 15272 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_158
timestamp 1649977179
transform 1 0 15640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_194
timestamp 1649977179
transform 1 0 18952 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_202
timestamp 1649977179
transform 1 0 19688 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_208
timestamp 1649977179
transform 1 0 20240 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp 1649977179
transform 1 0 21344 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_7
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_35
timestamp 1649977179
transform 1 0 4324 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_123
timestamp 1649977179
transform 1 0 12420 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_152
timestamp 1649977179
transform 1 0 15088 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_190 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18584 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_6_200
timestamp 1649977179
transform 1 0 19504 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_212
timestamp 1649977179
transform 1 0 20608 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_220
timestamp 1649977179
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_73
timestamp 1649977179
transform 1 0 7820 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_83
timestamp 1649977179
transform 1 0 8740 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_192
timestamp 1649977179
transform 1 0 18768 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_204
timestamp 1649977179
transform 1 0 19872 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_216
timestamp 1649977179
transform 1 0 20976 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_9
timestamp 1649977179
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_129
timestamp 1649977179
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_66
timestamp 1649977179
transform 1 0 7176 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_87
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_158
timestamp 1649977179
transform 1 0 15640 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1649977179
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 1649977179
transform 1 0 4600 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_100
timestamp 1649977179
transform 1 0 10304 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1649977179
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_152
timestamp 1649977179
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_170
timestamp 1649977179
transform 1 0 16744 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_182
timestamp 1649977179
transform 1 0 17848 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1649977179
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_68
timestamp 1649977179
transform 1 0 7360 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_82
timestamp 1649977179
transform 1 0 8648 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_101
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_122
timestamp 1649977179
transform 1 0 12328 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_158
timestamp 1649977179
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_6
timestamp 1649977179
transform 1 0 1656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_70
timestamp 1649977179
transform 1 0 7544 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_127
timestamp 1649977179
transform 1 0 12788 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_167
timestamp 1649977179
transform 1 0 16468 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_179
timestamp 1649977179
transform 1 0 17572 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_191
timestamp 1649977179
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_45
timestamp 1649977179
transform 1 0 5244 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_62
timestamp 1649977179
transform 1 0 6808 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_107
timestamp 1649977179
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_122
timestamp 1649977179
transform 1 0 12328 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_134
timestamp 1649977179
transform 1 0 13432 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_146
timestamp 1649977179
transform 1 0 14536 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp 1649977179
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_50
timestamp 1649977179
transform 1 0 5704 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1649977179
transform 1 0 9660 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_99
timestamp 1649977179
transform 1 0 10212 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_102
timestamp 1649977179
transform 1 0 10488 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_152
timestamp 1649977179
transform 1 0 15088 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_164
timestamp 1649977179
transform 1 0 16192 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_176
timestamp 1649977179
transform 1 0 17296 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_188
timestamp 1649977179
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_73
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_79
timestamp 1649977179
transform 1 0 8372 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_98
timestamp 1649977179
transform 1 0 10120 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_108
timestamp 1649977179
transform 1 0 11040 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_115
timestamp 1649977179
transform 1 0 11684 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_119
timestamp 1649977179
transform 1 0 12052 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_157
timestamp 1649977179
transform 1 0 15548 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 1649977179
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_37
timestamp 1649977179
transform 1 0 4508 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_120
timestamp 1649977179
transform 1 0 12144 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_143
timestamp 1649977179
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_164
timestamp 1649977179
transform 1 0 16192 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_176
timestamp 1649977179
transform 1 0 17296 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_188
timestamp 1649977179
transform 1 0 18400 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_71
timestamp 1649977179
transform 1 0 7636 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_138
timestamp 1649977179
transform 1 0 13800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_142
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_31
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_50
timestamp 1649977179
transform 1 0 5704 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_68
timestamp 1649977179
transform 1 0 7360 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_136
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_167
timestamp 1649977179
transform 1 0 16468 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_179
timestamp 1649977179
transform 1 0 17572 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1649977179
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_84
timestamp 1649977179
transform 1 0 8832 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_104
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1649977179
transform 1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_142
timestamp 1649977179
transform 1 0 14168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_6
timestamp 1649977179
transform 1 0 1656 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_33
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_87
timestamp 1649977179
transform 1 0 9108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 1649977179
transform 1 0 9384 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1649977179
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_162
timestamp 1649977179
transform 1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_181
timestamp 1649977179
transform 1 0 17756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1649977179
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_14
timestamp 1649977179
transform 1 0 2392 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_99
timestamp 1649977179
transform 1 0 10212 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_115
timestamp 1649977179
transform 1 0 11684 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 1649977179
transform 1 0 12420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_140
timestamp 1649977179
transform 1 0 13984 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_146
timestamp 1649977179
transform 1 0 14536 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_156
timestamp 1649977179
transform 1 0 15456 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_162
timestamp 1649977179
transform 1 0 16008 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_35
timestamp 1649977179
transform 1 0 4324 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_47
timestamp 1649977179
transform 1 0 5428 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1649977179
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_90
timestamp 1649977179
transform 1 0 9384 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_100
timestamp 1649977179
transform 1 0 10304 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_112
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_122
timestamp 1649977179
transform 1 0 12328 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_128
timestamp 1649977179
transform 1 0 12880 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_145
timestamp 1649977179
transform 1 0 14444 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_171
timestamp 1649977179
transform 1 0 16836 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_183
timestamp 1649977179
transform 1 0 17940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_76
timestamp 1649977179
transform 1 0 8096 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_158
timestamp 1649977179
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 1649977179
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_40
timestamp 1649977179
transform 1 0 4784 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_44
timestamp 1649977179
transform 1 0 5152 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_92
timestamp 1649977179
transform 1 0 9568 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_100
timestamp 1649977179
transform 1 0 10304 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1649977179
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_26
timestamp 1649977179
transform 1 0 3496 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_46
timestamp 1649977179
transform 1 0 5336 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_122
timestamp 1649977179
transform 1 0 12328 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_139
timestamp 1649977179
transform 1 0 13892 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_151
timestamp 1649977179
transform 1 0 14996 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_163
timestamp 1649977179
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_87
timestamp 1649977179
transform 1 0 9108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_123
timestamp 1649977179
transform 1 0 12420 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1649977179
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_149
timestamp 1649977179
transform 1 0 14812 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_161
timestamp 1649977179
transform 1 0 15916 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_173
timestamp 1649977179
transform 1 0 17020 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_185
timestamp 1649977179
transform 1 0 18124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1649977179
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_11
timestamp 1649977179
transform 1 0 2116 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_127
timestamp 1649977179
transform 1 0 12788 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_134
timestamp 1649977179
transform 1 0 13432 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_146
timestamp 1649977179
transform 1 0 14536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_158
timestamp 1649977179
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1649977179
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_61
timestamp 1649977179
transform 1 0 6716 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_108
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_142
timestamp 1649977179
transform 1 0 14168 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_154
timestamp 1649977179
transform 1 0 15272 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1649977179
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_38
timestamp 1649977179
transform 1 0 4600 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_43
timestamp 1649977179
transform 1 0 5060 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_79
timestamp 1649977179
transform 1 0 8372 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_151
timestamp 1649977179
transform 1 0 14996 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_163
timestamp 1649977179
transform 1 0 16100 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_175
timestamp 1649977179
transform 1 0 17204 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1649977179
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_98
timestamp 1649977179
transform 1 0 10120 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 1649977179
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_183
timestamp 1649977179
transform 1 0 17940 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_194
timestamp 1649977179
transform 1 0 18952 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_206
timestamp 1649977179
transform 1 0 20056 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_218
timestamp 1649977179
transform 1 0 21160 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_222
timestamp 1649977179
transform 1 0 21528 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_23
timestamp 1649977179
transform 1 0 3220 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_48
timestamp 1649977179
transform 1 0 5520 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1649977179
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_200
timestamp 1649977179
transform 1 0 19504 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_206
timestamp 1649977179
transform 1 0 20056 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_212
timestamp 1649977179
transform 1 0 20608 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_65
timestamp 1649977179
transform 1 0 7084 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_135
timestamp 1649977179
transform 1 0 13524 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_145
timestamp 1649977179
transform 1 0 14444 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_150
timestamp 1649977179
transform 1 0 14904 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_155
timestamp 1649977179
transform 1 0 15364 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_160
timestamp 1649977179
transform 1 0 15824 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_185
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_190
timestamp 1649977179
transform 1 0 18584 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_195
timestamp 1649977179
transform 1 0 19044 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_210
timestamp 1649977179
transform 1 0 20424 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_215
timestamp 1649977179
transform 1 0 20884 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _066_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1649977179
transform 1 0 2116 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1649977179
transform 1 0 1840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1649977179
transform 1 0 1840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform 1 0 2392 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform 1 0 1840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform 1 0 2116 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform 1 0 1840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform 1 0 2944 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform 1 0 3220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform 1 0 2392 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform 1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform -1 0 2944 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform 1 0 3220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform 1 0 6624 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform 1 0 3128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform -1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform -1 0 13708 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform -1 0 15732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform 1 0 15732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform -1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform -1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform -1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform -1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform -1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform -1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 19320 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform -1 0 19780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform -1 0 20240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform -1 0 20700 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform -1 0 16560 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform -1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform -1 0 13616 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform -1 0 13616 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform -1 0 13892 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1649977179
transform -1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 14904 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1649977179
transform -1 0 15180 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1649977179
transform -1 0 15456 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1649977179
transform -1 0 15916 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1649977179
transform -1 0 16192 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1649977179
transform -1 0 17204 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1649977179
transform -1 0 17756 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1649977179
transform -1 0 18032 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1649977179
transform -1 0 18308 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1649977179
transform -1 0 18584 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1649977179
transform -1 0 13340 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1649977179
transform -1 0 19504 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1649977179
transform -1 0 19872 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1649977179
transform -1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1649977179
transform -1 0 14628 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1649977179
transform -1 0 13892 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11408 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 10396 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 10396 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8832 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1649977179
transform 1 0 10672 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1649977179
transform 1 0 15732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1649977179
transform 1 0 3496 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1649977179
transform -1 0 16284 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1649977179
transform 1 0 2944 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1649977179
transform -1 0 2944 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1649977179
transform 1 0 9752 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1649977179
transform 1 0 6992 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1649977179
transform 1 0 6624 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1649977179
transform 1 0 15732 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1649977179
transform 1 0 5244 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1649977179
transform -1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1649977179
transform 1 0 7912 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1649977179
transform 1 0 13892 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1649977179
transform 1 0 7912 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1649977179
transform 1 0 13524 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1649977179
transform 1 0 8832 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1649977179
transform -1 0 8832 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1649977179
transform 1 0 12052 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1649977179
transform 1 0 5520 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1649977179
transform -1 0 2116 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1649977179
transform 1 0 12604 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1649977179
transform 1 0 15548 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1649977179
transform 1 0 7176 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1649977179
transform 1 0 18032 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1649977179
transform -1 0 5980 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1649977179
transform -1 0 6256 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1649977179
transform 1 0 1472 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1649977179
transform -1 0 2116 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1649977179
transform 1 0 5428 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1649977179
transform -1 0 5336 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1649977179
transform -1 0 8188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1649977179
transform -1 0 2116 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 8372 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 7360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 3680 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 3680 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform 1 0 21344 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 21344 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 2208 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 1932 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform -1 0 1656 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 3588 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 4784 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 5244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform -1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 4324 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 1932 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform -1 0 1932 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 10028 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input34
timestamp 1649977179
transform -1 0 10580 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1649977179
transform -1 0 9660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1649977179
transform -1 0 11040 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1649977179
transform -1 0 12420 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input40
timestamp 1649977179
transform -1 0 13340 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform 1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform 1 0 7544 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform 1 0 4692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1649977179
transform -1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1649977179
transform -1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform -1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform -1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1649977179
transform -1 0 8832 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform -1 0 2760 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1649977179
transform -1 0 8832 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform 1 0 8924 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1649977179
transform -1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1649977179
transform -1 0 10764 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input56
timestamp 1649977179
transform -1 0 10580 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform 1 0 9200 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1649977179
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1649977179
transform 1 0 12420 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input60
timestamp 1649977179
transform -1 0 13156 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform 1 0 12788 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1649977179
transform -1 0 5060 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1649977179
transform -1 0 3680 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1649977179
transform -1 0 3680 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1649977179
transform -1 0 5060 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1649977179
transform 1 0 5888 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input70
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input71
timestamp 1649977179
transform -1 0 7084 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1649977179
transform 1 0 6164 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1649977179
transform -1 0 3220 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1649977179
transform 1 0 1564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input77
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input79
timestamp 1649977179
transform -1 0 2300 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp 1649977179
transform -1 0 3220 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input81
timestamp 1649977179
transform -1 0 2300 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1649977179
transform -1 0 3220 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input83
timestamp 1649977179
transform -1 0 3036 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1649977179
transform -1 0 3220 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input85
timestamp 1649977179
transform -1 0 4692 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1649977179
transform -1 0 2760 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1649977179
transform 1 0 21344 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13708 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9568 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10396 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10028 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8556 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4784 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6164 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7268 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7360 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9200 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11040 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12512 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13984 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12512 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 13340 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12696 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14168 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15272 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15640 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18584 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3312 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 1840 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2392 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3404 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 2944 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 3312 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3588 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 2852 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 1932 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3128 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 1932 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3220 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6164 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 6256 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4784 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4784 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4600 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8372 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5244 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4048 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5520 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3680 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4048 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 5520 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7820 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 3864 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4968 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6440 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6900 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8372 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9844 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13248 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10580 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12420 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10396 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10120 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8556 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8372 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4600 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4048 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6256 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 6624 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4232 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6164 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17756 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9384 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4784 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 5888 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7360 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9200 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11960 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12328 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9844 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12420 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16008 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 15732 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16192 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10672 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12144 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 14536 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7176 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10120 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9200 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12328 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform -1 0 11500 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform -1 0 11408 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 11408 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 10120 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l2_in_3__175 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 10304 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1649977179
transform -1 0 10856 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 10948 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10120 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1649977179
transform -1 0 10672 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7912 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7544 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8096 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1649977179
transform -1 0 5428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_3.mux_l2_in_3__178
timestamp 1649977179
transform 1 0 8188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1649977179
transform -1 0 6164 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7636 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6716 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10580 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10580 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1649977179
transform -1 0 7360 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1649977179
transform -1 0 7912 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_4_
timestamp 1649977179
transform -1 0 8096 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_5_
timestamp 1649977179
transform 1 0 8096 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_6_
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7912 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1649977179
transform -1 0 8740 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l2_in_3__180
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 9752 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 9752 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 9752 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1649977179
transform -1 0 12880 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13432 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14260 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 13432 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_3__181
timestamp 1649977179
transform -1 0 13984 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 15640 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13708 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1649977179
transform -1 0 14536 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform -1 0 12788 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13892 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_17.mux_l1_in_3__176
timestamp 1649977179
transform -1 0 14536 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_3_
timestamp 1649977179
transform -1 0 14904 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14812 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14904 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15732 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15640 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18124 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1649977179
transform -1 0 12604 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13800 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16560 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l2_in_1__177
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17296 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17572 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_33.mux_l2_in_1__179
timestamp 1649977179
transform 1 0 4140 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3312 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3588 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3680 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2392 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_1.mux_l1_in_3__182
timestamp 1649977179
transform 1 0 3220 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1649977179
transform -1 0 2392 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2760 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2024 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 1932 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1932 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 4508 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2576 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_3.mux_l1_in_3__159
timestamp 1649977179
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 2852 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2576 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2760 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3772 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4416 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_5.mux_l1_in_3__165
timestamp 1649977179
transform 1 0 3220 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1649977179
transform -1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2852 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 4416 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 2944 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6256 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5428 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_7.mux_l1_in_3__166
timestamp 1649977179
transform -1 0 6256 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_3_
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1649977179
transform -1 0 4692 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4692 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4784 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_9.mux_l2_in_1__167
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5336 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7636 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7360 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_11.mux_l2_in_1__183
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5060 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2392 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5244 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4416 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_13.mux_l2_in_1__184
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4048 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3220 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8188 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7360 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_15.mux_l2_in_1__185
timestamp 1649977179
transform 1 0 7820 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6532 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8188 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_17.mux_l1_in_1__153
timestamp 1649977179
transform -1 0 3864 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1649977179
transform -1 0 4784 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4048 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2116 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7452 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_19.mux_l1_in_1__154
timestamp 1649977179
transform -1 0 6900 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6808 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2944 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9568 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_21.mux_l1_in_1__155
timestamp 1649977179
transform 1 0 9752 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_1_
timestamp 1649977179
transform -1 0 9752 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9016 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11592 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_23.mux_l1_in_1__156
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11224 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10304 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3496 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11684 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10580 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_25.mux_l1_in_1__157
timestamp 1649977179
transform 1 0 11132 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10580 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10488 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9844 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_29.mux_l2_in_0__158
timestamp 1649977179
transform -1 0 8924 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 8372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7268 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_31.mux_l2_in_0__160
timestamp 1649977179
transform -1 0 3312 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6440 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2300 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_33.mux_l2_in_0__161
timestamp 1649977179
transform 1 0 9476 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2668 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5612 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5060 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_35.mux_l2_in_0__162
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2944 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4416 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_37.mux_l2_in_0__163
timestamp 1649977179
transform -1 0 3036 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2484 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3864 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_39.mux_l2_in_0__164
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3036 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3128 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8004 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9384 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12788 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7728 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8004 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 5060 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_0.mux_l2_in_3__168
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5428 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7084 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 5888 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 7360 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13064 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9568 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9660 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10488 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 12788 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1649977179
transform -1 0 13616 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_2.mux_l2_in_3__170
timestamp 1649977179
transform -1 0 11960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10396 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12788 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 12788 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12788 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11500 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10304 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 10580 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_3_
timestamp 1649977179
transform -1 0 9844 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_4_
timestamp 1649977179
transform 1 0 14628 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_5_
timestamp 1649977179
transform -1 0 13800 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_6_
timestamp 1649977179
transform -1 0 13800 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11224 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 11224 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13800 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_4.mux_l2_in_3__173
timestamp 1649977179
transform -1 0 12696 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1649977179
transform -1 0 13616 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 13616 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13432 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16008 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15456 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15824 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 15088 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_8.mux_l2_in_3__174
timestamp 1649977179
transform -1 0 14720 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1649977179
transform -1 0 15364 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15088 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 15732 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14260 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14812 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12144 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13064 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_16.mux_l1_in_3__169
timestamp 1649977179
transform 1 0 11776 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_3_
timestamp 1649977179
transform -1 0 12236 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12328 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13064 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15272 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8740 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10212 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1649977179
transform -1 0 6624 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_24.mux_l1_in_3__171
timestamp 1649977179
transform 1 0 7360 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_3_
timestamp 1649977179
transform -1 0 6256 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8464 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7084 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8556 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16928 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9292 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9200 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1649977179
transform -1 0 10028 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9568 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10120 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_32.mux_l2_in_1__172
timestamp 1649977179
transform -1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10396 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18952 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output88 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 2484 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 2116 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 2116 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 2852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 2852 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform 1 0 3220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 2116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 2116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 2484 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform -1 0 2116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform 1 0 18032 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform 1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform 1 0 20424 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform 1 0 20884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1649977179
transform 1 0 21252 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform 1 0 21252 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform 1 0 20884 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform -1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform -1 0 15640 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform 1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform -1 0 13524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform 1 0 18216 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1649977179
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1649977179
transform 1 0 20056 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1649977179
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1649977179
transform 1 0 20976 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1649977179
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1649977179
transform 1 0 20884 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1649977179
transform 1 0 13616 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1649977179
transform 1 0 14536 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1649977179
transform 1 0 15456 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1649977179
transform 1 0 17388 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17480 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater149
timestamp 1649977179
transform -1 0 11316 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater150
timestamp 1649977179
transform 1 0 13616 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater151
timestamp 1649977179
transform -1 0 8832 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater152
timestamp 1649977179
transform -1 0 9108 0 -1 7616
box -38 -48 406 592
<< labels >>
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 0 nsew ground input
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 0 nsew ground input
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 0 nsew ground input
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 1 nsew power input
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 1 nsew power input
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 1 nsew power input
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 1 nsew power input
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 2 nsew signal input
rlabel metal2 s 662 0 718 800 6 bottom_left_grid_pin_43_
port 3 nsew signal input
rlabel metal2 s 1122 0 1178 800 6 bottom_left_grid_pin_44_
port 4 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 bottom_left_grid_pin_45_
port 5 nsew signal input
rlabel metal2 s 2042 0 2098 800 6 bottom_left_grid_pin_46_
port 6 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 bottom_left_grid_pin_47_
port 7 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 bottom_left_grid_pin_48_
port 8 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 bottom_left_grid_pin_49_
port 9 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 bottom_right_grid_pin_1_
port 10 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 ccff_head
port 11 nsew signal input
rlabel metal3 s 22200 17144 23000 17264 6 ccff_tail
port 12 nsew signal tristate
rlabel metal3 s 0 3952 800 4072 6 chanx_left_in[0]
port 13 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 chanx_left_in[10]
port 14 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 chanx_left_in[11]
port 15 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[12]
port 16 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 chanx_left_in[13]
port 17 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 chanx_left_in[14]
port 18 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 chanx_left_in[15]
port 19 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 chanx_left_in[16]
port 20 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 chanx_left_in[17]
port 21 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 chanx_left_in[18]
port 22 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 chanx_left_in[19]
port 23 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[1]
port 24 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 chanx_left_in[2]
port 25 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 chanx_left_in[3]
port 26 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 chanx_left_in[4]
port 27 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 chanx_left_in[5]
port 28 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 chanx_left_in[6]
port 29 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 chanx_left_in[7]
port 30 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 chanx_left_in[8]
port 31 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 chanx_left_in[9]
port 32 nsew signal input
rlabel metal3 s 0 13472 800 13592 6 chanx_left_out[0]
port 33 nsew signal tristate
rlabel metal3 s 0 18232 800 18352 6 chanx_left_out[10]
port 34 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[11]
port 35 nsew signal tristate
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[12]
port 36 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[13]
port 37 nsew signal tristate
rlabel metal3 s 0 20136 800 20256 6 chanx_left_out[14]
port 38 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[15]
port 39 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 chanx_left_out[16]
port 40 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[17]
port 41 nsew signal tristate
rlabel metal3 s 0 22040 800 22160 6 chanx_left_out[18]
port 42 nsew signal tristate
rlabel metal3 s 0 22584 800 22704 6 chanx_left_out[19]
port 43 nsew signal tristate
rlabel metal3 s 0 14016 800 14136 6 chanx_left_out[1]
port 44 nsew signal tristate
rlabel metal3 s 0 14424 800 14544 6 chanx_left_out[2]
port 45 nsew signal tristate
rlabel metal3 s 0 14968 800 15088 6 chanx_left_out[3]
port 46 nsew signal tristate
rlabel metal3 s 0 15376 800 15496 6 chanx_left_out[4]
port 47 nsew signal tristate
rlabel metal3 s 0 15920 800 16040 6 chanx_left_out[5]
port 48 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 chanx_left_out[6]
port 49 nsew signal tristate
rlabel metal3 s 0 16872 800 16992 6 chanx_left_out[7]
port 50 nsew signal tristate
rlabel metal3 s 0 17280 800 17400 6 chanx_left_out[8]
port 51 nsew signal tristate
rlabel metal3 s 0 17824 800 17944 6 chanx_left_out[9]
port 52 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 chany_bottom_in[0]
port 53 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[10]
port 54 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 chany_bottom_in[11]
port 55 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[12]
port 56 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[13]
port 57 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[14]
port 58 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 chany_bottom_in[15]
port 59 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[16]
port 60 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[17]
port 61 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_in[18]
port 62 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 chany_bottom_in[19]
port 63 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 chany_bottom_in[1]
port 64 nsew signal input
rlabel metal2 s 4894 0 4950 800 6 chany_bottom_in[2]
port 65 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 chany_bottom_in[3]
port 66 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 chany_bottom_in[4]
port 67 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 chany_bottom_in[5]
port 68 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 chany_bottom_in[6]
port 69 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 chany_bottom_in[7]
port 70 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[8]
port 71 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[9]
port 72 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[0]
port 73 nsew signal tristate
rlabel metal2 s 17958 0 18014 800 6 chany_bottom_out[10]
port 74 nsew signal tristate
rlabel metal2 s 18418 0 18474 800 6 chany_bottom_out[11]
port 75 nsew signal tristate
rlabel metal2 s 18970 0 19026 800 6 chany_bottom_out[12]
port 76 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 chany_bottom_out[13]
port 77 nsew signal tristate
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_out[14]
port 78 nsew signal tristate
rlabel metal2 s 20350 0 20406 800 6 chany_bottom_out[15]
port 79 nsew signal tristate
rlabel metal2 s 20810 0 20866 800 6 chany_bottom_out[16]
port 80 nsew signal tristate
rlabel metal2 s 21270 0 21326 800 6 chany_bottom_out[17]
port 81 nsew signal tristate
rlabel metal2 s 21730 0 21786 800 6 chany_bottom_out[18]
port 82 nsew signal tristate
rlabel metal2 s 22190 0 22246 800 6 chany_bottom_out[19]
port 83 nsew signal tristate
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_out[1]
port 84 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 chany_bottom_out[2]
port 85 nsew signal tristate
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_out[3]
port 86 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_out[4]
port 87 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_out[5]
port 88 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 chany_bottom_out[6]
port 89 nsew signal tristate
rlabel metal2 s 16578 0 16634 800 6 chany_bottom_out[7]
port 90 nsew signal tristate
rlabel metal2 s 17038 0 17094 800 6 chany_bottom_out[8]
port 91 nsew signal tristate
rlabel metal2 s 17498 0 17554 800 6 chany_bottom_out[9]
port 92 nsew signal tristate
rlabel metal2 s 3882 22200 3938 23000 6 chany_top_in[0]
port 93 nsew signal input
rlabel metal2 s 8482 22200 8538 23000 6 chany_top_in[10]
port 94 nsew signal input
rlabel metal2 s 8942 22200 8998 23000 6 chany_top_in[11]
port 95 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[12]
port 96 nsew signal input
rlabel metal2 s 9862 22200 9918 23000 6 chany_top_in[13]
port 97 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[14]
port 98 nsew signal input
rlabel metal2 s 10782 22200 10838 23000 6 chany_top_in[15]
port 99 nsew signal input
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_in[16]
port 100 nsew signal input
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_in[17]
port 101 nsew signal input
rlabel metal2 s 12162 22200 12218 23000 6 chany_top_in[18]
port 102 nsew signal input
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_in[19]
port 103 nsew signal input
rlabel metal2 s 4342 22200 4398 23000 6 chany_top_in[1]
port 104 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[2]
port 105 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[3]
port 106 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 chany_top_in[4]
port 107 nsew signal input
rlabel metal2 s 6182 22200 6238 23000 6 chany_top_in[5]
port 108 nsew signal input
rlabel metal2 s 6642 22200 6698 23000 6 chany_top_in[6]
port 109 nsew signal input
rlabel metal2 s 7102 22200 7158 23000 6 chany_top_in[7]
port 110 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[8]
port 111 nsew signal input
rlabel metal2 s 8022 22200 8078 23000 6 chany_top_in[9]
port 112 nsew signal input
rlabel metal2 s 13082 22200 13138 23000 6 chany_top_out[0]
port 113 nsew signal tristate
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 114 nsew signal tristate
rlabel metal2 s 18142 22200 18198 23000 6 chany_top_out[11]
port 115 nsew signal tristate
rlabel metal2 s 18602 22200 18658 23000 6 chany_top_out[12]
port 116 nsew signal tristate
rlabel metal2 s 19062 22200 19118 23000 6 chany_top_out[13]
port 117 nsew signal tristate
rlabel metal2 s 19522 22200 19578 23000 6 chany_top_out[14]
port 118 nsew signal tristate
rlabel metal2 s 19982 22200 20038 23000 6 chany_top_out[15]
port 119 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[16]
port 120 nsew signal tristate
rlabel metal2 s 20902 22200 20958 23000 6 chany_top_out[17]
port 121 nsew signal tristate
rlabel metal2 s 21362 22200 21418 23000 6 chany_top_out[18]
port 122 nsew signal tristate
rlabel metal2 s 21822 22200 21878 23000 6 chany_top_out[19]
port 123 nsew signal tristate
rlabel metal2 s 13542 22200 13598 23000 6 chany_top_out[1]
port 124 nsew signal tristate
rlabel metal2 s 14002 22200 14058 23000 6 chany_top_out[2]
port 125 nsew signal tristate
rlabel metal2 s 14462 22200 14518 23000 6 chany_top_out[3]
port 126 nsew signal tristate
rlabel metal2 s 14922 22200 14978 23000 6 chany_top_out[4]
port 127 nsew signal tristate
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[5]
port 128 nsew signal tristate
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[6]
port 129 nsew signal tristate
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[7]
port 130 nsew signal tristate
rlabel metal2 s 16762 22200 16818 23000 6 chany_top_out[8]
port 131 nsew signal tristate
rlabel metal2 s 17222 22200 17278 23000 6 chany_top_out[9]
port 132 nsew signal tristate
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 133 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 134 nsew signal input
rlabel metal3 s 0 1096 800 1216 6 left_bottom_grid_pin_36_
port 135 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_37_
port 136 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 left_bottom_grid_pin_38_
port 137 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_39_
port 138 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 left_bottom_grid_pin_40_
port 139 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 140 nsew signal input
rlabel metal2 s 22282 22200 22338 23000 6 prog_clk_0_N_in
port 141 nsew signal input
rlabel metal2 s 202 22200 258 23000 6 top_left_grid_pin_42_
port 142 nsew signal input
rlabel metal2 s 662 22200 718 23000 6 top_left_grid_pin_43_
port 143 nsew signal input
rlabel metal2 s 1122 22200 1178 23000 6 top_left_grid_pin_44_
port 144 nsew signal input
rlabel metal2 s 1582 22200 1638 23000 6 top_left_grid_pin_45_
port 145 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_46_
port 146 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 top_left_grid_pin_47_
port 147 nsew signal input
rlabel metal2 s 2962 22200 3018 23000 6 top_left_grid_pin_48_
port 148 nsew signal input
rlabel metal2 s 3422 22200 3478 23000 6 top_left_grid_pin_49_
port 149 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 top_right_grid_pin_1_
port 150 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
