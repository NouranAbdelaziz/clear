magic
tech sky130A
magscale 1 2
timestamp 1650892240
<< obsli1 >>
rect 1104 2159 21896 20689
<< obsm1 >>
rect 290 2128 22710 20720
<< metal2 >>
rect 294 22200 350 23000
rect 846 22200 902 23000
rect 1398 22200 1454 23000
rect 1950 22200 2006 23000
rect 2502 22200 2558 23000
rect 3054 22200 3110 23000
rect 3606 22200 3662 23000
rect 4158 22200 4214 23000
rect 4710 22200 4766 23000
rect 5262 22200 5318 23000
rect 5814 22200 5870 23000
rect 6458 22200 6514 23000
rect 7010 22200 7066 23000
rect 7562 22200 7618 23000
rect 8114 22200 8170 23000
rect 8666 22200 8722 23000
rect 9218 22200 9274 23000
rect 9770 22200 9826 23000
rect 10322 22200 10378 23000
rect 10874 22200 10930 23000
rect 11426 22200 11482 23000
rect 12070 22200 12126 23000
rect 12622 22200 12678 23000
rect 13174 22200 13230 23000
rect 13726 22200 13782 23000
rect 14278 22200 14334 23000
rect 14830 22200 14886 23000
rect 15382 22200 15438 23000
rect 15934 22200 15990 23000
rect 16486 22200 16542 23000
rect 17038 22200 17094 23000
rect 17682 22200 17738 23000
rect 18234 22200 18290 23000
rect 18786 22200 18842 23000
rect 19338 22200 19394 23000
rect 19890 22200 19946 23000
rect 20442 22200 20498 23000
rect 20994 22200 21050 23000
rect 21546 22200 21602 23000
rect 22098 22200 22154 23000
rect 22650 22200 22706 23000
<< obsm2 >>
rect 406 22144 790 22681
rect 958 22144 1342 22681
rect 1510 22144 1894 22681
rect 2062 22144 2446 22681
rect 2614 22144 2998 22681
rect 3166 22144 3550 22681
rect 3718 22144 4102 22681
rect 4270 22144 4654 22681
rect 4822 22144 5206 22681
rect 5374 22144 5758 22681
rect 5926 22144 6402 22681
rect 6570 22144 6954 22681
rect 7122 22144 7506 22681
rect 7674 22144 8058 22681
rect 8226 22144 8610 22681
rect 8778 22144 9162 22681
rect 9330 22144 9714 22681
rect 9882 22144 10266 22681
rect 10434 22144 10818 22681
rect 10986 22144 11370 22681
rect 11538 22144 12014 22681
rect 12182 22144 12566 22681
rect 12734 22144 13118 22681
rect 13286 22144 13670 22681
rect 13838 22144 14222 22681
rect 14390 22144 14774 22681
rect 14942 22144 15326 22681
rect 15494 22144 15878 22681
rect 16046 22144 16430 22681
rect 16598 22144 16982 22681
rect 17150 22144 17626 22681
rect 17794 22144 18178 22681
rect 18346 22144 18730 22681
rect 18898 22144 19282 22681
rect 19450 22144 19834 22681
rect 20002 22144 20386 22681
rect 20554 22144 20938 22681
rect 21106 22144 21490 22681
rect 21658 22144 22042 22681
rect 22210 22144 22594 22681
rect 296 167 22704 22144
<< metal3 >>
rect 22200 22584 23000 22704
rect 22200 22176 23000 22296
rect 22200 21632 23000 21752
rect 22200 21224 23000 21344
rect 22200 20816 23000 20936
rect 22200 20272 23000 20392
rect 22200 19864 23000 19984
rect 22200 19320 23000 19440
rect 22200 18912 23000 19032
rect 22200 18504 23000 18624
rect 22200 17960 23000 18080
rect 22200 17552 23000 17672
rect 0 17144 800 17264
rect 22200 17144 23000 17264
rect 22200 16600 23000 16720
rect 22200 16192 23000 16312
rect 22200 15648 23000 15768
rect 22200 15240 23000 15360
rect 22200 14832 23000 14952
rect 22200 14288 23000 14408
rect 22200 13880 23000 14000
rect 22200 13472 23000 13592
rect 22200 12928 23000 13048
rect 22200 12520 23000 12640
rect 22200 11976 23000 12096
rect 22200 11568 23000 11688
rect 22200 11160 23000 11280
rect 22200 10616 23000 10736
rect 22200 10208 23000 10328
rect 22200 9664 23000 9784
rect 22200 9256 23000 9376
rect 22200 8848 23000 8968
rect 22200 8304 23000 8424
rect 22200 7896 23000 8016
rect 22200 7488 23000 7608
rect 22200 6944 23000 7064
rect 22200 6536 23000 6656
rect 22200 5992 23000 6112
rect 0 5720 800 5840
rect 22200 5584 23000 5704
rect 22200 5176 23000 5296
rect 22200 4632 23000 4752
rect 22200 4224 23000 4344
rect 22200 3816 23000 3936
rect 22200 3272 23000 3392
rect 22200 2864 23000 2984
rect 22200 2320 23000 2440
rect 22200 1912 23000 2032
rect 22200 1504 23000 1624
rect 22200 960 23000 1080
rect 22200 552 23000 672
rect 22200 144 23000 264
<< obsm3 >>
rect 800 22504 22120 22677
rect 800 22376 22200 22504
rect 800 22096 22120 22376
rect 800 21832 22200 22096
rect 800 21552 22120 21832
rect 800 21424 22200 21552
rect 800 21144 22120 21424
rect 800 21016 22200 21144
rect 800 20736 22120 21016
rect 800 20472 22200 20736
rect 800 20192 22120 20472
rect 800 20064 22200 20192
rect 800 19784 22120 20064
rect 800 19520 22200 19784
rect 800 19240 22120 19520
rect 800 19112 22200 19240
rect 800 18832 22120 19112
rect 800 18704 22200 18832
rect 800 18424 22120 18704
rect 800 18160 22200 18424
rect 800 17880 22120 18160
rect 800 17752 22200 17880
rect 800 17472 22120 17752
rect 800 17344 22200 17472
rect 880 17064 22120 17344
rect 800 16800 22200 17064
rect 800 16520 22120 16800
rect 800 16392 22200 16520
rect 800 16112 22120 16392
rect 800 15848 22200 16112
rect 800 15568 22120 15848
rect 800 15440 22200 15568
rect 800 15160 22120 15440
rect 800 15032 22200 15160
rect 800 14752 22120 15032
rect 800 14488 22200 14752
rect 800 14208 22120 14488
rect 800 14080 22200 14208
rect 800 13800 22120 14080
rect 800 13672 22200 13800
rect 800 13392 22120 13672
rect 800 13128 22200 13392
rect 800 12848 22120 13128
rect 800 12720 22200 12848
rect 800 12440 22120 12720
rect 800 12176 22200 12440
rect 800 11896 22120 12176
rect 800 11768 22200 11896
rect 800 11488 22120 11768
rect 800 11360 22200 11488
rect 800 11080 22120 11360
rect 800 10816 22200 11080
rect 800 10536 22120 10816
rect 800 10408 22200 10536
rect 800 10128 22120 10408
rect 800 9864 22200 10128
rect 800 9584 22120 9864
rect 800 9456 22200 9584
rect 800 9176 22120 9456
rect 800 9048 22200 9176
rect 800 8768 22120 9048
rect 800 8504 22200 8768
rect 800 8224 22120 8504
rect 800 8096 22200 8224
rect 800 7816 22120 8096
rect 800 7688 22200 7816
rect 800 7408 22120 7688
rect 800 7144 22200 7408
rect 800 6864 22120 7144
rect 800 6736 22200 6864
rect 800 6456 22120 6736
rect 800 6192 22200 6456
rect 800 5920 22120 6192
rect 880 5912 22120 5920
rect 880 5784 22200 5912
rect 880 5640 22120 5784
rect 800 5504 22120 5640
rect 800 5376 22200 5504
rect 800 5096 22120 5376
rect 800 4832 22200 5096
rect 800 4552 22120 4832
rect 800 4424 22200 4552
rect 800 4144 22120 4424
rect 800 4016 22200 4144
rect 800 3736 22120 4016
rect 800 3472 22200 3736
rect 800 3192 22120 3472
rect 800 3064 22200 3192
rect 800 2784 22120 3064
rect 800 2520 22200 2784
rect 800 2240 22120 2520
rect 800 2112 22200 2240
rect 800 1832 22120 2112
rect 800 1704 22200 1832
rect 800 1424 22120 1704
rect 800 1160 22200 1424
rect 800 880 22120 1160
rect 800 752 22200 880
rect 800 472 22120 752
rect 800 344 22200 472
rect 800 171 22120 344
<< metal4 >>
rect 3543 2128 3863 20720
rect 6142 2128 6462 20720
rect 8741 2128 9061 20720
rect 11340 2128 11660 20720
rect 13939 2128 14259 20720
rect 16538 2128 16858 20720
rect 19137 2128 19457 20720
<< obsm4 >>
rect 18643 5339 18893 19549
<< labels >>
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 1 nsew ground input
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 1 nsew ground input
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 1 nsew ground input
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 2 nsew power input
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 2 nsew power input
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 2 nsew power input
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 2 nsew power input
rlabel metal3 s 0 5720 800 5840 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 ccff_tail
port 4 nsew signal output
rlabel metal3 s 22200 4224 23000 4344 6 chanx_right_in[0]
port 5 nsew signal input
rlabel metal3 s 22200 8848 23000 8968 6 chanx_right_in[10]
port 6 nsew signal input
rlabel metal3 s 22200 9256 23000 9376 6 chanx_right_in[11]
port 7 nsew signal input
rlabel metal3 s 22200 9664 23000 9784 6 chanx_right_in[12]
port 8 nsew signal input
rlabel metal3 s 22200 10208 23000 10328 6 chanx_right_in[13]
port 9 nsew signal input
rlabel metal3 s 22200 10616 23000 10736 6 chanx_right_in[14]
port 10 nsew signal input
rlabel metal3 s 22200 11160 23000 11280 6 chanx_right_in[15]
port 11 nsew signal input
rlabel metal3 s 22200 11568 23000 11688 6 chanx_right_in[16]
port 12 nsew signal input
rlabel metal3 s 22200 11976 23000 12096 6 chanx_right_in[17]
port 13 nsew signal input
rlabel metal3 s 22200 12520 23000 12640 6 chanx_right_in[18]
port 14 nsew signal input
rlabel metal3 s 22200 12928 23000 13048 6 chanx_right_in[19]
port 15 nsew signal input
rlabel metal3 s 22200 4632 23000 4752 6 chanx_right_in[1]
port 16 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[2]
port 17 nsew signal input
rlabel metal3 s 22200 5584 23000 5704 6 chanx_right_in[3]
port 18 nsew signal input
rlabel metal3 s 22200 5992 23000 6112 6 chanx_right_in[4]
port 19 nsew signal input
rlabel metal3 s 22200 6536 23000 6656 6 chanx_right_in[5]
port 20 nsew signal input
rlabel metal3 s 22200 6944 23000 7064 6 chanx_right_in[6]
port 21 nsew signal input
rlabel metal3 s 22200 7488 23000 7608 6 chanx_right_in[7]
port 22 nsew signal input
rlabel metal3 s 22200 7896 23000 8016 6 chanx_right_in[8]
port 23 nsew signal input
rlabel metal3 s 22200 8304 23000 8424 6 chanx_right_in[9]
port 24 nsew signal input
rlabel metal3 s 22200 13472 23000 13592 6 chanx_right_out[0]
port 25 nsew signal output
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[10]
port 26 nsew signal output
rlabel metal3 s 22200 18504 23000 18624 6 chanx_right_out[11]
port 27 nsew signal output
rlabel metal3 s 22200 18912 23000 19032 6 chanx_right_out[12]
port 28 nsew signal output
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[13]
port 29 nsew signal output
rlabel metal3 s 22200 19864 23000 19984 6 chanx_right_out[14]
port 30 nsew signal output
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[15]
port 31 nsew signal output
rlabel metal3 s 22200 20816 23000 20936 6 chanx_right_out[16]
port 32 nsew signal output
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[17]
port 33 nsew signal output
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[18]
port 34 nsew signal output
rlabel metal3 s 22200 22176 23000 22296 6 chanx_right_out[19]
port 35 nsew signal output
rlabel metal3 s 22200 13880 23000 14000 6 chanx_right_out[1]
port 36 nsew signal output
rlabel metal3 s 22200 14288 23000 14408 6 chanx_right_out[2]
port 37 nsew signal output
rlabel metal3 s 22200 14832 23000 14952 6 chanx_right_out[3]
port 38 nsew signal output
rlabel metal3 s 22200 15240 23000 15360 6 chanx_right_out[4]
port 39 nsew signal output
rlabel metal3 s 22200 15648 23000 15768 6 chanx_right_out[5]
port 40 nsew signal output
rlabel metal3 s 22200 16192 23000 16312 6 chanx_right_out[6]
port 41 nsew signal output
rlabel metal3 s 22200 16600 23000 16720 6 chanx_right_out[7]
port 42 nsew signal output
rlabel metal3 s 22200 17144 23000 17264 6 chanx_right_out[8]
port 43 nsew signal output
rlabel metal3 s 22200 17552 23000 17672 6 chanx_right_out[9]
port 44 nsew signal output
rlabel metal2 s 846 22200 902 23000 6 chany_top_in[0]
port 45 nsew signal input
rlabel metal2 s 6458 22200 6514 23000 6 chany_top_in[10]
port 46 nsew signal input
rlabel metal2 s 7010 22200 7066 23000 6 chany_top_in[11]
port 47 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[12]
port 48 nsew signal input
rlabel metal2 s 8114 22200 8170 23000 6 chany_top_in[13]
port 49 nsew signal input
rlabel metal2 s 8666 22200 8722 23000 6 chany_top_in[14]
port 50 nsew signal input
rlabel metal2 s 9218 22200 9274 23000 6 chany_top_in[15]
port 51 nsew signal input
rlabel metal2 s 9770 22200 9826 23000 6 chany_top_in[16]
port 52 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[17]
port 53 nsew signal input
rlabel metal2 s 10874 22200 10930 23000 6 chany_top_in[18]
port 54 nsew signal input
rlabel metal2 s 11426 22200 11482 23000 6 chany_top_in[19]
port 55 nsew signal input
rlabel metal2 s 1398 22200 1454 23000 6 chany_top_in[1]
port 56 nsew signal input
rlabel metal2 s 1950 22200 2006 23000 6 chany_top_in[2]
port 57 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 chany_top_in[3]
port 58 nsew signal input
rlabel metal2 s 3054 22200 3110 23000 6 chany_top_in[4]
port 59 nsew signal input
rlabel metal2 s 3606 22200 3662 23000 6 chany_top_in[5]
port 60 nsew signal input
rlabel metal2 s 4158 22200 4214 23000 6 chany_top_in[6]
port 61 nsew signal input
rlabel metal2 s 4710 22200 4766 23000 6 chany_top_in[7]
port 62 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[8]
port 63 nsew signal input
rlabel metal2 s 5814 22200 5870 23000 6 chany_top_in[9]
port 64 nsew signal input
rlabel metal2 s 12070 22200 12126 23000 6 chany_top_out[0]
port 65 nsew signal output
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 66 nsew signal output
rlabel metal2 s 18234 22200 18290 23000 6 chany_top_out[11]
port 67 nsew signal output
rlabel metal2 s 18786 22200 18842 23000 6 chany_top_out[12]
port 68 nsew signal output
rlabel metal2 s 19338 22200 19394 23000 6 chany_top_out[13]
port 69 nsew signal output
rlabel metal2 s 19890 22200 19946 23000 6 chany_top_out[14]
port 70 nsew signal output
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[15]
port 71 nsew signal output
rlabel metal2 s 20994 22200 21050 23000 6 chany_top_out[16]
port 72 nsew signal output
rlabel metal2 s 21546 22200 21602 23000 6 chany_top_out[17]
port 73 nsew signal output
rlabel metal2 s 22098 22200 22154 23000 6 chany_top_out[18]
port 74 nsew signal output
rlabel metal2 s 22650 22200 22706 23000 6 chany_top_out[19]
port 75 nsew signal output
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_out[1]
port 76 nsew signal output
rlabel metal2 s 13174 22200 13230 23000 6 chany_top_out[2]
port 77 nsew signal output
rlabel metal2 s 13726 22200 13782 23000 6 chany_top_out[3]
port 78 nsew signal output
rlabel metal2 s 14278 22200 14334 23000 6 chany_top_out[4]
port 79 nsew signal output
rlabel metal2 s 14830 22200 14886 23000 6 chany_top_out[5]
port 80 nsew signal output
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[6]
port 81 nsew signal output
rlabel metal2 s 15934 22200 15990 23000 6 chany_top_out[7]
port 82 nsew signal output
rlabel metal2 s 16486 22200 16542 23000 6 chany_top_out[8]
port 83 nsew signal output
rlabel metal2 s 17038 22200 17094 23000 6 chany_top_out[9]
port 84 nsew signal output
rlabel metal3 s 22200 22584 23000 22704 6 prog_clk_0_E_in
port 85 nsew signal input
rlabel metal3 s 22200 2320 23000 2440 6 right_bottom_grid_pin_11_
port 86 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_13_
port 87 nsew signal input
rlabel metal3 s 22200 3272 23000 3392 6 right_bottom_grid_pin_15_
port 88 nsew signal input
rlabel metal3 s 22200 3816 23000 3936 6 right_bottom_grid_pin_17_
port 89 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_1_
port 90 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_3_
port 91 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_5_
port 92 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_7_
port 93 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_9_
port 94 nsew signal input
rlabel metal2 s 294 22200 350 23000 6 top_left_grid_pin_1_
port 95 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 923478
string GDS_FILE /home/karim/work/ef/clear-harden/openlane/sb_0__0_/runs/22_04_25_15_09/results/signoff/sb_0__0_.magic.gds
string GDS_START 94790
<< end >>

