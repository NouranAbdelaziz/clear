VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tie_array
  CLASS BLOCK ;
  FOREIGN tie_array ;
  ORIGIN 0.000 0.000 ;
  SIZE 60.000 BY 70.000 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 16.960 10.640 18.560 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 29.200 10.640 30.800 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 41.440 10.640 43.040 57.360 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 10.840 10.640 12.440 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.080 10.640 24.680 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 35.320 10.640 36.920 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.560 10.640 49.160 57.360 ;
    END
  END VPWR
  PIN x[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END x[0]
  PIN x[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 0.000 11.410 4.000 ;
    END
  END x[1]
  PIN x[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END x[2]
  PIN x[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END x[3]
  PIN x[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 0.000 33.950 4.000 ;
    END
  END x[4]
  PIN x[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END x[5]
  PIN x[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END x[6]
  PIN x[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END x[7]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 54.280 57.205 ;
      LAYER met1 ;
        RECT 3.750 10.640 56.050 57.360 ;
      LAYER met2 ;
        RECT 3.780 4.280 56.020 57.360 ;
        RECT 4.330 4.000 10.850 4.280 ;
        RECT 11.690 4.000 18.210 4.280 ;
        RECT 19.050 4.000 25.570 4.280 ;
        RECT 26.410 4.000 33.390 4.280 ;
        RECT 34.230 4.000 40.750 4.280 ;
        RECT 41.590 4.000 48.110 4.280 ;
        RECT 48.950 4.000 55.470 4.280 ;
      LAYER met3 ;
        RECT 10.840 10.715 49.160 57.285 ;
  END
END tie_array
END LIBRARY

